//
// by teak gui
//
// Generated on: Tue Oct 14 13:30:34 BST 2014
//


`timescale 1ns/1ps

// tko31m32_1nm1b0_2apt1o0w1bi0w31b TeakO [
//     (1,TeakOConstant 1 0),
//     (2,TeakOAppend 1 [(1,0+:1),(0,0+:31)])] [One 31,One 32]
module tko31m32_1nm1b0_2apt1o0w1bi0w31b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [30:0] i_0r0;
  input [30:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [30:0] gocomp_0;
  wire [10:0] simp331_0;
  wire tech34_int;
  wire tech35_int;
  wire tech36_int;
  wire tech37_int;
  wire tech38_int;
  wire tech39_int;
  wire tech40_int;
  wire tech41_int;
  wire tech42_int;
  wire tech43_int;
  wire [3:0] simp332_0;
  wire tech46_int;
  wire tech47_int;
  wire tech48_int;
  wire [1:0] simp333_0;
  wire tech51_int;
  wire termf_1;
  wire termt_1;
  OR2EHD I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2EHD I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2EHD I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2EHD I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2EHD I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2EHD I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2EHD I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2EHD I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2EHD I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2EHD I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2EHD I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2EHD I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2EHD I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2EHD I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2EHD I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2EHD I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2EHD I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2EHD I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2EHD I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2EHD I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2EHD I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2EHD I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2EHD I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2EHD I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2EHD I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2EHD I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2EHD I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2EHD I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2EHD I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2EHD I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2EHD I30 (gocomp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  AO222EHD I31 (tech34_int, gocomp_0[0:0], gocomp_0[1:1], tech34_int, gocomp_0[0:0], tech34_int, gocomp_0[1:1]);
  AO222EHD I32 (simp331_0[0:0], tech34_int, gocomp_0[2:2], simp331_0[0:0], tech34_int, simp331_0[0:0], gocomp_0[2:2]);
  AO222EHD I33 (tech35_int, gocomp_0[3:3], gocomp_0[4:4], tech35_int, gocomp_0[3:3], tech35_int, gocomp_0[4:4]);
  AO222EHD I34 (simp331_0[1:1], tech35_int, gocomp_0[5:5], simp331_0[1:1], tech35_int, simp331_0[1:1], gocomp_0[5:5]);
  AO222EHD I35 (tech36_int, gocomp_0[6:6], gocomp_0[7:7], tech36_int, gocomp_0[6:6], tech36_int, gocomp_0[7:7]);
  AO222EHD I36 (simp331_0[2:2], tech36_int, gocomp_0[8:8], simp331_0[2:2], tech36_int, simp331_0[2:2], gocomp_0[8:8]);
  AO222EHD I37 (tech37_int, gocomp_0[9:9], gocomp_0[10:10], tech37_int, gocomp_0[9:9], tech37_int, gocomp_0[10:10]);
  AO222EHD I38 (simp331_0[3:3], tech37_int, gocomp_0[11:11], simp331_0[3:3], tech37_int, simp331_0[3:3], gocomp_0[11:11]);
  AO222EHD I39 (tech38_int, gocomp_0[12:12], gocomp_0[13:13], tech38_int, gocomp_0[12:12], tech38_int, gocomp_0[13:13]);
  AO222EHD I40 (simp331_0[4:4], tech38_int, gocomp_0[14:14], simp331_0[4:4], tech38_int, simp331_0[4:4], gocomp_0[14:14]);
  AO222EHD I41 (tech39_int, gocomp_0[15:15], gocomp_0[16:16], tech39_int, gocomp_0[15:15], tech39_int, gocomp_0[16:16]);
  AO222EHD I42 (simp331_0[5:5], tech39_int, gocomp_0[17:17], simp331_0[5:5], tech39_int, simp331_0[5:5], gocomp_0[17:17]);
  AO222EHD I43 (tech40_int, gocomp_0[18:18], gocomp_0[19:19], tech40_int, gocomp_0[18:18], tech40_int, gocomp_0[19:19]);
  AO222EHD I44 (simp331_0[6:6], tech40_int, gocomp_0[20:20], simp331_0[6:6], tech40_int, simp331_0[6:6], gocomp_0[20:20]);
  AO222EHD I45 (tech41_int, gocomp_0[21:21], gocomp_0[22:22], tech41_int, gocomp_0[21:21], tech41_int, gocomp_0[22:22]);
  AO222EHD I46 (simp331_0[7:7], tech41_int, gocomp_0[23:23], simp331_0[7:7], tech41_int, simp331_0[7:7], gocomp_0[23:23]);
  AO222EHD I47 (tech42_int, gocomp_0[24:24], gocomp_0[25:25], tech42_int, gocomp_0[24:24], tech42_int, gocomp_0[25:25]);
  AO222EHD I48 (simp331_0[8:8], tech42_int, gocomp_0[26:26], simp331_0[8:8], tech42_int, simp331_0[8:8], gocomp_0[26:26]);
  AO222EHD I49 (tech43_int, gocomp_0[27:27], gocomp_0[28:28], tech43_int, gocomp_0[27:27], tech43_int, gocomp_0[28:28]);
  AO222EHD I50 (simp331_0[9:9], tech43_int, gocomp_0[29:29], simp331_0[9:9], tech43_int, simp331_0[9:9], gocomp_0[29:29]);
  BUFEHD I51 (simp331_0[10:10], gocomp_0[30:30]);
  AO222EHD I52 (tech46_int, simp331_0[0:0], simp331_0[1:1], tech46_int, simp331_0[0:0], tech46_int, simp331_0[1:1]);
  AO222EHD I53 (simp332_0[0:0], tech46_int, simp331_0[2:2], simp332_0[0:0], tech46_int, simp332_0[0:0], simp331_0[2:2]);
  AO222EHD I54 (tech47_int, simp331_0[3:3], simp331_0[4:4], tech47_int, simp331_0[3:3], tech47_int, simp331_0[4:4]);
  AO222EHD I55 (simp332_0[1:1], tech47_int, simp331_0[5:5], simp332_0[1:1], tech47_int, simp332_0[1:1], simp331_0[5:5]);
  AO222EHD I56 (tech48_int, simp331_0[6:6], simp331_0[7:7], tech48_int, simp331_0[6:6], tech48_int, simp331_0[7:7]);
  AO222EHD I57 (simp332_0[2:2], tech48_int, simp331_0[8:8], simp332_0[2:2], tech48_int, simp332_0[2:2], simp331_0[8:8]);
  AO222EHD I58 (simp332_0[3:3], simp331_0[9:9], simp331_0[10:10], simp332_0[3:3], simp331_0[9:9], simp332_0[3:3], simp331_0[10:10]);
  AO222EHD I59 (tech51_int, simp332_0[0:0], simp332_0[1:1], tech51_int, simp332_0[0:0], tech51_int, simp332_0[1:1]);
  AO222EHD I60 (simp333_0[0:0], tech51_int, simp332_0[2:2], simp333_0[0:0], tech51_int, simp333_0[0:0], simp332_0[2:2]);
  BUFEHD I61 (simp333_0[1:1], simp332_0[3:3]);
  AO222EHD I62 (go_0, simp333_0[0:0], simp333_0[1:1], go_0, simp333_0[0:0], go_0, simp333_0[1:1]);
  BUFEHD I63 (termf_1, go_0);
  TIE0DND I64 (termt_1);
  BUFEHD I65 (o_0r0[0:0], termf_1);
  BUFEHD I66 (o_0r0[1:1], i_0r0[0:0]);
  BUFEHD I67 (o_0r0[2:2], i_0r0[1:1]);
  BUFEHD I68 (o_0r0[3:3], i_0r0[2:2]);
  BUFEHD I69 (o_0r0[4:4], i_0r0[3:3]);
  BUFEHD I70 (o_0r0[5:5], i_0r0[4:4]);
  BUFEHD I71 (o_0r0[6:6], i_0r0[5:5]);
  BUFEHD I72 (o_0r0[7:7], i_0r0[6:6]);
  BUFEHD I73 (o_0r0[8:8], i_0r0[7:7]);
  BUFEHD I74 (o_0r0[9:9], i_0r0[8:8]);
  BUFEHD I75 (o_0r0[10:10], i_0r0[9:9]);
  BUFEHD I76 (o_0r0[11:11], i_0r0[10:10]);
  BUFEHD I77 (o_0r0[12:12], i_0r0[11:11]);
  BUFEHD I78 (o_0r0[13:13], i_0r0[12:12]);
  BUFEHD I79 (o_0r0[14:14], i_0r0[13:13]);
  BUFEHD I80 (o_0r0[15:15], i_0r0[14:14]);
  BUFEHD I81 (o_0r0[16:16], i_0r0[15:15]);
  BUFEHD I82 (o_0r0[17:17], i_0r0[16:16]);
  BUFEHD I83 (o_0r0[18:18], i_0r0[17:17]);
  BUFEHD I84 (o_0r0[19:19], i_0r0[18:18]);
  BUFEHD I85 (o_0r0[20:20], i_0r0[19:19]);
  BUFEHD I86 (o_0r0[21:21], i_0r0[20:20]);
  BUFEHD I87 (o_0r0[22:22], i_0r0[21:21]);
  BUFEHD I88 (o_0r0[23:23], i_0r0[22:22]);
  BUFEHD I89 (o_0r0[24:24], i_0r0[23:23]);
  BUFEHD I90 (o_0r0[25:25], i_0r0[24:24]);
  BUFEHD I91 (o_0r0[26:26], i_0r0[25:25]);
  BUFEHD I92 (o_0r0[27:27], i_0r0[26:26]);
  BUFEHD I93 (o_0r0[28:28], i_0r0[27:27]);
  BUFEHD I94 (o_0r0[29:29], i_0r0[28:28]);
  BUFEHD I95 (o_0r0[30:30], i_0r0[29:29]);
  BUFEHD I96 (o_0r0[31:31], i_0r0[30:30]);
  BUFEHD I97 (o_0r1[0:0], termt_1);
  BUFEHD I98 (o_0r1[1:1], i_0r1[0:0]);
  BUFEHD I99 (o_0r1[2:2], i_0r1[1:1]);
  BUFEHD I100 (o_0r1[3:3], i_0r1[2:2]);
  BUFEHD I101 (o_0r1[4:4], i_0r1[3:3]);
  BUFEHD I102 (o_0r1[5:5], i_0r1[4:4]);
  BUFEHD I103 (o_0r1[6:6], i_0r1[5:5]);
  BUFEHD I104 (o_0r1[7:7], i_0r1[6:6]);
  BUFEHD I105 (o_0r1[8:8], i_0r1[7:7]);
  BUFEHD I106 (o_0r1[9:9], i_0r1[8:8]);
  BUFEHD I107 (o_0r1[10:10], i_0r1[9:9]);
  BUFEHD I108 (o_0r1[11:11], i_0r1[10:10]);
  BUFEHD I109 (o_0r1[12:12], i_0r1[11:11]);
  BUFEHD I110 (o_0r1[13:13], i_0r1[12:12]);
  BUFEHD I111 (o_0r1[14:14], i_0r1[13:13]);
  BUFEHD I112 (o_0r1[15:15], i_0r1[14:14]);
  BUFEHD I113 (o_0r1[16:16], i_0r1[15:15]);
  BUFEHD I114 (o_0r1[17:17], i_0r1[16:16]);
  BUFEHD I115 (o_0r1[18:18], i_0r1[17:17]);
  BUFEHD I116 (o_0r1[19:19], i_0r1[18:18]);
  BUFEHD I117 (o_0r1[20:20], i_0r1[19:19]);
  BUFEHD I118 (o_0r1[21:21], i_0r1[20:20]);
  BUFEHD I119 (o_0r1[22:22], i_0r1[21:21]);
  BUFEHD I120 (o_0r1[23:23], i_0r1[22:22]);
  BUFEHD I121 (o_0r1[24:24], i_0r1[23:23]);
  BUFEHD I122 (o_0r1[25:25], i_0r1[24:24]);
  BUFEHD I123 (o_0r1[26:26], i_0r1[25:25]);
  BUFEHD I124 (o_0r1[27:27], i_0r1[26:26]);
  BUFEHD I125 (o_0r1[28:28], i_0r1[27:27]);
  BUFEHD I126 (o_0r1[29:29], i_0r1[28:28]);
  BUFEHD I127 (o_0r1[30:30], i_0r1[29:29]);
  BUFEHD I128 (o_0r1[31:31], i_0r1[30:30]);
  BUFEHD I129 (i_0a, o_0a);
endmodule

// tko31m32_1nm1b0_2api0w31bt1o0w1b TeakO [
//     (1,TeakOConstant 1 0),
//     (2,TeakOAppend 1 [(0,0+:31),(1,0+:1)])] [One 31,One 32]
module tko31m32_1nm1b0_2api0w31bt1o0w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [30:0] i_0r0;
  input [30:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [30:0] gocomp_0;
  wire [10:0] simp331_0;
  wire tech34_int;
  wire tech35_int;
  wire tech36_int;
  wire tech37_int;
  wire tech38_int;
  wire tech39_int;
  wire tech40_int;
  wire tech41_int;
  wire tech42_int;
  wire tech43_int;
  wire [3:0] simp332_0;
  wire tech46_int;
  wire tech47_int;
  wire tech48_int;
  wire [1:0] simp333_0;
  wire tech51_int;
  wire termf_1;
  wire termt_1;
  OR2EHD I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2EHD I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2EHD I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2EHD I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2EHD I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2EHD I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2EHD I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2EHD I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2EHD I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2EHD I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2EHD I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2EHD I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2EHD I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2EHD I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2EHD I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2EHD I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2EHD I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2EHD I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2EHD I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2EHD I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2EHD I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2EHD I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2EHD I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2EHD I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2EHD I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2EHD I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2EHD I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2EHD I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2EHD I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2EHD I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2EHD I30 (gocomp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  AO222EHD I31 (tech34_int, gocomp_0[0:0], gocomp_0[1:1], tech34_int, gocomp_0[0:0], tech34_int, gocomp_0[1:1]);
  AO222EHD I32 (simp331_0[0:0], tech34_int, gocomp_0[2:2], simp331_0[0:0], tech34_int, simp331_0[0:0], gocomp_0[2:2]);
  AO222EHD I33 (tech35_int, gocomp_0[3:3], gocomp_0[4:4], tech35_int, gocomp_0[3:3], tech35_int, gocomp_0[4:4]);
  AO222EHD I34 (simp331_0[1:1], tech35_int, gocomp_0[5:5], simp331_0[1:1], tech35_int, simp331_0[1:1], gocomp_0[5:5]);
  AO222EHD I35 (tech36_int, gocomp_0[6:6], gocomp_0[7:7], tech36_int, gocomp_0[6:6], tech36_int, gocomp_0[7:7]);
  AO222EHD I36 (simp331_0[2:2], tech36_int, gocomp_0[8:8], simp331_0[2:2], tech36_int, simp331_0[2:2], gocomp_0[8:8]);
  AO222EHD I37 (tech37_int, gocomp_0[9:9], gocomp_0[10:10], tech37_int, gocomp_0[9:9], tech37_int, gocomp_0[10:10]);
  AO222EHD I38 (simp331_0[3:3], tech37_int, gocomp_0[11:11], simp331_0[3:3], tech37_int, simp331_0[3:3], gocomp_0[11:11]);
  AO222EHD I39 (tech38_int, gocomp_0[12:12], gocomp_0[13:13], tech38_int, gocomp_0[12:12], tech38_int, gocomp_0[13:13]);
  AO222EHD I40 (simp331_0[4:4], tech38_int, gocomp_0[14:14], simp331_0[4:4], tech38_int, simp331_0[4:4], gocomp_0[14:14]);
  AO222EHD I41 (tech39_int, gocomp_0[15:15], gocomp_0[16:16], tech39_int, gocomp_0[15:15], tech39_int, gocomp_0[16:16]);
  AO222EHD I42 (simp331_0[5:5], tech39_int, gocomp_0[17:17], simp331_0[5:5], tech39_int, simp331_0[5:5], gocomp_0[17:17]);
  AO222EHD I43 (tech40_int, gocomp_0[18:18], gocomp_0[19:19], tech40_int, gocomp_0[18:18], tech40_int, gocomp_0[19:19]);
  AO222EHD I44 (simp331_0[6:6], tech40_int, gocomp_0[20:20], simp331_0[6:6], tech40_int, simp331_0[6:6], gocomp_0[20:20]);
  AO222EHD I45 (tech41_int, gocomp_0[21:21], gocomp_0[22:22], tech41_int, gocomp_0[21:21], tech41_int, gocomp_0[22:22]);
  AO222EHD I46 (simp331_0[7:7], tech41_int, gocomp_0[23:23], simp331_0[7:7], tech41_int, simp331_0[7:7], gocomp_0[23:23]);
  AO222EHD I47 (tech42_int, gocomp_0[24:24], gocomp_0[25:25], tech42_int, gocomp_0[24:24], tech42_int, gocomp_0[25:25]);
  AO222EHD I48 (simp331_0[8:8], tech42_int, gocomp_0[26:26], simp331_0[8:8], tech42_int, simp331_0[8:8], gocomp_0[26:26]);
  AO222EHD I49 (tech43_int, gocomp_0[27:27], gocomp_0[28:28], tech43_int, gocomp_0[27:27], tech43_int, gocomp_0[28:28]);
  AO222EHD I50 (simp331_0[9:9], tech43_int, gocomp_0[29:29], simp331_0[9:9], tech43_int, simp331_0[9:9], gocomp_0[29:29]);
  BUFEHD I51 (simp331_0[10:10], gocomp_0[30:30]);
  AO222EHD I52 (tech46_int, simp331_0[0:0], simp331_0[1:1], tech46_int, simp331_0[0:0], tech46_int, simp331_0[1:1]);
  AO222EHD I53 (simp332_0[0:0], tech46_int, simp331_0[2:2], simp332_0[0:0], tech46_int, simp332_0[0:0], simp331_0[2:2]);
  AO222EHD I54 (tech47_int, simp331_0[3:3], simp331_0[4:4], tech47_int, simp331_0[3:3], tech47_int, simp331_0[4:4]);
  AO222EHD I55 (simp332_0[1:1], tech47_int, simp331_0[5:5], simp332_0[1:1], tech47_int, simp332_0[1:1], simp331_0[5:5]);
  AO222EHD I56 (tech48_int, simp331_0[6:6], simp331_0[7:7], tech48_int, simp331_0[6:6], tech48_int, simp331_0[7:7]);
  AO222EHD I57 (simp332_0[2:2], tech48_int, simp331_0[8:8], simp332_0[2:2], tech48_int, simp332_0[2:2], simp331_0[8:8]);
  AO222EHD I58 (simp332_0[3:3], simp331_0[9:9], simp331_0[10:10], simp332_0[3:3], simp331_0[9:9], simp332_0[3:3], simp331_0[10:10]);
  AO222EHD I59 (tech51_int, simp332_0[0:0], simp332_0[1:1], tech51_int, simp332_0[0:0], tech51_int, simp332_0[1:1]);
  AO222EHD I60 (simp333_0[0:0], tech51_int, simp332_0[2:2], simp333_0[0:0], tech51_int, simp333_0[0:0], simp332_0[2:2]);
  BUFEHD I61 (simp333_0[1:1], simp332_0[3:3]);
  AO222EHD I62 (go_0, simp333_0[0:0], simp333_0[1:1], go_0, simp333_0[0:0], go_0, simp333_0[1:1]);
  BUFEHD I63 (termf_1, go_0);
  TIE0DND I64 (termt_1);
  BUFEHD I65 (o_0r0[0:0], i_0r0[0:0]);
  BUFEHD I66 (o_0r0[1:1], i_0r0[1:1]);
  BUFEHD I67 (o_0r0[2:2], i_0r0[2:2]);
  BUFEHD I68 (o_0r0[3:3], i_0r0[3:3]);
  BUFEHD I69 (o_0r0[4:4], i_0r0[4:4]);
  BUFEHD I70 (o_0r0[5:5], i_0r0[5:5]);
  BUFEHD I71 (o_0r0[6:6], i_0r0[6:6]);
  BUFEHD I72 (o_0r0[7:7], i_0r0[7:7]);
  BUFEHD I73 (o_0r0[8:8], i_0r0[8:8]);
  BUFEHD I74 (o_0r0[9:9], i_0r0[9:9]);
  BUFEHD I75 (o_0r0[10:10], i_0r0[10:10]);
  BUFEHD I76 (o_0r0[11:11], i_0r0[11:11]);
  BUFEHD I77 (o_0r0[12:12], i_0r0[12:12]);
  BUFEHD I78 (o_0r0[13:13], i_0r0[13:13]);
  BUFEHD I79 (o_0r0[14:14], i_0r0[14:14]);
  BUFEHD I80 (o_0r0[15:15], i_0r0[15:15]);
  BUFEHD I81 (o_0r0[16:16], i_0r0[16:16]);
  BUFEHD I82 (o_0r0[17:17], i_0r0[17:17]);
  BUFEHD I83 (o_0r0[18:18], i_0r0[18:18]);
  BUFEHD I84 (o_0r0[19:19], i_0r0[19:19]);
  BUFEHD I85 (o_0r0[20:20], i_0r0[20:20]);
  BUFEHD I86 (o_0r0[21:21], i_0r0[21:21]);
  BUFEHD I87 (o_0r0[22:22], i_0r0[22:22]);
  BUFEHD I88 (o_0r0[23:23], i_0r0[23:23]);
  BUFEHD I89 (o_0r0[24:24], i_0r0[24:24]);
  BUFEHD I90 (o_0r0[25:25], i_0r0[25:25]);
  BUFEHD I91 (o_0r0[26:26], i_0r0[26:26]);
  BUFEHD I92 (o_0r0[27:27], i_0r0[27:27]);
  BUFEHD I93 (o_0r0[28:28], i_0r0[28:28]);
  BUFEHD I94 (o_0r0[29:29], i_0r0[29:29]);
  BUFEHD I95 (o_0r0[30:30], i_0r0[30:30]);
  BUFEHD I96 (o_0r0[31:31], termf_1);
  BUFEHD I97 (o_0r1[0:0], i_0r1[0:0]);
  BUFEHD I98 (o_0r1[1:1], i_0r1[1:1]);
  BUFEHD I99 (o_0r1[2:2], i_0r1[2:2]);
  BUFEHD I100 (o_0r1[3:3], i_0r1[3:3]);
  BUFEHD I101 (o_0r1[4:4], i_0r1[4:4]);
  BUFEHD I102 (o_0r1[5:5], i_0r1[5:5]);
  BUFEHD I103 (o_0r1[6:6], i_0r1[6:6]);
  BUFEHD I104 (o_0r1[7:7], i_0r1[7:7]);
  BUFEHD I105 (o_0r1[8:8], i_0r1[8:8]);
  BUFEHD I106 (o_0r1[9:9], i_0r1[9:9]);
  BUFEHD I107 (o_0r1[10:10], i_0r1[10:10]);
  BUFEHD I108 (o_0r1[11:11], i_0r1[11:11]);
  BUFEHD I109 (o_0r1[12:12], i_0r1[12:12]);
  BUFEHD I110 (o_0r1[13:13], i_0r1[13:13]);
  BUFEHD I111 (o_0r1[14:14], i_0r1[14:14]);
  BUFEHD I112 (o_0r1[15:15], i_0r1[15:15]);
  BUFEHD I113 (o_0r1[16:16], i_0r1[16:16]);
  BUFEHD I114 (o_0r1[17:17], i_0r1[17:17]);
  BUFEHD I115 (o_0r1[18:18], i_0r1[18:18]);
  BUFEHD I116 (o_0r1[19:19], i_0r1[19:19]);
  BUFEHD I117 (o_0r1[20:20], i_0r1[20:20]);
  BUFEHD I118 (o_0r1[21:21], i_0r1[21:21]);
  BUFEHD I119 (o_0r1[22:22], i_0r1[22:22]);
  BUFEHD I120 (o_0r1[23:23], i_0r1[23:23]);
  BUFEHD I121 (o_0r1[24:24], i_0r1[24:24]);
  BUFEHD I122 (o_0r1[25:25], i_0r1[25:25]);
  BUFEHD I123 (o_0r1[26:26], i_0r1[26:26]);
  BUFEHD I124 (o_0r1[27:27], i_0r1[27:27]);
  BUFEHD I125 (o_0r1[28:28], i_0r1[28:28]);
  BUFEHD I126 (o_0r1[29:29], i_0r1[29:29]);
  BUFEHD I127 (o_0r1[30:30], i_0r1[30:30]);
  BUFEHD I128 (o_0r1[31:31], termt_1);
  BUFEHD I129 (i_0a, o_0a);
endmodule

// tko31m32_1nm1b1_2api0w31bt1o0w1b TeakO [
//     (1,TeakOConstant 1 1),
//     (2,TeakOAppend 1 [(0,0+:31),(1,0+:1)])] [One 31,One 32]
module tko31m32_1nm1b1_2api0w31bt1o0w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [30:0] i_0r0;
  input [30:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [30:0] gocomp_0;
  wire [10:0] simp331_0;
  wire tech34_int;
  wire tech35_int;
  wire tech36_int;
  wire tech37_int;
  wire tech38_int;
  wire tech39_int;
  wire tech40_int;
  wire tech41_int;
  wire tech42_int;
  wire tech43_int;
  wire [3:0] simp332_0;
  wire tech46_int;
  wire tech47_int;
  wire tech48_int;
  wire [1:0] simp333_0;
  wire tech51_int;
  wire termf_1;
  wire termt_1;
  OR2EHD I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2EHD I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2EHD I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2EHD I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2EHD I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2EHD I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2EHD I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2EHD I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2EHD I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2EHD I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2EHD I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2EHD I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2EHD I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2EHD I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2EHD I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2EHD I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2EHD I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2EHD I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2EHD I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2EHD I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2EHD I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2EHD I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2EHD I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2EHD I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2EHD I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2EHD I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2EHD I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2EHD I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2EHD I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2EHD I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2EHD I30 (gocomp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  AO222EHD I31 (tech34_int, gocomp_0[0:0], gocomp_0[1:1], tech34_int, gocomp_0[0:0], tech34_int, gocomp_0[1:1]);
  AO222EHD I32 (simp331_0[0:0], tech34_int, gocomp_0[2:2], simp331_0[0:0], tech34_int, simp331_0[0:0], gocomp_0[2:2]);
  AO222EHD I33 (tech35_int, gocomp_0[3:3], gocomp_0[4:4], tech35_int, gocomp_0[3:3], tech35_int, gocomp_0[4:4]);
  AO222EHD I34 (simp331_0[1:1], tech35_int, gocomp_0[5:5], simp331_0[1:1], tech35_int, simp331_0[1:1], gocomp_0[5:5]);
  AO222EHD I35 (tech36_int, gocomp_0[6:6], gocomp_0[7:7], tech36_int, gocomp_0[6:6], tech36_int, gocomp_0[7:7]);
  AO222EHD I36 (simp331_0[2:2], tech36_int, gocomp_0[8:8], simp331_0[2:2], tech36_int, simp331_0[2:2], gocomp_0[8:8]);
  AO222EHD I37 (tech37_int, gocomp_0[9:9], gocomp_0[10:10], tech37_int, gocomp_0[9:9], tech37_int, gocomp_0[10:10]);
  AO222EHD I38 (simp331_0[3:3], tech37_int, gocomp_0[11:11], simp331_0[3:3], tech37_int, simp331_0[3:3], gocomp_0[11:11]);
  AO222EHD I39 (tech38_int, gocomp_0[12:12], gocomp_0[13:13], tech38_int, gocomp_0[12:12], tech38_int, gocomp_0[13:13]);
  AO222EHD I40 (simp331_0[4:4], tech38_int, gocomp_0[14:14], simp331_0[4:4], tech38_int, simp331_0[4:4], gocomp_0[14:14]);
  AO222EHD I41 (tech39_int, gocomp_0[15:15], gocomp_0[16:16], tech39_int, gocomp_0[15:15], tech39_int, gocomp_0[16:16]);
  AO222EHD I42 (simp331_0[5:5], tech39_int, gocomp_0[17:17], simp331_0[5:5], tech39_int, simp331_0[5:5], gocomp_0[17:17]);
  AO222EHD I43 (tech40_int, gocomp_0[18:18], gocomp_0[19:19], tech40_int, gocomp_0[18:18], tech40_int, gocomp_0[19:19]);
  AO222EHD I44 (simp331_0[6:6], tech40_int, gocomp_0[20:20], simp331_0[6:6], tech40_int, simp331_0[6:6], gocomp_0[20:20]);
  AO222EHD I45 (tech41_int, gocomp_0[21:21], gocomp_0[22:22], tech41_int, gocomp_0[21:21], tech41_int, gocomp_0[22:22]);
  AO222EHD I46 (simp331_0[7:7], tech41_int, gocomp_0[23:23], simp331_0[7:7], tech41_int, simp331_0[7:7], gocomp_0[23:23]);
  AO222EHD I47 (tech42_int, gocomp_0[24:24], gocomp_0[25:25], tech42_int, gocomp_0[24:24], tech42_int, gocomp_0[25:25]);
  AO222EHD I48 (simp331_0[8:8], tech42_int, gocomp_0[26:26], simp331_0[8:8], tech42_int, simp331_0[8:8], gocomp_0[26:26]);
  AO222EHD I49 (tech43_int, gocomp_0[27:27], gocomp_0[28:28], tech43_int, gocomp_0[27:27], tech43_int, gocomp_0[28:28]);
  AO222EHD I50 (simp331_0[9:9], tech43_int, gocomp_0[29:29], simp331_0[9:9], tech43_int, simp331_0[9:9], gocomp_0[29:29]);
  BUFEHD I51 (simp331_0[10:10], gocomp_0[30:30]);
  AO222EHD I52 (tech46_int, simp331_0[0:0], simp331_0[1:1], tech46_int, simp331_0[0:0], tech46_int, simp331_0[1:1]);
  AO222EHD I53 (simp332_0[0:0], tech46_int, simp331_0[2:2], simp332_0[0:0], tech46_int, simp332_0[0:0], simp331_0[2:2]);
  AO222EHD I54 (tech47_int, simp331_0[3:3], simp331_0[4:4], tech47_int, simp331_0[3:3], tech47_int, simp331_0[4:4]);
  AO222EHD I55 (simp332_0[1:1], tech47_int, simp331_0[5:5], simp332_0[1:1], tech47_int, simp332_0[1:1], simp331_0[5:5]);
  AO222EHD I56 (tech48_int, simp331_0[6:6], simp331_0[7:7], tech48_int, simp331_0[6:6], tech48_int, simp331_0[7:7]);
  AO222EHD I57 (simp332_0[2:2], tech48_int, simp331_0[8:8], simp332_0[2:2], tech48_int, simp332_0[2:2], simp331_0[8:8]);
  AO222EHD I58 (simp332_0[3:3], simp331_0[9:9], simp331_0[10:10], simp332_0[3:3], simp331_0[9:9], simp332_0[3:3], simp331_0[10:10]);
  AO222EHD I59 (tech51_int, simp332_0[0:0], simp332_0[1:1], tech51_int, simp332_0[0:0], tech51_int, simp332_0[1:1]);
  AO222EHD I60 (simp333_0[0:0], tech51_int, simp332_0[2:2], simp333_0[0:0], tech51_int, simp333_0[0:0], simp332_0[2:2]);
  BUFEHD I61 (simp333_0[1:1], simp332_0[3:3]);
  AO222EHD I62 (go_0, simp333_0[0:0], simp333_0[1:1], go_0, simp333_0[0:0], go_0, simp333_0[1:1]);
  BUFEHD I63 (termt_1, go_0);
  TIE0DND I64 (termf_1);
  BUFEHD I65 (o_0r0[0:0], i_0r0[0:0]);
  BUFEHD I66 (o_0r0[1:1], i_0r0[1:1]);
  BUFEHD I67 (o_0r0[2:2], i_0r0[2:2]);
  BUFEHD I68 (o_0r0[3:3], i_0r0[3:3]);
  BUFEHD I69 (o_0r0[4:4], i_0r0[4:4]);
  BUFEHD I70 (o_0r0[5:5], i_0r0[5:5]);
  BUFEHD I71 (o_0r0[6:6], i_0r0[6:6]);
  BUFEHD I72 (o_0r0[7:7], i_0r0[7:7]);
  BUFEHD I73 (o_0r0[8:8], i_0r0[8:8]);
  BUFEHD I74 (o_0r0[9:9], i_0r0[9:9]);
  BUFEHD I75 (o_0r0[10:10], i_0r0[10:10]);
  BUFEHD I76 (o_0r0[11:11], i_0r0[11:11]);
  BUFEHD I77 (o_0r0[12:12], i_0r0[12:12]);
  BUFEHD I78 (o_0r0[13:13], i_0r0[13:13]);
  BUFEHD I79 (o_0r0[14:14], i_0r0[14:14]);
  BUFEHD I80 (o_0r0[15:15], i_0r0[15:15]);
  BUFEHD I81 (o_0r0[16:16], i_0r0[16:16]);
  BUFEHD I82 (o_0r0[17:17], i_0r0[17:17]);
  BUFEHD I83 (o_0r0[18:18], i_0r0[18:18]);
  BUFEHD I84 (o_0r0[19:19], i_0r0[19:19]);
  BUFEHD I85 (o_0r0[20:20], i_0r0[20:20]);
  BUFEHD I86 (o_0r0[21:21], i_0r0[21:21]);
  BUFEHD I87 (o_0r0[22:22], i_0r0[22:22]);
  BUFEHD I88 (o_0r0[23:23], i_0r0[23:23]);
  BUFEHD I89 (o_0r0[24:24], i_0r0[24:24]);
  BUFEHD I90 (o_0r0[25:25], i_0r0[25:25]);
  BUFEHD I91 (o_0r0[26:26], i_0r0[26:26]);
  BUFEHD I92 (o_0r0[27:27], i_0r0[27:27]);
  BUFEHD I93 (o_0r0[28:28], i_0r0[28:28]);
  BUFEHD I94 (o_0r0[29:29], i_0r0[29:29]);
  BUFEHD I95 (o_0r0[30:30], i_0r0[30:30]);
  BUFEHD I96 (o_0r0[31:31], termf_1);
  BUFEHD I97 (o_0r1[0:0], i_0r1[0:0]);
  BUFEHD I98 (o_0r1[1:1], i_0r1[1:1]);
  BUFEHD I99 (o_0r1[2:2], i_0r1[2:2]);
  BUFEHD I100 (o_0r1[3:3], i_0r1[3:3]);
  BUFEHD I101 (o_0r1[4:4], i_0r1[4:4]);
  BUFEHD I102 (o_0r1[5:5], i_0r1[5:5]);
  BUFEHD I103 (o_0r1[6:6], i_0r1[6:6]);
  BUFEHD I104 (o_0r1[7:7], i_0r1[7:7]);
  BUFEHD I105 (o_0r1[8:8], i_0r1[8:8]);
  BUFEHD I106 (o_0r1[9:9], i_0r1[9:9]);
  BUFEHD I107 (o_0r1[10:10], i_0r1[10:10]);
  BUFEHD I108 (o_0r1[11:11], i_0r1[11:11]);
  BUFEHD I109 (o_0r1[12:12], i_0r1[12:12]);
  BUFEHD I110 (o_0r1[13:13], i_0r1[13:13]);
  BUFEHD I111 (o_0r1[14:14], i_0r1[14:14]);
  BUFEHD I112 (o_0r1[15:15], i_0r1[15:15]);
  BUFEHD I113 (o_0r1[16:16], i_0r1[16:16]);
  BUFEHD I114 (o_0r1[17:17], i_0r1[17:17]);
  BUFEHD I115 (o_0r1[18:18], i_0r1[18:18]);
  BUFEHD I116 (o_0r1[19:19], i_0r1[19:19]);
  BUFEHD I117 (o_0r1[20:20], i_0r1[20:20]);
  BUFEHD I118 (o_0r1[21:21], i_0r1[21:21]);
  BUFEHD I119 (o_0r1[22:22], i_0r1[22:22]);
  BUFEHD I120 (o_0r1[23:23], i_0r1[23:23]);
  BUFEHD I121 (o_0r1[24:24], i_0r1[24:24]);
  BUFEHD I122 (o_0r1[25:25], i_0r1[25:25]);
  BUFEHD I123 (o_0r1[26:26], i_0r1[26:26]);
  BUFEHD I124 (o_0r1[27:27], i_0r1[27:27]);
  BUFEHD I125 (o_0r1[28:28], i_0r1[28:28]);
  BUFEHD I126 (o_0r1[29:29], i_0r1[29:29]);
  BUFEHD I127 (o_0r1[30:30], i_0r1[30:30]);
  BUFEHD I128 (o_0r1[31:31], termt_1);
  BUFEHD I129 (i_0a, o_0a);
endmodule

// tkvi32_wo0w32_ro0w32o0w31o1w31o1w31 TeakV "i" 32 [] [0] [0,0,1,1] [Many [32],Many [0],Many [0,0,0,0]
//   ,Many [32,31,31,31]]
module tkvi32_wo0w32_ro0w32o0w31o1w31o1w31 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [30:0] rd_1r0;
  output [30:0] rd_1r1;
  input rd_1a;
  output [30:0] rd_2r0;
  output [30:0] rd_2r1;
  input rd_2a;
  output [30:0] rd_3r0;
  output [30:0] rd_3r1;
  input rd_3a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire tech239_int;
  wire tech240_int;
  wire tech241_int;
  wire tech242_int;
  wire tech243_int;
  wire tech244_int;
  wire tech245_int;
  wire tech246_int;
  wire tech247_int;
  wire tech248_int;
  wire [3:0] simp2382_0;
  wire tech251_int;
  wire tech252_int;
  wire tech253_int;
  wire [1:0] simp2383_0;
  wire tech256_int;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire tech428_int;
  wire tech429_int;
  wire tech430_int;
  wire tech431_int;
  wire tech432_int;
  wire tech433_int;
  wire tech434_int;
  wire tech435_int;
  wire tech436_int;
  wire tech437_int;
  wire tech438_int;
  wire [3:0] simp4072_0;
  wire tech440_int;
  wire tech441_int;
  wire tech442_int;
  wire [1:0] simp4073_0;
  wire tech445_int;
  wire [2:0] simp6581_0;
  INVHHD I0 (nreset_0, reset);
  AN2EHD I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AN2EHD I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AN2EHD I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AN2EHD I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AN2EHD I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AN2EHD I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AN2EHD I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AN2EHD I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AN2EHD I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AN2EHD I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AN2EHD I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AN2EHD I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AN2EHD I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AN2EHD I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AN2EHD I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AN2EHD I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AN2EHD I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AN2EHD I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AN2EHD I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AN2EHD I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AN2EHD I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AN2EHD I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AN2EHD I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AN2EHD I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AN2EHD I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AN2EHD I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AN2EHD I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AN2EHD I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AN2EHD I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AN2EHD I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AN2EHD I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AN2EHD I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AN2EHD I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AN2EHD I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AN2EHD I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AN2EHD I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AN2EHD I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AN2EHD I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AN2EHD I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AN2EHD I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AN2EHD I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AN2EHD I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AN2EHD I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AN2EHD I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AN2EHD I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AN2EHD I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AN2EHD I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AN2EHD I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AN2EHD I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AN2EHD I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AN2EHD I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AN2EHD I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AN2EHD I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AN2EHD I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AN2EHD I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AN2EHD I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AN2EHD I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AN2EHD I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AN2EHD I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AN2EHD I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AN2EHD I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AN2EHD I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AN2EHD I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AN2EHD I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AN2EHD I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AN2EHD I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AN2EHD I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AN2EHD I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AN2EHD I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AN2EHD I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AN2EHD I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AN2EHD I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AN2EHD I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AN2EHD I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AN2EHD I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AN2EHD I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AN2EHD I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AN2EHD I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AN2EHD I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AN2EHD I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AN2EHD I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AN2EHD I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AN2EHD I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AN2EHD I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AN2EHD I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AN2EHD I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AN2EHD I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AN2EHD I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AN2EHD I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AN2EHD I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AN2EHD I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AN2EHD I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AN2EHD I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AN2EHD I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AN2EHD I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AN2EHD I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NR2EHD I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NR2EHD I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NR2EHD I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NR2EHD I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NR2EHD I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NR2EHD I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NR2EHD I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NR2EHD I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NR2EHD I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NR2EHD I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NR2EHD I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NR2EHD I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NR2EHD I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NR2EHD I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NR2EHD I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NR2EHD I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NR2EHD I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NR2EHD I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NR2EHD I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NR2EHD I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NR2EHD I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NR2EHD I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NR2EHD I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NR2EHD I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NR2EHD I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NR2EHD I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NR2EHD I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NR2EHD I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NR2EHD I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NR2EHD I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NR2EHD I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NR2EHD I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NR3EHD I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NR3EHD I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NR3EHD I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NR3EHD I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NR3EHD I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NR3EHD I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NR3EHD I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NR3EHD I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NR3EHD I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NR3EHD I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NR3EHD I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NR3EHD I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NR3EHD I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NR3EHD I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NR3EHD I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NR3EHD I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NR3EHD I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NR3EHD I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NR3EHD I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NR3EHD I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NR3EHD I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NR3EHD I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NR3EHD I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NR3EHD I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NR3EHD I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NR3EHD I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NR3EHD I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NR3EHD I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NR3EHD I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NR3EHD I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NR3EHD I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NR3EHD I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22EHD I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22EHD I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22EHD I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22EHD I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22EHD I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22EHD I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22EHD I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22EHD I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22EHD I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22EHD I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22EHD I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22EHD I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22EHD I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22EHD I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22EHD I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22EHD I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22EHD I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22EHD I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22EHD I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22EHD I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22EHD I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22EHD I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22EHD I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22EHD I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22EHD I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22EHD I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22EHD I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22EHD I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22EHD I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22EHD I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22EHD I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22EHD I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2EHD I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2EHD I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2EHD I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2EHD I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2EHD I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2EHD I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2EHD I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2EHD I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2EHD I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2EHD I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2EHD I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2EHD I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2EHD I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2EHD I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2EHD I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2EHD I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2EHD I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2EHD I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2EHD I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2EHD I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2EHD I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2EHD I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2EHD I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2EHD I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2EHD I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2EHD I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2EHD I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2EHD I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2EHD I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2EHD I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2EHD I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2EHD I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  AO222EHD I225 (tech239_int, comp0_0[0:0], comp0_0[1:1], tech239_int, comp0_0[0:0], tech239_int, comp0_0[1:1]);
  AO222EHD I226 (simp2381_0[0:0], tech239_int, comp0_0[2:2], simp2381_0[0:0], tech239_int, simp2381_0[0:0], comp0_0[2:2]);
  AO222EHD I227 (tech240_int, comp0_0[3:3], comp0_0[4:4], tech240_int, comp0_0[3:3], tech240_int, comp0_0[4:4]);
  AO222EHD I228 (simp2381_0[1:1], tech240_int, comp0_0[5:5], simp2381_0[1:1], tech240_int, simp2381_0[1:1], comp0_0[5:5]);
  AO222EHD I229 (tech241_int, comp0_0[6:6], comp0_0[7:7], tech241_int, comp0_0[6:6], tech241_int, comp0_0[7:7]);
  AO222EHD I230 (simp2381_0[2:2], tech241_int, comp0_0[8:8], simp2381_0[2:2], tech241_int, simp2381_0[2:2], comp0_0[8:8]);
  AO222EHD I231 (tech242_int, comp0_0[9:9], comp0_0[10:10], tech242_int, comp0_0[9:9], tech242_int, comp0_0[10:10]);
  AO222EHD I232 (simp2381_0[3:3], tech242_int, comp0_0[11:11], simp2381_0[3:3], tech242_int, simp2381_0[3:3], comp0_0[11:11]);
  AO222EHD I233 (tech243_int, comp0_0[12:12], comp0_0[13:13], tech243_int, comp0_0[12:12], tech243_int, comp0_0[13:13]);
  AO222EHD I234 (simp2381_0[4:4], tech243_int, comp0_0[14:14], simp2381_0[4:4], tech243_int, simp2381_0[4:4], comp0_0[14:14]);
  AO222EHD I235 (tech244_int, comp0_0[15:15], comp0_0[16:16], tech244_int, comp0_0[15:15], tech244_int, comp0_0[16:16]);
  AO222EHD I236 (simp2381_0[5:5], tech244_int, comp0_0[17:17], simp2381_0[5:5], tech244_int, simp2381_0[5:5], comp0_0[17:17]);
  AO222EHD I237 (tech245_int, comp0_0[18:18], comp0_0[19:19], tech245_int, comp0_0[18:18], tech245_int, comp0_0[19:19]);
  AO222EHD I238 (simp2381_0[6:6], tech245_int, comp0_0[20:20], simp2381_0[6:6], tech245_int, simp2381_0[6:6], comp0_0[20:20]);
  AO222EHD I239 (tech246_int, comp0_0[21:21], comp0_0[22:22], tech246_int, comp0_0[21:21], tech246_int, comp0_0[22:22]);
  AO222EHD I240 (simp2381_0[7:7], tech246_int, comp0_0[23:23], simp2381_0[7:7], tech246_int, simp2381_0[7:7], comp0_0[23:23]);
  AO222EHD I241 (tech247_int, comp0_0[24:24], comp0_0[25:25], tech247_int, comp0_0[24:24], tech247_int, comp0_0[25:25]);
  AO222EHD I242 (simp2381_0[8:8], tech247_int, comp0_0[26:26], simp2381_0[8:8], tech247_int, simp2381_0[8:8], comp0_0[26:26]);
  AO222EHD I243 (tech248_int, comp0_0[27:27], comp0_0[28:28], tech248_int, comp0_0[27:27], tech248_int, comp0_0[28:28]);
  AO222EHD I244 (simp2381_0[9:9], tech248_int, comp0_0[29:29], simp2381_0[9:9], tech248_int, simp2381_0[9:9], comp0_0[29:29]);
  AO222EHD I245 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31], simp2381_0[10:10], comp0_0[30:30], simp2381_0[10:10], comp0_0[31:31]);
  AO222EHD I246 (tech251_int, simp2381_0[0:0], simp2381_0[1:1], tech251_int, simp2381_0[0:0], tech251_int, simp2381_0[1:1]);
  AO222EHD I247 (simp2382_0[0:0], tech251_int, simp2381_0[2:2], simp2382_0[0:0], tech251_int, simp2382_0[0:0], simp2381_0[2:2]);
  AO222EHD I248 (tech252_int, simp2381_0[3:3], simp2381_0[4:4], tech252_int, simp2381_0[3:3], tech252_int, simp2381_0[4:4]);
  AO222EHD I249 (simp2382_0[1:1], tech252_int, simp2381_0[5:5], simp2382_0[1:1], tech252_int, simp2382_0[1:1], simp2381_0[5:5]);
  AO222EHD I250 (tech253_int, simp2381_0[6:6], simp2381_0[7:7], tech253_int, simp2381_0[6:6], tech253_int, simp2381_0[7:7]);
  AO222EHD I251 (simp2382_0[2:2], tech253_int, simp2381_0[8:8], simp2382_0[2:2], tech253_int, simp2382_0[2:2], simp2381_0[8:8]);
  AO222EHD I252 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10], simp2382_0[3:3], simp2381_0[9:9], simp2382_0[3:3], simp2381_0[10:10]);
  AO222EHD I253 (tech256_int, simp2382_0[0:0], simp2382_0[1:1], tech256_int, simp2382_0[0:0], tech256_int, simp2382_0[1:1]);
  AO222EHD I254 (simp2383_0[0:0], tech256_int, simp2382_0[2:2], simp2383_0[0:0], tech256_int, simp2383_0[0:0], simp2382_0[2:2]);
  BUFEHD I255 (simp2383_0[1:1], simp2382_0[3:3]);
  AO222EHD I256 (wc_0, simp2383_0[0:0], simp2383_0[1:1], wc_0, simp2383_0[0:0], wc_0, simp2383_0[1:1]);
  AN2EHD I257 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AN2EHD I258 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AN2EHD I259 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AN2EHD I260 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AN2EHD I261 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AN2EHD I262 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AN2EHD I263 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AN2EHD I264 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AN2EHD I265 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AN2EHD I266 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AN2EHD I267 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AN2EHD I268 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AN2EHD I269 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AN2EHD I270 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AN2EHD I271 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AN2EHD I272 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AN2EHD I273 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AN2EHD I274 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AN2EHD I275 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AN2EHD I276 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AN2EHD I277 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AN2EHD I278 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AN2EHD I279 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AN2EHD I280 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AN2EHD I281 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AN2EHD I282 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AN2EHD I283 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AN2EHD I284 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AN2EHD I285 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AN2EHD I286 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AN2EHD I287 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AN2EHD I288 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AN2EHD I289 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AN2EHD I290 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AN2EHD I291 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AN2EHD I292 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AN2EHD I293 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AN2EHD I294 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AN2EHD I295 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AN2EHD I296 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AN2EHD I297 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AN2EHD I298 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AN2EHD I299 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AN2EHD I300 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AN2EHD I301 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AN2EHD I302 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AN2EHD I303 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AN2EHD I304 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AN2EHD I305 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AN2EHD I306 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AN2EHD I307 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AN2EHD I308 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AN2EHD I309 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AN2EHD I310 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AN2EHD I311 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AN2EHD I312 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AN2EHD I313 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AN2EHD I314 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AN2EHD I315 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AN2EHD I316 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AN2EHD I317 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AN2EHD I318 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AN2EHD I319 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AN2EHD I320 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFEHD I321 (conwigc_0, wc_0);
  AO12EHD I322 (conwig_0, conwigc_0, conwigc_0, conwigcanw_0);
  NR2EHD I323 (conwigcanw_0, anyread_0, conwig_0);
  BUFEHD I324 (wf_0[0:0], conwgif_0[0:0]);
  BUFEHD I325 (wt_0[0:0], conwgit_0[0:0]);
  BUFEHD I326 (wenr_0[0:0], wc_0);
  BUFEHD I327 (wf_0[1:1], conwgif_0[1:1]);
  BUFEHD I328 (wt_0[1:1], conwgit_0[1:1]);
  BUFEHD I329 (wenr_0[1:1], wc_0);
  BUFEHD I330 (wf_0[2:2], conwgif_0[2:2]);
  BUFEHD I331 (wt_0[2:2], conwgit_0[2:2]);
  BUFEHD I332 (wenr_0[2:2], wc_0);
  BUFEHD I333 (wf_0[3:3], conwgif_0[3:3]);
  BUFEHD I334 (wt_0[3:3], conwgit_0[3:3]);
  BUFEHD I335 (wenr_0[3:3], wc_0);
  BUFEHD I336 (wf_0[4:4], conwgif_0[4:4]);
  BUFEHD I337 (wt_0[4:4], conwgit_0[4:4]);
  BUFEHD I338 (wenr_0[4:4], wc_0);
  BUFEHD I339 (wf_0[5:5], conwgif_0[5:5]);
  BUFEHD I340 (wt_0[5:5], conwgit_0[5:5]);
  BUFEHD I341 (wenr_0[5:5], wc_0);
  BUFEHD I342 (wf_0[6:6], conwgif_0[6:6]);
  BUFEHD I343 (wt_0[6:6], conwgit_0[6:6]);
  BUFEHD I344 (wenr_0[6:6], wc_0);
  BUFEHD I345 (wf_0[7:7], conwgif_0[7:7]);
  BUFEHD I346 (wt_0[7:7], conwgit_0[7:7]);
  BUFEHD I347 (wenr_0[7:7], wc_0);
  BUFEHD I348 (wf_0[8:8], conwgif_0[8:8]);
  BUFEHD I349 (wt_0[8:8], conwgit_0[8:8]);
  BUFEHD I350 (wenr_0[8:8], wc_0);
  BUFEHD I351 (wf_0[9:9], conwgif_0[9:9]);
  BUFEHD I352 (wt_0[9:9], conwgit_0[9:9]);
  BUFEHD I353 (wenr_0[9:9], wc_0);
  BUFEHD I354 (wf_0[10:10], conwgif_0[10:10]);
  BUFEHD I355 (wt_0[10:10], conwgit_0[10:10]);
  BUFEHD I356 (wenr_0[10:10], wc_0);
  BUFEHD I357 (wf_0[11:11], conwgif_0[11:11]);
  BUFEHD I358 (wt_0[11:11], conwgit_0[11:11]);
  BUFEHD I359 (wenr_0[11:11], wc_0);
  BUFEHD I360 (wf_0[12:12], conwgif_0[12:12]);
  BUFEHD I361 (wt_0[12:12], conwgit_0[12:12]);
  BUFEHD I362 (wenr_0[12:12], wc_0);
  BUFEHD I363 (wf_0[13:13], conwgif_0[13:13]);
  BUFEHD I364 (wt_0[13:13], conwgit_0[13:13]);
  BUFEHD I365 (wenr_0[13:13], wc_0);
  BUFEHD I366 (wf_0[14:14], conwgif_0[14:14]);
  BUFEHD I367 (wt_0[14:14], conwgit_0[14:14]);
  BUFEHD I368 (wenr_0[14:14], wc_0);
  BUFEHD I369 (wf_0[15:15], conwgif_0[15:15]);
  BUFEHD I370 (wt_0[15:15], conwgit_0[15:15]);
  BUFEHD I371 (wenr_0[15:15], wc_0);
  BUFEHD I372 (wf_0[16:16], conwgif_0[16:16]);
  BUFEHD I373 (wt_0[16:16], conwgit_0[16:16]);
  BUFEHD I374 (wenr_0[16:16], wc_0);
  BUFEHD I375 (wf_0[17:17], conwgif_0[17:17]);
  BUFEHD I376 (wt_0[17:17], conwgit_0[17:17]);
  BUFEHD I377 (wenr_0[17:17], wc_0);
  BUFEHD I378 (wf_0[18:18], conwgif_0[18:18]);
  BUFEHD I379 (wt_0[18:18], conwgit_0[18:18]);
  BUFEHD I380 (wenr_0[18:18], wc_0);
  BUFEHD I381 (wf_0[19:19], conwgif_0[19:19]);
  BUFEHD I382 (wt_0[19:19], conwgit_0[19:19]);
  BUFEHD I383 (wenr_0[19:19], wc_0);
  BUFEHD I384 (wf_0[20:20], conwgif_0[20:20]);
  BUFEHD I385 (wt_0[20:20], conwgit_0[20:20]);
  BUFEHD I386 (wenr_0[20:20], wc_0);
  BUFEHD I387 (wf_0[21:21], conwgif_0[21:21]);
  BUFEHD I388 (wt_0[21:21], conwgit_0[21:21]);
  BUFEHD I389 (wenr_0[21:21], wc_0);
  BUFEHD I390 (wf_0[22:22], conwgif_0[22:22]);
  BUFEHD I391 (wt_0[22:22], conwgit_0[22:22]);
  BUFEHD I392 (wenr_0[22:22], wc_0);
  BUFEHD I393 (wf_0[23:23], conwgif_0[23:23]);
  BUFEHD I394 (wt_0[23:23], conwgit_0[23:23]);
  BUFEHD I395 (wenr_0[23:23], wc_0);
  BUFEHD I396 (wf_0[24:24], conwgif_0[24:24]);
  BUFEHD I397 (wt_0[24:24], conwgit_0[24:24]);
  BUFEHD I398 (wenr_0[24:24], wc_0);
  BUFEHD I399 (wf_0[25:25], conwgif_0[25:25]);
  BUFEHD I400 (wt_0[25:25], conwgit_0[25:25]);
  BUFEHD I401 (wenr_0[25:25], wc_0);
  BUFEHD I402 (wf_0[26:26], conwgif_0[26:26]);
  BUFEHD I403 (wt_0[26:26], conwgit_0[26:26]);
  BUFEHD I404 (wenr_0[26:26], wc_0);
  BUFEHD I405 (wf_0[27:27], conwgif_0[27:27]);
  BUFEHD I406 (wt_0[27:27], conwgit_0[27:27]);
  BUFEHD I407 (wenr_0[27:27], wc_0);
  BUFEHD I408 (wf_0[28:28], conwgif_0[28:28]);
  BUFEHD I409 (wt_0[28:28], conwgit_0[28:28]);
  BUFEHD I410 (wenr_0[28:28], wc_0);
  BUFEHD I411 (wf_0[29:29], conwgif_0[29:29]);
  BUFEHD I412 (wt_0[29:29], conwgit_0[29:29]);
  BUFEHD I413 (wenr_0[29:29], wc_0);
  BUFEHD I414 (wf_0[30:30], conwgif_0[30:30]);
  BUFEHD I415 (wt_0[30:30], conwgit_0[30:30]);
  BUFEHD I416 (wenr_0[30:30], wc_0);
  BUFEHD I417 (wf_0[31:31], conwgif_0[31:31]);
  BUFEHD I418 (wt_0[31:31], conwgit_0[31:31]);
  BUFEHD I419 (wenr_0[31:31], wc_0);
  AO222EHD I420 (tech428_int, conwig_0, wacks_0[0:0], tech428_int, conwig_0, tech428_int, wacks_0[0:0]);
  AO222EHD I421 (simp4071_0[0:0], tech428_int, wacks_0[1:1], simp4071_0[0:0], tech428_int, simp4071_0[0:0], wacks_0[1:1]);
  AO222EHD I422 (tech429_int, wacks_0[2:2], wacks_0[3:3], tech429_int, wacks_0[2:2], tech429_int, wacks_0[3:3]);
  AO222EHD I423 (simp4071_0[1:1], tech429_int, wacks_0[4:4], simp4071_0[1:1], tech429_int, simp4071_0[1:1], wacks_0[4:4]);
  AO222EHD I424 (tech430_int, wacks_0[5:5], wacks_0[6:6], tech430_int, wacks_0[5:5], tech430_int, wacks_0[6:6]);
  AO222EHD I425 (simp4071_0[2:2], tech430_int, wacks_0[7:7], simp4071_0[2:2], tech430_int, simp4071_0[2:2], wacks_0[7:7]);
  AO222EHD I426 (tech431_int, wacks_0[8:8], wacks_0[9:9], tech431_int, wacks_0[8:8], tech431_int, wacks_0[9:9]);
  AO222EHD I427 (simp4071_0[3:3], tech431_int, wacks_0[10:10], simp4071_0[3:3], tech431_int, simp4071_0[3:3], wacks_0[10:10]);
  AO222EHD I428 (tech432_int, wacks_0[11:11], wacks_0[12:12], tech432_int, wacks_0[11:11], tech432_int, wacks_0[12:12]);
  AO222EHD I429 (simp4071_0[4:4], tech432_int, wacks_0[13:13], simp4071_0[4:4], tech432_int, simp4071_0[4:4], wacks_0[13:13]);
  AO222EHD I430 (tech433_int, wacks_0[14:14], wacks_0[15:15], tech433_int, wacks_0[14:14], tech433_int, wacks_0[15:15]);
  AO222EHD I431 (simp4071_0[5:5], tech433_int, wacks_0[16:16], simp4071_0[5:5], tech433_int, simp4071_0[5:5], wacks_0[16:16]);
  AO222EHD I432 (tech434_int, wacks_0[17:17], wacks_0[18:18], tech434_int, wacks_0[17:17], tech434_int, wacks_0[18:18]);
  AO222EHD I433 (simp4071_0[6:6], tech434_int, wacks_0[19:19], simp4071_0[6:6], tech434_int, simp4071_0[6:6], wacks_0[19:19]);
  AO222EHD I434 (tech435_int, wacks_0[20:20], wacks_0[21:21], tech435_int, wacks_0[20:20], tech435_int, wacks_0[21:21]);
  AO222EHD I435 (simp4071_0[7:7], tech435_int, wacks_0[22:22], simp4071_0[7:7], tech435_int, simp4071_0[7:7], wacks_0[22:22]);
  AO222EHD I436 (tech436_int, wacks_0[23:23], wacks_0[24:24], tech436_int, wacks_0[23:23], tech436_int, wacks_0[24:24]);
  AO222EHD I437 (simp4071_0[8:8], tech436_int, wacks_0[25:25], simp4071_0[8:8], tech436_int, simp4071_0[8:8], wacks_0[25:25]);
  AO222EHD I438 (tech437_int, wacks_0[26:26], wacks_0[27:27], tech437_int, wacks_0[26:26], tech437_int, wacks_0[27:27]);
  AO222EHD I439 (simp4071_0[9:9], tech437_int, wacks_0[28:28], simp4071_0[9:9], tech437_int, simp4071_0[9:9], wacks_0[28:28]);
  AO222EHD I440 (tech438_int, wacks_0[29:29], wacks_0[30:30], tech438_int, wacks_0[29:29], tech438_int, wacks_0[30:30]);
  AO222EHD I441 (simp4071_0[10:10], tech438_int, wacks_0[31:31], simp4071_0[10:10], tech438_int, simp4071_0[10:10], wacks_0[31:31]);
  AO222EHD I442 (tech440_int, simp4071_0[0:0], simp4071_0[1:1], tech440_int, simp4071_0[0:0], tech440_int, simp4071_0[1:1]);
  AO222EHD I443 (simp4072_0[0:0], tech440_int, simp4071_0[2:2], simp4072_0[0:0], tech440_int, simp4072_0[0:0], simp4071_0[2:2]);
  AO222EHD I444 (tech441_int, simp4071_0[3:3], simp4071_0[4:4], tech441_int, simp4071_0[3:3], tech441_int, simp4071_0[4:4]);
  AO222EHD I445 (simp4072_0[1:1], tech441_int, simp4071_0[5:5], simp4072_0[1:1], tech441_int, simp4072_0[1:1], simp4071_0[5:5]);
  AO222EHD I446 (tech442_int, simp4071_0[6:6], simp4071_0[7:7], tech442_int, simp4071_0[6:6], tech442_int, simp4071_0[7:7]);
  AO222EHD I447 (simp4072_0[2:2], tech442_int, simp4071_0[8:8], simp4072_0[2:2], tech442_int, simp4072_0[2:2], simp4071_0[8:8]);
  AO222EHD I448 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10], simp4072_0[3:3], simp4071_0[9:9], simp4072_0[3:3], simp4071_0[10:10]);
  AO222EHD I449 (tech445_int, simp4072_0[0:0], simp4072_0[1:1], tech445_int, simp4072_0[0:0], tech445_int, simp4072_0[1:1]);
  AO222EHD I450 (simp4073_0[0:0], tech445_int, simp4072_0[2:2], simp4073_0[0:0], tech445_int, simp4073_0[0:0], simp4072_0[2:2]);
  BUFEHD I451 (simp4073_0[1:1], simp4072_0[3:3]);
  AO222EHD I452 (wd_0r, simp4073_0[0:0], simp4073_0[1:1], wd_0r, simp4073_0[0:0], wd_0r, simp4073_0[1:1]);
  AN2EHD I453 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AN2EHD I454 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AN2EHD I455 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AN2EHD I456 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AN2EHD I457 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AN2EHD I458 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AN2EHD I459 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AN2EHD I460 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AN2EHD I461 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AN2EHD I462 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AN2EHD I463 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AN2EHD I464 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AN2EHD I465 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AN2EHD I466 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AN2EHD I467 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AN2EHD I468 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AN2EHD I469 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AN2EHD I470 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AN2EHD I471 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AN2EHD I472 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AN2EHD I473 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AN2EHD I474 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AN2EHD I475 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AN2EHD I476 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AN2EHD I477 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AN2EHD I478 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AN2EHD I479 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AN2EHD I480 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AN2EHD I481 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AN2EHD I482 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AN2EHD I483 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AN2EHD I484 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AN2EHD I485 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AN2EHD I486 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AN2EHD I487 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AN2EHD I488 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AN2EHD I489 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AN2EHD I490 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AN2EHD I491 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AN2EHD I492 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AN2EHD I493 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AN2EHD I494 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AN2EHD I495 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AN2EHD I496 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AN2EHD I497 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AN2EHD I498 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AN2EHD I499 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AN2EHD I500 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AN2EHD I501 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AN2EHD I502 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AN2EHD I503 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AN2EHD I504 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AN2EHD I505 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AN2EHD I506 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AN2EHD I507 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AN2EHD I508 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AN2EHD I509 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AN2EHD I510 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AN2EHD I511 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AN2EHD I512 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AN2EHD I513 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AN2EHD I514 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AN2EHD I515 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AN2EHD I516 (rd_2r0[0:0], df_0[1:1], rg_2r);
  AN2EHD I517 (rd_2r0[1:1], df_0[2:2], rg_2r);
  AN2EHD I518 (rd_2r0[2:2], df_0[3:3], rg_2r);
  AN2EHD I519 (rd_2r0[3:3], df_0[4:4], rg_2r);
  AN2EHD I520 (rd_2r0[4:4], df_0[5:5], rg_2r);
  AN2EHD I521 (rd_2r0[5:5], df_0[6:6], rg_2r);
  AN2EHD I522 (rd_2r0[6:6], df_0[7:7], rg_2r);
  AN2EHD I523 (rd_2r0[7:7], df_0[8:8], rg_2r);
  AN2EHD I524 (rd_2r0[8:8], df_0[9:9], rg_2r);
  AN2EHD I525 (rd_2r0[9:9], df_0[10:10], rg_2r);
  AN2EHD I526 (rd_2r0[10:10], df_0[11:11], rg_2r);
  AN2EHD I527 (rd_2r0[11:11], df_0[12:12], rg_2r);
  AN2EHD I528 (rd_2r0[12:12], df_0[13:13], rg_2r);
  AN2EHD I529 (rd_2r0[13:13], df_0[14:14], rg_2r);
  AN2EHD I530 (rd_2r0[14:14], df_0[15:15], rg_2r);
  AN2EHD I531 (rd_2r0[15:15], df_0[16:16], rg_2r);
  AN2EHD I532 (rd_2r0[16:16], df_0[17:17], rg_2r);
  AN2EHD I533 (rd_2r0[17:17], df_0[18:18], rg_2r);
  AN2EHD I534 (rd_2r0[18:18], df_0[19:19], rg_2r);
  AN2EHD I535 (rd_2r0[19:19], df_0[20:20], rg_2r);
  AN2EHD I536 (rd_2r0[20:20], df_0[21:21], rg_2r);
  AN2EHD I537 (rd_2r0[21:21], df_0[22:22], rg_2r);
  AN2EHD I538 (rd_2r0[22:22], df_0[23:23], rg_2r);
  AN2EHD I539 (rd_2r0[23:23], df_0[24:24], rg_2r);
  AN2EHD I540 (rd_2r0[24:24], df_0[25:25], rg_2r);
  AN2EHD I541 (rd_2r0[25:25], df_0[26:26], rg_2r);
  AN2EHD I542 (rd_2r0[26:26], df_0[27:27], rg_2r);
  AN2EHD I543 (rd_2r0[27:27], df_0[28:28], rg_2r);
  AN2EHD I544 (rd_2r0[28:28], df_0[29:29], rg_2r);
  AN2EHD I545 (rd_2r0[29:29], df_0[30:30], rg_2r);
  AN2EHD I546 (rd_2r0[30:30], df_0[31:31], rg_2r);
  AN2EHD I547 (rd_3r0[0:0], df_0[1:1], rg_3r);
  AN2EHD I548 (rd_3r0[1:1], df_0[2:2], rg_3r);
  AN2EHD I549 (rd_3r0[2:2], df_0[3:3], rg_3r);
  AN2EHD I550 (rd_3r0[3:3], df_0[4:4], rg_3r);
  AN2EHD I551 (rd_3r0[4:4], df_0[5:5], rg_3r);
  AN2EHD I552 (rd_3r0[5:5], df_0[6:6], rg_3r);
  AN2EHD I553 (rd_3r0[6:6], df_0[7:7], rg_3r);
  AN2EHD I554 (rd_3r0[7:7], df_0[8:8], rg_3r);
  AN2EHD I555 (rd_3r0[8:8], df_0[9:9], rg_3r);
  AN2EHD I556 (rd_3r0[9:9], df_0[10:10], rg_3r);
  AN2EHD I557 (rd_3r0[10:10], df_0[11:11], rg_3r);
  AN2EHD I558 (rd_3r0[11:11], df_0[12:12], rg_3r);
  AN2EHD I559 (rd_3r0[12:12], df_0[13:13], rg_3r);
  AN2EHD I560 (rd_3r0[13:13], df_0[14:14], rg_3r);
  AN2EHD I561 (rd_3r0[14:14], df_0[15:15], rg_3r);
  AN2EHD I562 (rd_3r0[15:15], df_0[16:16], rg_3r);
  AN2EHD I563 (rd_3r0[16:16], df_0[17:17], rg_3r);
  AN2EHD I564 (rd_3r0[17:17], df_0[18:18], rg_3r);
  AN2EHD I565 (rd_3r0[18:18], df_0[19:19], rg_3r);
  AN2EHD I566 (rd_3r0[19:19], df_0[20:20], rg_3r);
  AN2EHD I567 (rd_3r0[20:20], df_0[21:21], rg_3r);
  AN2EHD I568 (rd_3r0[21:21], df_0[22:22], rg_3r);
  AN2EHD I569 (rd_3r0[22:22], df_0[23:23], rg_3r);
  AN2EHD I570 (rd_3r0[23:23], df_0[24:24], rg_3r);
  AN2EHD I571 (rd_3r0[24:24], df_0[25:25], rg_3r);
  AN2EHD I572 (rd_3r0[25:25], df_0[26:26], rg_3r);
  AN2EHD I573 (rd_3r0[26:26], df_0[27:27], rg_3r);
  AN2EHD I574 (rd_3r0[27:27], df_0[28:28], rg_3r);
  AN2EHD I575 (rd_3r0[28:28], df_0[29:29], rg_3r);
  AN2EHD I576 (rd_3r0[29:29], df_0[30:30], rg_3r);
  AN2EHD I577 (rd_3r0[30:30], df_0[31:31], rg_3r);
  AN2EHD I578 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AN2EHD I579 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AN2EHD I580 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AN2EHD I581 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AN2EHD I582 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AN2EHD I583 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AN2EHD I584 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AN2EHD I585 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AN2EHD I586 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AN2EHD I587 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AN2EHD I588 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AN2EHD I589 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AN2EHD I590 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AN2EHD I591 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AN2EHD I592 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AN2EHD I593 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AN2EHD I594 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AN2EHD I595 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AN2EHD I596 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AN2EHD I597 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AN2EHD I598 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AN2EHD I599 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AN2EHD I600 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AN2EHD I601 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AN2EHD I602 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AN2EHD I603 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AN2EHD I604 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AN2EHD I605 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AN2EHD I606 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AN2EHD I607 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AN2EHD I608 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AN2EHD I609 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AN2EHD I610 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AN2EHD I611 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AN2EHD I612 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AN2EHD I613 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AN2EHD I614 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AN2EHD I615 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AN2EHD I616 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AN2EHD I617 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AN2EHD I618 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AN2EHD I619 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AN2EHD I620 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AN2EHD I621 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AN2EHD I622 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AN2EHD I623 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AN2EHD I624 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AN2EHD I625 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AN2EHD I626 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AN2EHD I627 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AN2EHD I628 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AN2EHD I629 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AN2EHD I630 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AN2EHD I631 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AN2EHD I632 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AN2EHD I633 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AN2EHD I634 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AN2EHD I635 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AN2EHD I636 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AN2EHD I637 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AN2EHD I638 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AN2EHD I639 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AN2EHD I640 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AN2EHD I641 (rd_2r1[0:0], dt_0[1:1], rg_2r);
  AN2EHD I642 (rd_2r1[1:1], dt_0[2:2], rg_2r);
  AN2EHD I643 (rd_2r1[2:2], dt_0[3:3], rg_2r);
  AN2EHD I644 (rd_2r1[3:3], dt_0[4:4], rg_2r);
  AN2EHD I645 (rd_2r1[4:4], dt_0[5:5], rg_2r);
  AN2EHD I646 (rd_2r1[5:5], dt_0[6:6], rg_2r);
  AN2EHD I647 (rd_2r1[6:6], dt_0[7:7], rg_2r);
  AN2EHD I648 (rd_2r1[7:7], dt_0[8:8], rg_2r);
  AN2EHD I649 (rd_2r1[8:8], dt_0[9:9], rg_2r);
  AN2EHD I650 (rd_2r1[9:9], dt_0[10:10], rg_2r);
  AN2EHD I651 (rd_2r1[10:10], dt_0[11:11], rg_2r);
  AN2EHD I652 (rd_2r1[11:11], dt_0[12:12], rg_2r);
  AN2EHD I653 (rd_2r1[12:12], dt_0[13:13], rg_2r);
  AN2EHD I654 (rd_2r1[13:13], dt_0[14:14], rg_2r);
  AN2EHD I655 (rd_2r1[14:14], dt_0[15:15], rg_2r);
  AN2EHD I656 (rd_2r1[15:15], dt_0[16:16], rg_2r);
  AN2EHD I657 (rd_2r1[16:16], dt_0[17:17], rg_2r);
  AN2EHD I658 (rd_2r1[17:17], dt_0[18:18], rg_2r);
  AN2EHD I659 (rd_2r1[18:18], dt_0[19:19], rg_2r);
  AN2EHD I660 (rd_2r1[19:19], dt_0[20:20], rg_2r);
  AN2EHD I661 (rd_2r1[20:20], dt_0[21:21], rg_2r);
  AN2EHD I662 (rd_2r1[21:21], dt_0[22:22], rg_2r);
  AN2EHD I663 (rd_2r1[22:22], dt_0[23:23], rg_2r);
  AN2EHD I664 (rd_2r1[23:23], dt_0[24:24], rg_2r);
  AN2EHD I665 (rd_2r1[24:24], dt_0[25:25], rg_2r);
  AN2EHD I666 (rd_2r1[25:25], dt_0[26:26], rg_2r);
  AN2EHD I667 (rd_2r1[26:26], dt_0[27:27], rg_2r);
  AN2EHD I668 (rd_2r1[27:27], dt_0[28:28], rg_2r);
  AN2EHD I669 (rd_2r1[28:28], dt_0[29:29], rg_2r);
  AN2EHD I670 (rd_2r1[29:29], dt_0[30:30], rg_2r);
  AN2EHD I671 (rd_2r1[30:30], dt_0[31:31], rg_2r);
  AN2EHD I672 (rd_3r1[0:0], dt_0[1:1], rg_3r);
  AN2EHD I673 (rd_3r1[1:1], dt_0[2:2], rg_3r);
  AN2EHD I674 (rd_3r1[2:2], dt_0[3:3], rg_3r);
  AN2EHD I675 (rd_3r1[3:3], dt_0[4:4], rg_3r);
  AN2EHD I676 (rd_3r1[4:4], dt_0[5:5], rg_3r);
  AN2EHD I677 (rd_3r1[5:5], dt_0[6:6], rg_3r);
  AN2EHD I678 (rd_3r1[6:6], dt_0[7:7], rg_3r);
  AN2EHD I679 (rd_3r1[7:7], dt_0[8:8], rg_3r);
  AN2EHD I680 (rd_3r1[8:8], dt_0[9:9], rg_3r);
  AN2EHD I681 (rd_3r1[9:9], dt_0[10:10], rg_3r);
  AN2EHD I682 (rd_3r1[10:10], dt_0[11:11], rg_3r);
  AN2EHD I683 (rd_3r1[11:11], dt_0[12:12], rg_3r);
  AN2EHD I684 (rd_3r1[12:12], dt_0[13:13], rg_3r);
  AN2EHD I685 (rd_3r1[13:13], dt_0[14:14], rg_3r);
  AN2EHD I686 (rd_3r1[14:14], dt_0[15:15], rg_3r);
  AN2EHD I687 (rd_3r1[15:15], dt_0[16:16], rg_3r);
  AN2EHD I688 (rd_3r1[16:16], dt_0[17:17], rg_3r);
  AN2EHD I689 (rd_3r1[17:17], dt_0[18:18], rg_3r);
  AN2EHD I690 (rd_3r1[18:18], dt_0[19:19], rg_3r);
  AN2EHD I691 (rd_3r1[19:19], dt_0[20:20], rg_3r);
  AN2EHD I692 (rd_3r1[20:20], dt_0[21:21], rg_3r);
  AN2EHD I693 (rd_3r1[21:21], dt_0[22:22], rg_3r);
  AN2EHD I694 (rd_3r1[22:22], dt_0[23:23], rg_3r);
  AN2EHD I695 (rd_3r1[23:23], dt_0[24:24], rg_3r);
  AN2EHD I696 (rd_3r1[24:24], dt_0[25:25], rg_3r);
  AN2EHD I697 (rd_3r1[25:25], dt_0[26:26], rg_3r);
  AN2EHD I698 (rd_3r1[26:26], dt_0[27:27], rg_3r);
  AN2EHD I699 (rd_3r1[27:27], dt_0[28:28], rg_3r);
  AN2EHD I700 (rd_3r1[28:28], dt_0[29:29], rg_3r);
  AN2EHD I701 (rd_3r1[29:29], dt_0[30:30], rg_3r);
  AN2EHD I702 (rd_3r1[30:30], dt_0[31:31], rg_3r);
  NR3EHD I703 (simp6581_0[0:0], rg_0r, rg_1r, rg_2r);
  NR3EHD I704 (simp6581_0[1:1], rg_3r, rg_0a, rg_1a);
  NR2EHD I705 (simp6581_0[2:2], rg_2a, rg_3a);
  ND3EHD I706 (anyread_0, simp6581_0[0:0], simp6581_0[1:1], simp6581_0[2:2]);
  BUFEHD I707 (wg_0a, wd_0a);
  BUFEHD I708 (rg_0a, rd_0a);
  BUFEHD I709 (rg_1a, rd_1a);
  BUFEHD I710 (rg_2a, rd_2a);
  BUFEHD I711 (rg_3a, rd_3a);
endmodule

// tko30m32_1nm2b0_2apt1o0w2bi0w30b TeakO [
//     (1,TeakOConstant 2 0),
//     (2,TeakOAppend 1 [(1,0+:2),(0,0+:30)])] [One 30,One 32]
module tko30m32_1nm2b0_2apt1o0w2bi0w30b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [29:0] i_0r0;
  input [29:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [29:0] gocomp_0;
  wire [9:0] simp321_0;
  wire tech33_int;
  wire tech34_int;
  wire tech35_int;
  wire tech36_int;
  wire tech37_int;
  wire tech38_int;
  wire tech39_int;
  wire tech40_int;
  wire tech41_int;
  wire tech42_int;
  wire [3:0] simp322_0;
  wire tech44_int;
  wire tech45_int;
  wire tech46_int;
  wire [1:0] simp323_0;
  wire tech49_int;
  wire [1:0] termf_1;
  wire [1:0] termt_1;
  OR2EHD I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2EHD I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2EHD I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2EHD I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2EHD I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2EHD I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2EHD I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2EHD I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2EHD I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2EHD I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2EHD I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2EHD I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2EHD I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2EHD I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2EHD I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2EHD I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2EHD I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2EHD I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2EHD I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2EHD I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2EHD I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2EHD I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2EHD I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2EHD I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2EHD I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2EHD I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2EHD I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2EHD I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2EHD I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2EHD I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  AO222EHD I30 (tech33_int, gocomp_0[0:0], gocomp_0[1:1], tech33_int, gocomp_0[0:0], tech33_int, gocomp_0[1:1]);
  AO222EHD I31 (simp321_0[0:0], tech33_int, gocomp_0[2:2], simp321_0[0:0], tech33_int, simp321_0[0:0], gocomp_0[2:2]);
  AO222EHD I32 (tech34_int, gocomp_0[3:3], gocomp_0[4:4], tech34_int, gocomp_0[3:3], tech34_int, gocomp_0[4:4]);
  AO222EHD I33 (simp321_0[1:1], tech34_int, gocomp_0[5:5], simp321_0[1:1], tech34_int, simp321_0[1:1], gocomp_0[5:5]);
  AO222EHD I34 (tech35_int, gocomp_0[6:6], gocomp_0[7:7], tech35_int, gocomp_0[6:6], tech35_int, gocomp_0[7:7]);
  AO222EHD I35 (simp321_0[2:2], tech35_int, gocomp_0[8:8], simp321_0[2:2], tech35_int, simp321_0[2:2], gocomp_0[8:8]);
  AO222EHD I36 (tech36_int, gocomp_0[9:9], gocomp_0[10:10], tech36_int, gocomp_0[9:9], tech36_int, gocomp_0[10:10]);
  AO222EHD I37 (simp321_0[3:3], tech36_int, gocomp_0[11:11], simp321_0[3:3], tech36_int, simp321_0[3:3], gocomp_0[11:11]);
  AO222EHD I38 (tech37_int, gocomp_0[12:12], gocomp_0[13:13], tech37_int, gocomp_0[12:12], tech37_int, gocomp_0[13:13]);
  AO222EHD I39 (simp321_0[4:4], tech37_int, gocomp_0[14:14], simp321_0[4:4], tech37_int, simp321_0[4:4], gocomp_0[14:14]);
  AO222EHD I40 (tech38_int, gocomp_0[15:15], gocomp_0[16:16], tech38_int, gocomp_0[15:15], tech38_int, gocomp_0[16:16]);
  AO222EHD I41 (simp321_0[5:5], tech38_int, gocomp_0[17:17], simp321_0[5:5], tech38_int, simp321_0[5:5], gocomp_0[17:17]);
  AO222EHD I42 (tech39_int, gocomp_0[18:18], gocomp_0[19:19], tech39_int, gocomp_0[18:18], tech39_int, gocomp_0[19:19]);
  AO222EHD I43 (simp321_0[6:6], tech39_int, gocomp_0[20:20], simp321_0[6:6], tech39_int, simp321_0[6:6], gocomp_0[20:20]);
  AO222EHD I44 (tech40_int, gocomp_0[21:21], gocomp_0[22:22], tech40_int, gocomp_0[21:21], tech40_int, gocomp_0[22:22]);
  AO222EHD I45 (simp321_0[7:7], tech40_int, gocomp_0[23:23], simp321_0[7:7], tech40_int, simp321_0[7:7], gocomp_0[23:23]);
  AO222EHD I46 (tech41_int, gocomp_0[24:24], gocomp_0[25:25], tech41_int, gocomp_0[24:24], tech41_int, gocomp_0[25:25]);
  AO222EHD I47 (simp321_0[8:8], tech41_int, gocomp_0[26:26], simp321_0[8:8], tech41_int, simp321_0[8:8], gocomp_0[26:26]);
  AO222EHD I48 (tech42_int, gocomp_0[27:27], gocomp_0[28:28], tech42_int, gocomp_0[27:27], tech42_int, gocomp_0[28:28]);
  AO222EHD I49 (simp321_0[9:9], tech42_int, gocomp_0[29:29], simp321_0[9:9], tech42_int, simp321_0[9:9], gocomp_0[29:29]);
  AO222EHD I50 (tech44_int, simp321_0[0:0], simp321_0[1:1], tech44_int, simp321_0[0:0], tech44_int, simp321_0[1:1]);
  AO222EHD I51 (simp322_0[0:0], tech44_int, simp321_0[2:2], simp322_0[0:0], tech44_int, simp322_0[0:0], simp321_0[2:2]);
  AO222EHD I52 (tech45_int, simp321_0[3:3], simp321_0[4:4], tech45_int, simp321_0[3:3], tech45_int, simp321_0[4:4]);
  AO222EHD I53 (simp322_0[1:1], tech45_int, simp321_0[5:5], simp322_0[1:1], tech45_int, simp322_0[1:1], simp321_0[5:5]);
  AO222EHD I54 (tech46_int, simp321_0[6:6], simp321_0[7:7], tech46_int, simp321_0[6:6], tech46_int, simp321_0[7:7]);
  AO222EHD I55 (simp322_0[2:2], tech46_int, simp321_0[8:8], simp322_0[2:2], tech46_int, simp322_0[2:2], simp321_0[8:8]);
  BUFEHD I56 (simp322_0[3:3], simp321_0[9:9]);
  AO222EHD I57 (tech49_int, simp322_0[0:0], simp322_0[1:1], tech49_int, simp322_0[0:0], tech49_int, simp322_0[1:1]);
  AO222EHD I58 (simp323_0[0:0], tech49_int, simp322_0[2:2], simp323_0[0:0], tech49_int, simp323_0[0:0], simp322_0[2:2]);
  BUFEHD I59 (simp323_0[1:1], simp322_0[3:3]);
  AO222EHD I60 (go_0, simp323_0[0:0], simp323_0[1:1], go_0, simp323_0[0:0], go_0, simp323_0[1:1]);
  BUFEHD I61 (termf_1[0:0], go_0);
  BUFEHD I62 (termf_1[1:1], go_0);
  TIE0DND I63 (termt_1[0:0]);
  TIE0DND I64 (termt_1[1:1]);
  BUFEHD I65 (o_0r0[0:0], termf_1[0:0]);
  BUFEHD I66 (o_0r0[1:1], termf_1[1:1]);
  BUFEHD I67 (o_0r0[2:2], i_0r0[0:0]);
  BUFEHD I68 (o_0r0[3:3], i_0r0[1:1]);
  BUFEHD I69 (o_0r0[4:4], i_0r0[2:2]);
  BUFEHD I70 (o_0r0[5:5], i_0r0[3:3]);
  BUFEHD I71 (o_0r0[6:6], i_0r0[4:4]);
  BUFEHD I72 (o_0r0[7:7], i_0r0[5:5]);
  BUFEHD I73 (o_0r0[8:8], i_0r0[6:6]);
  BUFEHD I74 (o_0r0[9:9], i_0r0[7:7]);
  BUFEHD I75 (o_0r0[10:10], i_0r0[8:8]);
  BUFEHD I76 (o_0r0[11:11], i_0r0[9:9]);
  BUFEHD I77 (o_0r0[12:12], i_0r0[10:10]);
  BUFEHD I78 (o_0r0[13:13], i_0r0[11:11]);
  BUFEHD I79 (o_0r0[14:14], i_0r0[12:12]);
  BUFEHD I80 (o_0r0[15:15], i_0r0[13:13]);
  BUFEHD I81 (o_0r0[16:16], i_0r0[14:14]);
  BUFEHD I82 (o_0r0[17:17], i_0r0[15:15]);
  BUFEHD I83 (o_0r0[18:18], i_0r0[16:16]);
  BUFEHD I84 (o_0r0[19:19], i_0r0[17:17]);
  BUFEHD I85 (o_0r0[20:20], i_0r0[18:18]);
  BUFEHD I86 (o_0r0[21:21], i_0r0[19:19]);
  BUFEHD I87 (o_0r0[22:22], i_0r0[20:20]);
  BUFEHD I88 (o_0r0[23:23], i_0r0[21:21]);
  BUFEHD I89 (o_0r0[24:24], i_0r0[22:22]);
  BUFEHD I90 (o_0r0[25:25], i_0r0[23:23]);
  BUFEHD I91 (o_0r0[26:26], i_0r0[24:24]);
  BUFEHD I92 (o_0r0[27:27], i_0r0[25:25]);
  BUFEHD I93 (o_0r0[28:28], i_0r0[26:26]);
  BUFEHD I94 (o_0r0[29:29], i_0r0[27:27]);
  BUFEHD I95 (o_0r0[30:30], i_0r0[28:28]);
  BUFEHD I96 (o_0r0[31:31], i_0r0[29:29]);
  BUFEHD I97 (o_0r1[0:0], termt_1[0:0]);
  BUFEHD I98 (o_0r1[1:1], termt_1[1:1]);
  BUFEHD I99 (o_0r1[2:2], i_0r1[0:0]);
  BUFEHD I100 (o_0r1[3:3], i_0r1[1:1]);
  BUFEHD I101 (o_0r1[4:4], i_0r1[2:2]);
  BUFEHD I102 (o_0r1[5:5], i_0r1[3:3]);
  BUFEHD I103 (o_0r1[6:6], i_0r1[4:4]);
  BUFEHD I104 (o_0r1[7:7], i_0r1[5:5]);
  BUFEHD I105 (o_0r1[8:8], i_0r1[6:6]);
  BUFEHD I106 (o_0r1[9:9], i_0r1[7:7]);
  BUFEHD I107 (o_0r1[10:10], i_0r1[8:8]);
  BUFEHD I108 (o_0r1[11:11], i_0r1[9:9]);
  BUFEHD I109 (o_0r1[12:12], i_0r1[10:10]);
  BUFEHD I110 (o_0r1[13:13], i_0r1[11:11]);
  BUFEHD I111 (o_0r1[14:14], i_0r1[12:12]);
  BUFEHD I112 (o_0r1[15:15], i_0r1[13:13]);
  BUFEHD I113 (o_0r1[16:16], i_0r1[14:14]);
  BUFEHD I114 (o_0r1[17:17], i_0r1[15:15]);
  BUFEHD I115 (o_0r1[18:18], i_0r1[16:16]);
  BUFEHD I116 (o_0r1[19:19], i_0r1[17:17]);
  BUFEHD I117 (o_0r1[20:20], i_0r1[18:18]);
  BUFEHD I118 (o_0r1[21:21], i_0r1[19:19]);
  BUFEHD I119 (o_0r1[22:22], i_0r1[20:20]);
  BUFEHD I120 (o_0r1[23:23], i_0r1[21:21]);
  BUFEHD I121 (o_0r1[24:24], i_0r1[22:22]);
  BUFEHD I122 (o_0r1[25:25], i_0r1[23:23]);
  BUFEHD I123 (o_0r1[26:26], i_0r1[24:24]);
  BUFEHD I124 (o_0r1[27:27], i_0r1[25:25]);
  BUFEHD I125 (o_0r1[28:28], i_0r1[26:26]);
  BUFEHD I126 (o_0r1[29:29], i_0r1[27:27]);
  BUFEHD I127 (o_0r1[30:30], i_0r1[28:28]);
  BUFEHD I128 (o_0r1[31:31], i_0r1[29:29]);
  BUFEHD I129 (i_0a, o_0a);
endmodule

// tko30m32_1nm2b0_2api0w30bt1o0w2b TeakO [
//     (1,TeakOConstant 2 0),
//     (2,TeakOAppend 1 [(0,0+:30),(1,0+:2)])] [One 30,One 32]
module tko30m32_1nm2b0_2api0w30bt1o0w2b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [29:0] i_0r0;
  input [29:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [29:0] gocomp_0;
  wire [9:0] simp321_0;
  wire tech33_int;
  wire tech34_int;
  wire tech35_int;
  wire tech36_int;
  wire tech37_int;
  wire tech38_int;
  wire tech39_int;
  wire tech40_int;
  wire tech41_int;
  wire tech42_int;
  wire [3:0] simp322_0;
  wire tech44_int;
  wire tech45_int;
  wire tech46_int;
  wire [1:0] simp323_0;
  wire tech49_int;
  wire [1:0] termf_1;
  wire [1:0] termt_1;
  OR2EHD I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2EHD I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2EHD I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2EHD I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2EHD I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2EHD I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2EHD I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2EHD I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2EHD I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2EHD I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2EHD I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2EHD I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2EHD I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2EHD I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2EHD I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2EHD I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2EHD I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2EHD I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2EHD I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2EHD I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2EHD I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2EHD I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2EHD I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2EHD I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2EHD I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2EHD I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2EHD I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2EHD I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2EHD I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2EHD I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  AO222EHD I30 (tech33_int, gocomp_0[0:0], gocomp_0[1:1], tech33_int, gocomp_0[0:0], tech33_int, gocomp_0[1:1]);
  AO222EHD I31 (simp321_0[0:0], tech33_int, gocomp_0[2:2], simp321_0[0:0], tech33_int, simp321_0[0:0], gocomp_0[2:2]);
  AO222EHD I32 (tech34_int, gocomp_0[3:3], gocomp_0[4:4], tech34_int, gocomp_0[3:3], tech34_int, gocomp_0[4:4]);
  AO222EHD I33 (simp321_0[1:1], tech34_int, gocomp_0[5:5], simp321_0[1:1], tech34_int, simp321_0[1:1], gocomp_0[5:5]);
  AO222EHD I34 (tech35_int, gocomp_0[6:6], gocomp_0[7:7], tech35_int, gocomp_0[6:6], tech35_int, gocomp_0[7:7]);
  AO222EHD I35 (simp321_0[2:2], tech35_int, gocomp_0[8:8], simp321_0[2:2], tech35_int, simp321_0[2:2], gocomp_0[8:8]);
  AO222EHD I36 (tech36_int, gocomp_0[9:9], gocomp_0[10:10], tech36_int, gocomp_0[9:9], tech36_int, gocomp_0[10:10]);
  AO222EHD I37 (simp321_0[3:3], tech36_int, gocomp_0[11:11], simp321_0[3:3], tech36_int, simp321_0[3:3], gocomp_0[11:11]);
  AO222EHD I38 (tech37_int, gocomp_0[12:12], gocomp_0[13:13], tech37_int, gocomp_0[12:12], tech37_int, gocomp_0[13:13]);
  AO222EHD I39 (simp321_0[4:4], tech37_int, gocomp_0[14:14], simp321_0[4:4], tech37_int, simp321_0[4:4], gocomp_0[14:14]);
  AO222EHD I40 (tech38_int, gocomp_0[15:15], gocomp_0[16:16], tech38_int, gocomp_0[15:15], tech38_int, gocomp_0[16:16]);
  AO222EHD I41 (simp321_0[5:5], tech38_int, gocomp_0[17:17], simp321_0[5:5], tech38_int, simp321_0[5:5], gocomp_0[17:17]);
  AO222EHD I42 (tech39_int, gocomp_0[18:18], gocomp_0[19:19], tech39_int, gocomp_0[18:18], tech39_int, gocomp_0[19:19]);
  AO222EHD I43 (simp321_0[6:6], tech39_int, gocomp_0[20:20], simp321_0[6:6], tech39_int, simp321_0[6:6], gocomp_0[20:20]);
  AO222EHD I44 (tech40_int, gocomp_0[21:21], gocomp_0[22:22], tech40_int, gocomp_0[21:21], tech40_int, gocomp_0[22:22]);
  AO222EHD I45 (simp321_0[7:7], tech40_int, gocomp_0[23:23], simp321_0[7:7], tech40_int, simp321_0[7:7], gocomp_0[23:23]);
  AO222EHD I46 (tech41_int, gocomp_0[24:24], gocomp_0[25:25], tech41_int, gocomp_0[24:24], tech41_int, gocomp_0[25:25]);
  AO222EHD I47 (simp321_0[8:8], tech41_int, gocomp_0[26:26], simp321_0[8:8], tech41_int, simp321_0[8:8], gocomp_0[26:26]);
  AO222EHD I48 (tech42_int, gocomp_0[27:27], gocomp_0[28:28], tech42_int, gocomp_0[27:27], tech42_int, gocomp_0[28:28]);
  AO222EHD I49 (simp321_0[9:9], tech42_int, gocomp_0[29:29], simp321_0[9:9], tech42_int, simp321_0[9:9], gocomp_0[29:29]);
  AO222EHD I50 (tech44_int, simp321_0[0:0], simp321_0[1:1], tech44_int, simp321_0[0:0], tech44_int, simp321_0[1:1]);
  AO222EHD I51 (simp322_0[0:0], tech44_int, simp321_0[2:2], simp322_0[0:0], tech44_int, simp322_0[0:0], simp321_0[2:2]);
  AO222EHD I52 (tech45_int, simp321_0[3:3], simp321_0[4:4], tech45_int, simp321_0[3:3], tech45_int, simp321_0[4:4]);
  AO222EHD I53 (simp322_0[1:1], tech45_int, simp321_0[5:5], simp322_0[1:1], tech45_int, simp322_0[1:1], simp321_0[5:5]);
  AO222EHD I54 (tech46_int, simp321_0[6:6], simp321_0[7:7], tech46_int, simp321_0[6:6], tech46_int, simp321_0[7:7]);
  AO222EHD I55 (simp322_0[2:2], tech46_int, simp321_0[8:8], simp322_0[2:2], tech46_int, simp322_0[2:2], simp321_0[8:8]);
  BUFEHD I56 (simp322_0[3:3], simp321_0[9:9]);
  AO222EHD I57 (tech49_int, simp322_0[0:0], simp322_0[1:1], tech49_int, simp322_0[0:0], tech49_int, simp322_0[1:1]);
  AO222EHD I58 (simp323_0[0:0], tech49_int, simp322_0[2:2], simp323_0[0:0], tech49_int, simp323_0[0:0], simp322_0[2:2]);
  BUFEHD I59 (simp323_0[1:1], simp322_0[3:3]);
  AO222EHD I60 (go_0, simp323_0[0:0], simp323_0[1:1], go_0, simp323_0[0:0], go_0, simp323_0[1:1]);
  BUFEHD I61 (termf_1[0:0], go_0);
  BUFEHD I62 (termf_1[1:1], go_0);
  TIE0DND I63 (termt_1[0:0]);
  TIE0DND I64 (termt_1[1:1]);
  BUFEHD I65 (o_0r0[0:0], i_0r0[0:0]);
  BUFEHD I66 (o_0r0[1:1], i_0r0[1:1]);
  BUFEHD I67 (o_0r0[2:2], i_0r0[2:2]);
  BUFEHD I68 (o_0r0[3:3], i_0r0[3:3]);
  BUFEHD I69 (o_0r0[4:4], i_0r0[4:4]);
  BUFEHD I70 (o_0r0[5:5], i_0r0[5:5]);
  BUFEHD I71 (o_0r0[6:6], i_0r0[6:6]);
  BUFEHD I72 (o_0r0[7:7], i_0r0[7:7]);
  BUFEHD I73 (o_0r0[8:8], i_0r0[8:8]);
  BUFEHD I74 (o_0r0[9:9], i_0r0[9:9]);
  BUFEHD I75 (o_0r0[10:10], i_0r0[10:10]);
  BUFEHD I76 (o_0r0[11:11], i_0r0[11:11]);
  BUFEHD I77 (o_0r0[12:12], i_0r0[12:12]);
  BUFEHD I78 (o_0r0[13:13], i_0r0[13:13]);
  BUFEHD I79 (o_0r0[14:14], i_0r0[14:14]);
  BUFEHD I80 (o_0r0[15:15], i_0r0[15:15]);
  BUFEHD I81 (o_0r0[16:16], i_0r0[16:16]);
  BUFEHD I82 (o_0r0[17:17], i_0r0[17:17]);
  BUFEHD I83 (o_0r0[18:18], i_0r0[18:18]);
  BUFEHD I84 (o_0r0[19:19], i_0r0[19:19]);
  BUFEHD I85 (o_0r0[20:20], i_0r0[20:20]);
  BUFEHD I86 (o_0r0[21:21], i_0r0[21:21]);
  BUFEHD I87 (o_0r0[22:22], i_0r0[22:22]);
  BUFEHD I88 (o_0r0[23:23], i_0r0[23:23]);
  BUFEHD I89 (o_0r0[24:24], i_0r0[24:24]);
  BUFEHD I90 (o_0r0[25:25], i_0r0[25:25]);
  BUFEHD I91 (o_0r0[26:26], i_0r0[26:26]);
  BUFEHD I92 (o_0r0[27:27], i_0r0[27:27]);
  BUFEHD I93 (o_0r0[28:28], i_0r0[28:28]);
  BUFEHD I94 (o_0r0[29:29], i_0r0[29:29]);
  BUFEHD I95 (o_0r0[30:30], termf_1[0:0]);
  BUFEHD I96 (o_0r0[31:31], termf_1[1:1]);
  BUFEHD I97 (o_0r1[0:0], i_0r1[0:0]);
  BUFEHD I98 (o_0r1[1:1], i_0r1[1:1]);
  BUFEHD I99 (o_0r1[2:2], i_0r1[2:2]);
  BUFEHD I100 (o_0r1[3:3], i_0r1[3:3]);
  BUFEHD I101 (o_0r1[4:4], i_0r1[4:4]);
  BUFEHD I102 (o_0r1[5:5], i_0r1[5:5]);
  BUFEHD I103 (o_0r1[6:6], i_0r1[6:6]);
  BUFEHD I104 (o_0r1[7:7], i_0r1[7:7]);
  BUFEHD I105 (o_0r1[8:8], i_0r1[8:8]);
  BUFEHD I106 (o_0r1[9:9], i_0r1[9:9]);
  BUFEHD I107 (o_0r1[10:10], i_0r1[10:10]);
  BUFEHD I108 (o_0r1[11:11], i_0r1[11:11]);
  BUFEHD I109 (o_0r1[12:12], i_0r1[12:12]);
  BUFEHD I110 (o_0r1[13:13], i_0r1[13:13]);
  BUFEHD I111 (o_0r1[14:14], i_0r1[14:14]);
  BUFEHD I112 (o_0r1[15:15], i_0r1[15:15]);
  BUFEHD I113 (o_0r1[16:16], i_0r1[16:16]);
  BUFEHD I114 (o_0r1[17:17], i_0r1[17:17]);
  BUFEHD I115 (o_0r1[18:18], i_0r1[18:18]);
  BUFEHD I116 (o_0r1[19:19], i_0r1[19:19]);
  BUFEHD I117 (o_0r1[20:20], i_0r1[20:20]);
  BUFEHD I118 (o_0r1[21:21], i_0r1[21:21]);
  BUFEHD I119 (o_0r1[22:22], i_0r1[22:22]);
  BUFEHD I120 (o_0r1[23:23], i_0r1[23:23]);
  BUFEHD I121 (o_0r1[24:24], i_0r1[24:24]);
  BUFEHD I122 (o_0r1[25:25], i_0r1[25:25]);
  BUFEHD I123 (o_0r1[26:26], i_0r1[26:26]);
  BUFEHD I124 (o_0r1[27:27], i_0r1[27:27]);
  BUFEHD I125 (o_0r1[28:28], i_0r1[28:28]);
  BUFEHD I126 (o_0r1[29:29], i_0r1[29:29]);
  BUFEHD I127 (o_0r1[30:30], termt_1[0:0]);
  BUFEHD I128 (o_0r1[31:31], termt_1[1:1]);
  BUFEHD I129 (i_0a, o_0a);
endmodule

// tko30m32_1nm2b3_2api0w30bt1o0w2b TeakO [
//     (1,TeakOConstant 2 3),
//     (2,TeakOAppend 1 [(0,0+:30),(1,0+:2)])] [One 30,One 32]
module tko30m32_1nm2b3_2api0w30bt1o0w2b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [29:0] i_0r0;
  input [29:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [29:0] gocomp_0;
  wire [9:0] simp321_0;
  wire tech33_int;
  wire tech34_int;
  wire tech35_int;
  wire tech36_int;
  wire tech37_int;
  wire tech38_int;
  wire tech39_int;
  wire tech40_int;
  wire tech41_int;
  wire tech42_int;
  wire [3:0] simp322_0;
  wire tech44_int;
  wire tech45_int;
  wire tech46_int;
  wire [1:0] simp323_0;
  wire tech49_int;
  wire [1:0] termf_1;
  wire [1:0] termt_1;
  OR2EHD I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2EHD I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2EHD I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2EHD I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2EHD I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2EHD I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2EHD I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2EHD I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2EHD I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2EHD I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2EHD I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2EHD I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2EHD I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2EHD I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2EHD I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2EHD I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2EHD I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2EHD I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2EHD I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2EHD I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2EHD I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2EHD I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2EHD I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2EHD I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2EHD I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2EHD I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2EHD I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2EHD I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2EHD I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2EHD I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  AO222EHD I30 (tech33_int, gocomp_0[0:0], gocomp_0[1:1], tech33_int, gocomp_0[0:0], tech33_int, gocomp_0[1:1]);
  AO222EHD I31 (simp321_0[0:0], tech33_int, gocomp_0[2:2], simp321_0[0:0], tech33_int, simp321_0[0:0], gocomp_0[2:2]);
  AO222EHD I32 (tech34_int, gocomp_0[3:3], gocomp_0[4:4], tech34_int, gocomp_0[3:3], tech34_int, gocomp_0[4:4]);
  AO222EHD I33 (simp321_0[1:1], tech34_int, gocomp_0[5:5], simp321_0[1:1], tech34_int, simp321_0[1:1], gocomp_0[5:5]);
  AO222EHD I34 (tech35_int, gocomp_0[6:6], gocomp_0[7:7], tech35_int, gocomp_0[6:6], tech35_int, gocomp_0[7:7]);
  AO222EHD I35 (simp321_0[2:2], tech35_int, gocomp_0[8:8], simp321_0[2:2], tech35_int, simp321_0[2:2], gocomp_0[8:8]);
  AO222EHD I36 (tech36_int, gocomp_0[9:9], gocomp_0[10:10], tech36_int, gocomp_0[9:9], tech36_int, gocomp_0[10:10]);
  AO222EHD I37 (simp321_0[3:3], tech36_int, gocomp_0[11:11], simp321_0[3:3], tech36_int, simp321_0[3:3], gocomp_0[11:11]);
  AO222EHD I38 (tech37_int, gocomp_0[12:12], gocomp_0[13:13], tech37_int, gocomp_0[12:12], tech37_int, gocomp_0[13:13]);
  AO222EHD I39 (simp321_0[4:4], tech37_int, gocomp_0[14:14], simp321_0[4:4], tech37_int, simp321_0[4:4], gocomp_0[14:14]);
  AO222EHD I40 (tech38_int, gocomp_0[15:15], gocomp_0[16:16], tech38_int, gocomp_0[15:15], tech38_int, gocomp_0[16:16]);
  AO222EHD I41 (simp321_0[5:5], tech38_int, gocomp_0[17:17], simp321_0[5:5], tech38_int, simp321_0[5:5], gocomp_0[17:17]);
  AO222EHD I42 (tech39_int, gocomp_0[18:18], gocomp_0[19:19], tech39_int, gocomp_0[18:18], tech39_int, gocomp_0[19:19]);
  AO222EHD I43 (simp321_0[6:6], tech39_int, gocomp_0[20:20], simp321_0[6:6], tech39_int, simp321_0[6:6], gocomp_0[20:20]);
  AO222EHD I44 (tech40_int, gocomp_0[21:21], gocomp_0[22:22], tech40_int, gocomp_0[21:21], tech40_int, gocomp_0[22:22]);
  AO222EHD I45 (simp321_0[7:7], tech40_int, gocomp_0[23:23], simp321_0[7:7], tech40_int, simp321_0[7:7], gocomp_0[23:23]);
  AO222EHD I46 (tech41_int, gocomp_0[24:24], gocomp_0[25:25], tech41_int, gocomp_0[24:24], tech41_int, gocomp_0[25:25]);
  AO222EHD I47 (simp321_0[8:8], tech41_int, gocomp_0[26:26], simp321_0[8:8], tech41_int, simp321_0[8:8], gocomp_0[26:26]);
  AO222EHD I48 (tech42_int, gocomp_0[27:27], gocomp_0[28:28], tech42_int, gocomp_0[27:27], tech42_int, gocomp_0[28:28]);
  AO222EHD I49 (simp321_0[9:9], tech42_int, gocomp_0[29:29], simp321_0[9:9], tech42_int, simp321_0[9:9], gocomp_0[29:29]);
  AO222EHD I50 (tech44_int, simp321_0[0:0], simp321_0[1:1], tech44_int, simp321_0[0:0], tech44_int, simp321_0[1:1]);
  AO222EHD I51 (simp322_0[0:0], tech44_int, simp321_0[2:2], simp322_0[0:0], tech44_int, simp322_0[0:0], simp321_0[2:2]);
  AO222EHD I52 (tech45_int, simp321_0[3:3], simp321_0[4:4], tech45_int, simp321_0[3:3], tech45_int, simp321_0[4:4]);
  AO222EHD I53 (simp322_0[1:1], tech45_int, simp321_0[5:5], simp322_0[1:1], tech45_int, simp322_0[1:1], simp321_0[5:5]);
  AO222EHD I54 (tech46_int, simp321_0[6:6], simp321_0[7:7], tech46_int, simp321_0[6:6], tech46_int, simp321_0[7:7]);
  AO222EHD I55 (simp322_0[2:2], tech46_int, simp321_0[8:8], simp322_0[2:2], tech46_int, simp322_0[2:2], simp321_0[8:8]);
  BUFEHD I56 (simp322_0[3:3], simp321_0[9:9]);
  AO222EHD I57 (tech49_int, simp322_0[0:0], simp322_0[1:1], tech49_int, simp322_0[0:0], tech49_int, simp322_0[1:1]);
  AO222EHD I58 (simp323_0[0:0], tech49_int, simp322_0[2:2], simp323_0[0:0], tech49_int, simp323_0[0:0], simp322_0[2:2]);
  BUFEHD I59 (simp323_0[1:1], simp322_0[3:3]);
  AO222EHD I60 (go_0, simp323_0[0:0], simp323_0[1:1], go_0, simp323_0[0:0], go_0, simp323_0[1:1]);
  BUFEHD I61 (termt_1[0:0], go_0);
  BUFEHD I62 (termt_1[1:1], go_0);
  TIE0DND I63 (termf_1[0:0]);
  TIE0DND I64 (termf_1[1:1]);
  BUFEHD I65 (o_0r0[0:0], i_0r0[0:0]);
  BUFEHD I66 (o_0r0[1:1], i_0r0[1:1]);
  BUFEHD I67 (o_0r0[2:2], i_0r0[2:2]);
  BUFEHD I68 (o_0r0[3:3], i_0r0[3:3]);
  BUFEHD I69 (o_0r0[4:4], i_0r0[4:4]);
  BUFEHD I70 (o_0r0[5:5], i_0r0[5:5]);
  BUFEHD I71 (o_0r0[6:6], i_0r0[6:6]);
  BUFEHD I72 (o_0r0[7:7], i_0r0[7:7]);
  BUFEHD I73 (o_0r0[8:8], i_0r0[8:8]);
  BUFEHD I74 (o_0r0[9:9], i_0r0[9:9]);
  BUFEHD I75 (o_0r0[10:10], i_0r0[10:10]);
  BUFEHD I76 (o_0r0[11:11], i_0r0[11:11]);
  BUFEHD I77 (o_0r0[12:12], i_0r0[12:12]);
  BUFEHD I78 (o_0r0[13:13], i_0r0[13:13]);
  BUFEHD I79 (o_0r0[14:14], i_0r0[14:14]);
  BUFEHD I80 (o_0r0[15:15], i_0r0[15:15]);
  BUFEHD I81 (o_0r0[16:16], i_0r0[16:16]);
  BUFEHD I82 (o_0r0[17:17], i_0r0[17:17]);
  BUFEHD I83 (o_0r0[18:18], i_0r0[18:18]);
  BUFEHD I84 (o_0r0[19:19], i_0r0[19:19]);
  BUFEHD I85 (o_0r0[20:20], i_0r0[20:20]);
  BUFEHD I86 (o_0r0[21:21], i_0r0[21:21]);
  BUFEHD I87 (o_0r0[22:22], i_0r0[22:22]);
  BUFEHD I88 (o_0r0[23:23], i_0r0[23:23]);
  BUFEHD I89 (o_0r0[24:24], i_0r0[24:24]);
  BUFEHD I90 (o_0r0[25:25], i_0r0[25:25]);
  BUFEHD I91 (o_0r0[26:26], i_0r0[26:26]);
  BUFEHD I92 (o_0r0[27:27], i_0r0[27:27]);
  BUFEHD I93 (o_0r0[28:28], i_0r0[28:28]);
  BUFEHD I94 (o_0r0[29:29], i_0r0[29:29]);
  BUFEHD I95 (o_0r0[30:30], termf_1[0:0]);
  BUFEHD I96 (o_0r0[31:31], termf_1[1:1]);
  BUFEHD I97 (o_0r1[0:0], i_0r1[0:0]);
  BUFEHD I98 (o_0r1[1:1], i_0r1[1:1]);
  BUFEHD I99 (o_0r1[2:2], i_0r1[2:2]);
  BUFEHD I100 (o_0r1[3:3], i_0r1[3:3]);
  BUFEHD I101 (o_0r1[4:4], i_0r1[4:4]);
  BUFEHD I102 (o_0r1[5:5], i_0r1[5:5]);
  BUFEHD I103 (o_0r1[6:6], i_0r1[6:6]);
  BUFEHD I104 (o_0r1[7:7], i_0r1[7:7]);
  BUFEHD I105 (o_0r1[8:8], i_0r1[8:8]);
  BUFEHD I106 (o_0r1[9:9], i_0r1[9:9]);
  BUFEHD I107 (o_0r1[10:10], i_0r1[10:10]);
  BUFEHD I108 (o_0r1[11:11], i_0r1[11:11]);
  BUFEHD I109 (o_0r1[12:12], i_0r1[12:12]);
  BUFEHD I110 (o_0r1[13:13], i_0r1[13:13]);
  BUFEHD I111 (o_0r1[14:14], i_0r1[14:14]);
  BUFEHD I112 (o_0r1[15:15], i_0r1[15:15]);
  BUFEHD I113 (o_0r1[16:16], i_0r1[16:16]);
  BUFEHD I114 (o_0r1[17:17], i_0r1[17:17]);
  BUFEHD I115 (o_0r1[18:18], i_0r1[18:18]);
  BUFEHD I116 (o_0r1[19:19], i_0r1[19:19]);
  BUFEHD I117 (o_0r1[20:20], i_0r1[20:20]);
  BUFEHD I118 (o_0r1[21:21], i_0r1[21:21]);
  BUFEHD I119 (o_0r1[22:22], i_0r1[22:22]);
  BUFEHD I120 (o_0r1[23:23], i_0r1[23:23]);
  BUFEHD I121 (o_0r1[24:24], i_0r1[24:24]);
  BUFEHD I122 (o_0r1[25:25], i_0r1[25:25]);
  BUFEHD I123 (o_0r1[26:26], i_0r1[26:26]);
  BUFEHD I124 (o_0r1[27:27], i_0r1[27:27]);
  BUFEHD I125 (o_0r1[28:28], i_0r1[28:28]);
  BUFEHD I126 (o_0r1[29:29], i_0r1[29:29]);
  BUFEHD I127 (o_0r1[30:30], termt_1[0:0]);
  BUFEHD I128 (o_0r1[31:31], termt_1[1:1]);
  BUFEHD I129 (i_0a, o_0a);
endmodule

// tkvi32_wo0w32_ro0w32o0w30o2w30o2w30 TeakV "i" 32 [] [0] [0,0,2,2] [Many [32],Many [0],Many [0,0,0,0]
//   ,Many [32,30,30,30]]
module tkvi32_wo0w32_ro0w32o0w30o2w30o2w30 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [29:0] rd_1r0;
  output [29:0] rd_1r1;
  input rd_1a;
  output [29:0] rd_2r0;
  output [29:0] rd_2r1;
  input rd_2a;
  output [29:0] rd_3r0;
  output [29:0] rd_3r1;
  input rd_3a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire tech239_int;
  wire tech240_int;
  wire tech241_int;
  wire tech242_int;
  wire tech243_int;
  wire tech244_int;
  wire tech245_int;
  wire tech246_int;
  wire tech247_int;
  wire tech248_int;
  wire [3:0] simp2382_0;
  wire tech251_int;
  wire tech252_int;
  wire tech253_int;
  wire [1:0] simp2383_0;
  wire tech256_int;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire tech428_int;
  wire tech429_int;
  wire tech430_int;
  wire tech431_int;
  wire tech432_int;
  wire tech433_int;
  wire tech434_int;
  wire tech435_int;
  wire tech436_int;
  wire tech437_int;
  wire tech438_int;
  wire [3:0] simp4072_0;
  wire tech440_int;
  wire tech441_int;
  wire tech442_int;
  wire [1:0] simp4073_0;
  wire tech445_int;
  wire [2:0] simp6521_0;
  INVHHD I0 (nreset_0, reset);
  AN2EHD I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AN2EHD I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AN2EHD I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AN2EHD I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AN2EHD I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AN2EHD I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AN2EHD I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AN2EHD I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AN2EHD I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AN2EHD I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AN2EHD I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AN2EHD I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AN2EHD I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AN2EHD I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AN2EHD I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AN2EHD I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AN2EHD I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AN2EHD I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AN2EHD I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AN2EHD I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AN2EHD I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AN2EHD I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AN2EHD I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AN2EHD I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AN2EHD I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AN2EHD I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AN2EHD I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AN2EHD I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AN2EHD I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AN2EHD I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AN2EHD I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AN2EHD I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AN2EHD I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AN2EHD I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AN2EHD I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AN2EHD I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AN2EHD I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AN2EHD I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AN2EHD I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AN2EHD I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AN2EHD I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AN2EHD I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AN2EHD I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AN2EHD I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AN2EHD I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AN2EHD I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AN2EHD I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AN2EHD I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AN2EHD I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AN2EHD I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AN2EHD I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AN2EHD I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AN2EHD I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AN2EHD I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AN2EHD I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AN2EHD I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AN2EHD I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AN2EHD I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AN2EHD I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AN2EHD I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AN2EHD I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AN2EHD I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AN2EHD I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AN2EHD I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AN2EHD I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AN2EHD I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AN2EHD I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AN2EHD I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AN2EHD I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AN2EHD I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AN2EHD I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AN2EHD I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AN2EHD I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AN2EHD I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AN2EHD I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AN2EHD I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AN2EHD I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AN2EHD I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AN2EHD I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AN2EHD I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AN2EHD I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AN2EHD I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AN2EHD I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AN2EHD I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AN2EHD I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AN2EHD I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AN2EHD I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AN2EHD I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AN2EHD I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AN2EHD I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AN2EHD I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AN2EHD I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AN2EHD I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AN2EHD I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AN2EHD I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AN2EHD I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NR2EHD I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NR2EHD I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NR2EHD I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NR2EHD I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NR2EHD I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NR2EHD I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NR2EHD I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NR2EHD I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NR2EHD I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NR2EHD I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NR2EHD I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NR2EHD I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NR2EHD I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NR2EHD I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NR2EHD I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NR2EHD I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NR2EHD I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NR2EHD I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NR2EHD I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NR2EHD I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NR2EHD I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NR2EHD I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NR2EHD I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NR2EHD I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NR2EHD I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NR2EHD I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NR2EHD I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NR2EHD I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NR2EHD I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NR2EHD I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NR2EHD I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NR2EHD I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NR3EHD I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NR3EHD I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NR3EHD I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NR3EHD I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NR3EHD I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NR3EHD I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NR3EHD I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NR3EHD I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NR3EHD I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NR3EHD I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NR3EHD I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NR3EHD I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NR3EHD I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NR3EHD I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NR3EHD I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NR3EHD I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NR3EHD I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NR3EHD I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NR3EHD I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NR3EHD I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NR3EHD I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NR3EHD I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NR3EHD I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NR3EHD I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NR3EHD I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NR3EHD I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NR3EHD I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NR3EHD I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NR3EHD I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NR3EHD I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NR3EHD I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NR3EHD I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22EHD I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22EHD I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22EHD I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22EHD I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22EHD I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22EHD I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22EHD I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22EHD I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22EHD I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22EHD I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22EHD I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22EHD I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22EHD I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22EHD I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22EHD I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22EHD I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22EHD I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22EHD I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22EHD I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22EHD I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22EHD I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22EHD I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22EHD I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22EHD I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22EHD I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22EHD I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22EHD I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22EHD I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22EHD I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22EHD I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22EHD I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22EHD I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2EHD I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2EHD I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2EHD I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2EHD I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2EHD I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2EHD I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2EHD I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2EHD I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2EHD I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2EHD I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2EHD I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2EHD I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2EHD I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2EHD I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2EHD I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2EHD I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2EHD I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2EHD I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2EHD I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2EHD I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2EHD I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2EHD I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2EHD I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2EHD I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2EHD I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2EHD I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2EHD I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2EHD I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2EHD I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2EHD I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2EHD I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2EHD I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  AO222EHD I225 (tech239_int, comp0_0[0:0], comp0_0[1:1], tech239_int, comp0_0[0:0], tech239_int, comp0_0[1:1]);
  AO222EHD I226 (simp2381_0[0:0], tech239_int, comp0_0[2:2], simp2381_0[0:0], tech239_int, simp2381_0[0:0], comp0_0[2:2]);
  AO222EHD I227 (tech240_int, comp0_0[3:3], comp0_0[4:4], tech240_int, comp0_0[3:3], tech240_int, comp0_0[4:4]);
  AO222EHD I228 (simp2381_0[1:1], tech240_int, comp0_0[5:5], simp2381_0[1:1], tech240_int, simp2381_0[1:1], comp0_0[5:5]);
  AO222EHD I229 (tech241_int, comp0_0[6:6], comp0_0[7:7], tech241_int, comp0_0[6:6], tech241_int, comp0_0[7:7]);
  AO222EHD I230 (simp2381_0[2:2], tech241_int, comp0_0[8:8], simp2381_0[2:2], tech241_int, simp2381_0[2:2], comp0_0[8:8]);
  AO222EHD I231 (tech242_int, comp0_0[9:9], comp0_0[10:10], tech242_int, comp0_0[9:9], tech242_int, comp0_0[10:10]);
  AO222EHD I232 (simp2381_0[3:3], tech242_int, comp0_0[11:11], simp2381_0[3:3], tech242_int, simp2381_0[3:3], comp0_0[11:11]);
  AO222EHD I233 (tech243_int, comp0_0[12:12], comp0_0[13:13], tech243_int, comp0_0[12:12], tech243_int, comp0_0[13:13]);
  AO222EHD I234 (simp2381_0[4:4], tech243_int, comp0_0[14:14], simp2381_0[4:4], tech243_int, simp2381_0[4:4], comp0_0[14:14]);
  AO222EHD I235 (tech244_int, comp0_0[15:15], comp0_0[16:16], tech244_int, comp0_0[15:15], tech244_int, comp0_0[16:16]);
  AO222EHD I236 (simp2381_0[5:5], tech244_int, comp0_0[17:17], simp2381_0[5:5], tech244_int, simp2381_0[5:5], comp0_0[17:17]);
  AO222EHD I237 (tech245_int, comp0_0[18:18], comp0_0[19:19], tech245_int, comp0_0[18:18], tech245_int, comp0_0[19:19]);
  AO222EHD I238 (simp2381_0[6:6], tech245_int, comp0_0[20:20], simp2381_0[6:6], tech245_int, simp2381_0[6:6], comp0_0[20:20]);
  AO222EHD I239 (tech246_int, comp0_0[21:21], comp0_0[22:22], tech246_int, comp0_0[21:21], tech246_int, comp0_0[22:22]);
  AO222EHD I240 (simp2381_0[7:7], tech246_int, comp0_0[23:23], simp2381_0[7:7], tech246_int, simp2381_0[7:7], comp0_0[23:23]);
  AO222EHD I241 (tech247_int, comp0_0[24:24], comp0_0[25:25], tech247_int, comp0_0[24:24], tech247_int, comp0_0[25:25]);
  AO222EHD I242 (simp2381_0[8:8], tech247_int, comp0_0[26:26], simp2381_0[8:8], tech247_int, simp2381_0[8:8], comp0_0[26:26]);
  AO222EHD I243 (tech248_int, comp0_0[27:27], comp0_0[28:28], tech248_int, comp0_0[27:27], tech248_int, comp0_0[28:28]);
  AO222EHD I244 (simp2381_0[9:9], tech248_int, comp0_0[29:29], simp2381_0[9:9], tech248_int, simp2381_0[9:9], comp0_0[29:29]);
  AO222EHD I245 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31], simp2381_0[10:10], comp0_0[30:30], simp2381_0[10:10], comp0_0[31:31]);
  AO222EHD I246 (tech251_int, simp2381_0[0:0], simp2381_0[1:1], tech251_int, simp2381_0[0:0], tech251_int, simp2381_0[1:1]);
  AO222EHD I247 (simp2382_0[0:0], tech251_int, simp2381_0[2:2], simp2382_0[0:0], tech251_int, simp2382_0[0:0], simp2381_0[2:2]);
  AO222EHD I248 (tech252_int, simp2381_0[3:3], simp2381_0[4:4], tech252_int, simp2381_0[3:3], tech252_int, simp2381_0[4:4]);
  AO222EHD I249 (simp2382_0[1:1], tech252_int, simp2381_0[5:5], simp2382_0[1:1], tech252_int, simp2382_0[1:1], simp2381_0[5:5]);
  AO222EHD I250 (tech253_int, simp2381_0[6:6], simp2381_0[7:7], tech253_int, simp2381_0[6:6], tech253_int, simp2381_0[7:7]);
  AO222EHD I251 (simp2382_0[2:2], tech253_int, simp2381_0[8:8], simp2382_0[2:2], tech253_int, simp2382_0[2:2], simp2381_0[8:8]);
  AO222EHD I252 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10], simp2382_0[3:3], simp2381_0[9:9], simp2382_0[3:3], simp2381_0[10:10]);
  AO222EHD I253 (tech256_int, simp2382_0[0:0], simp2382_0[1:1], tech256_int, simp2382_0[0:0], tech256_int, simp2382_0[1:1]);
  AO222EHD I254 (simp2383_0[0:0], tech256_int, simp2382_0[2:2], simp2383_0[0:0], tech256_int, simp2383_0[0:0], simp2382_0[2:2]);
  BUFEHD I255 (simp2383_0[1:1], simp2382_0[3:3]);
  AO222EHD I256 (wc_0, simp2383_0[0:0], simp2383_0[1:1], wc_0, simp2383_0[0:0], wc_0, simp2383_0[1:1]);
  AN2EHD I257 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AN2EHD I258 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AN2EHD I259 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AN2EHD I260 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AN2EHD I261 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AN2EHD I262 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AN2EHD I263 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AN2EHD I264 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AN2EHD I265 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AN2EHD I266 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AN2EHD I267 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AN2EHD I268 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AN2EHD I269 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AN2EHD I270 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AN2EHD I271 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AN2EHD I272 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AN2EHD I273 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AN2EHD I274 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AN2EHD I275 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AN2EHD I276 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AN2EHD I277 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AN2EHD I278 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AN2EHD I279 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AN2EHD I280 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AN2EHD I281 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AN2EHD I282 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AN2EHD I283 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AN2EHD I284 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AN2EHD I285 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AN2EHD I286 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AN2EHD I287 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AN2EHD I288 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AN2EHD I289 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AN2EHD I290 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AN2EHD I291 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AN2EHD I292 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AN2EHD I293 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AN2EHD I294 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AN2EHD I295 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AN2EHD I296 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AN2EHD I297 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AN2EHD I298 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AN2EHD I299 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AN2EHD I300 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AN2EHD I301 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AN2EHD I302 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AN2EHD I303 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AN2EHD I304 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AN2EHD I305 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AN2EHD I306 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AN2EHD I307 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AN2EHD I308 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AN2EHD I309 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AN2EHD I310 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AN2EHD I311 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AN2EHD I312 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AN2EHD I313 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AN2EHD I314 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AN2EHD I315 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AN2EHD I316 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AN2EHD I317 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AN2EHD I318 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AN2EHD I319 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AN2EHD I320 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFEHD I321 (conwigc_0, wc_0);
  AO12EHD I322 (conwig_0, conwigc_0, conwigc_0, conwigcanw_0);
  NR2EHD I323 (conwigcanw_0, anyread_0, conwig_0);
  BUFEHD I324 (wf_0[0:0], conwgif_0[0:0]);
  BUFEHD I325 (wt_0[0:0], conwgit_0[0:0]);
  BUFEHD I326 (wenr_0[0:0], wc_0);
  BUFEHD I327 (wf_0[1:1], conwgif_0[1:1]);
  BUFEHD I328 (wt_0[1:1], conwgit_0[1:1]);
  BUFEHD I329 (wenr_0[1:1], wc_0);
  BUFEHD I330 (wf_0[2:2], conwgif_0[2:2]);
  BUFEHD I331 (wt_0[2:2], conwgit_0[2:2]);
  BUFEHD I332 (wenr_0[2:2], wc_0);
  BUFEHD I333 (wf_0[3:3], conwgif_0[3:3]);
  BUFEHD I334 (wt_0[3:3], conwgit_0[3:3]);
  BUFEHD I335 (wenr_0[3:3], wc_0);
  BUFEHD I336 (wf_0[4:4], conwgif_0[4:4]);
  BUFEHD I337 (wt_0[4:4], conwgit_0[4:4]);
  BUFEHD I338 (wenr_0[4:4], wc_0);
  BUFEHD I339 (wf_0[5:5], conwgif_0[5:5]);
  BUFEHD I340 (wt_0[5:5], conwgit_0[5:5]);
  BUFEHD I341 (wenr_0[5:5], wc_0);
  BUFEHD I342 (wf_0[6:6], conwgif_0[6:6]);
  BUFEHD I343 (wt_0[6:6], conwgit_0[6:6]);
  BUFEHD I344 (wenr_0[6:6], wc_0);
  BUFEHD I345 (wf_0[7:7], conwgif_0[7:7]);
  BUFEHD I346 (wt_0[7:7], conwgit_0[7:7]);
  BUFEHD I347 (wenr_0[7:7], wc_0);
  BUFEHD I348 (wf_0[8:8], conwgif_0[8:8]);
  BUFEHD I349 (wt_0[8:8], conwgit_0[8:8]);
  BUFEHD I350 (wenr_0[8:8], wc_0);
  BUFEHD I351 (wf_0[9:9], conwgif_0[9:9]);
  BUFEHD I352 (wt_0[9:9], conwgit_0[9:9]);
  BUFEHD I353 (wenr_0[9:9], wc_0);
  BUFEHD I354 (wf_0[10:10], conwgif_0[10:10]);
  BUFEHD I355 (wt_0[10:10], conwgit_0[10:10]);
  BUFEHD I356 (wenr_0[10:10], wc_0);
  BUFEHD I357 (wf_0[11:11], conwgif_0[11:11]);
  BUFEHD I358 (wt_0[11:11], conwgit_0[11:11]);
  BUFEHD I359 (wenr_0[11:11], wc_0);
  BUFEHD I360 (wf_0[12:12], conwgif_0[12:12]);
  BUFEHD I361 (wt_0[12:12], conwgit_0[12:12]);
  BUFEHD I362 (wenr_0[12:12], wc_0);
  BUFEHD I363 (wf_0[13:13], conwgif_0[13:13]);
  BUFEHD I364 (wt_0[13:13], conwgit_0[13:13]);
  BUFEHD I365 (wenr_0[13:13], wc_0);
  BUFEHD I366 (wf_0[14:14], conwgif_0[14:14]);
  BUFEHD I367 (wt_0[14:14], conwgit_0[14:14]);
  BUFEHD I368 (wenr_0[14:14], wc_0);
  BUFEHD I369 (wf_0[15:15], conwgif_0[15:15]);
  BUFEHD I370 (wt_0[15:15], conwgit_0[15:15]);
  BUFEHD I371 (wenr_0[15:15], wc_0);
  BUFEHD I372 (wf_0[16:16], conwgif_0[16:16]);
  BUFEHD I373 (wt_0[16:16], conwgit_0[16:16]);
  BUFEHD I374 (wenr_0[16:16], wc_0);
  BUFEHD I375 (wf_0[17:17], conwgif_0[17:17]);
  BUFEHD I376 (wt_0[17:17], conwgit_0[17:17]);
  BUFEHD I377 (wenr_0[17:17], wc_0);
  BUFEHD I378 (wf_0[18:18], conwgif_0[18:18]);
  BUFEHD I379 (wt_0[18:18], conwgit_0[18:18]);
  BUFEHD I380 (wenr_0[18:18], wc_0);
  BUFEHD I381 (wf_0[19:19], conwgif_0[19:19]);
  BUFEHD I382 (wt_0[19:19], conwgit_0[19:19]);
  BUFEHD I383 (wenr_0[19:19], wc_0);
  BUFEHD I384 (wf_0[20:20], conwgif_0[20:20]);
  BUFEHD I385 (wt_0[20:20], conwgit_0[20:20]);
  BUFEHD I386 (wenr_0[20:20], wc_0);
  BUFEHD I387 (wf_0[21:21], conwgif_0[21:21]);
  BUFEHD I388 (wt_0[21:21], conwgit_0[21:21]);
  BUFEHD I389 (wenr_0[21:21], wc_0);
  BUFEHD I390 (wf_0[22:22], conwgif_0[22:22]);
  BUFEHD I391 (wt_0[22:22], conwgit_0[22:22]);
  BUFEHD I392 (wenr_0[22:22], wc_0);
  BUFEHD I393 (wf_0[23:23], conwgif_0[23:23]);
  BUFEHD I394 (wt_0[23:23], conwgit_0[23:23]);
  BUFEHD I395 (wenr_0[23:23], wc_0);
  BUFEHD I396 (wf_0[24:24], conwgif_0[24:24]);
  BUFEHD I397 (wt_0[24:24], conwgit_0[24:24]);
  BUFEHD I398 (wenr_0[24:24], wc_0);
  BUFEHD I399 (wf_0[25:25], conwgif_0[25:25]);
  BUFEHD I400 (wt_0[25:25], conwgit_0[25:25]);
  BUFEHD I401 (wenr_0[25:25], wc_0);
  BUFEHD I402 (wf_0[26:26], conwgif_0[26:26]);
  BUFEHD I403 (wt_0[26:26], conwgit_0[26:26]);
  BUFEHD I404 (wenr_0[26:26], wc_0);
  BUFEHD I405 (wf_0[27:27], conwgif_0[27:27]);
  BUFEHD I406 (wt_0[27:27], conwgit_0[27:27]);
  BUFEHD I407 (wenr_0[27:27], wc_0);
  BUFEHD I408 (wf_0[28:28], conwgif_0[28:28]);
  BUFEHD I409 (wt_0[28:28], conwgit_0[28:28]);
  BUFEHD I410 (wenr_0[28:28], wc_0);
  BUFEHD I411 (wf_0[29:29], conwgif_0[29:29]);
  BUFEHD I412 (wt_0[29:29], conwgit_0[29:29]);
  BUFEHD I413 (wenr_0[29:29], wc_0);
  BUFEHD I414 (wf_0[30:30], conwgif_0[30:30]);
  BUFEHD I415 (wt_0[30:30], conwgit_0[30:30]);
  BUFEHD I416 (wenr_0[30:30], wc_0);
  BUFEHD I417 (wf_0[31:31], conwgif_0[31:31]);
  BUFEHD I418 (wt_0[31:31], conwgit_0[31:31]);
  BUFEHD I419 (wenr_0[31:31], wc_0);
  AO222EHD I420 (tech428_int, conwig_0, wacks_0[0:0], tech428_int, conwig_0, tech428_int, wacks_0[0:0]);
  AO222EHD I421 (simp4071_0[0:0], tech428_int, wacks_0[1:1], simp4071_0[0:0], tech428_int, simp4071_0[0:0], wacks_0[1:1]);
  AO222EHD I422 (tech429_int, wacks_0[2:2], wacks_0[3:3], tech429_int, wacks_0[2:2], tech429_int, wacks_0[3:3]);
  AO222EHD I423 (simp4071_0[1:1], tech429_int, wacks_0[4:4], simp4071_0[1:1], tech429_int, simp4071_0[1:1], wacks_0[4:4]);
  AO222EHD I424 (tech430_int, wacks_0[5:5], wacks_0[6:6], tech430_int, wacks_0[5:5], tech430_int, wacks_0[6:6]);
  AO222EHD I425 (simp4071_0[2:2], tech430_int, wacks_0[7:7], simp4071_0[2:2], tech430_int, simp4071_0[2:2], wacks_0[7:7]);
  AO222EHD I426 (tech431_int, wacks_0[8:8], wacks_0[9:9], tech431_int, wacks_0[8:8], tech431_int, wacks_0[9:9]);
  AO222EHD I427 (simp4071_0[3:3], tech431_int, wacks_0[10:10], simp4071_0[3:3], tech431_int, simp4071_0[3:3], wacks_0[10:10]);
  AO222EHD I428 (tech432_int, wacks_0[11:11], wacks_0[12:12], tech432_int, wacks_0[11:11], tech432_int, wacks_0[12:12]);
  AO222EHD I429 (simp4071_0[4:4], tech432_int, wacks_0[13:13], simp4071_0[4:4], tech432_int, simp4071_0[4:4], wacks_0[13:13]);
  AO222EHD I430 (tech433_int, wacks_0[14:14], wacks_0[15:15], tech433_int, wacks_0[14:14], tech433_int, wacks_0[15:15]);
  AO222EHD I431 (simp4071_0[5:5], tech433_int, wacks_0[16:16], simp4071_0[5:5], tech433_int, simp4071_0[5:5], wacks_0[16:16]);
  AO222EHD I432 (tech434_int, wacks_0[17:17], wacks_0[18:18], tech434_int, wacks_0[17:17], tech434_int, wacks_0[18:18]);
  AO222EHD I433 (simp4071_0[6:6], tech434_int, wacks_0[19:19], simp4071_0[6:6], tech434_int, simp4071_0[6:6], wacks_0[19:19]);
  AO222EHD I434 (tech435_int, wacks_0[20:20], wacks_0[21:21], tech435_int, wacks_0[20:20], tech435_int, wacks_0[21:21]);
  AO222EHD I435 (simp4071_0[7:7], tech435_int, wacks_0[22:22], simp4071_0[7:7], tech435_int, simp4071_0[7:7], wacks_0[22:22]);
  AO222EHD I436 (tech436_int, wacks_0[23:23], wacks_0[24:24], tech436_int, wacks_0[23:23], tech436_int, wacks_0[24:24]);
  AO222EHD I437 (simp4071_0[8:8], tech436_int, wacks_0[25:25], simp4071_0[8:8], tech436_int, simp4071_0[8:8], wacks_0[25:25]);
  AO222EHD I438 (tech437_int, wacks_0[26:26], wacks_0[27:27], tech437_int, wacks_0[26:26], tech437_int, wacks_0[27:27]);
  AO222EHD I439 (simp4071_0[9:9], tech437_int, wacks_0[28:28], simp4071_0[9:9], tech437_int, simp4071_0[9:9], wacks_0[28:28]);
  AO222EHD I440 (tech438_int, wacks_0[29:29], wacks_0[30:30], tech438_int, wacks_0[29:29], tech438_int, wacks_0[30:30]);
  AO222EHD I441 (simp4071_0[10:10], tech438_int, wacks_0[31:31], simp4071_0[10:10], tech438_int, simp4071_0[10:10], wacks_0[31:31]);
  AO222EHD I442 (tech440_int, simp4071_0[0:0], simp4071_0[1:1], tech440_int, simp4071_0[0:0], tech440_int, simp4071_0[1:1]);
  AO222EHD I443 (simp4072_0[0:0], tech440_int, simp4071_0[2:2], simp4072_0[0:0], tech440_int, simp4072_0[0:0], simp4071_0[2:2]);
  AO222EHD I444 (tech441_int, simp4071_0[3:3], simp4071_0[4:4], tech441_int, simp4071_0[3:3], tech441_int, simp4071_0[4:4]);
  AO222EHD I445 (simp4072_0[1:1], tech441_int, simp4071_0[5:5], simp4072_0[1:1], tech441_int, simp4072_0[1:1], simp4071_0[5:5]);
  AO222EHD I446 (tech442_int, simp4071_0[6:6], simp4071_0[7:7], tech442_int, simp4071_0[6:6], tech442_int, simp4071_0[7:7]);
  AO222EHD I447 (simp4072_0[2:2], tech442_int, simp4071_0[8:8], simp4072_0[2:2], tech442_int, simp4072_0[2:2], simp4071_0[8:8]);
  AO222EHD I448 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10], simp4072_0[3:3], simp4071_0[9:9], simp4072_0[3:3], simp4071_0[10:10]);
  AO222EHD I449 (tech445_int, simp4072_0[0:0], simp4072_0[1:1], tech445_int, simp4072_0[0:0], tech445_int, simp4072_0[1:1]);
  AO222EHD I450 (simp4073_0[0:0], tech445_int, simp4072_0[2:2], simp4073_0[0:0], tech445_int, simp4073_0[0:0], simp4072_0[2:2]);
  BUFEHD I451 (simp4073_0[1:1], simp4072_0[3:3]);
  AO222EHD I452 (wd_0r, simp4073_0[0:0], simp4073_0[1:1], wd_0r, simp4073_0[0:0], wd_0r, simp4073_0[1:1]);
  AN2EHD I453 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AN2EHD I454 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AN2EHD I455 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AN2EHD I456 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AN2EHD I457 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AN2EHD I458 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AN2EHD I459 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AN2EHD I460 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AN2EHD I461 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AN2EHD I462 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AN2EHD I463 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AN2EHD I464 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AN2EHD I465 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AN2EHD I466 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AN2EHD I467 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AN2EHD I468 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AN2EHD I469 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AN2EHD I470 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AN2EHD I471 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AN2EHD I472 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AN2EHD I473 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AN2EHD I474 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AN2EHD I475 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AN2EHD I476 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AN2EHD I477 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AN2EHD I478 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AN2EHD I479 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AN2EHD I480 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AN2EHD I481 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AN2EHD I482 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AN2EHD I483 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AN2EHD I484 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AN2EHD I485 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AN2EHD I486 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AN2EHD I487 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AN2EHD I488 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AN2EHD I489 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AN2EHD I490 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AN2EHD I491 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AN2EHD I492 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AN2EHD I493 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AN2EHD I494 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AN2EHD I495 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AN2EHD I496 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AN2EHD I497 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AN2EHD I498 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AN2EHD I499 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AN2EHD I500 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AN2EHD I501 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AN2EHD I502 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AN2EHD I503 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AN2EHD I504 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AN2EHD I505 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AN2EHD I506 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AN2EHD I507 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AN2EHD I508 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AN2EHD I509 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AN2EHD I510 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AN2EHD I511 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AN2EHD I512 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AN2EHD I513 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AN2EHD I514 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AN2EHD I515 (rd_2r0[0:0], df_0[2:2], rg_2r);
  AN2EHD I516 (rd_2r0[1:1], df_0[3:3], rg_2r);
  AN2EHD I517 (rd_2r0[2:2], df_0[4:4], rg_2r);
  AN2EHD I518 (rd_2r0[3:3], df_0[5:5], rg_2r);
  AN2EHD I519 (rd_2r0[4:4], df_0[6:6], rg_2r);
  AN2EHD I520 (rd_2r0[5:5], df_0[7:7], rg_2r);
  AN2EHD I521 (rd_2r0[6:6], df_0[8:8], rg_2r);
  AN2EHD I522 (rd_2r0[7:7], df_0[9:9], rg_2r);
  AN2EHD I523 (rd_2r0[8:8], df_0[10:10], rg_2r);
  AN2EHD I524 (rd_2r0[9:9], df_0[11:11], rg_2r);
  AN2EHD I525 (rd_2r0[10:10], df_0[12:12], rg_2r);
  AN2EHD I526 (rd_2r0[11:11], df_0[13:13], rg_2r);
  AN2EHD I527 (rd_2r0[12:12], df_0[14:14], rg_2r);
  AN2EHD I528 (rd_2r0[13:13], df_0[15:15], rg_2r);
  AN2EHD I529 (rd_2r0[14:14], df_0[16:16], rg_2r);
  AN2EHD I530 (rd_2r0[15:15], df_0[17:17], rg_2r);
  AN2EHD I531 (rd_2r0[16:16], df_0[18:18], rg_2r);
  AN2EHD I532 (rd_2r0[17:17], df_0[19:19], rg_2r);
  AN2EHD I533 (rd_2r0[18:18], df_0[20:20], rg_2r);
  AN2EHD I534 (rd_2r0[19:19], df_0[21:21], rg_2r);
  AN2EHD I535 (rd_2r0[20:20], df_0[22:22], rg_2r);
  AN2EHD I536 (rd_2r0[21:21], df_0[23:23], rg_2r);
  AN2EHD I537 (rd_2r0[22:22], df_0[24:24], rg_2r);
  AN2EHD I538 (rd_2r0[23:23], df_0[25:25], rg_2r);
  AN2EHD I539 (rd_2r0[24:24], df_0[26:26], rg_2r);
  AN2EHD I540 (rd_2r0[25:25], df_0[27:27], rg_2r);
  AN2EHD I541 (rd_2r0[26:26], df_0[28:28], rg_2r);
  AN2EHD I542 (rd_2r0[27:27], df_0[29:29], rg_2r);
  AN2EHD I543 (rd_2r0[28:28], df_0[30:30], rg_2r);
  AN2EHD I544 (rd_2r0[29:29], df_0[31:31], rg_2r);
  AN2EHD I545 (rd_3r0[0:0], df_0[2:2], rg_3r);
  AN2EHD I546 (rd_3r0[1:1], df_0[3:3], rg_3r);
  AN2EHD I547 (rd_3r0[2:2], df_0[4:4], rg_3r);
  AN2EHD I548 (rd_3r0[3:3], df_0[5:5], rg_3r);
  AN2EHD I549 (rd_3r0[4:4], df_0[6:6], rg_3r);
  AN2EHD I550 (rd_3r0[5:5], df_0[7:7], rg_3r);
  AN2EHD I551 (rd_3r0[6:6], df_0[8:8], rg_3r);
  AN2EHD I552 (rd_3r0[7:7], df_0[9:9], rg_3r);
  AN2EHD I553 (rd_3r0[8:8], df_0[10:10], rg_3r);
  AN2EHD I554 (rd_3r0[9:9], df_0[11:11], rg_3r);
  AN2EHD I555 (rd_3r0[10:10], df_0[12:12], rg_3r);
  AN2EHD I556 (rd_3r0[11:11], df_0[13:13], rg_3r);
  AN2EHD I557 (rd_3r0[12:12], df_0[14:14], rg_3r);
  AN2EHD I558 (rd_3r0[13:13], df_0[15:15], rg_3r);
  AN2EHD I559 (rd_3r0[14:14], df_0[16:16], rg_3r);
  AN2EHD I560 (rd_3r0[15:15], df_0[17:17], rg_3r);
  AN2EHD I561 (rd_3r0[16:16], df_0[18:18], rg_3r);
  AN2EHD I562 (rd_3r0[17:17], df_0[19:19], rg_3r);
  AN2EHD I563 (rd_3r0[18:18], df_0[20:20], rg_3r);
  AN2EHD I564 (rd_3r0[19:19], df_0[21:21], rg_3r);
  AN2EHD I565 (rd_3r0[20:20], df_0[22:22], rg_3r);
  AN2EHD I566 (rd_3r0[21:21], df_0[23:23], rg_3r);
  AN2EHD I567 (rd_3r0[22:22], df_0[24:24], rg_3r);
  AN2EHD I568 (rd_3r0[23:23], df_0[25:25], rg_3r);
  AN2EHD I569 (rd_3r0[24:24], df_0[26:26], rg_3r);
  AN2EHD I570 (rd_3r0[25:25], df_0[27:27], rg_3r);
  AN2EHD I571 (rd_3r0[26:26], df_0[28:28], rg_3r);
  AN2EHD I572 (rd_3r0[27:27], df_0[29:29], rg_3r);
  AN2EHD I573 (rd_3r0[28:28], df_0[30:30], rg_3r);
  AN2EHD I574 (rd_3r0[29:29], df_0[31:31], rg_3r);
  AN2EHD I575 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AN2EHD I576 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AN2EHD I577 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AN2EHD I578 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AN2EHD I579 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AN2EHD I580 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AN2EHD I581 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AN2EHD I582 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AN2EHD I583 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AN2EHD I584 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AN2EHD I585 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AN2EHD I586 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AN2EHD I587 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AN2EHD I588 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AN2EHD I589 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AN2EHD I590 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AN2EHD I591 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AN2EHD I592 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AN2EHD I593 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AN2EHD I594 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AN2EHD I595 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AN2EHD I596 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AN2EHD I597 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AN2EHD I598 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AN2EHD I599 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AN2EHD I600 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AN2EHD I601 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AN2EHD I602 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AN2EHD I603 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AN2EHD I604 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AN2EHD I605 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AN2EHD I606 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AN2EHD I607 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AN2EHD I608 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AN2EHD I609 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AN2EHD I610 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AN2EHD I611 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AN2EHD I612 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AN2EHD I613 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AN2EHD I614 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AN2EHD I615 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AN2EHD I616 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AN2EHD I617 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AN2EHD I618 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AN2EHD I619 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AN2EHD I620 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AN2EHD I621 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AN2EHD I622 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AN2EHD I623 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AN2EHD I624 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AN2EHD I625 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AN2EHD I626 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AN2EHD I627 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AN2EHD I628 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AN2EHD I629 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AN2EHD I630 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AN2EHD I631 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AN2EHD I632 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AN2EHD I633 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AN2EHD I634 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AN2EHD I635 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AN2EHD I636 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AN2EHD I637 (rd_2r1[0:0], dt_0[2:2], rg_2r);
  AN2EHD I638 (rd_2r1[1:1], dt_0[3:3], rg_2r);
  AN2EHD I639 (rd_2r1[2:2], dt_0[4:4], rg_2r);
  AN2EHD I640 (rd_2r1[3:3], dt_0[5:5], rg_2r);
  AN2EHD I641 (rd_2r1[4:4], dt_0[6:6], rg_2r);
  AN2EHD I642 (rd_2r1[5:5], dt_0[7:7], rg_2r);
  AN2EHD I643 (rd_2r1[6:6], dt_0[8:8], rg_2r);
  AN2EHD I644 (rd_2r1[7:7], dt_0[9:9], rg_2r);
  AN2EHD I645 (rd_2r1[8:8], dt_0[10:10], rg_2r);
  AN2EHD I646 (rd_2r1[9:9], dt_0[11:11], rg_2r);
  AN2EHD I647 (rd_2r1[10:10], dt_0[12:12], rg_2r);
  AN2EHD I648 (rd_2r1[11:11], dt_0[13:13], rg_2r);
  AN2EHD I649 (rd_2r1[12:12], dt_0[14:14], rg_2r);
  AN2EHD I650 (rd_2r1[13:13], dt_0[15:15], rg_2r);
  AN2EHD I651 (rd_2r1[14:14], dt_0[16:16], rg_2r);
  AN2EHD I652 (rd_2r1[15:15], dt_0[17:17], rg_2r);
  AN2EHD I653 (rd_2r1[16:16], dt_0[18:18], rg_2r);
  AN2EHD I654 (rd_2r1[17:17], dt_0[19:19], rg_2r);
  AN2EHD I655 (rd_2r1[18:18], dt_0[20:20], rg_2r);
  AN2EHD I656 (rd_2r1[19:19], dt_0[21:21], rg_2r);
  AN2EHD I657 (rd_2r1[20:20], dt_0[22:22], rg_2r);
  AN2EHD I658 (rd_2r1[21:21], dt_0[23:23], rg_2r);
  AN2EHD I659 (rd_2r1[22:22], dt_0[24:24], rg_2r);
  AN2EHD I660 (rd_2r1[23:23], dt_0[25:25], rg_2r);
  AN2EHD I661 (rd_2r1[24:24], dt_0[26:26], rg_2r);
  AN2EHD I662 (rd_2r1[25:25], dt_0[27:27], rg_2r);
  AN2EHD I663 (rd_2r1[26:26], dt_0[28:28], rg_2r);
  AN2EHD I664 (rd_2r1[27:27], dt_0[29:29], rg_2r);
  AN2EHD I665 (rd_2r1[28:28], dt_0[30:30], rg_2r);
  AN2EHD I666 (rd_2r1[29:29], dt_0[31:31], rg_2r);
  AN2EHD I667 (rd_3r1[0:0], dt_0[2:2], rg_3r);
  AN2EHD I668 (rd_3r1[1:1], dt_0[3:3], rg_3r);
  AN2EHD I669 (rd_3r1[2:2], dt_0[4:4], rg_3r);
  AN2EHD I670 (rd_3r1[3:3], dt_0[5:5], rg_3r);
  AN2EHD I671 (rd_3r1[4:4], dt_0[6:6], rg_3r);
  AN2EHD I672 (rd_3r1[5:5], dt_0[7:7], rg_3r);
  AN2EHD I673 (rd_3r1[6:6], dt_0[8:8], rg_3r);
  AN2EHD I674 (rd_3r1[7:7], dt_0[9:9], rg_3r);
  AN2EHD I675 (rd_3r1[8:8], dt_0[10:10], rg_3r);
  AN2EHD I676 (rd_3r1[9:9], dt_0[11:11], rg_3r);
  AN2EHD I677 (rd_3r1[10:10], dt_0[12:12], rg_3r);
  AN2EHD I678 (rd_3r1[11:11], dt_0[13:13], rg_3r);
  AN2EHD I679 (rd_3r1[12:12], dt_0[14:14], rg_3r);
  AN2EHD I680 (rd_3r1[13:13], dt_0[15:15], rg_3r);
  AN2EHD I681 (rd_3r1[14:14], dt_0[16:16], rg_3r);
  AN2EHD I682 (rd_3r1[15:15], dt_0[17:17], rg_3r);
  AN2EHD I683 (rd_3r1[16:16], dt_0[18:18], rg_3r);
  AN2EHD I684 (rd_3r1[17:17], dt_0[19:19], rg_3r);
  AN2EHD I685 (rd_3r1[18:18], dt_0[20:20], rg_3r);
  AN2EHD I686 (rd_3r1[19:19], dt_0[21:21], rg_3r);
  AN2EHD I687 (rd_3r1[20:20], dt_0[22:22], rg_3r);
  AN2EHD I688 (rd_3r1[21:21], dt_0[23:23], rg_3r);
  AN2EHD I689 (rd_3r1[22:22], dt_0[24:24], rg_3r);
  AN2EHD I690 (rd_3r1[23:23], dt_0[25:25], rg_3r);
  AN2EHD I691 (rd_3r1[24:24], dt_0[26:26], rg_3r);
  AN2EHD I692 (rd_3r1[25:25], dt_0[27:27], rg_3r);
  AN2EHD I693 (rd_3r1[26:26], dt_0[28:28], rg_3r);
  AN2EHD I694 (rd_3r1[27:27], dt_0[29:29], rg_3r);
  AN2EHD I695 (rd_3r1[28:28], dt_0[30:30], rg_3r);
  AN2EHD I696 (rd_3r1[29:29], dt_0[31:31], rg_3r);
  NR3EHD I697 (simp6521_0[0:0], rg_0r, rg_1r, rg_2r);
  NR3EHD I698 (simp6521_0[1:1], rg_3r, rg_0a, rg_1a);
  NR2EHD I699 (simp6521_0[2:2], rg_2a, rg_3a);
  ND3EHD I700 (anyread_0, simp6521_0[0:0], simp6521_0[1:1], simp6521_0[2:2]);
  BUFEHD I701 (wg_0a, wd_0a);
  BUFEHD I702 (rg_0a, rd_0a);
  BUFEHD I703 (rg_1a, rd_1a);
  BUFEHD I704 (rg_2a, rd_2a);
  BUFEHD I705 (rg_3a, rd_3a);
endmodule

// tkj0m0_0_0 TeakJ [Many [0,0,0],One 0]
module tkj0m0_0_0 (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  output o_0r;
  input o_0a;
  input reset;
  wire tech0_int;
  AO222EHD I0 (tech0_int, i_0r, i_1r, tech0_int, i_0r, tech0_int, i_1r);
  AO222EHD I1 (o_0r, tech0_int, i_2r, o_0r, tech0_int, o_0r, i_2r);
  BUFEHD I2 (i_0a, o_0a);
  BUFEHD I3 (i_1a, o_0a);
  BUFEHD I4 (i_2a, o_0a);
endmodule

// tkm4x32b TeakM [Many [32,32,32,32],One 32]
module tkm4x32b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  input [31:0] i_2r0;
  input [31:0] i_2r1;
  output i_2a;
  input [31:0] i_3r0;
  input [31:0] i_3r1;
  output i_3a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire [31:0] gfint_0;
  wire [31:0] gfint_1;
  wire [31:0] gfint_2;
  wire [31:0] gfint_3;
  wire [31:0] gtint_0;
  wire [31:0] gtint_1;
  wire [31:0] gtint_2;
  wire [31:0] gtint_3;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire icomp_3;
  wire nchosen_0;
  wire [1:0] simp181_0;
  wire [1:0] simp191_0;
  wire [1:0] simp201_0;
  wire [1:0] simp211_0;
  wire [1:0] simp221_0;
  wire [1:0] simp231_0;
  wire [1:0] simp241_0;
  wire [1:0] simp251_0;
  wire [1:0] simp261_0;
  wire [1:0] simp271_0;
  wire [1:0] simp281_0;
  wire [1:0] simp291_0;
  wire [1:0] simp301_0;
  wire [1:0] simp311_0;
  wire [1:0] simp321_0;
  wire [1:0] simp331_0;
  wire [1:0] simp341_0;
  wire [1:0] simp351_0;
  wire [1:0] simp361_0;
  wire [1:0] simp371_0;
  wire [1:0] simp381_0;
  wire [1:0] simp391_0;
  wire [1:0] simp401_0;
  wire [1:0] simp411_0;
  wire [1:0] simp421_0;
  wire [1:0] simp431_0;
  wire [1:0] simp441_0;
  wire [1:0] simp451_0;
  wire [1:0] simp461_0;
  wire [1:0] simp471_0;
  wire [1:0] simp481_0;
  wire [1:0] simp491_0;
  wire [1:0] simp501_0;
  wire [1:0] simp511_0;
  wire [1:0] simp521_0;
  wire [1:0] simp531_0;
  wire [1:0] simp541_0;
  wire [1:0] simp551_0;
  wire [1:0] simp561_0;
  wire [1:0] simp571_0;
  wire [1:0] simp581_0;
  wire [1:0] simp591_0;
  wire [1:0] simp601_0;
  wire [1:0] simp611_0;
  wire [1:0] simp621_0;
  wire [1:0] simp631_0;
  wire [1:0] simp641_0;
  wire [1:0] simp651_0;
  wire [1:0] simp661_0;
  wire [1:0] simp671_0;
  wire [1:0] simp681_0;
  wire [1:0] simp691_0;
  wire [1:0] simp701_0;
  wire [1:0] simp711_0;
  wire [1:0] simp721_0;
  wire [1:0] simp731_0;
  wire [1:0] simp741_0;
  wire [1:0] simp751_0;
  wire [1:0] simp761_0;
  wire [1:0] simp771_0;
  wire [1:0] simp781_0;
  wire [1:0] simp791_0;
  wire [1:0] simp801_0;
  wire [1:0] simp811_0;
  wire [31:0] comp0_0;
  wire [10:0] simp3711_0;
  wire tech564_int;
  wire tech565_int;
  wire tech566_int;
  wire tech567_int;
  wire tech568_int;
  wire tech569_int;
  wire tech570_int;
  wire tech571_int;
  wire tech572_int;
  wire tech573_int;
  wire [3:0] simp3712_0;
  wire tech576_int;
  wire tech577_int;
  wire tech578_int;
  wire [1:0] simp3713_0;
  wire tech581_int;
  wire [31:0] comp1_0;
  wire [10:0] simp4051_0;
  wire tech618_int;
  wire tech619_int;
  wire tech620_int;
  wire tech621_int;
  wire tech622_int;
  wire tech623_int;
  wire tech624_int;
  wire tech625_int;
  wire tech626_int;
  wire tech627_int;
  wire [3:0] simp4052_0;
  wire tech630_int;
  wire tech631_int;
  wire tech632_int;
  wire [1:0] simp4053_0;
  wire tech635_int;
  wire [31:0] comp2_0;
  wire [10:0] simp4391_0;
  wire tech672_int;
  wire tech673_int;
  wire tech674_int;
  wire tech675_int;
  wire tech676_int;
  wire tech677_int;
  wire tech678_int;
  wire tech679_int;
  wire tech680_int;
  wire tech681_int;
  wire [3:0] simp4392_0;
  wire tech684_int;
  wire tech685_int;
  wire tech686_int;
  wire [1:0] simp4393_0;
  wire tech689_int;
  wire [31:0] comp3_0;
  wire [10:0] simp4731_0;
  wire tech726_int;
  wire tech727_int;
  wire tech728_int;
  wire tech729_int;
  wire tech730_int;
  wire tech731_int;
  wire tech732_int;
  wire tech733_int;
  wire tech734_int;
  wire tech735_int;
  wire [3:0] simp4732_0;
  wire tech738_int;
  wire tech739_int;
  wire tech740_int;
  wire [1:0] simp4733_0;
  wire tech743_int;
  wire tech746_oint;
  wire tech747_oint;
  wire tech748_oint;
  wire tech749_oint;
  wire [1:0] simp4781_0;
  wire tech755_oint;
  wire tech756_oint;
  wire tech757_oint;
  wire tech758_oint;
  NR3EHD I0 (simp181_0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  INVHHD I1 (simp181_0[1:1], gfint_3[0:0]);
  ND2HHD I2 (o_0r0[0:0], simp181_0[0:0], simp181_0[1:1]);
  NR3EHD I3 (simp191_0[0:0], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  INVHHD I4 (simp191_0[1:1], gfint_3[1:1]);
  ND2HHD I5 (o_0r0[1:1], simp191_0[0:0], simp191_0[1:1]);
  NR3EHD I6 (simp201_0[0:0], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  INVHHD I7 (simp201_0[1:1], gfint_3[2:2]);
  ND2HHD I8 (o_0r0[2:2], simp201_0[0:0], simp201_0[1:1]);
  NR3EHD I9 (simp211_0[0:0], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  INVHHD I10 (simp211_0[1:1], gfint_3[3:3]);
  ND2HHD I11 (o_0r0[3:3], simp211_0[0:0], simp211_0[1:1]);
  NR3EHD I12 (simp221_0[0:0], gfint_0[4:4], gfint_1[4:4], gfint_2[4:4]);
  INVHHD I13 (simp221_0[1:1], gfint_3[4:4]);
  ND2HHD I14 (o_0r0[4:4], simp221_0[0:0], simp221_0[1:1]);
  NR3EHD I15 (simp231_0[0:0], gfint_0[5:5], gfint_1[5:5], gfint_2[5:5]);
  INVHHD I16 (simp231_0[1:1], gfint_3[5:5]);
  ND2HHD I17 (o_0r0[5:5], simp231_0[0:0], simp231_0[1:1]);
  NR3EHD I18 (simp241_0[0:0], gfint_0[6:6], gfint_1[6:6], gfint_2[6:6]);
  INVHHD I19 (simp241_0[1:1], gfint_3[6:6]);
  ND2HHD I20 (o_0r0[6:6], simp241_0[0:0], simp241_0[1:1]);
  NR3EHD I21 (simp251_0[0:0], gfint_0[7:7], gfint_1[7:7], gfint_2[7:7]);
  INVHHD I22 (simp251_0[1:1], gfint_3[7:7]);
  ND2HHD I23 (o_0r0[7:7], simp251_0[0:0], simp251_0[1:1]);
  NR3EHD I24 (simp261_0[0:0], gfint_0[8:8], gfint_1[8:8], gfint_2[8:8]);
  INVHHD I25 (simp261_0[1:1], gfint_3[8:8]);
  ND2HHD I26 (o_0r0[8:8], simp261_0[0:0], simp261_0[1:1]);
  NR3EHD I27 (simp271_0[0:0], gfint_0[9:9], gfint_1[9:9], gfint_2[9:9]);
  INVHHD I28 (simp271_0[1:1], gfint_3[9:9]);
  ND2HHD I29 (o_0r0[9:9], simp271_0[0:0], simp271_0[1:1]);
  NR3EHD I30 (simp281_0[0:0], gfint_0[10:10], gfint_1[10:10], gfint_2[10:10]);
  INVHHD I31 (simp281_0[1:1], gfint_3[10:10]);
  ND2HHD I32 (o_0r0[10:10], simp281_0[0:0], simp281_0[1:1]);
  NR3EHD I33 (simp291_0[0:0], gfint_0[11:11], gfint_1[11:11], gfint_2[11:11]);
  INVHHD I34 (simp291_0[1:1], gfint_3[11:11]);
  ND2HHD I35 (o_0r0[11:11], simp291_0[0:0], simp291_0[1:1]);
  NR3EHD I36 (simp301_0[0:0], gfint_0[12:12], gfint_1[12:12], gfint_2[12:12]);
  INVHHD I37 (simp301_0[1:1], gfint_3[12:12]);
  ND2HHD I38 (o_0r0[12:12], simp301_0[0:0], simp301_0[1:1]);
  NR3EHD I39 (simp311_0[0:0], gfint_0[13:13], gfint_1[13:13], gfint_2[13:13]);
  INVHHD I40 (simp311_0[1:1], gfint_3[13:13]);
  ND2HHD I41 (o_0r0[13:13], simp311_0[0:0], simp311_0[1:1]);
  NR3EHD I42 (simp321_0[0:0], gfint_0[14:14], gfint_1[14:14], gfint_2[14:14]);
  INVHHD I43 (simp321_0[1:1], gfint_3[14:14]);
  ND2HHD I44 (o_0r0[14:14], simp321_0[0:0], simp321_0[1:1]);
  NR3EHD I45 (simp331_0[0:0], gfint_0[15:15], gfint_1[15:15], gfint_2[15:15]);
  INVHHD I46 (simp331_0[1:1], gfint_3[15:15]);
  ND2HHD I47 (o_0r0[15:15], simp331_0[0:0], simp331_0[1:1]);
  NR3EHD I48 (simp341_0[0:0], gfint_0[16:16], gfint_1[16:16], gfint_2[16:16]);
  INVHHD I49 (simp341_0[1:1], gfint_3[16:16]);
  ND2HHD I50 (o_0r0[16:16], simp341_0[0:0], simp341_0[1:1]);
  NR3EHD I51 (simp351_0[0:0], gfint_0[17:17], gfint_1[17:17], gfint_2[17:17]);
  INVHHD I52 (simp351_0[1:1], gfint_3[17:17]);
  ND2HHD I53 (o_0r0[17:17], simp351_0[0:0], simp351_0[1:1]);
  NR3EHD I54 (simp361_0[0:0], gfint_0[18:18], gfint_1[18:18], gfint_2[18:18]);
  INVHHD I55 (simp361_0[1:1], gfint_3[18:18]);
  ND2HHD I56 (o_0r0[18:18], simp361_0[0:0], simp361_0[1:1]);
  NR3EHD I57 (simp371_0[0:0], gfint_0[19:19], gfint_1[19:19], gfint_2[19:19]);
  INVHHD I58 (simp371_0[1:1], gfint_3[19:19]);
  ND2HHD I59 (o_0r0[19:19], simp371_0[0:0], simp371_0[1:1]);
  NR3EHD I60 (simp381_0[0:0], gfint_0[20:20], gfint_1[20:20], gfint_2[20:20]);
  INVHHD I61 (simp381_0[1:1], gfint_3[20:20]);
  ND2HHD I62 (o_0r0[20:20], simp381_0[0:0], simp381_0[1:1]);
  NR3EHD I63 (simp391_0[0:0], gfint_0[21:21], gfint_1[21:21], gfint_2[21:21]);
  INVHHD I64 (simp391_0[1:1], gfint_3[21:21]);
  ND2HHD I65 (o_0r0[21:21], simp391_0[0:0], simp391_0[1:1]);
  NR3EHD I66 (simp401_0[0:0], gfint_0[22:22], gfint_1[22:22], gfint_2[22:22]);
  INVHHD I67 (simp401_0[1:1], gfint_3[22:22]);
  ND2HHD I68 (o_0r0[22:22], simp401_0[0:0], simp401_0[1:1]);
  NR3EHD I69 (simp411_0[0:0], gfint_0[23:23], gfint_1[23:23], gfint_2[23:23]);
  INVHHD I70 (simp411_0[1:1], gfint_3[23:23]);
  ND2HHD I71 (o_0r0[23:23], simp411_0[0:0], simp411_0[1:1]);
  NR3EHD I72 (simp421_0[0:0], gfint_0[24:24], gfint_1[24:24], gfint_2[24:24]);
  INVHHD I73 (simp421_0[1:1], gfint_3[24:24]);
  ND2HHD I74 (o_0r0[24:24], simp421_0[0:0], simp421_0[1:1]);
  NR3EHD I75 (simp431_0[0:0], gfint_0[25:25], gfint_1[25:25], gfint_2[25:25]);
  INVHHD I76 (simp431_0[1:1], gfint_3[25:25]);
  ND2HHD I77 (o_0r0[25:25], simp431_0[0:0], simp431_0[1:1]);
  NR3EHD I78 (simp441_0[0:0], gfint_0[26:26], gfint_1[26:26], gfint_2[26:26]);
  INVHHD I79 (simp441_0[1:1], gfint_3[26:26]);
  ND2HHD I80 (o_0r0[26:26], simp441_0[0:0], simp441_0[1:1]);
  NR3EHD I81 (simp451_0[0:0], gfint_0[27:27], gfint_1[27:27], gfint_2[27:27]);
  INVHHD I82 (simp451_0[1:1], gfint_3[27:27]);
  ND2HHD I83 (o_0r0[27:27], simp451_0[0:0], simp451_0[1:1]);
  NR3EHD I84 (simp461_0[0:0], gfint_0[28:28], gfint_1[28:28], gfint_2[28:28]);
  INVHHD I85 (simp461_0[1:1], gfint_3[28:28]);
  ND2HHD I86 (o_0r0[28:28], simp461_0[0:0], simp461_0[1:1]);
  NR3EHD I87 (simp471_0[0:0], gfint_0[29:29], gfint_1[29:29], gfint_2[29:29]);
  INVHHD I88 (simp471_0[1:1], gfint_3[29:29]);
  ND2HHD I89 (o_0r0[29:29], simp471_0[0:0], simp471_0[1:1]);
  NR3EHD I90 (simp481_0[0:0], gfint_0[30:30], gfint_1[30:30], gfint_2[30:30]);
  INVHHD I91 (simp481_0[1:1], gfint_3[30:30]);
  ND2HHD I92 (o_0r0[30:30], simp481_0[0:0], simp481_0[1:1]);
  NR3EHD I93 (simp491_0[0:0], gfint_0[31:31], gfint_1[31:31], gfint_2[31:31]);
  INVHHD I94 (simp491_0[1:1], gfint_3[31:31]);
  ND2HHD I95 (o_0r0[31:31], simp491_0[0:0], simp491_0[1:1]);
  NR3EHD I96 (simp501_0[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  INVHHD I97 (simp501_0[1:1], gtint_3[0:0]);
  ND2HHD I98 (o_0r1[0:0], simp501_0[0:0], simp501_0[1:1]);
  NR3EHD I99 (simp511_0[0:0], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  INVHHD I100 (simp511_0[1:1], gtint_3[1:1]);
  ND2HHD I101 (o_0r1[1:1], simp511_0[0:0], simp511_0[1:1]);
  NR3EHD I102 (simp521_0[0:0], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  INVHHD I103 (simp521_0[1:1], gtint_3[2:2]);
  ND2HHD I104 (o_0r1[2:2], simp521_0[0:0], simp521_0[1:1]);
  NR3EHD I105 (simp531_0[0:0], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  INVHHD I106 (simp531_0[1:1], gtint_3[3:3]);
  ND2HHD I107 (o_0r1[3:3], simp531_0[0:0], simp531_0[1:1]);
  NR3EHD I108 (simp541_0[0:0], gtint_0[4:4], gtint_1[4:4], gtint_2[4:4]);
  INVHHD I109 (simp541_0[1:1], gtint_3[4:4]);
  ND2HHD I110 (o_0r1[4:4], simp541_0[0:0], simp541_0[1:1]);
  NR3EHD I111 (simp551_0[0:0], gtint_0[5:5], gtint_1[5:5], gtint_2[5:5]);
  INVHHD I112 (simp551_0[1:1], gtint_3[5:5]);
  ND2HHD I113 (o_0r1[5:5], simp551_0[0:0], simp551_0[1:1]);
  NR3EHD I114 (simp561_0[0:0], gtint_0[6:6], gtint_1[6:6], gtint_2[6:6]);
  INVHHD I115 (simp561_0[1:1], gtint_3[6:6]);
  ND2HHD I116 (o_0r1[6:6], simp561_0[0:0], simp561_0[1:1]);
  NR3EHD I117 (simp571_0[0:0], gtint_0[7:7], gtint_1[7:7], gtint_2[7:7]);
  INVHHD I118 (simp571_0[1:1], gtint_3[7:7]);
  ND2HHD I119 (o_0r1[7:7], simp571_0[0:0], simp571_0[1:1]);
  NR3EHD I120 (simp581_0[0:0], gtint_0[8:8], gtint_1[8:8], gtint_2[8:8]);
  INVHHD I121 (simp581_0[1:1], gtint_3[8:8]);
  ND2HHD I122 (o_0r1[8:8], simp581_0[0:0], simp581_0[1:1]);
  NR3EHD I123 (simp591_0[0:0], gtint_0[9:9], gtint_1[9:9], gtint_2[9:9]);
  INVHHD I124 (simp591_0[1:1], gtint_3[9:9]);
  ND2HHD I125 (o_0r1[9:9], simp591_0[0:0], simp591_0[1:1]);
  NR3EHD I126 (simp601_0[0:0], gtint_0[10:10], gtint_1[10:10], gtint_2[10:10]);
  INVHHD I127 (simp601_0[1:1], gtint_3[10:10]);
  ND2HHD I128 (o_0r1[10:10], simp601_0[0:0], simp601_0[1:1]);
  NR3EHD I129 (simp611_0[0:0], gtint_0[11:11], gtint_1[11:11], gtint_2[11:11]);
  INVHHD I130 (simp611_0[1:1], gtint_3[11:11]);
  ND2HHD I131 (o_0r1[11:11], simp611_0[0:0], simp611_0[1:1]);
  NR3EHD I132 (simp621_0[0:0], gtint_0[12:12], gtint_1[12:12], gtint_2[12:12]);
  INVHHD I133 (simp621_0[1:1], gtint_3[12:12]);
  ND2HHD I134 (o_0r1[12:12], simp621_0[0:0], simp621_0[1:1]);
  NR3EHD I135 (simp631_0[0:0], gtint_0[13:13], gtint_1[13:13], gtint_2[13:13]);
  INVHHD I136 (simp631_0[1:1], gtint_3[13:13]);
  ND2HHD I137 (o_0r1[13:13], simp631_0[0:0], simp631_0[1:1]);
  NR3EHD I138 (simp641_0[0:0], gtint_0[14:14], gtint_1[14:14], gtint_2[14:14]);
  INVHHD I139 (simp641_0[1:1], gtint_3[14:14]);
  ND2HHD I140 (o_0r1[14:14], simp641_0[0:0], simp641_0[1:1]);
  NR3EHD I141 (simp651_0[0:0], gtint_0[15:15], gtint_1[15:15], gtint_2[15:15]);
  INVHHD I142 (simp651_0[1:1], gtint_3[15:15]);
  ND2HHD I143 (o_0r1[15:15], simp651_0[0:0], simp651_0[1:1]);
  NR3EHD I144 (simp661_0[0:0], gtint_0[16:16], gtint_1[16:16], gtint_2[16:16]);
  INVHHD I145 (simp661_0[1:1], gtint_3[16:16]);
  ND2HHD I146 (o_0r1[16:16], simp661_0[0:0], simp661_0[1:1]);
  NR3EHD I147 (simp671_0[0:0], gtint_0[17:17], gtint_1[17:17], gtint_2[17:17]);
  INVHHD I148 (simp671_0[1:1], gtint_3[17:17]);
  ND2HHD I149 (o_0r1[17:17], simp671_0[0:0], simp671_0[1:1]);
  NR3EHD I150 (simp681_0[0:0], gtint_0[18:18], gtint_1[18:18], gtint_2[18:18]);
  INVHHD I151 (simp681_0[1:1], gtint_3[18:18]);
  ND2HHD I152 (o_0r1[18:18], simp681_0[0:0], simp681_0[1:1]);
  NR3EHD I153 (simp691_0[0:0], gtint_0[19:19], gtint_1[19:19], gtint_2[19:19]);
  INVHHD I154 (simp691_0[1:1], gtint_3[19:19]);
  ND2HHD I155 (o_0r1[19:19], simp691_0[0:0], simp691_0[1:1]);
  NR3EHD I156 (simp701_0[0:0], gtint_0[20:20], gtint_1[20:20], gtint_2[20:20]);
  INVHHD I157 (simp701_0[1:1], gtint_3[20:20]);
  ND2HHD I158 (o_0r1[20:20], simp701_0[0:0], simp701_0[1:1]);
  NR3EHD I159 (simp711_0[0:0], gtint_0[21:21], gtint_1[21:21], gtint_2[21:21]);
  INVHHD I160 (simp711_0[1:1], gtint_3[21:21]);
  ND2HHD I161 (o_0r1[21:21], simp711_0[0:0], simp711_0[1:1]);
  NR3EHD I162 (simp721_0[0:0], gtint_0[22:22], gtint_1[22:22], gtint_2[22:22]);
  INVHHD I163 (simp721_0[1:1], gtint_3[22:22]);
  ND2HHD I164 (o_0r1[22:22], simp721_0[0:0], simp721_0[1:1]);
  NR3EHD I165 (simp731_0[0:0], gtint_0[23:23], gtint_1[23:23], gtint_2[23:23]);
  INVHHD I166 (simp731_0[1:1], gtint_3[23:23]);
  ND2HHD I167 (o_0r1[23:23], simp731_0[0:0], simp731_0[1:1]);
  NR3EHD I168 (simp741_0[0:0], gtint_0[24:24], gtint_1[24:24], gtint_2[24:24]);
  INVHHD I169 (simp741_0[1:1], gtint_3[24:24]);
  ND2HHD I170 (o_0r1[24:24], simp741_0[0:0], simp741_0[1:1]);
  NR3EHD I171 (simp751_0[0:0], gtint_0[25:25], gtint_1[25:25], gtint_2[25:25]);
  INVHHD I172 (simp751_0[1:1], gtint_3[25:25]);
  ND2HHD I173 (o_0r1[25:25], simp751_0[0:0], simp751_0[1:1]);
  NR3EHD I174 (simp761_0[0:0], gtint_0[26:26], gtint_1[26:26], gtint_2[26:26]);
  INVHHD I175 (simp761_0[1:1], gtint_3[26:26]);
  ND2HHD I176 (o_0r1[26:26], simp761_0[0:0], simp761_0[1:1]);
  NR3EHD I177 (simp771_0[0:0], gtint_0[27:27], gtint_1[27:27], gtint_2[27:27]);
  INVHHD I178 (simp771_0[1:1], gtint_3[27:27]);
  ND2HHD I179 (o_0r1[27:27], simp771_0[0:0], simp771_0[1:1]);
  NR3EHD I180 (simp781_0[0:0], gtint_0[28:28], gtint_1[28:28], gtint_2[28:28]);
  INVHHD I181 (simp781_0[1:1], gtint_3[28:28]);
  ND2HHD I182 (o_0r1[28:28], simp781_0[0:0], simp781_0[1:1]);
  NR3EHD I183 (simp791_0[0:0], gtint_0[29:29], gtint_1[29:29], gtint_2[29:29]);
  INVHHD I184 (simp791_0[1:1], gtint_3[29:29]);
  ND2HHD I185 (o_0r1[29:29], simp791_0[0:0], simp791_0[1:1]);
  NR3EHD I186 (simp801_0[0:0], gtint_0[30:30], gtint_1[30:30], gtint_2[30:30]);
  INVHHD I187 (simp801_0[1:1], gtint_3[30:30]);
  ND2HHD I188 (o_0r1[30:30], simp801_0[0:0], simp801_0[1:1]);
  NR3EHD I189 (simp811_0[0:0], gtint_0[31:31], gtint_1[31:31], gtint_2[31:31]);
  INVHHD I190 (simp811_0[1:1], gtint_3[31:31]);
  ND2HHD I191 (o_0r1[31:31], simp811_0[0:0], simp811_0[1:1]);
  AN2EHD I192 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AN2EHD I193 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AN2EHD I194 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AN2EHD I195 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AN2EHD I196 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AN2EHD I197 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AN2EHD I198 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AN2EHD I199 (gtint_0[7:7], choice_0, i_0r1[7:7]);
  AN2EHD I200 (gtint_0[8:8], choice_0, i_0r1[8:8]);
  AN2EHD I201 (gtint_0[9:9], choice_0, i_0r1[9:9]);
  AN2EHD I202 (gtint_0[10:10], choice_0, i_0r1[10:10]);
  AN2EHD I203 (gtint_0[11:11], choice_0, i_0r1[11:11]);
  AN2EHD I204 (gtint_0[12:12], choice_0, i_0r1[12:12]);
  AN2EHD I205 (gtint_0[13:13], choice_0, i_0r1[13:13]);
  AN2EHD I206 (gtint_0[14:14], choice_0, i_0r1[14:14]);
  AN2EHD I207 (gtint_0[15:15], choice_0, i_0r1[15:15]);
  AN2EHD I208 (gtint_0[16:16], choice_0, i_0r1[16:16]);
  AN2EHD I209 (gtint_0[17:17], choice_0, i_0r1[17:17]);
  AN2EHD I210 (gtint_0[18:18], choice_0, i_0r1[18:18]);
  AN2EHD I211 (gtint_0[19:19], choice_0, i_0r1[19:19]);
  AN2EHD I212 (gtint_0[20:20], choice_0, i_0r1[20:20]);
  AN2EHD I213 (gtint_0[21:21], choice_0, i_0r1[21:21]);
  AN2EHD I214 (gtint_0[22:22], choice_0, i_0r1[22:22]);
  AN2EHD I215 (gtint_0[23:23], choice_0, i_0r1[23:23]);
  AN2EHD I216 (gtint_0[24:24], choice_0, i_0r1[24:24]);
  AN2EHD I217 (gtint_0[25:25], choice_0, i_0r1[25:25]);
  AN2EHD I218 (gtint_0[26:26], choice_0, i_0r1[26:26]);
  AN2EHD I219 (gtint_0[27:27], choice_0, i_0r1[27:27]);
  AN2EHD I220 (gtint_0[28:28], choice_0, i_0r1[28:28]);
  AN2EHD I221 (gtint_0[29:29], choice_0, i_0r1[29:29]);
  AN2EHD I222 (gtint_0[30:30], choice_0, i_0r1[30:30]);
  AN2EHD I223 (gtint_0[31:31], choice_0, i_0r1[31:31]);
  AN2EHD I224 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AN2EHD I225 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AN2EHD I226 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AN2EHD I227 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AN2EHD I228 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AN2EHD I229 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AN2EHD I230 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AN2EHD I231 (gtint_1[7:7], choice_1, i_1r1[7:7]);
  AN2EHD I232 (gtint_1[8:8], choice_1, i_1r1[8:8]);
  AN2EHD I233 (gtint_1[9:9], choice_1, i_1r1[9:9]);
  AN2EHD I234 (gtint_1[10:10], choice_1, i_1r1[10:10]);
  AN2EHD I235 (gtint_1[11:11], choice_1, i_1r1[11:11]);
  AN2EHD I236 (gtint_1[12:12], choice_1, i_1r1[12:12]);
  AN2EHD I237 (gtint_1[13:13], choice_1, i_1r1[13:13]);
  AN2EHD I238 (gtint_1[14:14], choice_1, i_1r1[14:14]);
  AN2EHD I239 (gtint_1[15:15], choice_1, i_1r1[15:15]);
  AN2EHD I240 (gtint_1[16:16], choice_1, i_1r1[16:16]);
  AN2EHD I241 (gtint_1[17:17], choice_1, i_1r1[17:17]);
  AN2EHD I242 (gtint_1[18:18], choice_1, i_1r1[18:18]);
  AN2EHD I243 (gtint_1[19:19], choice_1, i_1r1[19:19]);
  AN2EHD I244 (gtint_1[20:20], choice_1, i_1r1[20:20]);
  AN2EHD I245 (gtint_1[21:21], choice_1, i_1r1[21:21]);
  AN2EHD I246 (gtint_1[22:22], choice_1, i_1r1[22:22]);
  AN2EHD I247 (gtint_1[23:23], choice_1, i_1r1[23:23]);
  AN2EHD I248 (gtint_1[24:24], choice_1, i_1r1[24:24]);
  AN2EHD I249 (gtint_1[25:25], choice_1, i_1r1[25:25]);
  AN2EHD I250 (gtint_1[26:26], choice_1, i_1r1[26:26]);
  AN2EHD I251 (gtint_1[27:27], choice_1, i_1r1[27:27]);
  AN2EHD I252 (gtint_1[28:28], choice_1, i_1r1[28:28]);
  AN2EHD I253 (gtint_1[29:29], choice_1, i_1r1[29:29]);
  AN2EHD I254 (gtint_1[30:30], choice_1, i_1r1[30:30]);
  AN2EHD I255 (gtint_1[31:31], choice_1, i_1r1[31:31]);
  AN2EHD I256 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AN2EHD I257 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AN2EHD I258 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AN2EHD I259 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AN2EHD I260 (gtint_2[4:4], choice_2, i_2r1[4:4]);
  AN2EHD I261 (gtint_2[5:5], choice_2, i_2r1[5:5]);
  AN2EHD I262 (gtint_2[6:6], choice_2, i_2r1[6:6]);
  AN2EHD I263 (gtint_2[7:7], choice_2, i_2r1[7:7]);
  AN2EHD I264 (gtint_2[8:8], choice_2, i_2r1[8:8]);
  AN2EHD I265 (gtint_2[9:9], choice_2, i_2r1[9:9]);
  AN2EHD I266 (gtint_2[10:10], choice_2, i_2r1[10:10]);
  AN2EHD I267 (gtint_2[11:11], choice_2, i_2r1[11:11]);
  AN2EHD I268 (gtint_2[12:12], choice_2, i_2r1[12:12]);
  AN2EHD I269 (gtint_2[13:13], choice_2, i_2r1[13:13]);
  AN2EHD I270 (gtint_2[14:14], choice_2, i_2r1[14:14]);
  AN2EHD I271 (gtint_2[15:15], choice_2, i_2r1[15:15]);
  AN2EHD I272 (gtint_2[16:16], choice_2, i_2r1[16:16]);
  AN2EHD I273 (gtint_2[17:17], choice_2, i_2r1[17:17]);
  AN2EHD I274 (gtint_2[18:18], choice_2, i_2r1[18:18]);
  AN2EHD I275 (gtint_2[19:19], choice_2, i_2r1[19:19]);
  AN2EHD I276 (gtint_2[20:20], choice_2, i_2r1[20:20]);
  AN2EHD I277 (gtint_2[21:21], choice_2, i_2r1[21:21]);
  AN2EHD I278 (gtint_2[22:22], choice_2, i_2r1[22:22]);
  AN2EHD I279 (gtint_2[23:23], choice_2, i_2r1[23:23]);
  AN2EHD I280 (gtint_2[24:24], choice_2, i_2r1[24:24]);
  AN2EHD I281 (gtint_2[25:25], choice_2, i_2r1[25:25]);
  AN2EHD I282 (gtint_2[26:26], choice_2, i_2r1[26:26]);
  AN2EHD I283 (gtint_2[27:27], choice_2, i_2r1[27:27]);
  AN2EHD I284 (gtint_2[28:28], choice_2, i_2r1[28:28]);
  AN2EHD I285 (gtint_2[29:29], choice_2, i_2r1[29:29]);
  AN2EHD I286 (gtint_2[30:30], choice_2, i_2r1[30:30]);
  AN2EHD I287 (gtint_2[31:31], choice_2, i_2r1[31:31]);
  AN2EHD I288 (gtint_3[0:0], choice_3, i_3r1[0:0]);
  AN2EHD I289 (gtint_3[1:1], choice_3, i_3r1[1:1]);
  AN2EHD I290 (gtint_3[2:2], choice_3, i_3r1[2:2]);
  AN2EHD I291 (gtint_3[3:3], choice_3, i_3r1[3:3]);
  AN2EHD I292 (gtint_3[4:4], choice_3, i_3r1[4:4]);
  AN2EHD I293 (gtint_3[5:5], choice_3, i_3r1[5:5]);
  AN2EHD I294 (gtint_3[6:6], choice_3, i_3r1[6:6]);
  AN2EHD I295 (gtint_3[7:7], choice_3, i_3r1[7:7]);
  AN2EHD I296 (gtint_3[8:8], choice_3, i_3r1[8:8]);
  AN2EHD I297 (gtint_3[9:9], choice_3, i_3r1[9:9]);
  AN2EHD I298 (gtint_3[10:10], choice_3, i_3r1[10:10]);
  AN2EHD I299 (gtint_3[11:11], choice_3, i_3r1[11:11]);
  AN2EHD I300 (gtint_3[12:12], choice_3, i_3r1[12:12]);
  AN2EHD I301 (gtint_3[13:13], choice_3, i_3r1[13:13]);
  AN2EHD I302 (gtint_3[14:14], choice_3, i_3r1[14:14]);
  AN2EHD I303 (gtint_3[15:15], choice_3, i_3r1[15:15]);
  AN2EHD I304 (gtint_3[16:16], choice_3, i_3r1[16:16]);
  AN2EHD I305 (gtint_3[17:17], choice_3, i_3r1[17:17]);
  AN2EHD I306 (gtint_3[18:18], choice_3, i_3r1[18:18]);
  AN2EHD I307 (gtint_3[19:19], choice_3, i_3r1[19:19]);
  AN2EHD I308 (gtint_3[20:20], choice_3, i_3r1[20:20]);
  AN2EHD I309 (gtint_3[21:21], choice_3, i_3r1[21:21]);
  AN2EHD I310 (gtint_3[22:22], choice_3, i_3r1[22:22]);
  AN2EHD I311 (gtint_3[23:23], choice_3, i_3r1[23:23]);
  AN2EHD I312 (gtint_3[24:24], choice_3, i_3r1[24:24]);
  AN2EHD I313 (gtint_3[25:25], choice_3, i_3r1[25:25]);
  AN2EHD I314 (gtint_3[26:26], choice_3, i_3r1[26:26]);
  AN2EHD I315 (gtint_3[27:27], choice_3, i_3r1[27:27]);
  AN2EHD I316 (gtint_3[28:28], choice_3, i_3r1[28:28]);
  AN2EHD I317 (gtint_3[29:29], choice_3, i_3r1[29:29]);
  AN2EHD I318 (gtint_3[30:30], choice_3, i_3r1[30:30]);
  AN2EHD I319 (gtint_3[31:31], choice_3, i_3r1[31:31]);
  AN2EHD I320 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AN2EHD I321 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AN2EHD I322 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AN2EHD I323 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AN2EHD I324 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AN2EHD I325 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AN2EHD I326 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AN2EHD I327 (gfint_0[7:7], choice_0, i_0r0[7:7]);
  AN2EHD I328 (gfint_0[8:8], choice_0, i_0r0[8:8]);
  AN2EHD I329 (gfint_0[9:9], choice_0, i_0r0[9:9]);
  AN2EHD I330 (gfint_0[10:10], choice_0, i_0r0[10:10]);
  AN2EHD I331 (gfint_0[11:11], choice_0, i_0r0[11:11]);
  AN2EHD I332 (gfint_0[12:12], choice_0, i_0r0[12:12]);
  AN2EHD I333 (gfint_0[13:13], choice_0, i_0r0[13:13]);
  AN2EHD I334 (gfint_0[14:14], choice_0, i_0r0[14:14]);
  AN2EHD I335 (gfint_0[15:15], choice_0, i_0r0[15:15]);
  AN2EHD I336 (gfint_0[16:16], choice_0, i_0r0[16:16]);
  AN2EHD I337 (gfint_0[17:17], choice_0, i_0r0[17:17]);
  AN2EHD I338 (gfint_0[18:18], choice_0, i_0r0[18:18]);
  AN2EHD I339 (gfint_0[19:19], choice_0, i_0r0[19:19]);
  AN2EHD I340 (gfint_0[20:20], choice_0, i_0r0[20:20]);
  AN2EHD I341 (gfint_0[21:21], choice_0, i_0r0[21:21]);
  AN2EHD I342 (gfint_0[22:22], choice_0, i_0r0[22:22]);
  AN2EHD I343 (gfint_0[23:23], choice_0, i_0r0[23:23]);
  AN2EHD I344 (gfint_0[24:24], choice_0, i_0r0[24:24]);
  AN2EHD I345 (gfint_0[25:25], choice_0, i_0r0[25:25]);
  AN2EHD I346 (gfint_0[26:26], choice_0, i_0r0[26:26]);
  AN2EHD I347 (gfint_0[27:27], choice_0, i_0r0[27:27]);
  AN2EHD I348 (gfint_0[28:28], choice_0, i_0r0[28:28]);
  AN2EHD I349 (gfint_0[29:29], choice_0, i_0r0[29:29]);
  AN2EHD I350 (gfint_0[30:30], choice_0, i_0r0[30:30]);
  AN2EHD I351 (gfint_0[31:31], choice_0, i_0r0[31:31]);
  AN2EHD I352 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AN2EHD I353 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AN2EHD I354 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AN2EHD I355 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AN2EHD I356 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AN2EHD I357 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AN2EHD I358 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AN2EHD I359 (gfint_1[7:7], choice_1, i_1r0[7:7]);
  AN2EHD I360 (gfint_1[8:8], choice_1, i_1r0[8:8]);
  AN2EHD I361 (gfint_1[9:9], choice_1, i_1r0[9:9]);
  AN2EHD I362 (gfint_1[10:10], choice_1, i_1r0[10:10]);
  AN2EHD I363 (gfint_1[11:11], choice_1, i_1r0[11:11]);
  AN2EHD I364 (gfint_1[12:12], choice_1, i_1r0[12:12]);
  AN2EHD I365 (gfint_1[13:13], choice_1, i_1r0[13:13]);
  AN2EHD I366 (gfint_1[14:14], choice_1, i_1r0[14:14]);
  AN2EHD I367 (gfint_1[15:15], choice_1, i_1r0[15:15]);
  AN2EHD I368 (gfint_1[16:16], choice_1, i_1r0[16:16]);
  AN2EHD I369 (gfint_1[17:17], choice_1, i_1r0[17:17]);
  AN2EHD I370 (gfint_1[18:18], choice_1, i_1r0[18:18]);
  AN2EHD I371 (gfint_1[19:19], choice_1, i_1r0[19:19]);
  AN2EHD I372 (gfint_1[20:20], choice_1, i_1r0[20:20]);
  AN2EHD I373 (gfint_1[21:21], choice_1, i_1r0[21:21]);
  AN2EHD I374 (gfint_1[22:22], choice_1, i_1r0[22:22]);
  AN2EHD I375 (gfint_1[23:23], choice_1, i_1r0[23:23]);
  AN2EHD I376 (gfint_1[24:24], choice_1, i_1r0[24:24]);
  AN2EHD I377 (gfint_1[25:25], choice_1, i_1r0[25:25]);
  AN2EHD I378 (gfint_1[26:26], choice_1, i_1r0[26:26]);
  AN2EHD I379 (gfint_1[27:27], choice_1, i_1r0[27:27]);
  AN2EHD I380 (gfint_1[28:28], choice_1, i_1r0[28:28]);
  AN2EHD I381 (gfint_1[29:29], choice_1, i_1r0[29:29]);
  AN2EHD I382 (gfint_1[30:30], choice_1, i_1r0[30:30]);
  AN2EHD I383 (gfint_1[31:31], choice_1, i_1r0[31:31]);
  AN2EHD I384 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AN2EHD I385 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AN2EHD I386 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AN2EHD I387 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AN2EHD I388 (gfint_2[4:4], choice_2, i_2r0[4:4]);
  AN2EHD I389 (gfint_2[5:5], choice_2, i_2r0[5:5]);
  AN2EHD I390 (gfint_2[6:6], choice_2, i_2r0[6:6]);
  AN2EHD I391 (gfint_2[7:7], choice_2, i_2r0[7:7]);
  AN2EHD I392 (gfint_2[8:8], choice_2, i_2r0[8:8]);
  AN2EHD I393 (gfint_2[9:9], choice_2, i_2r0[9:9]);
  AN2EHD I394 (gfint_2[10:10], choice_2, i_2r0[10:10]);
  AN2EHD I395 (gfint_2[11:11], choice_2, i_2r0[11:11]);
  AN2EHD I396 (gfint_2[12:12], choice_2, i_2r0[12:12]);
  AN2EHD I397 (gfint_2[13:13], choice_2, i_2r0[13:13]);
  AN2EHD I398 (gfint_2[14:14], choice_2, i_2r0[14:14]);
  AN2EHD I399 (gfint_2[15:15], choice_2, i_2r0[15:15]);
  AN2EHD I400 (gfint_2[16:16], choice_2, i_2r0[16:16]);
  AN2EHD I401 (gfint_2[17:17], choice_2, i_2r0[17:17]);
  AN2EHD I402 (gfint_2[18:18], choice_2, i_2r0[18:18]);
  AN2EHD I403 (gfint_2[19:19], choice_2, i_2r0[19:19]);
  AN2EHD I404 (gfint_2[20:20], choice_2, i_2r0[20:20]);
  AN2EHD I405 (gfint_2[21:21], choice_2, i_2r0[21:21]);
  AN2EHD I406 (gfint_2[22:22], choice_2, i_2r0[22:22]);
  AN2EHD I407 (gfint_2[23:23], choice_2, i_2r0[23:23]);
  AN2EHD I408 (gfint_2[24:24], choice_2, i_2r0[24:24]);
  AN2EHD I409 (gfint_2[25:25], choice_2, i_2r0[25:25]);
  AN2EHD I410 (gfint_2[26:26], choice_2, i_2r0[26:26]);
  AN2EHD I411 (gfint_2[27:27], choice_2, i_2r0[27:27]);
  AN2EHD I412 (gfint_2[28:28], choice_2, i_2r0[28:28]);
  AN2EHD I413 (gfint_2[29:29], choice_2, i_2r0[29:29]);
  AN2EHD I414 (gfint_2[30:30], choice_2, i_2r0[30:30]);
  AN2EHD I415 (gfint_2[31:31], choice_2, i_2r0[31:31]);
  AN2EHD I416 (gfint_3[0:0], choice_3, i_3r0[0:0]);
  AN2EHD I417 (gfint_3[1:1], choice_3, i_3r0[1:1]);
  AN2EHD I418 (gfint_3[2:2], choice_3, i_3r0[2:2]);
  AN2EHD I419 (gfint_3[3:3], choice_3, i_3r0[3:3]);
  AN2EHD I420 (gfint_3[4:4], choice_3, i_3r0[4:4]);
  AN2EHD I421 (gfint_3[5:5], choice_3, i_3r0[5:5]);
  AN2EHD I422 (gfint_3[6:6], choice_3, i_3r0[6:6]);
  AN2EHD I423 (gfint_3[7:7], choice_3, i_3r0[7:7]);
  AN2EHD I424 (gfint_3[8:8], choice_3, i_3r0[8:8]);
  AN2EHD I425 (gfint_3[9:9], choice_3, i_3r0[9:9]);
  AN2EHD I426 (gfint_3[10:10], choice_3, i_3r0[10:10]);
  AN2EHD I427 (gfint_3[11:11], choice_3, i_3r0[11:11]);
  AN2EHD I428 (gfint_3[12:12], choice_3, i_3r0[12:12]);
  AN2EHD I429 (gfint_3[13:13], choice_3, i_3r0[13:13]);
  AN2EHD I430 (gfint_3[14:14], choice_3, i_3r0[14:14]);
  AN2EHD I431 (gfint_3[15:15], choice_3, i_3r0[15:15]);
  AN2EHD I432 (gfint_3[16:16], choice_3, i_3r0[16:16]);
  AN2EHD I433 (gfint_3[17:17], choice_3, i_3r0[17:17]);
  AN2EHD I434 (gfint_3[18:18], choice_3, i_3r0[18:18]);
  AN2EHD I435 (gfint_3[19:19], choice_3, i_3r0[19:19]);
  AN2EHD I436 (gfint_3[20:20], choice_3, i_3r0[20:20]);
  AN2EHD I437 (gfint_3[21:21], choice_3, i_3r0[21:21]);
  AN2EHD I438 (gfint_3[22:22], choice_3, i_3r0[22:22]);
  AN2EHD I439 (gfint_3[23:23], choice_3, i_3r0[23:23]);
  AN2EHD I440 (gfint_3[24:24], choice_3, i_3r0[24:24]);
  AN2EHD I441 (gfint_3[25:25], choice_3, i_3r0[25:25]);
  AN2EHD I442 (gfint_3[26:26], choice_3, i_3r0[26:26]);
  AN2EHD I443 (gfint_3[27:27], choice_3, i_3r0[27:27]);
  AN2EHD I444 (gfint_3[28:28], choice_3, i_3r0[28:28]);
  AN2EHD I445 (gfint_3[29:29], choice_3, i_3r0[29:29]);
  AN2EHD I446 (gfint_3[30:30], choice_3, i_3r0[30:30]);
  AN2EHD I447 (gfint_3[31:31], choice_3, i_3r0[31:31]);
  OR2EHD I448 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2EHD I449 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2EHD I450 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2EHD I451 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2EHD I452 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2EHD I453 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2EHD I454 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2EHD I455 (comp0_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2EHD I456 (comp0_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2EHD I457 (comp0_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2EHD I458 (comp0_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2EHD I459 (comp0_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2EHD I460 (comp0_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2EHD I461 (comp0_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2EHD I462 (comp0_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2EHD I463 (comp0_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2EHD I464 (comp0_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2EHD I465 (comp0_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2EHD I466 (comp0_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2EHD I467 (comp0_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2EHD I468 (comp0_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2EHD I469 (comp0_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2EHD I470 (comp0_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2EHD I471 (comp0_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2EHD I472 (comp0_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2EHD I473 (comp0_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2EHD I474 (comp0_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2EHD I475 (comp0_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2EHD I476 (comp0_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2EHD I477 (comp0_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2EHD I478 (comp0_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2EHD I479 (comp0_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  AO222EHD I480 (tech564_int, comp0_0[0:0], comp0_0[1:1], tech564_int, comp0_0[0:0], tech564_int, comp0_0[1:1]);
  AO222EHD I481 (simp3711_0[0:0], tech564_int, comp0_0[2:2], simp3711_0[0:0], tech564_int, simp3711_0[0:0], comp0_0[2:2]);
  AO222EHD I482 (tech565_int, comp0_0[3:3], comp0_0[4:4], tech565_int, comp0_0[3:3], tech565_int, comp0_0[4:4]);
  AO222EHD I483 (simp3711_0[1:1], tech565_int, comp0_0[5:5], simp3711_0[1:1], tech565_int, simp3711_0[1:1], comp0_0[5:5]);
  AO222EHD I484 (tech566_int, comp0_0[6:6], comp0_0[7:7], tech566_int, comp0_0[6:6], tech566_int, comp0_0[7:7]);
  AO222EHD I485 (simp3711_0[2:2], tech566_int, comp0_0[8:8], simp3711_0[2:2], tech566_int, simp3711_0[2:2], comp0_0[8:8]);
  AO222EHD I486 (tech567_int, comp0_0[9:9], comp0_0[10:10], tech567_int, comp0_0[9:9], tech567_int, comp0_0[10:10]);
  AO222EHD I487 (simp3711_0[3:3], tech567_int, comp0_0[11:11], simp3711_0[3:3], tech567_int, simp3711_0[3:3], comp0_0[11:11]);
  AO222EHD I488 (tech568_int, comp0_0[12:12], comp0_0[13:13], tech568_int, comp0_0[12:12], tech568_int, comp0_0[13:13]);
  AO222EHD I489 (simp3711_0[4:4], tech568_int, comp0_0[14:14], simp3711_0[4:4], tech568_int, simp3711_0[4:4], comp0_0[14:14]);
  AO222EHD I490 (tech569_int, comp0_0[15:15], comp0_0[16:16], tech569_int, comp0_0[15:15], tech569_int, comp0_0[16:16]);
  AO222EHD I491 (simp3711_0[5:5], tech569_int, comp0_0[17:17], simp3711_0[5:5], tech569_int, simp3711_0[5:5], comp0_0[17:17]);
  AO222EHD I492 (tech570_int, comp0_0[18:18], comp0_0[19:19], tech570_int, comp0_0[18:18], tech570_int, comp0_0[19:19]);
  AO222EHD I493 (simp3711_0[6:6], tech570_int, comp0_0[20:20], simp3711_0[6:6], tech570_int, simp3711_0[6:6], comp0_0[20:20]);
  AO222EHD I494 (tech571_int, comp0_0[21:21], comp0_0[22:22], tech571_int, comp0_0[21:21], tech571_int, comp0_0[22:22]);
  AO222EHD I495 (simp3711_0[7:7], tech571_int, comp0_0[23:23], simp3711_0[7:7], tech571_int, simp3711_0[7:7], comp0_0[23:23]);
  AO222EHD I496 (tech572_int, comp0_0[24:24], comp0_0[25:25], tech572_int, comp0_0[24:24], tech572_int, comp0_0[25:25]);
  AO222EHD I497 (simp3711_0[8:8], tech572_int, comp0_0[26:26], simp3711_0[8:8], tech572_int, simp3711_0[8:8], comp0_0[26:26]);
  AO222EHD I498 (tech573_int, comp0_0[27:27], comp0_0[28:28], tech573_int, comp0_0[27:27], tech573_int, comp0_0[28:28]);
  AO222EHD I499 (simp3711_0[9:9], tech573_int, comp0_0[29:29], simp3711_0[9:9], tech573_int, simp3711_0[9:9], comp0_0[29:29]);
  AO222EHD I500 (simp3711_0[10:10], comp0_0[30:30], comp0_0[31:31], simp3711_0[10:10], comp0_0[30:30], simp3711_0[10:10], comp0_0[31:31]);
  AO222EHD I501 (tech576_int, simp3711_0[0:0], simp3711_0[1:1], tech576_int, simp3711_0[0:0], tech576_int, simp3711_0[1:1]);
  AO222EHD I502 (simp3712_0[0:0], tech576_int, simp3711_0[2:2], simp3712_0[0:0], tech576_int, simp3712_0[0:0], simp3711_0[2:2]);
  AO222EHD I503 (tech577_int, simp3711_0[3:3], simp3711_0[4:4], tech577_int, simp3711_0[3:3], tech577_int, simp3711_0[4:4]);
  AO222EHD I504 (simp3712_0[1:1], tech577_int, simp3711_0[5:5], simp3712_0[1:1], tech577_int, simp3712_0[1:1], simp3711_0[5:5]);
  AO222EHD I505 (tech578_int, simp3711_0[6:6], simp3711_0[7:7], tech578_int, simp3711_0[6:6], tech578_int, simp3711_0[7:7]);
  AO222EHD I506 (simp3712_0[2:2], tech578_int, simp3711_0[8:8], simp3712_0[2:2], tech578_int, simp3712_0[2:2], simp3711_0[8:8]);
  AO222EHD I507 (simp3712_0[3:3], simp3711_0[9:9], simp3711_0[10:10], simp3712_0[3:3], simp3711_0[9:9], simp3712_0[3:3], simp3711_0[10:10]);
  AO222EHD I508 (tech581_int, simp3712_0[0:0], simp3712_0[1:1], tech581_int, simp3712_0[0:0], tech581_int, simp3712_0[1:1]);
  AO222EHD I509 (simp3713_0[0:0], tech581_int, simp3712_0[2:2], simp3713_0[0:0], tech581_int, simp3713_0[0:0], simp3712_0[2:2]);
  BUFEHD I510 (simp3713_0[1:1], simp3712_0[3:3]);
  AO222EHD I511 (icomp_0, simp3713_0[0:0], simp3713_0[1:1], icomp_0, simp3713_0[0:0], icomp_0, simp3713_0[1:1]);
  OR2EHD I512 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2EHD I513 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2EHD I514 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2EHD I515 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2EHD I516 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2EHD I517 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2EHD I518 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  OR2EHD I519 (comp1_0[7:7], i_1r0[7:7], i_1r1[7:7]);
  OR2EHD I520 (comp1_0[8:8], i_1r0[8:8], i_1r1[8:8]);
  OR2EHD I521 (comp1_0[9:9], i_1r0[9:9], i_1r1[9:9]);
  OR2EHD I522 (comp1_0[10:10], i_1r0[10:10], i_1r1[10:10]);
  OR2EHD I523 (comp1_0[11:11], i_1r0[11:11], i_1r1[11:11]);
  OR2EHD I524 (comp1_0[12:12], i_1r0[12:12], i_1r1[12:12]);
  OR2EHD I525 (comp1_0[13:13], i_1r0[13:13], i_1r1[13:13]);
  OR2EHD I526 (comp1_0[14:14], i_1r0[14:14], i_1r1[14:14]);
  OR2EHD I527 (comp1_0[15:15], i_1r0[15:15], i_1r1[15:15]);
  OR2EHD I528 (comp1_0[16:16], i_1r0[16:16], i_1r1[16:16]);
  OR2EHD I529 (comp1_0[17:17], i_1r0[17:17], i_1r1[17:17]);
  OR2EHD I530 (comp1_0[18:18], i_1r0[18:18], i_1r1[18:18]);
  OR2EHD I531 (comp1_0[19:19], i_1r0[19:19], i_1r1[19:19]);
  OR2EHD I532 (comp1_0[20:20], i_1r0[20:20], i_1r1[20:20]);
  OR2EHD I533 (comp1_0[21:21], i_1r0[21:21], i_1r1[21:21]);
  OR2EHD I534 (comp1_0[22:22], i_1r0[22:22], i_1r1[22:22]);
  OR2EHD I535 (comp1_0[23:23], i_1r0[23:23], i_1r1[23:23]);
  OR2EHD I536 (comp1_0[24:24], i_1r0[24:24], i_1r1[24:24]);
  OR2EHD I537 (comp1_0[25:25], i_1r0[25:25], i_1r1[25:25]);
  OR2EHD I538 (comp1_0[26:26], i_1r0[26:26], i_1r1[26:26]);
  OR2EHD I539 (comp1_0[27:27], i_1r0[27:27], i_1r1[27:27]);
  OR2EHD I540 (comp1_0[28:28], i_1r0[28:28], i_1r1[28:28]);
  OR2EHD I541 (comp1_0[29:29], i_1r0[29:29], i_1r1[29:29]);
  OR2EHD I542 (comp1_0[30:30], i_1r0[30:30], i_1r1[30:30]);
  OR2EHD I543 (comp1_0[31:31], i_1r0[31:31], i_1r1[31:31]);
  AO222EHD I544 (tech618_int, comp1_0[0:0], comp1_0[1:1], tech618_int, comp1_0[0:0], tech618_int, comp1_0[1:1]);
  AO222EHD I545 (simp4051_0[0:0], tech618_int, comp1_0[2:2], simp4051_0[0:0], tech618_int, simp4051_0[0:0], comp1_0[2:2]);
  AO222EHD I546 (tech619_int, comp1_0[3:3], comp1_0[4:4], tech619_int, comp1_0[3:3], tech619_int, comp1_0[4:4]);
  AO222EHD I547 (simp4051_0[1:1], tech619_int, comp1_0[5:5], simp4051_0[1:1], tech619_int, simp4051_0[1:1], comp1_0[5:5]);
  AO222EHD I548 (tech620_int, comp1_0[6:6], comp1_0[7:7], tech620_int, comp1_0[6:6], tech620_int, comp1_0[7:7]);
  AO222EHD I549 (simp4051_0[2:2], tech620_int, comp1_0[8:8], simp4051_0[2:2], tech620_int, simp4051_0[2:2], comp1_0[8:8]);
  AO222EHD I550 (tech621_int, comp1_0[9:9], comp1_0[10:10], tech621_int, comp1_0[9:9], tech621_int, comp1_0[10:10]);
  AO222EHD I551 (simp4051_0[3:3], tech621_int, comp1_0[11:11], simp4051_0[3:3], tech621_int, simp4051_0[3:3], comp1_0[11:11]);
  AO222EHD I552 (tech622_int, comp1_0[12:12], comp1_0[13:13], tech622_int, comp1_0[12:12], tech622_int, comp1_0[13:13]);
  AO222EHD I553 (simp4051_0[4:4], tech622_int, comp1_0[14:14], simp4051_0[4:4], tech622_int, simp4051_0[4:4], comp1_0[14:14]);
  AO222EHD I554 (tech623_int, comp1_0[15:15], comp1_0[16:16], tech623_int, comp1_0[15:15], tech623_int, comp1_0[16:16]);
  AO222EHD I555 (simp4051_0[5:5], tech623_int, comp1_0[17:17], simp4051_0[5:5], tech623_int, simp4051_0[5:5], comp1_0[17:17]);
  AO222EHD I556 (tech624_int, comp1_0[18:18], comp1_0[19:19], tech624_int, comp1_0[18:18], tech624_int, comp1_0[19:19]);
  AO222EHD I557 (simp4051_0[6:6], tech624_int, comp1_0[20:20], simp4051_0[6:6], tech624_int, simp4051_0[6:6], comp1_0[20:20]);
  AO222EHD I558 (tech625_int, comp1_0[21:21], comp1_0[22:22], tech625_int, comp1_0[21:21], tech625_int, comp1_0[22:22]);
  AO222EHD I559 (simp4051_0[7:7], tech625_int, comp1_0[23:23], simp4051_0[7:7], tech625_int, simp4051_0[7:7], comp1_0[23:23]);
  AO222EHD I560 (tech626_int, comp1_0[24:24], comp1_0[25:25], tech626_int, comp1_0[24:24], tech626_int, comp1_0[25:25]);
  AO222EHD I561 (simp4051_0[8:8], tech626_int, comp1_0[26:26], simp4051_0[8:8], tech626_int, simp4051_0[8:8], comp1_0[26:26]);
  AO222EHD I562 (tech627_int, comp1_0[27:27], comp1_0[28:28], tech627_int, comp1_0[27:27], tech627_int, comp1_0[28:28]);
  AO222EHD I563 (simp4051_0[9:9], tech627_int, comp1_0[29:29], simp4051_0[9:9], tech627_int, simp4051_0[9:9], comp1_0[29:29]);
  AO222EHD I564 (simp4051_0[10:10], comp1_0[30:30], comp1_0[31:31], simp4051_0[10:10], comp1_0[30:30], simp4051_0[10:10], comp1_0[31:31]);
  AO222EHD I565 (tech630_int, simp4051_0[0:0], simp4051_0[1:1], tech630_int, simp4051_0[0:0], tech630_int, simp4051_0[1:1]);
  AO222EHD I566 (simp4052_0[0:0], tech630_int, simp4051_0[2:2], simp4052_0[0:0], tech630_int, simp4052_0[0:0], simp4051_0[2:2]);
  AO222EHD I567 (tech631_int, simp4051_0[3:3], simp4051_0[4:4], tech631_int, simp4051_0[3:3], tech631_int, simp4051_0[4:4]);
  AO222EHD I568 (simp4052_0[1:1], tech631_int, simp4051_0[5:5], simp4052_0[1:1], tech631_int, simp4052_0[1:1], simp4051_0[5:5]);
  AO222EHD I569 (tech632_int, simp4051_0[6:6], simp4051_0[7:7], tech632_int, simp4051_0[6:6], tech632_int, simp4051_0[7:7]);
  AO222EHD I570 (simp4052_0[2:2], tech632_int, simp4051_0[8:8], simp4052_0[2:2], tech632_int, simp4052_0[2:2], simp4051_0[8:8]);
  AO222EHD I571 (simp4052_0[3:3], simp4051_0[9:9], simp4051_0[10:10], simp4052_0[3:3], simp4051_0[9:9], simp4052_0[3:3], simp4051_0[10:10]);
  AO222EHD I572 (tech635_int, simp4052_0[0:0], simp4052_0[1:1], tech635_int, simp4052_0[0:0], tech635_int, simp4052_0[1:1]);
  AO222EHD I573 (simp4053_0[0:0], tech635_int, simp4052_0[2:2], simp4053_0[0:0], tech635_int, simp4053_0[0:0], simp4052_0[2:2]);
  BUFEHD I574 (simp4053_0[1:1], simp4052_0[3:3]);
  AO222EHD I575 (icomp_1, simp4053_0[0:0], simp4053_0[1:1], icomp_1, simp4053_0[0:0], icomp_1, simp4053_0[1:1]);
  OR2EHD I576 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2EHD I577 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2EHD I578 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2EHD I579 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  OR2EHD I580 (comp2_0[4:4], i_2r0[4:4], i_2r1[4:4]);
  OR2EHD I581 (comp2_0[5:5], i_2r0[5:5], i_2r1[5:5]);
  OR2EHD I582 (comp2_0[6:6], i_2r0[6:6], i_2r1[6:6]);
  OR2EHD I583 (comp2_0[7:7], i_2r0[7:7], i_2r1[7:7]);
  OR2EHD I584 (comp2_0[8:8], i_2r0[8:8], i_2r1[8:8]);
  OR2EHD I585 (comp2_0[9:9], i_2r0[9:9], i_2r1[9:9]);
  OR2EHD I586 (comp2_0[10:10], i_2r0[10:10], i_2r1[10:10]);
  OR2EHD I587 (comp2_0[11:11], i_2r0[11:11], i_2r1[11:11]);
  OR2EHD I588 (comp2_0[12:12], i_2r0[12:12], i_2r1[12:12]);
  OR2EHD I589 (comp2_0[13:13], i_2r0[13:13], i_2r1[13:13]);
  OR2EHD I590 (comp2_0[14:14], i_2r0[14:14], i_2r1[14:14]);
  OR2EHD I591 (comp2_0[15:15], i_2r0[15:15], i_2r1[15:15]);
  OR2EHD I592 (comp2_0[16:16], i_2r0[16:16], i_2r1[16:16]);
  OR2EHD I593 (comp2_0[17:17], i_2r0[17:17], i_2r1[17:17]);
  OR2EHD I594 (comp2_0[18:18], i_2r0[18:18], i_2r1[18:18]);
  OR2EHD I595 (comp2_0[19:19], i_2r0[19:19], i_2r1[19:19]);
  OR2EHD I596 (comp2_0[20:20], i_2r0[20:20], i_2r1[20:20]);
  OR2EHD I597 (comp2_0[21:21], i_2r0[21:21], i_2r1[21:21]);
  OR2EHD I598 (comp2_0[22:22], i_2r0[22:22], i_2r1[22:22]);
  OR2EHD I599 (comp2_0[23:23], i_2r0[23:23], i_2r1[23:23]);
  OR2EHD I600 (comp2_0[24:24], i_2r0[24:24], i_2r1[24:24]);
  OR2EHD I601 (comp2_0[25:25], i_2r0[25:25], i_2r1[25:25]);
  OR2EHD I602 (comp2_0[26:26], i_2r0[26:26], i_2r1[26:26]);
  OR2EHD I603 (comp2_0[27:27], i_2r0[27:27], i_2r1[27:27]);
  OR2EHD I604 (comp2_0[28:28], i_2r0[28:28], i_2r1[28:28]);
  OR2EHD I605 (comp2_0[29:29], i_2r0[29:29], i_2r1[29:29]);
  OR2EHD I606 (comp2_0[30:30], i_2r0[30:30], i_2r1[30:30]);
  OR2EHD I607 (comp2_0[31:31], i_2r0[31:31], i_2r1[31:31]);
  AO222EHD I608 (tech672_int, comp2_0[0:0], comp2_0[1:1], tech672_int, comp2_0[0:0], tech672_int, comp2_0[1:1]);
  AO222EHD I609 (simp4391_0[0:0], tech672_int, comp2_0[2:2], simp4391_0[0:0], tech672_int, simp4391_0[0:0], comp2_0[2:2]);
  AO222EHD I610 (tech673_int, comp2_0[3:3], comp2_0[4:4], tech673_int, comp2_0[3:3], tech673_int, comp2_0[4:4]);
  AO222EHD I611 (simp4391_0[1:1], tech673_int, comp2_0[5:5], simp4391_0[1:1], tech673_int, simp4391_0[1:1], comp2_0[5:5]);
  AO222EHD I612 (tech674_int, comp2_0[6:6], comp2_0[7:7], tech674_int, comp2_0[6:6], tech674_int, comp2_0[7:7]);
  AO222EHD I613 (simp4391_0[2:2], tech674_int, comp2_0[8:8], simp4391_0[2:2], tech674_int, simp4391_0[2:2], comp2_0[8:8]);
  AO222EHD I614 (tech675_int, comp2_0[9:9], comp2_0[10:10], tech675_int, comp2_0[9:9], tech675_int, comp2_0[10:10]);
  AO222EHD I615 (simp4391_0[3:3], tech675_int, comp2_0[11:11], simp4391_0[3:3], tech675_int, simp4391_0[3:3], comp2_0[11:11]);
  AO222EHD I616 (tech676_int, comp2_0[12:12], comp2_0[13:13], tech676_int, comp2_0[12:12], tech676_int, comp2_0[13:13]);
  AO222EHD I617 (simp4391_0[4:4], tech676_int, comp2_0[14:14], simp4391_0[4:4], tech676_int, simp4391_0[4:4], comp2_0[14:14]);
  AO222EHD I618 (tech677_int, comp2_0[15:15], comp2_0[16:16], tech677_int, comp2_0[15:15], tech677_int, comp2_0[16:16]);
  AO222EHD I619 (simp4391_0[5:5], tech677_int, comp2_0[17:17], simp4391_0[5:5], tech677_int, simp4391_0[5:5], comp2_0[17:17]);
  AO222EHD I620 (tech678_int, comp2_0[18:18], comp2_0[19:19], tech678_int, comp2_0[18:18], tech678_int, comp2_0[19:19]);
  AO222EHD I621 (simp4391_0[6:6], tech678_int, comp2_0[20:20], simp4391_0[6:6], tech678_int, simp4391_0[6:6], comp2_0[20:20]);
  AO222EHD I622 (tech679_int, comp2_0[21:21], comp2_0[22:22], tech679_int, comp2_0[21:21], tech679_int, comp2_0[22:22]);
  AO222EHD I623 (simp4391_0[7:7], tech679_int, comp2_0[23:23], simp4391_0[7:7], tech679_int, simp4391_0[7:7], comp2_0[23:23]);
  AO222EHD I624 (tech680_int, comp2_0[24:24], comp2_0[25:25], tech680_int, comp2_0[24:24], tech680_int, comp2_0[25:25]);
  AO222EHD I625 (simp4391_0[8:8], tech680_int, comp2_0[26:26], simp4391_0[8:8], tech680_int, simp4391_0[8:8], comp2_0[26:26]);
  AO222EHD I626 (tech681_int, comp2_0[27:27], comp2_0[28:28], tech681_int, comp2_0[27:27], tech681_int, comp2_0[28:28]);
  AO222EHD I627 (simp4391_0[9:9], tech681_int, comp2_0[29:29], simp4391_0[9:9], tech681_int, simp4391_0[9:9], comp2_0[29:29]);
  AO222EHD I628 (simp4391_0[10:10], comp2_0[30:30], comp2_0[31:31], simp4391_0[10:10], comp2_0[30:30], simp4391_0[10:10], comp2_0[31:31]);
  AO222EHD I629 (tech684_int, simp4391_0[0:0], simp4391_0[1:1], tech684_int, simp4391_0[0:0], tech684_int, simp4391_0[1:1]);
  AO222EHD I630 (simp4392_0[0:0], tech684_int, simp4391_0[2:2], simp4392_0[0:0], tech684_int, simp4392_0[0:0], simp4391_0[2:2]);
  AO222EHD I631 (tech685_int, simp4391_0[3:3], simp4391_0[4:4], tech685_int, simp4391_0[3:3], tech685_int, simp4391_0[4:4]);
  AO222EHD I632 (simp4392_0[1:1], tech685_int, simp4391_0[5:5], simp4392_0[1:1], tech685_int, simp4392_0[1:1], simp4391_0[5:5]);
  AO222EHD I633 (tech686_int, simp4391_0[6:6], simp4391_0[7:7], tech686_int, simp4391_0[6:6], tech686_int, simp4391_0[7:7]);
  AO222EHD I634 (simp4392_0[2:2], tech686_int, simp4391_0[8:8], simp4392_0[2:2], tech686_int, simp4392_0[2:2], simp4391_0[8:8]);
  AO222EHD I635 (simp4392_0[3:3], simp4391_0[9:9], simp4391_0[10:10], simp4392_0[3:3], simp4391_0[9:9], simp4392_0[3:3], simp4391_0[10:10]);
  AO222EHD I636 (tech689_int, simp4392_0[0:0], simp4392_0[1:1], tech689_int, simp4392_0[0:0], tech689_int, simp4392_0[1:1]);
  AO222EHD I637 (simp4393_0[0:0], tech689_int, simp4392_0[2:2], simp4393_0[0:0], tech689_int, simp4393_0[0:0], simp4392_0[2:2]);
  BUFEHD I638 (simp4393_0[1:1], simp4392_0[3:3]);
  AO222EHD I639 (icomp_2, simp4393_0[0:0], simp4393_0[1:1], icomp_2, simp4393_0[0:0], icomp_2, simp4393_0[1:1]);
  OR2EHD I640 (comp3_0[0:0], i_3r0[0:0], i_3r1[0:0]);
  OR2EHD I641 (comp3_0[1:1], i_3r0[1:1], i_3r1[1:1]);
  OR2EHD I642 (comp3_0[2:2], i_3r0[2:2], i_3r1[2:2]);
  OR2EHD I643 (comp3_0[3:3], i_3r0[3:3], i_3r1[3:3]);
  OR2EHD I644 (comp3_0[4:4], i_3r0[4:4], i_3r1[4:4]);
  OR2EHD I645 (comp3_0[5:5], i_3r0[5:5], i_3r1[5:5]);
  OR2EHD I646 (comp3_0[6:6], i_3r0[6:6], i_3r1[6:6]);
  OR2EHD I647 (comp3_0[7:7], i_3r0[7:7], i_3r1[7:7]);
  OR2EHD I648 (comp3_0[8:8], i_3r0[8:8], i_3r1[8:8]);
  OR2EHD I649 (comp3_0[9:9], i_3r0[9:9], i_3r1[9:9]);
  OR2EHD I650 (comp3_0[10:10], i_3r0[10:10], i_3r1[10:10]);
  OR2EHD I651 (comp3_0[11:11], i_3r0[11:11], i_3r1[11:11]);
  OR2EHD I652 (comp3_0[12:12], i_3r0[12:12], i_3r1[12:12]);
  OR2EHD I653 (comp3_0[13:13], i_3r0[13:13], i_3r1[13:13]);
  OR2EHD I654 (comp3_0[14:14], i_3r0[14:14], i_3r1[14:14]);
  OR2EHD I655 (comp3_0[15:15], i_3r0[15:15], i_3r1[15:15]);
  OR2EHD I656 (comp3_0[16:16], i_3r0[16:16], i_3r1[16:16]);
  OR2EHD I657 (comp3_0[17:17], i_3r0[17:17], i_3r1[17:17]);
  OR2EHD I658 (comp3_0[18:18], i_3r0[18:18], i_3r1[18:18]);
  OR2EHD I659 (comp3_0[19:19], i_3r0[19:19], i_3r1[19:19]);
  OR2EHD I660 (comp3_0[20:20], i_3r0[20:20], i_3r1[20:20]);
  OR2EHD I661 (comp3_0[21:21], i_3r0[21:21], i_3r1[21:21]);
  OR2EHD I662 (comp3_0[22:22], i_3r0[22:22], i_3r1[22:22]);
  OR2EHD I663 (comp3_0[23:23], i_3r0[23:23], i_3r1[23:23]);
  OR2EHD I664 (comp3_0[24:24], i_3r0[24:24], i_3r1[24:24]);
  OR2EHD I665 (comp3_0[25:25], i_3r0[25:25], i_3r1[25:25]);
  OR2EHD I666 (comp3_0[26:26], i_3r0[26:26], i_3r1[26:26]);
  OR2EHD I667 (comp3_0[27:27], i_3r0[27:27], i_3r1[27:27]);
  OR2EHD I668 (comp3_0[28:28], i_3r0[28:28], i_3r1[28:28]);
  OR2EHD I669 (comp3_0[29:29], i_3r0[29:29], i_3r1[29:29]);
  OR2EHD I670 (comp3_0[30:30], i_3r0[30:30], i_3r1[30:30]);
  OR2EHD I671 (comp3_0[31:31], i_3r0[31:31], i_3r1[31:31]);
  AO222EHD I672 (tech726_int, comp3_0[0:0], comp3_0[1:1], tech726_int, comp3_0[0:0], tech726_int, comp3_0[1:1]);
  AO222EHD I673 (simp4731_0[0:0], tech726_int, comp3_0[2:2], simp4731_0[0:0], tech726_int, simp4731_0[0:0], comp3_0[2:2]);
  AO222EHD I674 (tech727_int, comp3_0[3:3], comp3_0[4:4], tech727_int, comp3_0[3:3], tech727_int, comp3_0[4:4]);
  AO222EHD I675 (simp4731_0[1:1], tech727_int, comp3_0[5:5], simp4731_0[1:1], tech727_int, simp4731_0[1:1], comp3_0[5:5]);
  AO222EHD I676 (tech728_int, comp3_0[6:6], comp3_0[7:7], tech728_int, comp3_0[6:6], tech728_int, comp3_0[7:7]);
  AO222EHD I677 (simp4731_0[2:2], tech728_int, comp3_0[8:8], simp4731_0[2:2], tech728_int, simp4731_0[2:2], comp3_0[8:8]);
  AO222EHD I678 (tech729_int, comp3_0[9:9], comp3_0[10:10], tech729_int, comp3_0[9:9], tech729_int, comp3_0[10:10]);
  AO222EHD I679 (simp4731_0[3:3], tech729_int, comp3_0[11:11], simp4731_0[3:3], tech729_int, simp4731_0[3:3], comp3_0[11:11]);
  AO222EHD I680 (tech730_int, comp3_0[12:12], comp3_0[13:13], tech730_int, comp3_0[12:12], tech730_int, comp3_0[13:13]);
  AO222EHD I681 (simp4731_0[4:4], tech730_int, comp3_0[14:14], simp4731_0[4:4], tech730_int, simp4731_0[4:4], comp3_0[14:14]);
  AO222EHD I682 (tech731_int, comp3_0[15:15], comp3_0[16:16], tech731_int, comp3_0[15:15], tech731_int, comp3_0[16:16]);
  AO222EHD I683 (simp4731_0[5:5], tech731_int, comp3_0[17:17], simp4731_0[5:5], tech731_int, simp4731_0[5:5], comp3_0[17:17]);
  AO222EHD I684 (tech732_int, comp3_0[18:18], comp3_0[19:19], tech732_int, comp3_0[18:18], tech732_int, comp3_0[19:19]);
  AO222EHD I685 (simp4731_0[6:6], tech732_int, comp3_0[20:20], simp4731_0[6:6], tech732_int, simp4731_0[6:6], comp3_0[20:20]);
  AO222EHD I686 (tech733_int, comp3_0[21:21], comp3_0[22:22], tech733_int, comp3_0[21:21], tech733_int, comp3_0[22:22]);
  AO222EHD I687 (simp4731_0[7:7], tech733_int, comp3_0[23:23], simp4731_0[7:7], tech733_int, simp4731_0[7:7], comp3_0[23:23]);
  AO222EHD I688 (tech734_int, comp3_0[24:24], comp3_0[25:25], tech734_int, comp3_0[24:24], tech734_int, comp3_0[25:25]);
  AO222EHD I689 (simp4731_0[8:8], tech734_int, comp3_0[26:26], simp4731_0[8:8], tech734_int, simp4731_0[8:8], comp3_0[26:26]);
  AO222EHD I690 (tech735_int, comp3_0[27:27], comp3_0[28:28], tech735_int, comp3_0[27:27], tech735_int, comp3_0[28:28]);
  AO222EHD I691 (simp4731_0[9:9], tech735_int, comp3_0[29:29], simp4731_0[9:9], tech735_int, simp4731_0[9:9], comp3_0[29:29]);
  AO222EHD I692 (simp4731_0[10:10], comp3_0[30:30], comp3_0[31:31], simp4731_0[10:10], comp3_0[30:30], simp4731_0[10:10], comp3_0[31:31]);
  AO222EHD I693 (tech738_int, simp4731_0[0:0], simp4731_0[1:1], tech738_int, simp4731_0[0:0], tech738_int, simp4731_0[1:1]);
  AO222EHD I694 (simp4732_0[0:0], tech738_int, simp4731_0[2:2], simp4732_0[0:0], tech738_int, simp4732_0[0:0], simp4731_0[2:2]);
  AO222EHD I695 (tech739_int, simp4731_0[3:3], simp4731_0[4:4], tech739_int, simp4731_0[3:3], tech739_int, simp4731_0[4:4]);
  AO222EHD I696 (simp4732_0[1:1], tech739_int, simp4731_0[5:5], simp4732_0[1:1], tech739_int, simp4732_0[1:1], simp4731_0[5:5]);
  AO222EHD I697 (tech740_int, simp4731_0[6:6], simp4731_0[7:7], tech740_int, simp4731_0[6:6], tech740_int, simp4731_0[7:7]);
  AO222EHD I698 (simp4732_0[2:2], tech740_int, simp4731_0[8:8], simp4732_0[2:2], tech740_int, simp4732_0[2:2], simp4731_0[8:8]);
  AO222EHD I699 (simp4732_0[3:3], simp4731_0[9:9], simp4731_0[10:10], simp4732_0[3:3], simp4731_0[9:9], simp4732_0[3:3], simp4731_0[10:10]);
  AO222EHD I700 (tech743_int, simp4732_0[0:0], simp4732_0[1:1], tech743_int, simp4732_0[0:0], tech743_int, simp4732_0[1:1]);
  AO222EHD I701 (simp4733_0[0:0], tech743_int, simp4732_0[2:2], simp4733_0[0:0], tech743_int, simp4733_0[0:0], simp4732_0[2:2]);
  BUFEHD I702 (simp4733_0[1:1], simp4732_0[3:3]);
  AO222EHD I703 (icomp_3, simp4733_0[0:0], simp4733_0[1:1], icomp_3, simp4733_0[0:0], icomp_3, simp4733_0[1:1]);
  AO222EHD I704 (choice_0, icomp_0, nchosen_0, tech746_oint, icomp_0, tech746_oint, nchosen_0);
  AN2B1CHD I705 (tech746_oint, choice_0, reset);
  AO222EHD I706 (choice_1, icomp_1, nchosen_0, tech747_oint, icomp_1, tech747_oint, nchosen_0);
  AN2B1CHD I707 (tech747_oint, choice_1, reset);
  AO222EHD I708 (choice_2, icomp_2, nchosen_0, tech748_oint, icomp_2, tech748_oint, nchosen_0);
  AN2B1CHD I709 (tech748_oint, choice_2, reset);
  AO222EHD I710 (choice_3, icomp_3, nchosen_0, tech749_oint, icomp_3, tech749_oint, nchosen_0);
  AN2B1CHD I711 (tech749_oint, choice_3, reset);
  NR3EHD I712 (simp4781_0[0:0], choice_0, choice_1, choice_2);
  INVHHD I713 (simp4781_0[1:1], choice_3);
  ND2HHD I714 (anychoice_0, simp4781_0[0:0], simp4781_0[1:1]);
  NR2EHD I715 (nchosen_0, anychoice_0, o_0a);
  AO222EHD I716 (i_0a, choice_0, o_0a, tech755_oint, choice_0, tech755_oint, o_0a);
  AN2B1CHD I717 (tech755_oint, i_0a, reset);
  AO222EHD I718 (i_1a, choice_1, o_0a, tech756_oint, choice_1, tech756_oint, o_0a);
  AN2B1CHD I719 (tech756_oint, i_1a, reset);
  AO222EHD I720 (i_2a, choice_2, o_0a, tech757_oint, choice_2, tech757_oint, o_0a);
  AN2B1CHD I721 (tech757_oint, i_2a, reset);
  AO222EHD I722 (i_3a, choice_3, o_0a, tech758_oint, choice_3, tech758_oint, o_0a);
  AN2B1CHD I723 (tech758_oint, i_3a, reset);
endmodule

// tkj32m32_0 TeakJ [Many [32,0],One 32]
module tkj32m32_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [31:0] joinf_0;
  wire [31:0] joint_0;
  BUFEHD I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFEHD I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFEHD I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFEHD I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFEHD I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFEHD I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFEHD I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFEHD I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFEHD I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFEHD I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFEHD I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFEHD I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFEHD I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFEHD I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFEHD I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFEHD I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFEHD I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFEHD I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFEHD I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFEHD I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFEHD I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFEHD I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFEHD I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFEHD I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFEHD I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFEHD I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFEHD I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFEHD I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFEHD I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFEHD I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFEHD I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFEHD I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFEHD I32 (joint_0[0:0], i_0r1[0:0]);
  BUFEHD I33 (joint_0[1:1], i_0r1[1:1]);
  BUFEHD I34 (joint_0[2:2], i_0r1[2:2]);
  BUFEHD I35 (joint_0[3:3], i_0r1[3:3]);
  BUFEHD I36 (joint_0[4:4], i_0r1[4:4]);
  BUFEHD I37 (joint_0[5:5], i_0r1[5:5]);
  BUFEHD I38 (joint_0[6:6], i_0r1[6:6]);
  BUFEHD I39 (joint_0[7:7], i_0r1[7:7]);
  BUFEHD I40 (joint_0[8:8], i_0r1[8:8]);
  BUFEHD I41 (joint_0[9:9], i_0r1[9:9]);
  BUFEHD I42 (joint_0[10:10], i_0r1[10:10]);
  BUFEHD I43 (joint_0[11:11], i_0r1[11:11]);
  BUFEHD I44 (joint_0[12:12], i_0r1[12:12]);
  BUFEHD I45 (joint_0[13:13], i_0r1[13:13]);
  BUFEHD I46 (joint_0[14:14], i_0r1[14:14]);
  BUFEHD I47 (joint_0[15:15], i_0r1[15:15]);
  BUFEHD I48 (joint_0[16:16], i_0r1[16:16]);
  BUFEHD I49 (joint_0[17:17], i_0r1[17:17]);
  BUFEHD I50 (joint_0[18:18], i_0r1[18:18]);
  BUFEHD I51 (joint_0[19:19], i_0r1[19:19]);
  BUFEHD I52 (joint_0[20:20], i_0r1[20:20]);
  BUFEHD I53 (joint_0[21:21], i_0r1[21:21]);
  BUFEHD I54 (joint_0[22:22], i_0r1[22:22]);
  BUFEHD I55 (joint_0[23:23], i_0r1[23:23]);
  BUFEHD I56 (joint_0[24:24], i_0r1[24:24]);
  BUFEHD I57 (joint_0[25:25], i_0r1[25:25]);
  BUFEHD I58 (joint_0[26:26], i_0r1[26:26]);
  BUFEHD I59 (joint_0[27:27], i_0r1[27:27]);
  BUFEHD I60 (joint_0[28:28], i_0r1[28:28]);
  BUFEHD I61 (joint_0[29:29], i_0r1[29:29]);
  BUFEHD I62 (joint_0[30:30], i_0r1[30:30]);
  BUFEHD I63 (joint_0[31:31], i_0r1[31:31]);
  BUFEHD I64 (icomplete_0, i_1r);
  AO222EHD I65 (o_0r0[0:0], joinf_0[0:0], icomplete_0, o_0r0[0:0], joinf_0[0:0], o_0r0[0:0], icomplete_0);
  AO222EHD I66 (o_0r1[0:0], joint_0[0:0], icomplete_0, o_0r1[0:0], joint_0[0:0], o_0r1[0:0], icomplete_0);
  BUFEHD I67 (o_0r0[1:1], joinf_0[1:1]);
  BUFEHD I68 (o_0r0[2:2], joinf_0[2:2]);
  BUFEHD I69 (o_0r0[3:3], joinf_0[3:3]);
  BUFEHD I70 (o_0r0[4:4], joinf_0[4:4]);
  BUFEHD I71 (o_0r0[5:5], joinf_0[5:5]);
  BUFEHD I72 (o_0r0[6:6], joinf_0[6:6]);
  BUFEHD I73 (o_0r0[7:7], joinf_0[7:7]);
  BUFEHD I74 (o_0r0[8:8], joinf_0[8:8]);
  BUFEHD I75 (o_0r0[9:9], joinf_0[9:9]);
  BUFEHD I76 (o_0r0[10:10], joinf_0[10:10]);
  BUFEHD I77 (o_0r0[11:11], joinf_0[11:11]);
  BUFEHD I78 (o_0r0[12:12], joinf_0[12:12]);
  BUFEHD I79 (o_0r0[13:13], joinf_0[13:13]);
  BUFEHD I80 (o_0r0[14:14], joinf_0[14:14]);
  BUFEHD I81 (o_0r0[15:15], joinf_0[15:15]);
  BUFEHD I82 (o_0r0[16:16], joinf_0[16:16]);
  BUFEHD I83 (o_0r0[17:17], joinf_0[17:17]);
  BUFEHD I84 (o_0r0[18:18], joinf_0[18:18]);
  BUFEHD I85 (o_0r0[19:19], joinf_0[19:19]);
  BUFEHD I86 (o_0r0[20:20], joinf_0[20:20]);
  BUFEHD I87 (o_0r0[21:21], joinf_0[21:21]);
  BUFEHD I88 (o_0r0[22:22], joinf_0[22:22]);
  BUFEHD I89 (o_0r0[23:23], joinf_0[23:23]);
  BUFEHD I90 (o_0r0[24:24], joinf_0[24:24]);
  BUFEHD I91 (o_0r0[25:25], joinf_0[25:25]);
  BUFEHD I92 (o_0r0[26:26], joinf_0[26:26]);
  BUFEHD I93 (o_0r0[27:27], joinf_0[27:27]);
  BUFEHD I94 (o_0r0[28:28], joinf_0[28:28]);
  BUFEHD I95 (o_0r0[29:29], joinf_0[29:29]);
  BUFEHD I96 (o_0r0[30:30], joinf_0[30:30]);
  BUFEHD I97 (o_0r0[31:31], joinf_0[31:31]);
  BUFEHD I98 (o_0r1[1:1], joint_0[1:1]);
  BUFEHD I99 (o_0r1[2:2], joint_0[2:2]);
  BUFEHD I100 (o_0r1[3:3], joint_0[3:3]);
  BUFEHD I101 (o_0r1[4:4], joint_0[4:4]);
  BUFEHD I102 (o_0r1[5:5], joint_0[5:5]);
  BUFEHD I103 (o_0r1[6:6], joint_0[6:6]);
  BUFEHD I104 (o_0r1[7:7], joint_0[7:7]);
  BUFEHD I105 (o_0r1[8:8], joint_0[8:8]);
  BUFEHD I106 (o_0r1[9:9], joint_0[9:9]);
  BUFEHD I107 (o_0r1[10:10], joint_0[10:10]);
  BUFEHD I108 (o_0r1[11:11], joint_0[11:11]);
  BUFEHD I109 (o_0r1[12:12], joint_0[12:12]);
  BUFEHD I110 (o_0r1[13:13], joint_0[13:13]);
  BUFEHD I111 (o_0r1[14:14], joint_0[14:14]);
  BUFEHD I112 (o_0r1[15:15], joint_0[15:15]);
  BUFEHD I113 (o_0r1[16:16], joint_0[16:16]);
  BUFEHD I114 (o_0r1[17:17], joint_0[17:17]);
  BUFEHD I115 (o_0r1[18:18], joint_0[18:18]);
  BUFEHD I116 (o_0r1[19:19], joint_0[19:19]);
  BUFEHD I117 (o_0r1[20:20], joint_0[20:20]);
  BUFEHD I118 (o_0r1[21:21], joint_0[21:21]);
  BUFEHD I119 (o_0r1[22:22], joint_0[22:22]);
  BUFEHD I120 (o_0r1[23:23], joint_0[23:23]);
  BUFEHD I121 (o_0r1[24:24], joint_0[24:24]);
  BUFEHD I122 (o_0r1[25:25], joint_0[25:25]);
  BUFEHD I123 (o_0r1[26:26], joint_0[26:26]);
  BUFEHD I124 (o_0r1[27:27], joint_0[27:27]);
  BUFEHD I125 (o_0r1[28:28], joint_0[28:28]);
  BUFEHD I126 (o_0r1[29:29], joint_0[29:29]);
  BUFEHD I127 (o_0r1[30:30], joint_0[30:30]);
  BUFEHD I128 (o_0r1[31:31], joint_0[31:31]);
  BUFEHD I129 (i_0a, o_0a);
  BUFEHD I130 (i_1a, o_0a);
endmodule

// tkf32mo0w0_o0w32 TeakF [0,0] [One 32,Many [0,32]]
module tkf32mo0w0_o0w32 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [31:0] o_1r0;
  output [31:0] o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  wire tech69_int;
  OR2EHD I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFEHD I1 (acomplete_0, icomplete_0);
  BUFEHD I2 (o_1r0[0:0], i_0r0[0:0]);
  BUFEHD I3 (o_1r0[1:1], i_0r0[1:1]);
  BUFEHD I4 (o_1r0[2:2], i_0r0[2:2]);
  BUFEHD I5 (o_1r0[3:3], i_0r0[3:3]);
  BUFEHD I6 (o_1r0[4:4], i_0r0[4:4]);
  BUFEHD I7 (o_1r0[5:5], i_0r0[5:5]);
  BUFEHD I8 (o_1r0[6:6], i_0r0[6:6]);
  BUFEHD I9 (o_1r0[7:7], i_0r0[7:7]);
  BUFEHD I10 (o_1r0[8:8], i_0r0[8:8]);
  BUFEHD I11 (o_1r0[9:9], i_0r0[9:9]);
  BUFEHD I12 (o_1r0[10:10], i_0r0[10:10]);
  BUFEHD I13 (o_1r0[11:11], i_0r0[11:11]);
  BUFEHD I14 (o_1r0[12:12], i_0r0[12:12]);
  BUFEHD I15 (o_1r0[13:13], i_0r0[13:13]);
  BUFEHD I16 (o_1r0[14:14], i_0r0[14:14]);
  BUFEHD I17 (o_1r0[15:15], i_0r0[15:15]);
  BUFEHD I18 (o_1r0[16:16], i_0r0[16:16]);
  BUFEHD I19 (o_1r0[17:17], i_0r0[17:17]);
  BUFEHD I20 (o_1r0[18:18], i_0r0[18:18]);
  BUFEHD I21 (o_1r0[19:19], i_0r0[19:19]);
  BUFEHD I22 (o_1r0[20:20], i_0r0[20:20]);
  BUFEHD I23 (o_1r0[21:21], i_0r0[21:21]);
  BUFEHD I24 (o_1r0[22:22], i_0r0[22:22]);
  BUFEHD I25 (o_1r0[23:23], i_0r0[23:23]);
  BUFEHD I26 (o_1r0[24:24], i_0r0[24:24]);
  BUFEHD I27 (o_1r0[25:25], i_0r0[25:25]);
  BUFEHD I28 (o_1r0[26:26], i_0r0[26:26]);
  BUFEHD I29 (o_1r0[27:27], i_0r0[27:27]);
  BUFEHD I30 (o_1r0[28:28], i_0r0[28:28]);
  BUFEHD I31 (o_1r0[29:29], i_0r0[29:29]);
  BUFEHD I32 (o_1r0[30:30], i_0r0[30:30]);
  BUFEHD I33 (o_1r0[31:31], i_0r0[31:31]);
  BUFEHD I34 (o_1r1[0:0], i_0r1[0:0]);
  BUFEHD I35 (o_1r1[1:1], i_0r1[1:1]);
  BUFEHD I36 (o_1r1[2:2], i_0r1[2:2]);
  BUFEHD I37 (o_1r1[3:3], i_0r1[3:3]);
  BUFEHD I38 (o_1r1[4:4], i_0r1[4:4]);
  BUFEHD I39 (o_1r1[5:5], i_0r1[5:5]);
  BUFEHD I40 (o_1r1[6:6], i_0r1[6:6]);
  BUFEHD I41 (o_1r1[7:7], i_0r1[7:7]);
  BUFEHD I42 (o_1r1[8:8], i_0r1[8:8]);
  BUFEHD I43 (o_1r1[9:9], i_0r1[9:9]);
  BUFEHD I44 (o_1r1[10:10], i_0r1[10:10]);
  BUFEHD I45 (o_1r1[11:11], i_0r1[11:11]);
  BUFEHD I46 (o_1r1[12:12], i_0r1[12:12]);
  BUFEHD I47 (o_1r1[13:13], i_0r1[13:13]);
  BUFEHD I48 (o_1r1[14:14], i_0r1[14:14]);
  BUFEHD I49 (o_1r1[15:15], i_0r1[15:15]);
  BUFEHD I50 (o_1r1[16:16], i_0r1[16:16]);
  BUFEHD I51 (o_1r1[17:17], i_0r1[17:17]);
  BUFEHD I52 (o_1r1[18:18], i_0r1[18:18]);
  BUFEHD I53 (o_1r1[19:19], i_0r1[19:19]);
  BUFEHD I54 (o_1r1[20:20], i_0r1[20:20]);
  BUFEHD I55 (o_1r1[21:21], i_0r1[21:21]);
  BUFEHD I56 (o_1r1[22:22], i_0r1[22:22]);
  BUFEHD I57 (o_1r1[23:23], i_0r1[23:23]);
  BUFEHD I58 (o_1r1[24:24], i_0r1[24:24]);
  BUFEHD I59 (o_1r1[25:25], i_0r1[25:25]);
  BUFEHD I60 (o_1r1[26:26], i_0r1[26:26]);
  BUFEHD I61 (o_1r1[27:27], i_0r1[27:27]);
  BUFEHD I62 (o_1r1[28:28], i_0r1[28:28]);
  BUFEHD I63 (o_1r1[29:29], i_0r1[29:29]);
  BUFEHD I64 (o_1r1[30:30], i_0r1[30:30]);
  BUFEHD I65 (o_1r1[31:31], i_0r1[31:31]);
  BUFEHD I66 (o_0r, icomplete_0);
  AO222EHD I67 (tech69_int, acomplete_0, o_0a, tech69_int, acomplete_0, tech69_int, o_0a);
  AO222EHD I68 (i_0a, tech69_int, o_1a, i_0a, tech69_int, i_0a, o_1a);
endmodule

// tkj7m5_2_0 TeakJ [Many [5,2,0],One 7]
module tkj7m5_2_0 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r, i_2a, o_0r0, o_0r1, o_0a, reset);
  input [4:0] i_0r0;
  input [4:0] i_0r1;
  output i_0a;
  input [1:0] i_1r0;
  input [1:0] i_1r1;
  output i_1a;
  input i_2r;
  output i_2a;
  output [6:0] o_0r0;
  output [6:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [6:0] joinf_0;
  wire [6:0] joint_0;
  wire dcomplete_0;
  BUFEHD I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFEHD I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFEHD I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFEHD I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFEHD I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFEHD I5 (joinf_0[5:5], i_1r0[0:0]);
  BUFEHD I6 (joinf_0[6:6], i_1r0[1:1]);
  BUFEHD I7 (joint_0[0:0], i_0r1[0:0]);
  BUFEHD I8 (joint_0[1:1], i_0r1[1:1]);
  BUFEHD I9 (joint_0[2:2], i_0r1[2:2]);
  BUFEHD I10 (joint_0[3:3], i_0r1[3:3]);
  BUFEHD I11 (joint_0[4:4], i_0r1[4:4]);
  BUFEHD I12 (joint_0[5:5], i_1r1[0:0]);
  BUFEHD I13 (joint_0[6:6], i_1r1[1:1]);
  OR2EHD I14 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  AO222EHD I15 (icomplete_0, i_2r, dcomplete_0, icomplete_0, i_2r, icomplete_0, dcomplete_0);
  AO222EHD I16 (o_0r0[0:0], joinf_0[0:0], icomplete_0, o_0r0[0:0], joinf_0[0:0], o_0r0[0:0], icomplete_0);
  AO222EHD I17 (o_0r1[0:0], joint_0[0:0], icomplete_0, o_0r1[0:0], joint_0[0:0], o_0r1[0:0], icomplete_0);
  BUFEHD I18 (o_0r0[1:1], joinf_0[1:1]);
  BUFEHD I19 (o_0r0[2:2], joinf_0[2:2]);
  BUFEHD I20 (o_0r0[3:3], joinf_0[3:3]);
  BUFEHD I21 (o_0r0[4:4], joinf_0[4:4]);
  BUFEHD I22 (o_0r0[5:5], joinf_0[5:5]);
  BUFEHD I23 (o_0r0[6:6], joinf_0[6:6]);
  BUFEHD I24 (o_0r1[1:1], joint_0[1:1]);
  BUFEHD I25 (o_0r1[2:2], joint_0[2:2]);
  BUFEHD I26 (o_0r1[3:3], joint_0[3:3]);
  BUFEHD I27 (o_0r1[4:4], joint_0[4:4]);
  BUFEHD I28 (o_0r1[5:5], joint_0[5:5]);
  BUFEHD I29 (o_0r1[6:6], joint_0[6:6]);
  BUFEHD I30 (i_0a, o_0a);
  BUFEHD I31 (i_1a, o_0a);
  BUFEHD I32 (i_2a, o_0a);
endmodule

// tkvdistanceIshift7_wo0w7_ro5w2o5w2 TeakV "distanceI-shift" 7 [] [0] [5,5] [Many [7],Many [0],Many [0
//   ,0],Many [2,2]]
module tkvdistanceIshift7_wo0w7_ro5w2o5w2 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, reset);
  input [6:0] wg_0r0;
  input [6:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [1:0] rd_0r0;
  output [1:0] rd_0r1;
  input rd_0a;
  output [1:0] rd_1r0;
  output [1:0] rd_1r1;
  input rd_1a;
  input reset;
  wire [6:0] wf_0;
  wire [6:0] wt_0;
  wire [6:0] df_0;
  wire [6:0] dt_0;
  wire wc_0;
  wire [6:0] wacks_0;
  wire [6:0] wenr_0;
  wire [6:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [6:0] drlgf_0;
  wire [6:0] drlgt_0;
  wire [6:0] comp0_0;
  wire [2:0] simp631_0;
  wire tech64_int;
  wire tech65_int;
  wire tech67_int;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [6:0] conwgit_0;
  wire [6:0] conwgif_0;
  wire conwig_0;
  wire [2:0] simp1071_0;
  wire tech112_int;
  wire tech113_int;
  wire tech115_int;
  wire [1:0] simp1161_0;
  INVHHD I0 (nreset_0, reset);
  AN2EHD I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AN2EHD I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AN2EHD I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AN2EHD I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AN2EHD I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AN2EHD I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AN2EHD I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AN2EHD I8 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AN2EHD I9 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AN2EHD I10 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AN2EHD I11 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AN2EHD I12 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AN2EHD I13 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AN2EHD I14 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AN2EHD I15 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AN2EHD I16 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AN2EHD I17 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AN2EHD I18 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AN2EHD I19 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AN2EHD I20 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AN2EHD I21 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  NR2EHD I22 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NR2EHD I23 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NR2EHD I24 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NR2EHD I25 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NR2EHD I26 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NR2EHD I27 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NR2EHD I28 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NR3EHD I29 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NR3EHD I30 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NR3EHD I31 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NR3EHD I32 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NR3EHD I33 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NR3EHD I34 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NR3EHD I35 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  AO22EHD I36 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22EHD I37 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22EHD I38 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22EHD I39 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22EHD I40 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22EHD I41 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22EHD I42 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  OR2EHD I43 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2EHD I44 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2EHD I45 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2EHD I46 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2EHD I47 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2EHD I48 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2EHD I49 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  AO222EHD I50 (tech64_int, comp0_0[0:0], comp0_0[1:1], tech64_int, comp0_0[0:0], tech64_int, comp0_0[1:1]);
  AO222EHD I51 (simp631_0[0:0], tech64_int, comp0_0[2:2], simp631_0[0:0], tech64_int, simp631_0[0:0], comp0_0[2:2]);
  AO222EHD I52 (tech65_int, comp0_0[3:3], comp0_0[4:4], tech65_int, comp0_0[3:3], tech65_int, comp0_0[4:4]);
  AO222EHD I53 (simp631_0[1:1], tech65_int, comp0_0[5:5], simp631_0[1:1], tech65_int, simp631_0[1:1], comp0_0[5:5]);
  BUFEHD I54 (simp631_0[2:2], comp0_0[6:6]);
  AO222EHD I55 (tech67_int, simp631_0[0:0], simp631_0[1:1], tech67_int, simp631_0[0:0], tech67_int, simp631_0[1:1]);
  AO222EHD I56 (wc_0, tech67_int, simp631_0[2:2], wc_0, tech67_int, wc_0, simp631_0[2:2]);
  AN2EHD I57 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AN2EHD I58 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AN2EHD I59 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AN2EHD I60 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AN2EHD I61 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AN2EHD I62 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AN2EHD I63 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AN2EHD I64 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AN2EHD I65 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AN2EHD I66 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AN2EHD I67 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AN2EHD I68 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AN2EHD I69 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AN2EHD I70 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  BUFEHD I71 (conwigc_0, wc_0);
  AO12EHD I72 (conwig_0, conwigc_0, conwigc_0, conwigcanw_0);
  NR2EHD I73 (conwigcanw_0, anyread_0, conwig_0);
  BUFEHD I74 (wf_0[0:0], conwgif_0[0:0]);
  BUFEHD I75 (wt_0[0:0], conwgit_0[0:0]);
  BUFEHD I76 (wenr_0[0:0], wc_0);
  BUFEHD I77 (wf_0[1:1], conwgif_0[1:1]);
  BUFEHD I78 (wt_0[1:1], conwgit_0[1:1]);
  BUFEHD I79 (wenr_0[1:1], wc_0);
  BUFEHD I80 (wf_0[2:2], conwgif_0[2:2]);
  BUFEHD I81 (wt_0[2:2], conwgit_0[2:2]);
  BUFEHD I82 (wenr_0[2:2], wc_0);
  BUFEHD I83 (wf_0[3:3], conwgif_0[3:3]);
  BUFEHD I84 (wt_0[3:3], conwgit_0[3:3]);
  BUFEHD I85 (wenr_0[3:3], wc_0);
  BUFEHD I86 (wf_0[4:4], conwgif_0[4:4]);
  BUFEHD I87 (wt_0[4:4], conwgit_0[4:4]);
  BUFEHD I88 (wenr_0[4:4], wc_0);
  BUFEHD I89 (wf_0[5:5], conwgif_0[5:5]);
  BUFEHD I90 (wt_0[5:5], conwgit_0[5:5]);
  BUFEHD I91 (wenr_0[5:5], wc_0);
  BUFEHD I92 (wf_0[6:6], conwgif_0[6:6]);
  BUFEHD I93 (wt_0[6:6], conwgit_0[6:6]);
  BUFEHD I94 (wenr_0[6:6], wc_0);
  AO222EHD I95 (tech112_int, conwig_0, wacks_0[0:0], tech112_int, conwig_0, tech112_int, wacks_0[0:0]);
  AO222EHD I96 (simp1071_0[0:0], tech112_int, wacks_0[1:1], simp1071_0[0:0], tech112_int, simp1071_0[0:0], wacks_0[1:1]);
  AO222EHD I97 (tech113_int, wacks_0[2:2], wacks_0[3:3], tech113_int, wacks_0[2:2], tech113_int, wacks_0[3:3]);
  AO222EHD I98 (simp1071_0[1:1], tech113_int, wacks_0[4:4], simp1071_0[1:1], tech113_int, simp1071_0[1:1], wacks_0[4:4]);
  AO222EHD I99 (simp1071_0[2:2], wacks_0[5:5], wacks_0[6:6], simp1071_0[2:2], wacks_0[5:5], simp1071_0[2:2], wacks_0[6:6]);
  AO222EHD I100 (tech115_int, simp1071_0[0:0], simp1071_0[1:1], tech115_int, simp1071_0[0:0], tech115_int, simp1071_0[1:1]);
  AO222EHD I101 (wd_0r, tech115_int, simp1071_0[2:2], wd_0r, tech115_int, wd_0r, simp1071_0[2:2]);
  AN2EHD I102 (rd_0r0[0:0], df_0[5:5], rg_0r);
  AN2EHD I103 (rd_0r0[1:1], df_0[6:6], rg_0r);
  AN2EHD I104 (rd_1r0[0:0], df_0[5:5], rg_1r);
  AN2EHD I105 (rd_1r0[1:1], df_0[6:6], rg_1r);
  AN2EHD I106 (rd_0r1[0:0], dt_0[5:5], rg_0r);
  AN2EHD I107 (rd_0r1[1:1], dt_0[6:6], rg_0r);
  AN2EHD I108 (rd_1r1[0:0], dt_0[5:5], rg_1r);
  AN2EHD I109 (rd_1r1[1:1], dt_0[6:6], rg_1r);
  NR3EHD I110 (simp1161_0[0:0], rg_0r, rg_1r, rg_0a);
  INVHHD I111 (simp1161_0[1:1], rg_1a);
  ND2HHD I112 (anyread_0, simp1161_0[0:0], simp1161_0[1:1]);
  BUFEHD I113 (wg_0a, wd_0a);
  BUFEHD I114 (rg_0a, rd_0a);
  BUFEHD I115 (rg_1a, rd_1a);
endmodule

// tkf7mo0w7_o2w1_o1w1 TeakF [0,2,1] [One 7,Many [7,1,1]]
module tkf7mo0w7_o2w1_o1w1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r0, o_1r1, o_1a, o_2r0, o_2r1, o_2a, reset);
  input [6:0] i_0r0;
  input [6:0] i_0r1;
  output i_0a;
  output [6:0] o_0r0;
  output [6:0] o_0r1;
  input o_0a;
  output o_1r0;
  output o_1r1;
  input o_1a;
  output o_2r0;
  output o_2r1;
  input o_2a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  wire [1:0] simp231_0;
  wire tech23_int;
  OR2EHD I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFEHD I1 (acomplete_0, icomplete_0);
  BUFEHD I2 (o_0r0[0:0], i_0r0[0:0]);
  BUFEHD I3 (o_0r0[1:1], i_0r0[1:1]);
  BUFEHD I4 (o_0r0[2:2], i_0r0[2:2]);
  BUFEHD I5 (o_0r0[3:3], i_0r0[3:3]);
  BUFEHD I6 (o_0r0[4:4], i_0r0[4:4]);
  BUFEHD I7 (o_0r0[5:5], i_0r0[5:5]);
  BUFEHD I8 (o_0r0[6:6], i_0r0[6:6]);
  AO222EHD I9 (o_1r0, i_0r0[2:2], icomplete_0, o_1r0, i_0r0[2:2], o_1r0, icomplete_0);
  AO222EHD I10 (o_2r0, i_0r0[1:1], icomplete_0, o_2r0, i_0r0[1:1], o_2r0, icomplete_0);
  BUFEHD I11 (o_0r1[0:0], i_0r1[0:0]);
  BUFEHD I12 (o_0r1[1:1], i_0r1[1:1]);
  BUFEHD I13 (o_0r1[2:2], i_0r1[2:2]);
  BUFEHD I14 (o_0r1[3:3], i_0r1[3:3]);
  BUFEHD I15 (o_0r1[4:4], i_0r1[4:4]);
  BUFEHD I16 (o_0r1[5:5], i_0r1[5:5]);
  BUFEHD I17 (o_0r1[6:6], i_0r1[6:6]);
  AO222EHD I18 (o_1r1, i_0r1[2:2], icomplete_0, o_1r1, i_0r1[2:2], o_1r1, icomplete_0);
  AO222EHD I19 (o_2r1, i_0r1[1:1], icomplete_0, o_2r1, i_0r1[1:1], o_2r1, icomplete_0);
  AO222EHD I20 (tech23_int, acomplete_0, o_0a, tech23_int, acomplete_0, tech23_int, o_0a);
  AO222EHD I21 (simp231_0[0:0], tech23_int, o_1a, simp231_0[0:0], tech23_int, simp231_0[0:0], o_1a);
  BUFEHD I22 (simp231_0[1:1], o_2a);
  AO222EHD I23 (i_0a, simp231_0[0:0], simp231_0[1:1], i_0a, simp231_0[0:0], i_0a, simp231_0[1:1]);
endmodule

// tkj1m1_0 TeakJ [Many [1,0],One 1]
module tkj1m1_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire joinf_0;
  wire joint_0;
  BUFEHD I0 (joinf_0, i_0r0);
  BUFEHD I1 (joint_0, i_0r1);
  BUFEHD I2 (icomplete_0, i_1r);
  AO222EHD I3 (o_0r0, joinf_0, icomplete_0, o_0r0, joinf_0, o_0r0, icomplete_0);
  AO222EHD I4 (o_0r1, joint_0, icomplete_0, o_0r1, joint_0, o_0r1, icomplete_0);
  BUFEHD I5 (i_0a, o_0a);
  BUFEHD I6 (i_1a, o_0a);
endmodule

// tkf0mo0w0_o0w0 TeakF [0,0] [One 0,Many [0,0]]
module tkf0mo0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  BUFEHD I0 (o_0r, i_0r);
  BUFEHD I1 (o_1r, i_0r);
  AO222EHD I2 (i_0a, o_0a, o_1a, i_0a, o_0a, i_0a, o_1a);
endmodule

// tks2_o0w2_3o0w0_0c2o0w0_1o0w0 TeakS (0+:2) [([Imp 3 0],0),([Imp 0 2],0),([Imp 1 0],0)] [One 2,Many [
//   0,0,0]]
module tks2_o0w2_3o0w0_0c2o0w0_1o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire match2_0;
  wire [1:0] comp_0;
  BUFEHD I0 (sel_0, match0_0);
  AO222EHD I1 (match0_0, i_0r1[0:0], i_0r1[1:1], match0_0, i_0r1[0:0], match0_0, i_0r1[1:1]);
  BUFEHD I2 (sel_1, match1_0);
  BUFEHD I3 (match1_0, i_0r0[0:0]);
  BUFEHD I4 (sel_2, match2_0);
  AO222EHD I5 (match2_0, i_0r1[0:0], i_0r0[1:1], match2_0, i_0r1[0:0], match2_0, i_0r0[1:1]);
  AO222EHD I6 (gsel_0, sel_0, icomplete_0, gsel_0, sel_0, gsel_0, icomplete_0);
  AO222EHD I7 (gsel_1, sel_1, icomplete_0, gsel_1, sel_1, gsel_1, icomplete_0);
  AO222EHD I8 (gsel_2, sel_2, icomplete_0, gsel_2, sel_2, gsel_2, icomplete_0);
  OR2EHD I9 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2EHD I10 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  AO222EHD I11 (icomplete_0, comp_0[0:0], comp_0[1:1], icomplete_0, comp_0[0:0], icomplete_0, comp_0[1:1]);
  BUFEHD I12 (o_0r, gsel_0);
  BUFEHD I13 (o_1r, gsel_1);
  BUFEHD I14 (o_2r, gsel_2);
  OR3EHD I15 (oack_0, o_0a, o_1a, o_2a);
  AO222EHD I16 (i_0a, oack_0, icomplete_0, i_0a, oack_0, i_0a, icomplete_0);
endmodule

// tkf1mo0w1_o0w0 TeakF [0,0] [One 1,Many [1,0]]
module tkf1mo0w1_o0w0 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r, o_1a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  wire tech7_int;
  OR2EHD I0 (icomplete_0, i_0r0, i_0r1);
  BUFEHD I1 (acomplete_0, icomplete_0);
  BUFEHD I2 (o_0r0, i_0r0);
  BUFEHD I3 (o_0r1, i_0r1);
  BUFEHD I4 (o_1r, icomplete_0);
  AO222EHD I5 (tech7_int, acomplete_0, o_0a, tech7_int, acomplete_0, tech7_int, o_0a);
  AO222EHD I6 (i_0a, tech7_int, o_1a, i_0a, tech7_int, i_0a, o_1a);
endmodule

// tks1_o0w1_0o0w0_1o0w0 TeakS (0+:1) [([Imp 0 0],0),([Imp 1 0],0)] [One 1,Many [0,0]]
module tks1_o0w1_0o0w0_1o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire comp_0;
  BUFEHD I0 (sel_0, match0_0);
  BUFEHD I1 (match0_0, i_0r0);
  BUFEHD I2 (sel_1, match1_0);
  BUFEHD I3 (match1_0, i_0r1);
  AO222EHD I4 (gsel_0, sel_0, icomplete_0, gsel_0, sel_0, gsel_0, icomplete_0);
  AO222EHD I5 (gsel_1, sel_1, icomplete_0, gsel_1, sel_1, gsel_1, icomplete_0);
  OR2EHD I6 (comp_0, i_0r0, i_0r1);
  BUFEHD I7 (icomplete_0, comp_0);
  BUFEHD I8 (o_0r, gsel_0);
  BUFEHD I9 (o_1r, gsel_1);
  OR2EHD I10 (oack_0, o_0a, o_1a);
  AO222EHD I11 (i_0a, oack_0, icomplete_0, i_0a, oack_0, i_0a, icomplete_0);
endmodule

// tki TeakI [One 0,One 0]
module tki (i_0r, i_0a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  input reset;
  wire nreset_0;
  wire firsthsa_0;
  wire nfirsthsa_0;
  wire firsthsd_0;
  wire noa_0;
  INVHHD I0 (nreset_0, reset);
  INVHHD I1 (nfirsthsa_0, firsthsa_0);
  INVHHD I2 (noa_0, o_0a);
  AO22EHD I3 (o_0r, nreset_0, nfirsthsa_0, i_0r, firsthsd_0);
  AO12EHD I4 (firsthsa_0, nreset_0, nreset_0, o_0a);
  AO12EHD I5 (firsthsd_0, firsthsa_0, firsthsa_0, noa_0);
  AN2EHD I6 (i_0a, o_0a, firsthsd_0);
endmodule

// latch tkl0x3 width = 0, depth = 3
module tkl0x3 (i_0r, i_0a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  input reset;
  wire bf_0;
  wire ba_0;
  wire bb_0;
  wire tech3_oint;
  wire bof_0;
  wire boa_0;
  wire bob_0;
  wire tech9_oint;
  wire boo_0;
  wire tech13_oint;
  AO222EHD I0 (bf_0, i_0r, bb_0, tech3_oint, i_0r, tech3_oint, bb_0);
  AN2B1CHD I1 (tech3_oint, bf_0, reset);
  INVHHD I2 (bb_0, ba_0);
  BUFEHD I3 (i_0a, bf_0);
  AO222EHD I4 (bof_0, bf_0, bob_0, tech9_oint, bf_0, tech9_oint, bob_0);
  AN2B1CHD I5 (tech9_oint, bof_0, reset);
  INVHHD I6 (bob_0, boa_0);
  BUFEHD I7 (ba_0, bof_0);
  AO222EHD I8 (o_0r, bof_0, boo_0, tech13_oint, bof_0, tech13_oint, boo_0);
  AN2B1CHD I9 (tech13_oint, o_0r, reset);
  INVHHD I10 (boo_0, o_0a);
  BUFEHD I11 (boa_0, o_0r);
endmodule

module teak_Shifter (shift_0r0, shift_0r1, shift_0a, distanceI_0r0, distanceI_0r1, distanceI_0a, result_0r0, result_0r1, result_0a, arg_0r0, arg_0r1, arg_0a, reset);
  input [1:0] shift_0r0;
  input [1:0] shift_0r1;
  output shift_0a;
  input [4:0] distanceI_0r0;
  input [4:0] distanceI_0r1;
  output distanceI_0a;
  output [31:0] result_0r0;
  output [31:0] result_0r1;
  input result_0a;
  input [31:0] arg_0r0;
  input [31:0] arg_0r1;
  output arg_0a;
  input reset;
  wire L1_0r;
  wire L1_0a;
  wire [31:0] L35_0r0;
  wire [31:0] L35_0r1;
  wire L35_0a;
  wire L37_0r;
  wire L37_0a;
  wire L38_0r;
  wire L38_0a;
  wire [31:0] L72_0r0;
  wire [31:0] L72_0r1;
  wire L72_0a;
  wire L74_0r;
  wire L74_0a;
  wire L76P_0r;
  wire L76P_0a;
  wire L76A_0r;
  wire L76A_0a;
  wire [31:0] L78_0r0;
  wire [31:0] L78_0r1;
  wire L78_0a;
  wire [31:0] L80_0r0;
  wire [31:0] L80_0r1;
  wire L80_0a;
  wire [31:0] L82_0r0;
  wire [31:0] L82_0r1;
  wire L82_0a;
  wire [31:0] L84_0r0;
  wire [31:0] L84_0r1;
  wire L84_0a;
  wire [31:0] L87_0r0;
  wire [31:0] L87_0r1;
  wire L87_0a;
  wire L100_0r;
  wire L100_0a;
  wire [31:0] L106_0r0;
  wire [31:0] L106_0r1;
  wire L106_0a;
  wire [31:0] L108_0r0;
  wire [31:0] L108_0r1;
  wire L108_0a;
  wire [31:0] L110_0r0;
  wire [31:0] L110_0r1;
  wire L110_0a;
  wire [31:0] L112_0r0;
  wire [31:0] L112_0r1;
  wire L112_0a;
  wire [31:0] L113_0r0;
  wire [31:0] L113_0r1;
  wire L113_0a;
  wire L114_0r;
  wire L114_0a;
  wire [6:0] L129_0r0;
  wire [6:0] L129_0r1;
  wire L129_0a;
  wire [30:0] L137_0r0;
  wire [30:0] L137_0r1;
  wire L137_0a;
  wire [30:0] L138_0r0;
  wire [30:0] L138_0r1;
  wire L138_0a;
  wire [30:0] L139_0r0;
  wire [30:0] L139_0r1;
  wire L139_0a;
  wire [29:0] L140_0r0;
  wire [29:0] L140_0r1;
  wire L140_0a;
  wire [29:0] L141_0r0;
  wire [29:0] L141_0r1;
  wire L141_0a;
  wire [29:0] L142_0r0;
  wire [29:0] L142_0r1;
  wire L142_0a;
  wire L143_0r;
  wire L143_0a;
  wire L144_0r;
  wire L144_0a;
  wire L148_0r0;
  wire L148_0r1;
  wire L148_0a;
  wire L149_0r;
  wire L149_0a;
  wire [6:0] L151_0r0;
  wire [6:0] L151_0r1;
  wire L151_0a;
  wire L152_0r0;
  wire L152_0r1;
  wire L152_0a;
  wire L154_0r;
  wire L154_0a;
  wire L156_0r;
  wire L156_0a;
  wire L157_0r;
  wire L157_0a;
  wire L158_0r;
  wire L158_0a;
  wire L159_0r;
  wire L159_0a;
  wire L160_0r;
  wire L160_0a;
  wire L161_0r;
  wire L161_0a;
  wire L162_0r;
  wire L162_0a;
  wire [1:0] L175_0r0;
  wire [1:0] L175_0r1;
  wire L175_0a;
  wire [1:0] L181_0r0;
  wire [1:0] L181_0r1;
  wire L181_0a;
  wire L183_0r;
  wire L183_0a;
  wire L184_0r;
  wire L184_0a;
  wire L185_0r0;
  wire L185_0r1;
  wire L185_0a;
  wire L186_0r0;
  wire L186_0r1;
  wire L186_0a;
  wire L188_0r0;
  wire L188_0r1;
  wire L188_0a;
  wire L189_0r0;
  wire L189_0r1;
  wire L189_0a;
  tko31m32_1nm1b0_2apt1o0w1bi0w31b I0 (L137_0r0[30:0], L137_0r1[30:0], L137_0a, L108_0r0[31:0], L108_0r1[31:0], L108_0a, reset);
  tko31m32_1nm1b0_2api0w31bt1o0w1b I1 (L138_0r0[30:0], L138_0r1[30:0], L138_0a, L110_0r0[31:0], L110_0r1[31:0], L110_0a, reset);
  tko31m32_1nm1b1_2api0w31bt1o0w1b I2 (L139_0r0[30:0], L139_0r1[30:0], L139_0a, L112_0r0[31:0], L112_0r1[31:0], L112_0a, reset);
  tkvi32_wo0w32_ro0w32o0w31o1w31o1w31 I3 (L35_0r0[31:0], L35_0r1[31:0], L35_0a, L1_0r, L1_0a, L144_0r, L144_0a, L160_0r, L160_0a, L161_0r, L161_0a, L162_0r, L162_0a, L106_0r0[31:0], L106_0r1[31:0], L106_0a, L137_0r0[30:0], L137_0r1[30:0], L137_0a, L138_0r0[30:0], L138_0r1[30:0], L138_0a, L139_0r0[30:0], L139_0r1[30:0], L139_0a, reset);
  tko30m32_1nm2b0_2apt1o0w2bi0w30b I4 (L140_0r0[29:0], L140_0r1[29:0], L140_0a, L80_0r0[31:0], L80_0r1[31:0], L80_0a, reset);
  tko30m32_1nm2b0_2api0w30bt1o0w2b I5 (L141_0r0[29:0], L141_0r1[29:0], L141_0a, L82_0r0[31:0], L82_0r1[31:0], L82_0a, reset);
  tko30m32_1nm2b3_2api0w30bt1o0w2b I6 (L142_0r0[29:0], L142_0r1[29:0], L142_0a, L84_0r0[31:0], L84_0r1[31:0], L84_0a, reset);
  tkvi32_wo0w32_ro0w32o0w30o2w30o2w30 I7 (L72_0r0[31:0], L72_0r1[31:0], L72_0a, L38_0r, L38_0a, L143_0r, L143_0a, L157_0r, L157_0a, L158_0r, L158_0a, L159_0r, L159_0a, L78_0r0[31:0], L78_0r1[31:0], L78_0a, L140_0r0[29:0], L140_0r1[29:0], L140_0a, L141_0r0[29:0], L141_0r1[29:0], L141_0a, L142_0r0[29:0], L142_0r1[29:0], L142_0a, reset);
  tkj0m0_0_0 I8 (L114_0r, L114_0a, L156_0r, L156_0a, L154_0r, L154_0a, L76A_0r, L76A_0a, reset);
  tkm4x32b I9 (L78_0r0[31:0], L78_0r1[31:0], L78_0a, L80_0r0[31:0], L80_0r1[31:0], L80_0a, L82_0r0[31:0], L82_0r1[31:0], L82_0a, L84_0r0[31:0], L84_0r1[31:0], L84_0a, L87_0r0[31:0], L87_0r1[31:0], L87_0a, reset);
  tkj32m32_0 I10 (L87_0r0[31:0], L87_0r1[31:0], L87_0a, L37_0r, L37_0a, L35_0r0[31:0], L35_0r1[31:0], L35_0a, reset);
  tkm4x32b I11 (L106_0r0[31:0], L106_0r1[31:0], L106_0a, L108_0r0[31:0], L108_0r1[31:0], L108_0a, L110_0r0[31:0], L110_0r1[31:0], L110_0a, L112_0r0[31:0], L112_0r1[31:0], L112_0a, L113_0r0[31:0], L113_0r1[31:0], L113_0a, reset);
  tkf32mo0w0_o0w32 I12 (L113_0r0[31:0], L113_0r1[31:0], L113_0a, L114_0r, L114_0a, result_0r0[31:0], result_0r1[31:0], result_0a, reset);
  tkj32m32_0 I13 (arg_0r0[31:0], arg_0r1[31:0], arg_0a, L74_0r, L74_0a, L72_0r0[31:0], L72_0r1[31:0], L72_0a, reset);
  tkj7m5_2_0 I14 (distanceI_0r0[4:0], distanceI_0r1[4:0], distanceI_0a, shift_0r0[1:0], shift_0r1[1:0], shift_0a, L100_0r, L100_0a, L129_0r0[6:0], L129_0r1[6:0], L129_0a, reset);
  tkvdistanceIshift7_wo0w7_ro5w2o5w2 I15 (L151_0r0[6:0], L151_0r1[6:0], L151_0a, L149_0r, L149_0a, L183_0r, L183_0a, L184_0r, L184_0a, L175_0r0[1:0], L175_0r1[1:0], L175_0a, L181_0r0[1:0], L181_0r1[1:0], L181_0a, reset);
  tkf7mo0w7_o2w1_o1w1 I16 (L129_0r0[6:0], L129_0r1[6:0], L129_0a, L151_0r0[6:0], L151_0r1[6:0], L151_0a, L152_0r0, L152_0r1, L152_0a, L148_0r0, L148_0r1, L148_0a, reset);
  tkj1m1_0 I17 (L148_0r0, L148_0r1, L148_0a, L1_0r, L1_0a, L185_0r0, L185_0r1, L185_0a, reset);
  tkj1m1_0 I18 (L152_0r0, L152_0r1, L152_0a, L38_0r, L38_0a, L188_0r0, L188_0r1, L188_0a, reset);
  tkf0mo0w0_o0w0 I19 (L149_0r, L149_0a, L74_0r, L74_0a, L37_0r, L37_0a, reset);
  tks2_o0w2_3o0w0_0c2o0w0_1o0w0 I20 (L175_0r0[1:0], L175_0r1[1:0], L175_0a, L162_0r, L162_0a, L160_0r, L160_0a, L161_0r, L161_0a, reset);
  tks2_o0w2_3o0w0_0c2o0w0_1o0w0 I21 (L181_0r0[1:0], L181_0r1[1:0], L181_0a, L159_0r, L159_0a, L157_0r, L157_0a, L158_0r, L158_0a, reset);
  tkf1mo0w1_o0w0 I22 (L185_0r0, L185_0r1, L185_0a, L186_0r0, L186_0r1, L186_0a, L156_0r, L156_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I23 (L186_0r0, L186_0r1, L186_0a, L144_0r, L144_0a, L183_0r, L183_0a, reset);
  tkf1mo0w1_o0w0 I24 (L188_0r0, L188_0r1, L188_0a, L189_0r0, L189_0r1, L189_0a, L154_0r, L154_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I25 (L189_0r0, L189_0r1, L189_0a, L143_0r, L143_0a, L184_0r, L184_0a, reset);
  tki I26 (L76P_0r, L76P_0a, L100_0r, L100_0a, reset);
  tkl0x3 I27 (L76A_0r, L76A_0a, L76P_0r, L76P_0a, reset);
endmodule

// Netlist costs:
// teak_Shifter: AN2B1CHD*19 AN2EHD*1370 AO12EHD*5 AO222EHD*630 AO22EHD*72 BUFEHD*1076 INVHHD*140 ND2HHD*131 ND3EHD*2 NR2EHD*78 NR3EHD*206 OR2EHD*523 OR3EHD*2 TIE0DND*9
// tkf0mo0w0_o0w0: AO222EHD*1 BUFEHD*2
// tkf1mo0w1_o0w0: AO222EHD*2 BUFEHD*4 OR2EHD*1
// tkf32mo0w0_o0w32: AO222EHD*2 BUFEHD*66 OR2EHD*1
// tkf7mo0w7_o2w1_o1w1: AO222EHD*7 BUFEHD*16 OR2EHD*1
// tki: AN2EHD*1 AO12EHD*2 AO22EHD*1 INVHHD*3
// tkj0m0_0_0: AO222EHD*2 BUFEHD*3
// tkj1m1_0: AO222EHD*2 BUFEHD*5
// tkj32m32_0: AO222EHD*2 BUFEHD*129
// tkj7m5_2_0: AO222EHD*3 BUFEHD*29 OR2EHD*1
// tkl0x3: AN2B1CHD*3 AO222EHD*3 BUFEHD*3 INVHHD*3
// tkm4x32b: AN2B1CHD*8 AN2EHD*256 AO222EHD*132 BUFEHD*4 INVHHD*65 ND2HHD*65 NR2EHD*1 NR3EHD*65 OR2EHD*128
// tko30m32_1nm2b0_2api0w30bt1o0w2b: AO222EHD*29 BUFEHD*69 OR2EHD*30 TIE0DND*2
// tko30m32_1nm2b0_2apt1o0w2bi0w30b: AO222EHD*29 BUFEHD*69 OR2EHD*30 TIE0DND*2
// tko30m32_1nm2b3_2api0w30bt1o0w2b: AO222EHD*29 BUFEHD*69 OR2EHD*30 TIE0DND*2
// tko31m32_1nm1b0_2api0w31bt1o0w1b: AO222EHD*30 BUFEHD*68 OR2EHD*31 TIE0DND*1
// tko31m32_1nm1b0_2apt1o0w1bi0w31b: AO222EHD*30 BUFEHD*68 OR2EHD*31 TIE0DND*1
// tko31m32_1nm1b1_2api0w31bt1o0w1b: AO222EHD*30 BUFEHD*68 OR2EHD*31 TIE0DND*1
// tks1_o0w1_0o0w0_1o0w0: AO222EHD*3 BUFEHD*7 OR2EHD*2
// tks2_o0w2_3o0w0_0c2o0w0_1o0w0: AO222EHD*7 BUFEHD*7 OR2EHD*2 OR3EHD*1
// tkvdistanceIshift7_wo0w7_ro5w2o5w2: AN2EHD*43 AO12EHD*1 AO222EHD*13 AO22EHD*7 BUFEHD*26 INVHHD*2 ND2HHD*1 NR2EHD*8 NR3EHD*8 OR2EHD*7
// tkvi32_wo0w32_ro0w32o0w30o2w30o2w30: AN2EHD*404 AO12EHD*1 AO222EHD*63 AO22EHD*32 BUFEHD*104 INVHHD*1 ND3EHD*1 NR2EHD*34 NR3EHD*34 OR2EHD*32
// tkvi32_wo0w32_ro0w32o0w31o1w31o1w31: AN2EHD*410 AO12EHD*1 AO222EHD*63 AO22EHD*32 BUFEHD*104 INVHHD*1 ND3EHD*1 NR2EHD*34 NR3EHD*34 OR2EHD*32
