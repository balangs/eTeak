//
// from command: teak -v --gates --test-protocol -L -l before-i=3 -n shifter.teak -o shifter
//
// Generated on: Sun Sep  6 07:18:06 BST 2015
//


`timescale 1ns/1ps

// tko31m32_1nm1b0_2apt1o0w1bi0w31b TeakO [
//     (1,TeakOConstant 1 0),
//     (2,TeakOAppend 1 [(1,0+:1),(0,0+:31)])] [One 31,One 32]
module tko31m32_1nm1b0_2apt1o0w1bi0w31b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [30:0] i_0r0;
  input [30:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [30:0] gocomp_0;
  wire [10:0] simp331_0;
  wire [3:0] simp332_0;
  wire [1:0] simp333_0;
  wire termf_1;
  wire termt_1;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I30 (gocomp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  C3 I31 (simp331_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  C3 I32 (simp331_0[1:1], gocomp_0[3:3], gocomp_0[4:4], gocomp_0[5:5]);
  C3 I33 (simp331_0[2:2], gocomp_0[6:6], gocomp_0[7:7], gocomp_0[8:8]);
  C3 I34 (simp331_0[3:3], gocomp_0[9:9], gocomp_0[10:10], gocomp_0[11:11]);
  C3 I35 (simp331_0[4:4], gocomp_0[12:12], gocomp_0[13:13], gocomp_0[14:14]);
  C3 I36 (simp331_0[5:5], gocomp_0[15:15], gocomp_0[16:16], gocomp_0[17:17]);
  C3 I37 (simp331_0[6:6], gocomp_0[18:18], gocomp_0[19:19], gocomp_0[20:20]);
  C3 I38 (simp331_0[7:7], gocomp_0[21:21], gocomp_0[22:22], gocomp_0[23:23]);
  C3 I39 (simp331_0[8:8], gocomp_0[24:24], gocomp_0[25:25], gocomp_0[26:26]);
  C3 I40 (simp331_0[9:9], gocomp_0[27:27], gocomp_0[28:28], gocomp_0[29:29]);
  BUFF I41 (simp331_0[10:10], gocomp_0[30:30]);
  C3 I42 (simp332_0[0:0], simp331_0[0:0], simp331_0[1:1], simp331_0[2:2]);
  C3 I43 (simp332_0[1:1], simp331_0[3:3], simp331_0[4:4], simp331_0[5:5]);
  C3 I44 (simp332_0[2:2], simp331_0[6:6], simp331_0[7:7], simp331_0[8:8]);
  C2 I45 (simp332_0[3:3], simp331_0[9:9], simp331_0[10:10]);
  C3 I46 (simp333_0[0:0], simp332_0[0:0], simp332_0[1:1], simp332_0[2:2]);
  BUFF I47 (simp333_0[1:1], simp332_0[3:3]);
  C2 I48 (go_0, simp333_0[0:0], simp333_0[1:1]);
  BUFF I49 (termf_1, go_0);
  GND I50 (termt_1);
  BUFF I51 (o_0r0[0:0], termf_1);
  BUFF I52 (o_0r0[1:1], i_0r0[0:0]);
  BUFF I53 (o_0r0[2:2], i_0r0[1:1]);
  BUFF I54 (o_0r0[3:3], i_0r0[2:2]);
  BUFF I55 (o_0r0[4:4], i_0r0[3:3]);
  BUFF I56 (o_0r0[5:5], i_0r0[4:4]);
  BUFF I57 (o_0r0[6:6], i_0r0[5:5]);
  BUFF I58 (o_0r0[7:7], i_0r0[6:6]);
  BUFF I59 (o_0r0[8:8], i_0r0[7:7]);
  BUFF I60 (o_0r0[9:9], i_0r0[8:8]);
  BUFF I61 (o_0r0[10:10], i_0r0[9:9]);
  BUFF I62 (o_0r0[11:11], i_0r0[10:10]);
  BUFF I63 (o_0r0[12:12], i_0r0[11:11]);
  BUFF I64 (o_0r0[13:13], i_0r0[12:12]);
  BUFF I65 (o_0r0[14:14], i_0r0[13:13]);
  BUFF I66 (o_0r0[15:15], i_0r0[14:14]);
  BUFF I67 (o_0r0[16:16], i_0r0[15:15]);
  BUFF I68 (o_0r0[17:17], i_0r0[16:16]);
  BUFF I69 (o_0r0[18:18], i_0r0[17:17]);
  BUFF I70 (o_0r0[19:19], i_0r0[18:18]);
  BUFF I71 (o_0r0[20:20], i_0r0[19:19]);
  BUFF I72 (o_0r0[21:21], i_0r0[20:20]);
  BUFF I73 (o_0r0[22:22], i_0r0[21:21]);
  BUFF I74 (o_0r0[23:23], i_0r0[22:22]);
  BUFF I75 (o_0r0[24:24], i_0r0[23:23]);
  BUFF I76 (o_0r0[25:25], i_0r0[24:24]);
  BUFF I77 (o_0r0[26:26], i_0r0[25:25]);
  BUFF I78 (o_0r0[27:27], i_0r0[26:26]);
  BUFF I79 (o_0r0[28:28], i_0r0[27:27]);
  BUFF I80 (o_0r0[29:29], i_0r0[28:28]);
  BUFF I81 (o_0r0[30:30], i_0r0[29:29]);
  BUFF I82 (o_0r0[31:31], i_0r0[30:30]);
  BUFF I83 (o_0r1[0:0], termt_1);
  BUFF I84 (o_0r1[1:1], i_0r1[0:0]);
  BUFF I85 (o_0r1[2:2], i_0r1[1:1]);
  BUFF I86 (o_0r1[3:3], i_0r1[2:2]);
  BUFF I87 (o_0r1[4:4], i_0r1[3:3]);
  BUFF I88 (o_0r1[5:5], i_0r1[4:4]);
  BUFF I89 (o_0r1[6:6], i_0r1[5:5]);
  BUFF I90 (o_0r1[7:7], i_0r1[6:6]);
  BUFF I91 (o_0r1[8:8], i_0r1[7:7]);
  BUFF I92 (o_0r1[9:9], i_0r1[8:8]);
  BUFF I93 (o_0r1[10:10], i_0r1[9:9]);
  BUFF I94 (o_0r1[11:11], i_0r1[10:10]);
  BUFF I95 (o_0r1[12:12], i_0r1[11:11]);
  BUFF I96 (o_0r1[13:13], i_0r1[12:12]);
  BUFF I97 (o_0r1[14:14], i_0r1[13:13]);
  BUFF I98 (o_0r1[15:15], i_0r1[14:14]);
  BUFF I99 (o_0r1[16:16], i_0r1[15:15]);
  BUFF I100 (o_0r1[17:17], i_0r1[16:16]);
  BUFF I101 (o_0r1[18:18], i_0r1[17:17]);
  BUFF I102 (o_0r1[19:19], i_0r1[18:18]);
  BUFF I103 (o_0r1[20:20], i_0r1[19:19]);
  BUFF I104 (o_0r1[21:21], i_0r1[20:20]);
  BUFF I105 (o_0r1[22:22], i_0r1[21:21]);
  BUFF I106 (o_0r1[23:23], i_0r1[22:22]);
  BUFF I107 (o_0r1[24:24], i_0r1[23:23]);
  BUFF I108 (o_0r1[25:25], i_0r1[24:24]);
  BUFF I109 (o_0r1[26:26], i_0r1[25:25]);
  BUFF I110 (o_0r1[27:27], i_0r1[26:26]);
  BUFF I111 (o_0r1[28:28], i_0r1[27:27]);
  BUFF I112 (o_0r1[29:29], i_0r1[28:28]);
  BUFF I113 (o_0r1[30:30], i_0r1[29:29]);
  BUFF I114 (o_0r1[31:31], i_0r1[30:30]);
  BUFF I115 (i_0a, o_0a);
endmodule

// tko31m32_1nm1b0_2api0w31bt1o0w1b TeakO [
//     (1,TeakOConstant 1 0),
//     (2,TeakOAppend 1 [(0,0+:31),(1,0+:1)])] [One 31,One 32]
module tko31m32_1nm1b0_2api0w31bt1o0w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [30:0] i_0r0;
  input [30:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [30:0] gocomp_0;
  wire [10:0] simp331_0;
  wire [3:0] simp332_0;
  wire [1:0] simp333_0;
  wire termf_1;
  wire termt_1;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I30 (gocomp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  C3 I31 (simp331_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  C3 I32 (simp331_0[1:1], gocomp_0[3:3], gocomp_0[4:4], gocomp_0[5:5]);
  C3 I33 (simp331_0[2:2], gocomp_0[6:6], gocomp_0[7:7], gocomp_0[8:8]);
  C3 I34 (simp331_0[3:3], gocomp_0[9:9], gocomp_0[10:10], gocomp_0[11:11]);
  C3 I35 (simp331_0[4:4], gocomp_0[12:12], gocomp_0[13:13], gocomp_0[14:14]);
  C3 I36 (simp331_0[5:5], gocomp_0[15:15], gocomp_0[16:16], gocomp_0[17:17]);
  C3 I37 (simp331_0[6:6], gocomp_0[18:18], gocomp_0[19:19], gocomp_0[20:20]);
  C3 I38 (simp331_0[7:7], gocomp_0[21:21], gocomp_0[22:22], gocomp_0[23:23]);
  C3 I39 (simp331_0[8:8], gocomp_0[24:24], gocomp_0[25:25], gocomp_0[26:26]);
  C3 I40 (simp331_0[9:9], gocomp_0[27:27], gocomp_0[28:28], gocomp_0[29:29]);
  BUFF I41 (simp331_0[10:10], gocomp_0[30:30]);
  C3 I42 (simp332_0[0:0], simp331_0[0:0], simp331_0[1:1], simp331_0[2:2]);
  C3 I43 (simp332_0[1:1], simp331_0[3:3], simp331_0[4:4], simp331_0[5:5]);
  C3 I44 (simp332_0[2:2], simp331_0[6:6], simp331_0[7:7], simp331_0[8:8]);
  C2 I45 (simp332_0[3:3], simp331_0[9:9], simp331_0[10:10]);
  C3 I46 (simp333_0[0:0], simp332_0[0:0], simp332_0[1:1], simp332_0[2:2]);
  BUFF I47 (simp333_0[1:1], simp332_0[3:3]);
  C2 I48 (go_0, simp333_0[0:0], simp333_0[1:1]);
  BUFF I49 (termf_1, go_0);
  GND I50 (termt_1);
  BUFF I51 (o_0r0[0:0], i_0r0[0:0]);
  BUFF I52 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I53 (o_0r0[2:2], i_0r0[2:2]);
  BUFF I54 (o_0r0[3:3], i_0r0[3:3]);
  BUFF I55 (o_0r0[4:4], i_0r0[4:4]);
  BUFF I56 (o_0r0[5:5], i_0r0[5:5]);
  BUFF I57 (o_0r0[6:6], i_0r0[6:6]);
  BUFF I58 (o_0r0[7:7], i_0r0[7:7]);
  BUFF I59 (o_0r0[8:8], i_0r0[8:8]);
  BUFF I60 (o_0r0[9:9], i_0r0[9:9]);
  BUFF I61 (o_0r0[10:10], i_0r0[10:10]);
  BUFF I62 (o_0r0[11:11], i_0r0[11:11]);
  BUFF I63 (o_0r0[12:12], i_0r0[12:12]);
  BUFF I64 (o_0r0[13:13], i_0r0[13:13]);
  BUFF I65 (o_0r0[14:14], i_0r0[14:14]);
  BUFF I66 (o_0r0[15:15], i_0r0[15:15]);
  BUFF I67 (o_0r0[16:16], i_0r0[16:16]);
  BUFF I68 (o_0r0[17:17], i_0r0[17:17]);
  BUFF I69 (o_0r0[18:18], i_0r0[18:18]);
  BUFF I70 (o_0r0[19:19], i_0r0[19:19]);
  BUFF I71 (o_0r0[20:20], i_0r0[20:20]);
  BUFF I72 (o_0r0[21:21], i_0r0[21:21]);
  BUFF I73 (o_0r0[22:22], i_0r0[22:22]);
  BUFF I74 (o_0r0[23:23], i_0r0[23:23]);
  BUFF I75 (o_0r0[24:24], i_0r0[24:24]);
  BUFF I76 (o_0r0[25:25], i_0r0[25:25]);
  BUFF I77 (o_0r0[26:26], i_0r0[26:26]);
  BUFF I78 (o_0r0[27:27], i_0r0[27:27]);
  BUFF I79 (o_0r0[28:28], i_0r0[28:28]);
  BUFF I80 (o_0r0[29:29], i_0r0[29:29]);
  BUFF I81 (o_0r0[30:30], i_0r0[30:30]);
  BUFF I82 (o_0r0[31:31], termf_1);
  BUFF I83 (o_0r1[0:0], i_0r1[0:0]);
  BUFF I84 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I85 (o_0r1[2:2], i_0r1[2:2]);
  BUFF I86 (o_0r1[3:3], i_0r1[3:3]);
  BUFF I87 (o_0r1[4:4], i_0r1[4:4]);
  BUFF I88 (o_0r1[5:5], i_0r1[5:5]);
  BUFF I89 (o_0r1[6:6], i_0r1[6:6]);
  BUFF I90 (o_0r1[7:7], i_0r1[7:7]);
  BUFF I91 (o_0r1[8:8], i_0r1[8:8]);
  BUFF I92 (o_0r1[9:9], i_0r1[9:9]);
  BUFF I93 (o_0r1[10:10], i_0r1[10:10]);
  BUFF I94 (o_0r1[11:11], i_0r1[11:11]);
  BUFF I95 (o_0r1[12:12], i_0r1[12:12]);
  BUFF I96 (o_0r1[13:13], i_0r1[13:13]);
  BUFF I97 (o_0r1[14:14], i_0r1[14:14]);
  BUFF I98 (o_0r1[15:15], i_0r1[15:15]);
  BUFF I99 (o_0r1[16:16], i_0r1[16:16]);
  BUFF I100 (o_0r1[17:17], i_0r1[17:17]);
  BUFF I101 (o_0r1[18:18], i_0r1[18:18]);
  BUFF I102 (o_0r1[19:19], i_0r1[19:19]);
  BUFF I103 (o_0r1[20:20], i_0r1[20:20]);
  BUFF I104 (o_0r1[21:21], i_0r1[21:21]);
  BUFF I105 (o_0r1[22:22], i_0r1[22:22]);
  BUFF I106 (o_0r1[23:23], i_0r1[23:23]);
  BUFF I107 (o_0r1[24:24], i_0r1[24:24]);
  BUFF I108 (o_0r1[25:25], i_0r1[25:25]);
  BUFF I109 (o_0r1[26:26], i_0r1[26:26]);
  BUFF I110 (o_0r1[27:27], i_0r1[27:27]);
  BUFF I111 (o_0r1[28:28], i_0r1[28:28]);
  BUFF I112 (o_0r1[29:29], i_0r1[29:29]);
  BUFF I113 (o_0r1[30:30], i_0r1[30:30]);
  BUFF I114 (o_0r1[31:31], termt_1);
  BUFF I115 (i_0a, o_0a);
endmodule

// tko31m32_1nm1b1_2api0w31bt1o0w1b TeakO [
//     (1,TeakOConstant 1 1),
//     (2,TeakOAppend 1 [(0,0+:31),(1,0+:1)])] [One 31,One 32]
module tko31m32_1nm1b1_2api0w31bt1o0w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [30:0] i_0r0;
  input [30:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [30:0] gocomp_0;
  wire [10:0] simp331_0;
  wire [3:0] simp332_0;
  wire [1:0] simp333_0;
  wire termf_1;
  wire termt_1;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I30 (gocomp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  C3 I31 (simp331_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  C3 I32 (simp331_0[1:1], gocomp_0[3:3], gocomp_0[4:4], gocomp_0[5:5]);
  C3 I33 (simp331_0[2:2], gocomp_0[6:6], gocomp_0[7:7], gocomp_0[8:8]);
  C3 I34 (simp331_0[3:3], gocomp_0[9:9], gocomp_0[10:10], gocomp_0[11:11]);
  C3 I35 (simp331_0[4:4], gocomp_0[12:12], gocomp_0[13:13], gocomp_0[14:14]);
  C3 I36 (simp331_0[5:5], gocomp_0[15:15], gocomp_0[16:16], gocomp_0[17:17]);
  C3 I37 (simp331_0[6:6], gocomp_0[18:18], gocomp_0[19:19], gocomp_0[20:20]);
  C3 I38 (simp331_0[7:7], gocomp_0[21:21], gocomp_0[22:22], gocomp_0[23:23]);
  C3 I39 (simp331_0[8:8], gocomp_0[24:24], gocomp_0[25:25], gocomp_0[26:26]);
  C3 I40 (simp331_0[9:9], gocomp_0[27:27], gocomp_0[28:28], gocomp_0[29:29]);
  BUFF I41 (simp331_0[10:10], gocomp_0[30:30]);
  C3 I42 (simp332_0[0:0], simp331_0[0:0], simp331_0[1:1], simp331_0[2:2]);
  C3 I43 (simp332_0[1:1], simp331_0[3:3], simp331_0[4:4], simp331_0[5:5]);
  C3 I44 (simp332_0[2:2], simp331_0[6:6], simp331_0[7:7], simp331_0[8:8]);
  C2 I45 (simp332_0[3:3], simp331_0[9:9], simp331_0[10:10]);
  C3 I46 (simp333_0[0:0], simp332_0[0:0], simp332_0[1:1], simp332_0[2:2]);
  BUFF I47 (simp333_0[1:1], simp332_0[3:3]);
  C2 I48 (go_0, simp333_0[0:0], simp333_0[1:1]);
  BUFF I49 (termt_1, go_0);
  GND I50 (termf_1);
  BUFF I51 (o_0r0[0:0], i_0r0[0:0]);
  BUFF I52 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I53 (o_0r0[2:2], i_0r0[2:2]);
  BUFF I54 (o_0r0[3:3], i_0r0[3:3]);
  BUFF I55 (o_0r0[4:4], i_0r0[4:4]);
  BUFF I56 (o_0r0[5:5], i_0r0[5:5]);
  BUFF I57 (o_0r0[6:6], i_0r0[6:6]);
  BUFF I58 (o_0r0[7:7], i_0r0[7:7]);
  BUFF I59 (o_0r0[8:8], i_0r0[8:8]);
  BUFF I60 (o_0r0[9:9], i_0r0[9:9]);
  BUFF I61 (o_0r0[10:10], i_0r0[10:10]);
  BUFF I62 (o_0r0[11:11], i_0r0[11:11]);
  BUFF I63 (o_0r0[12:12], i_0r0[12:12]);
  BUFF I64 (o_0r0[13:13], i_0r0[13:13]);
  BUFF I65 (o_0r0[14:14], i_0r0[14:14]);
  BUFF I66 (o_0r0[15:15], i_0r0[15:15]);
  BUFF I67 (o_0r0[16:16], i_0r0[16:16]);
  BUFF I68 (o_0r0[17:17], i_0r0[17:17]);
  BUFF I69 (o_0r0[18:18], i_0r0[18:18]);
  BUFF I70 (o_0r0[19:19], i_0r0[19:19]);
  BUFF I71 (o_0r0[20:20], i_0r0[20:20]);
  BUFF I72 (o_0r0[21:21], i_0r0[21:21]);
  BUFF I73 (o_0r0[22:22], i_0r0[22:22]);
  BUFF I74 (o_0r0[23:23], i_0r0[23:23]);
  BUFF I75 (o_0r0[24:24], i_0r0[24:24]);
  BUFF I76 (o_0r0[25:25], i_0r0[25:25]);
  BUFF I77 (o_0r0[26:26], i_0r0[26:26]);
  BUFF I78 (o_0r0[27:27], i_0r0[27:27]);
  BUFF I79 (o_0r0[28:28], i_0r0[28:28]);
  BUFF I80 (o_0r0[29:29], i_0r0[29:29]);
  BUFF I81 (o_0r0[30:30], i_0r0[30:30]);
  BUFF I82 (o_0r0[31:31], termf_1);
  BUFF I83 (o_0r1[0:0], i_0r1[0:0]);
  BUFF I84 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I85 (o_0r1[2:2], i_0r1[2:2]);
  BUFF I86 (o_0r1[3:3], i_0r1[3:3]);
  BUFF I87 (o_0r1[4:4], i_0r1[4:4]);
  BUFF I88 (o_0r1[5:5], i_0r1[5:5]);
  BUFF I89 (o_0r1[6:6], i_0r1[6:6]);
  BUFF I90 (o_0r1[7:7], i_0r1[7:7]);
  BUFF I91 (o_0r1[8:8], i_0r1[8:8]);
  BUFF I92 (o_0r1[9:9], i_0r1[9:9]);
  BUFF I93 (o_0r1[10:10], i_0r1[10:10]);
  BUFF I94 (o_0r1[11:11], i_0r1[11:11]);
  BUFF I95 (o_0r1[12:12], i_0r1[12:12]);
  BUFF I96 (o_0r1[13:13], i_0r1[13:13]);
  BUFF I97 (o_0r1[14:14], i_0r1[14:14]);
  BUFF I98 (o_0r1[15:15], i_0r1[15:15]);
  BUFF I99 (o_0r1[16:16], i_0r1[16:16]);
  BUFF I100 (o_0r1[17:17], i_0r1[17:17]);
  BUFF I101 (o_0r1[18:18], i_0r1[18:18]);
  BUFF I102 (o_0r1[19:19], i_0r1[19:19]);
  BUFF I103 (o_0r1[20:20], i_0r1[20:20]);
  BUFF I104 (o_0r1[21:21], i_0r1[21:21]);
  BUFF I105 (o_0r1[22:22], i_0r1[22:22]);
  BUFF I106 (o_0r1[23:23], i_0r1[23:23]);
  BUFF I107 (o_0r1[24:24], i_0r1[24:24]);
  BUFF I108 (o_0r1[25:25], i_0r1[25:25]);
  BUFF I109 (o_0r1[26:26], i_0r1[26:26]);
  BUFF I110 (o_0r1[27:27], i_0r1[27:27]);
  BUFF I111 (o_0r1[28:28], i_0r1[28:28]);
  BUFF I112 (o_0r1[29:29], i_0r1[29:29]);
  BUFF I113 (o_0r1[30:30], i_0r1[30:30]);
  BUFF I114 (o_0r1[31:31], termt_1);
  BUFF I115 (i_0a, o_0a);
endmodule

// tkvi32_wo0w32_ro0w32o0w31o1w31o1w31 TeakV "i" 32 [] [0] [0,0,1,1] [Many [32],Many [0],Many [0,0,0,0]
//   ,Many [32,31,31,31]]
module tkvi32_wo0w32_ro0w32o0w31o1w31o1w31 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [30:0] rd_1r0;
  output [30:0] rd_1r1;
  input rd_1a;
  output [30:0] rd_2r0;
  output [30:0] rd_2r1;
  input rd_2a;
  output [30:0] rd_3r0;
  output [30:0] rd_3r1;
  input rd_3a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [2:0] simp6581_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_2r0[0:0], df_0[1:1], rg_2r);
  AND2 I488 (rd_2r0[1:1], df_0[2:2], rg_2r);
  AND2 I489 (rd_2r0[2:2], df_0[3:3], rg_2r);
  AND2 I490 (rd_2r0[3:3], df_0[4:4], rg_2r);
  AND2 I491 (rd_2r0[4:4], df_0[5:5], rg_2r);
  AND2 I492 (rd_2r0[5:5], df_0[6:6], rg_2r);
  AND2 I493 (rd_2r0[6:6], df_0[7:7], rg_2r);
  AND2 I494 (rd_2r0[7:7], df_0[8:8], rg_2r);
  AND2 I495 (rd_2r0[8:8], df_0[9:9], rg_2r);
  AND2 I496 (rd_2r0[9:9], df_0[10:10], rg_2r);
  AND2 I497 (rd_2r0[10:10], df_0[11:11], rg_2r);
  AND2 I498 (rd_2r0[11:11], df_0[12:12], rg_2r);
  AND2 I499 (rd_2r0[12:12], df_0[13:13], rg_2r);
  AND2 I500 (rd_2r0[13:13], df_0[14:14], rg_2r);
  AND2 I501 (rd_2r0[14:14], df_0[15:15], rg_2r);
  AND2 I502 (rd_2r0[15:15], df_0[16:16], rg_2r);
  AND2 I503 (rd_2r0[16:16], df_0[17:17], rg_2r);
  AND2 I504 (rd_2r0[17:17], df_0[18:18], rg_2r);
  AND2 I505 (rd_2r0[18:18], df_0[19:19], rg_2r);
  AND2 I506 (rd_2r0[19:19], df_0[20:20], rg_2r);
  AND2 I507 (rd_2r0[20:20], df_0[21:21], rg_2r);
  AND2 I508 (rd_2r0[21:21], df_0[22:22], rg_2r);
  AND2 I509 (rd_2r0[22:22], df_0[23:23], rg_2r);
  AND2 I510 (rd_2r0[23:23], df_0[24:24], rg_2r);
  AND2 I511 (rd_2r0[24:24], df_0[25:25], rg_2r);
  AND2 I512 (rd_2r0[25:25], df_0[26:26], rg_2r);
  AND2 I513 (rd_2r0[26:26], df_0[27:27], rg_2r);
  AND2 I514 (rd_2r0[27:27], df_0[28:28], rg_2r);
  AND2 I515 (rd_2r0[28:28], df_0[29:29], rg_2r);
  AND2 I516 (rd_2r0[29:29], df_0[30:30], rg_2r);
  AND2 I517 (rd_2r0[30:30], df_0[31:31], rg_2r);
  AND2 I518 (rd_3r0[0:0], df_0[1:1], rg_3r);
  AND2 I519 (rd_3r0[1:1], df_0[2:2], rg_3r);
  AND2 I520 (rd_3r0[2:2], df_0[3:3], rg_3r);
  AND2 I521 (rd_3r0[3:3], df_0[4:4], rg_3r);
  AND2 I522 (rd_3r0[4:4], df_0[5:5], rg_3r);
  AND2 I523 (rd_3r0[5:5], df_0[6:6], rg_3r);
  AND2 I524 (rd_3r0[6:6], df_0[7:7], rg_3r);
  AND2 I525 (rd_3r0[7:7], df_0[8:8], rg_3r);
  AND2 I526 (rd_3r0[8:8], df_0[9:9], rg_3r);
  AND2 I527 (rd_3r0[9:9], df_0[10:10], rg_3r);
  AND2 I528 (rd_3r0[10:10], df_0[11:11], rg_3r);
  AND2 I529 (rd_3r0[11:11], df_0[12:12], rg_3r);
  AND2 I530 (rd_3r0[12:12], df_0[13:13], rg_3r);
  AND2 I531 (rd_3r0[13:13], df_0[14:14], rg_3r);
  AND2 I532 (rd_3r0[14:14], df_0[15:15], rg_3r);
  AND2 I533 (rd_3r0[15:15], df_0[16:16], rg_3r);
  AND2 I534 (rd_3r0[16:16], df_0[17:17], rg_3r);
  AND2 I535 (rd_3r0[17:17], df_0[18:18], rg_3r);
  AND2 I536 (rd_3r0[18:18], df_0[19:19], rg_3r);
  AND2 I537 (rd_3r0[19:19], df_0[20:20], rg_3r);
  AND2 I538 (rd_3r0[20:20], df_0[21:21], rg_3r);
  AND2 I539 (rd_3r0[21:21], df_0[22:22], rg_3r);
  AND2 I540 (rd_3r0[22:22], df_0[23:23], rg_3r);
  AND2 I541 (rd_3r0[23:23], df_0[24:24], rg_3r);
  AND2 I542 (rd_3r0[24:24], df_0[25:25], rg_3r);
  AND2 I543 (rd_3r0[25:25], df_0[26:26], rg_3r);
  AND2 I544 (rd_3r0[26:26], df_0[27:27], rg_3r);
  AND2 I545 (rd_3r0[27:27], df_0[28:28], rg_3r);
  AND2 I546 (rd_3r0[28:28], df_0[29:29], rg_3r);
  AND2 I547 (rd_3r0[29:29], df_0[30:30], rg_3r);
  AND2 I548 (rd_3r0[30:30], df_0[31:31], rg_3r);
  AND2 I549 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I550 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I551 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I552 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I553 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I554 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I555 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I556 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I557 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I558 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I559 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I560 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I561 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I562 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I563 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I564 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I565 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I566 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I567 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I568 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I569 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I570 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I571 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I572 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I573 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I574 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I575 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I576 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I577 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I578 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I579 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I580 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I581 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I582 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I583 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I584 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I585 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I586 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I587 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I588 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I589 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I590 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I591 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I592 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I593 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I594 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I595 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I596 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I597 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I598 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I599 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I600 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I601 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I602 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I603 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I604 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I605 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I606 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I607 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I608 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I609 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I610 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I611 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I612 (rd_2r1[0:0], dt_0[1:1], rg_2r);
  AND2 I613 (rd_2r1[1:1], dt_0[2:2], rg_2r);
  AND2 I614 (rd_2r1[2:2], dt_0[3:3], rg_2r);
  AND2 I615 (rd_2r1[3:3], dt_0[4:4], rg_2r);
  AND2 I616 (rd_2r1[4:4], dt_0[5:5], rg_2r);
  AND2 I617 (rd_2r1[5:5], dt_0[6:6], rg_2r);
  AND2 I618 (rd_2r1[6:6], dt_0[7:7], rg_2r);
  AND2 I619 (rd_2r1[7:7], dt_0[8:8], rg_2r);
  AND2 I620 (rd_2r1[8:8], dt_0[9:9], rg_2r);
  AND2 I621 (rd_2r1[9:9], dt_0[10:10], rg_2r);
  AND2 I622 (rd_2r1[10:10], dt_0[11:11], rg_2r);
  AND2 I623 (rd_2r1[11:11], dt_0[12:12], rg_2r);
  AND2 I624 (rd_2r1[12:12], dt_0[13:13], rg_2r);
  AND2 I625 (rd_2r1[13:13], dt_0[14:14], rg_2r);
  AND2 I626 (rd_2r1[14:14], dt_0[15:15], rg_2r);
  AND2 I627 (rd_2r1[15:15], dt_0[16:16], rg_2r);
  AND2 I628 (rd_2r1[16:16], dt_0[17:17], rg_2r);
  AND2 I629 (rd_2r1[17:17], dt_0[18:18], rg_2r);
  AND2 I630 (rd_2r1[18:18], dt_0[19:19], rg_2r);
  AND2 I631 (rd_2r1[19:19], dt_0[20:20], rg_2r);
  AND2 I632 (rd_2r1[20:20], dt_0[21:21], rg_2r);
  AND2 I633 (rd_2r1[21:21], dt_0[22:22], rg_2r);
  AND2 I634 (rd_2r1[22:22], dt_0[23:23], rg_2r);
  AND2 I635 (rd_2r1[23:23], dt_0[24:24], rg_2r);
  AND2 I636 (rd_2r1[24:24], dt_0[25:25], rg_2r);
  AND2 I637 (rd_2r1[25:25], dt_0[26:26], rg_2r);
  AND2 I638 (rd_2r1[26:26], dt_0[27:27], rg_2r);
  AND2 I639 (rd_2r1[27:27], dt_0[28:28], rg_2r);
  AND2 I640 (rd_2r1[28:28], dt_0[29:29], rg_2r);
  AND2 I641 (rd_2r1[29:29], dt_0[30:30], rg_2r);
  AND2 I642 (rd_2r1[30:30], dt_0[31:31], rg_2r);
  AND2 I643 (rd_3r1[0:0], dt_0[1:1], rg_3r);
  AND2 I644 (rd_3r1[1:1], dt_0[2:2], rg_3r);
  AND2 I645 (rd_3r1[2:2], dt_0[3:3], rg_3r);
  AND2 I646 (rd_3r1[3:3], dt_0[4:4], rg_3r);
  AND2 I647 (rd_3r1[4:4], dt_0[5:5], rg_3r);
  AND2 I648 (rd_3r1[5:5], dt_0[6:6], rg_3r);
  AND2 I649 (rd_3r1[6:6], dt_0[7:7], rg_3r);
  AND2 I650 (rd_3r1[7:7], dt_0[8:8], rg_3r);
  AND2 I651 (rd_3r1[8:8], dt_0[9:9], rg_3r);
  AND2 I652 (rd_3r1[9:9], dt_0[10:10], rg_3r);
  AND2 I653 (rd_3r1[10:10], dt_0[11:11], rg_3r);
  AND2 I654 (rd_3r1[11:11], dt_0[12:12], rg_3r);
  AND2 I655 (rd_3r1[12:12], dt_0[13:13], rg_3r);
  AND2 I656 (rd_3r1[13:13], dt_0[14:14], rg_3r);
  AND2 I657 (rd_3r1[14:14], dt_0[15:15], rg_3r);
  AND2 I658 (rd_3r1[15:15], dt_0[16:16], rg_3r);
  AND2 I659 (rd_3r1[16:16], dt_0[17:17], rg_3r);
  AND2 I660 (rd_3r1[17:17], dt_0[18:18], rg_3r);
  AND2 I661 (rd_3r1[18:18], dt_0[19:19], rg_3r);
  AND2 I662 (rd_3r1[19:19], dt_0[20:20], rg_3r);
  AND2 I663 (rd_3r1[20:20], dt_0[21:21], rg_3r);
  AND2 I664 (rd_3r1[21:21], dt_0[22:22], rg_3r);
  AND2 I665 (rd_3r1[22:22], dt_0[23:23], rg_3r);
  AND2 I666 (rd_3r1[23:23], dt_0[24:24], rg_3r);
  AND2 I667 (rd_3r1[24:24], dt_0[25:25], rg_3r);
  AND2 I668 (rd_3r1[25:25], dt_0[26:26], rg_3r);
  AND2 I669 (rd_3r1[26:26], dt_0[27:27], rg_3r);
  AND2 I670 (rd_3r1[27:27], dt_0[28:28], rg_3r);
  AND2 I671 (rd_3r1[28:28], dt_0[29:29], rg_3r);
  AND2 I672 (rd_3r1[29:29], dt_0[30:30], rg_3r);
  AND2 I673 (rd_3r1[30:30], dt_0[31:31], rg_3r);
  NOR3 I674 (simp6581_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I675 (simp6581_0[1:1], rg_3r, rg_0a, rg_1a);
  NOR2 I676 (simp6581_0[2:2], rg_2a, rg_3a);
  NAND3 I677 (anyread_0, simp6581_0[0:0], simp6581_0[1:1], simp6581_0[2:2]);
  BUFF I678 (wg_0a, wd_0a);
  BUFF I679 (rg_0a, rd_0a);
  BUFF I680 (rg_1a, rd_1a);
  BUFF I681 (rg_2a, rd_2a);
  BUFF I682 (rg_3a, rd_3a);
endmodule

// tko30m32_1nm2b0_2apt1o0w2bi0w30b TeakO [
//     (1,TeakOConstant 2 0),
//     (2,TeakOAppend 1 [(1,0+:2),(0,0+:30)])] [One 30,One 32]
module tko30m32_1nm2b0_2apt1o0w2bi0w30b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [29:0] i_0r0;
  input [29:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [29:0] gocomp_0;
  wire [9:0] simp321_0;
  wire [3:0] simp322_0;
  wire [1:0] simp323_0;
  wire [1:0] termf_1;
  wire [1:0] termt_1;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  C3 I30 (simp321_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  C3 I31 (simp321_0[1:1], gocomp_0[3:3], gocomp_0[4:4], gocomp_0[5:5]);
  C3 I32 (simp321_0[2:2], gocomp_0[6:6], gocomp_0[7:7], gocomp_0[8:8]);
  C3 I33 (simp321_0[3:3], gocomp_0[9:9], gocomp_0[10:10], gocomp_0[11:11]);
  C3 I34 (simp321_0[4:4], gocomp_0[12:12], gocomp_0[13:13], gocomp_0[14:14]);
  C3 I35 (simp321_0[5:5], gocomp_0[15:15], gocomp_0[16:16], gocomp_0[17:17]);
  C3 I36 (simp321_0[6:6], gocomp_0[18:18], gocomp_0[19:19], gocomp_0[20:20]);
  C3 I37 (simp321_0[7:7], gocomp_0[21:21], gocomp_0[22:22], gocomp_0[23:23]);
  C3 I38 (simp321_0[8:8], gocomp_0[24:24], gocomp_0[25:25], gocomp_0[26:26]);
  C3 I39 (simp321_0[9:9], gocomp_0[27:27], gocomp_0[28:28], gocomp_0[29:29]);
  C3 I40 (simp322_0[0:0], simp321_0[0:0], simp321_0[1:1], simp321_0[2:2]);
  C3 I41 (simp322_0[1:1], simp321_0[3:3], simp321_0[4:4], simp321_0[5:5]);
  C3 I42 (simp322_0[2:2], simp321_0[6:6], simp321_0[7:7], simp321_0[8:8]);
  BUFF I43 (simp322_0[3:3], simp321_0[9:9]);
  C3 I44 (simp323_0[0:0], simp322_0[0:0], simp322_0[1:1], simp322_0[2:2]);
  BUFF I45 (simp323_0[1:1], simp322_0[3:3]);
  C2 I46 (go_0, simp323_0[0:0], simp323_0[1:1]);
  BUFF I47 (termf_1[0:0], go_0);
  BUFF I48 (termf_1[1:1], go_0);
  GND I49 (termt_1[0:0]);
  GND I50 (termt_1[1:1]);
  BUFF I51 (o_0r0[0:0], termf_1[0:0]);
  BUFF I52 (o_0r0[1:1], termf_1[1:1]);
  BUFF I53 (o_0r0[2:2], i_0r0[0:0]);
  BUFF I54 (o_0r0[3:3], i_0r0[1:1]);
  BUFF I55 (o_0r0[4:4], i_0r0[2:2]);
  BUFF I56 (o_0r0[5:5], i_0r0[3:3]);
  BUFF I57 (o_0r0[6:6], i_0r0[4:4]);
  BUFF I58 (o_0r0[7:7], i_0r0[5:5]);
  BUFF I59 (o_0r0[8:8], i_0r0[6:6]);
  BUFF I60 (o_0r0[9:9], i_0r0[7:7]);
  BUFF I61 (o_0r0[10:10], i_0r0[8:8]);
  BUFF I62 (o_0r0[11:11], i_0r0[9:9]);
  BUFF I63 (o_0r0[12:12], i_0r0[10:10]);
  BUFF I64 (o_0r0[13:13], i_0r0[11:11]);
  BUFF I65 (o_0r0[14:14], i_0r0[12:12]);
  BUFF I66 (o_0r0[15:15], i_0r0[13:13]);
  BUFF I67 (o_0r0[16:16], i_0r0[14:14]);
  BUFF I68 (o_0r0[17:17], i_0r0[15:15]);
  BUFF I69 (o_0r0[18:18], i_0r0[16:16]);
  BUFF I70 (o_0r0[19:19], i_0r0[17:17]);
  BUFF I71 (o_0r0[20:20], i_0r0[18:18]);
  BUFF I72 (o_0r0[21:21], i_0r0[19:19]);
  BUFF I73 (o_0r0[22:22], i_0r0[20:20]);
  BUFF I74 (o_0r0[23:23], i_0r0[21:21]);
  BUFF I75 (o_0r0[24:24], i_0r0[22:22]);
  BUFF I76 (o_0r0[25:25], i_0r0[23:23]);
  BUFF I77 (o_0r0[26:26], i_0r0[24:24]);
  BUFF I78 (o_0r0[27:27], i_0r0[25:25]);
  BUFF I79 (o_0r0[28:28], i_0r0[26:26]);
  BUFF I80 (o_0r0[29:29], i_0r0[27:27]);
  BUFF I81 (o_0r0[30:30], i_0r0[28:28]);
  BUFF I82 (o_0r0[31:31], i_0r0[29:29]);
  BUFF I83 (o_0r1[0:0], termt_1[0:0]);
  BUFF I84 (o_0r1[1:1], termt_1[1:1]);
  BUFF I85 (o_0r1[2:2], i_0r1[0:0]);
  BUFF I86 (o_0r1[3:3], i_0r1[1:1]);
  BUFF I87 (o_0r1[4:4], i_0r1[2:2]);
  BUFF I88 (o_0r1[5:5], i_0r1[3:3]);
  BUFF I89 (o_0r1[6:6], i_0r1[4:4]);
  BUFF I90 (o_0r1[7:7], i_0r1[5:5]);
  BUFF I91 (o_0r1[8:8], i_0r1[6:6]);
  BUFF I92 (o_0r1[9:9], i_0r1[7:7]);
  BUFF I93 (o_0r1[10:10], i_0r1[8:8]);
  BUFF I94 (o_0r1[11:11], i_0r1[9:9]);
  BUFF I95 (o_0r1[12:12], i_0r1[10:10]);
  BUFF I96 (o_0r1[13:13], i_0r1[11:11]);
  BUFF I97 (o_0r1[14:14], i_0r1[12:12]);
  BUFF I98 (o_0r1[15:15], i_0r1[13:13]);
  BUFF I99 (o_0r1[16:16], i_0r1[14:14]);
  BUFF I100 (o_0r1[17:17], i_0r1[15:15]);
  BUFF I101 (o_0r1[18:18], i_0r1[16:16]);
  BUFF I102 (o_0r1[19:19], i_0r1[17:17]);
  BUFF I103 (o_0r1[20:20], i_0r1[18:18]);
  BUFF I104 (o_0r1[21:21], i_0r1[19:19]);
  BUFF I105 (o_0r1[22:22], i_0r1[20:20]);
  BUFF I106 (o_0r1[23:23], i_0r1[21:21]);
  BUFF I107 (o_0r1[24:24], i_0r1[22:22]);
  BUFF I108 (o_0r1[25:25], i_0r1[23:23]);
  BUFF I109 (o_0r1[26:26], i_0r1[24:24]);
  BUFF I110 (o_0r1[27:27], i_0r1[25:25]);
  BUFF I111 (o_0r1[28:28], i_0r1[26:26]);
  BUFF I112 (o_0r1[29:29], i_0r1[27:27]);
  BUFF I113 (o_0r1[30:30], i_0r1[28:28]);
  BUFF I114 (o_0r1[31:31], i_0r1[29:29]);
  BUFF I115 (i_0a, o_0a);
endmodule

// tko30m32_1nm2b0_2api0w30bt1o0w2b TeakO [
//     (1,TeakOConstant 2 0),
//     (2,TeakOAppend 1 [(0,0+:30),(1,0+:2)])] [One 30,One 32]
module tko30m32_1nm2b0_2api0w30bt1o0w2b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [29:0] i_0r0;
  input [29:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [29:0] gocomp_0;
  wire [9:0] simp321_0;
  wire [3:0] simp322_0;
  wire [1:0] simp323_0;
  wire [1:0] termf_1;
  wire [1:0] termt_1;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  C3 I30 (simp321_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  C3 I31 (simp321_0[1:1], gocomp_0[3:3], gocomp_0[4:4], gocomp_0[5:5]);
  C3 I32 (simp321_0[2:2], gocomp_0[6:6], gocomp_0[7:7], gocomp_0[8:8]);
  C3 I33 (simp321_0[3:3], gocomp_0[9:9], gocomp_0[10:10], gocomp_0[11:11]);
  C3 I34 (simp321_0[4:4], gocomp_0[12:12], gocomp_0[13:13], gocomp_0[14:14]);
  C3 I35 (simp321_0[5:5], gocomp_0[15:15], gocomp_0[16:16], gocomp_0[17:17]);
  C3 I36 (simp321_0[6:6], gocomp_0[18:18], gocomp_0[19:19], gocomp_0[20:20]);
  C3 I37 (simp321_0[7:7], gocomp_0[21:21], gocomp_0[22:22], gocomp_0[23:23]);
  C3 I38 (simp321_0[8:8], gocomp_0[24:24], gocomp_0[25:25], gocomp_0[26:26]);
  C3 I39 (simp321_0[9:9], gocomp_0[27:27], gocomp_0[28:28], gocomp_0[29:29]);
  C3 I40 (simp322_0[0:0], simp321_0[0:0], simp321_0[1:1], simp321_0[2:2]);
  C3 I41 (simp322_0[1:1], simp321_0[3:3], simp321_0[4:4], simp321_0[5:5]);
  C3 I42 (simp322_0[2:2], simp321_0[6:6], simp321_0[7:7], simp321_0[8:8]);
  BUFF I43 (simp322_0[3:3], simp321_0[9:9]);
  C3 I44 (simp323_0[0:0], simp322_0[0:0], simp322_0[1:1], simp322_0[2:2]);
  BUFF I45 (simp323_0[1:1], simp322_0[3:3]);
  C2 I46 (go_0, simp323_0[0:0], simp323_0[1:1]);
  BUFF I47 (termf_1[0:0], go_0);
  BUFF I48 (termf_1[1:1], go_0);
  GND I49 (termt_1[0:0]);
  GND I50 (termt_1[1:1]);
  BUFF I51 (o_0r0[0:0], i_0r0[0:0]);
  BUFF I52 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I53 (o_0r0[2:2], i_0r0[2:2]);
  BUFF I54 (o_0r0[3:3], i_0r0[3:3]);
  BUFF I55 (o_0r0[4:4], i_0r0[4:4]);
  BUFF I56 (o_0r0[5:5], i_0r0[5:5]);
  BUFF I57 (o_0r0[6:6], i_0r0[6:6]);
  BUFF I58 (o_0r0[7:7], i_0r0[7:7]);
  BUFF I59 (o_0r0[8:8], i_0r0[8:8]);
  BUFF I60 (o_0r0[9:9], i_0r0[9:9]);
  BUFF I61 (o_0r0[10:10], i_0r0[10:10]);
  BUFF I62 (o_0r0[11:11], i_0r0[11:11]);
  BUFF I63 (o_0r0[12:12], i_0r0[12:12]);
  BUFF I64 (o_0r0[13:13], i_0r0[13:13]);
  BUFF I65 (o_0r0[14:14], i_0r0[14:14]);
  BUFF I66 (o_0r0[15:15], i_0r0[15:15]);
  BUFF I67 (o_0r0[16:16], i_0r0[16:16]);
  BUFF I68 (o_0r0[17:17], i_0r0[17:17]);
  BUFF I69 (o_0r0[18:18], i_0r0[18:18]);
  BUFF I70 (o_0r0[19:19], i_0r0[19:19]);
  BUFF I71 (o_0r0[20:20], i_0r0[20:20]);
  BUFF I72 (o_0r0[21:21], i_0r0[21:21]);
  BUFF I73 (o_0r0[22:22], i_0r0[22:22]);
  BUFF I74 (o_0r0[23:23], i_0r0[23:23]);
  BUFF I75 (o_0r0[24:24], i_0r0[24:24]);
  BUFF I76 (o_0r0[25:25], i_0r0[25:25]);
  BUFF I77 (o_0r0[26:26], i_0r0[26:26]);
  BUFF I78 (o_0r0[27:27], i_0r0[27:27]);
  BUFF I79 (o_0r0[28:28], i_0r0[28:28]);
  BUFF I80 (o_0r0[29:29], i_0r0[29:29]);
  BUFF I81 (o_0r0[30:30], termf_1[0:0]);
  BUFF I82 (o_0r0[31:31], termf_1[1:1]);
  BUFF I83 (o_0r1[0:0], i_0r1[0:0]);
  BUFF I84 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I85 (o_0r1[2:2], i_0r1[2:2]);
  BUFF I86 (o_0r1[3:3], i_0r1[3:3]);
  BUFF I87 (o_0r1[4:4], i_0r1[4:4]);
  BUFF I88 (o_0r1[5:5], i_0r1[5:5]);
  BUFF I89 (o_0r1[6:6], i_0r1[6:6]);
  BUFF I90 (o_0r1[7:7], i_0r1[7:7]);
  BUFF I91 (o_0r1[8:8], i_0r1[8:8]);
  BUFF I92 (o_0r1[9:9], i_0r1[9:9]);
  BUFF I93 (o_0r1[10:10], i_0r1[10:10]);
  BUFF I94 (o_0r1[11:11], i_0r1[11:11]);
  BUFF I95 (o_0r1[12:12], i_0r1[12:12]);
  BUFF I96 (o_0r1[13:13], i_0r1[13:13]);
  BUFF I97 (o_0r1[14:14], i_0r1[14:14]);
  BUFF I98 (o_0r1[15:15], i_0r1[15:15]);
  BUFF I99 (o_0r1[16:16], i_0r1[16:16]);
  BUFF I100 (o_0r1[17:17], i_0r1[17:17]);
  BUFF I101 (o_0r1[18:18], i_0r1[18:18]);
  BUFF I102 (o_0r1[19:19], i_0r1[19:19]);
  BUFF I103 (o_0r1[20:20], i_0r1[20:20]);
  BUFF I104 (o_0r1[21:21], i_0r1[21:21]);
  BUFF I105 (o_0r1[22:22], i_0r1[22:22]);
  BUFF I106 (o_0r1[23:23], i_0r1[23:23]);
  BUFF I107 (o_0r1[24:24], i_0r1[24:24]);
  BUFF I108 (o_0r1[25:25], i_0r1[25:25]);
  BUFF I109 (o_0r1[26:26], i_0r1[26:26]);
  BUFF I110 (o_0r1[27:27], i_0r1[27:27]);
  BUFF I111 (o_0r1[28:28], i_0r1[28:28]);
  BUFF I112 (o_0r1[29:29], i_0r1[29:29]);
  BUFF I113 (o_0r1[30:30], termt_1[0:0]);
  BUFF I114 (o_0r1[31:31], termt_1[1:1]);
  BUFF I115 (i_0a, o_0a);
endmodule

// tko30m32_1nm2b3_2api0w30bt1o0w2b TeakO [
//     (1,TeakOConstant 2 3),
//     (2,TeakOAppend 1 [(0,0+:30),(1,0+:2)])] [One 30,One 32]
module tko30m32_1nm2b3_2api0w30bt1o0w2b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [29:0] i_0r0;
  input [29:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [29:0] gocomp_0;
  wire [9:0] simp321_0;
  wire [3:0] simp322_0;
  wire [1:0] simp323_0;
  wire [1:0] termf_1;
  wire [1:0] termt_1;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  C3 I30 (simp321_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  C3 I31 (simp321_0[1:1], gocomp_0[3:3], gocomp_0[4:4], gocomp_0[5:5]);
  C3 I32 (simp321_0[2:2], gocomp_0[6:6], gocomp_0[7:7], gocomp_0[8:8]);
  C3 I33 (simp321_0[3:3], gocomp_0[9:9], gocomp_0[10:10], gocomp_0[11:11]);
  C3 I34 (simp321_0[4:4], gocomp_0[12:12], gocomp_0[13:13], gocomp_0[14:14]);
  C3 I35 (simp321_0[5:5], gocomp_0[15:15], gocomp_0[16:16], gocomp_0[17:17]);
  C3 I36 (simp321_0[6:6], gocomp_0[18:18], gocomp_0[19:19], gocomp_0[20:20]);
  C3 I37 (simp321_0[7:7], gocomp_0[21:21], gocomp_0[22:22], gocomp_0[23:23]);
  C3 I38 (simp321_0[8:8], gocomp_0[24:24], gocomp_0[25:25], gocomp_0[26:26]);
  C3 I39 (simp321_0[9:9], gocomp_0[27:27], gocomp_0[28:28], gocomp_0[29:29]);
  C3 I40 (simp322_0[0:0], simp321_0[0:0], simp321_0[1:1], simp321_0[2:2]);
  C3 I41 (simp322_0[1:1], simp321_0[3:3], simp321_0[4:4], simp321_0[5:5]);
  C3 I42 (simp322_0[2:2], simp321_0[6:6], simp321_0[7:7], simp321_0[8:8]);
  BUFF I43 (simp322_0[3:3], simp321_0[9:9]);
  C3 I44 (simp323_0[0:0], simp322_0[0:0], simp322_0[1:1], simp322_0[2:2]);
  BUFF I45 (simp323_0[1:1], simp322_0[3:3]);
  C2 I46 (go_0, simp323_0[0:0], simp323_0[1:1]);
  BUFF I47 (termt_1[0:0], go_0);
  BUFF I48 (termt_1[1:1], go_0);
  GND I49 (termf_1[0:0]);
  GND I50 (termf_1[1:1]);
  BUFF I51 (o_0r0[0:0], i_0r0[0:0]);
  BUFF I52 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I53 (o_0r0[2:2], i_0r0[2:2]);
  BUFF I54 (o_0r0[3:3], i_0r0[3:3]);
  BUFF I55 (o_0r0[4:4], i_0r0[4:4]);
  BUFF I56 (o_0r0[5:5], i_0r0[5:5]);
  BUFF I57 (o_0r0[6:6], i_0r0[6:6]);
  BUFF I58 (o_0r0[7:7], i_0r0[7:7]);
  BUFF I59 (o_0r0[8:8], i_0r0[8:8]);
  BUFF I60 (o_0r0[9:9], i_0r0[9:9]);
  BUFF I61 (o_0r0[10:10], i_0r0[10:10]);
  BUFF I62 (o_0r0[11:11], i_0r0[11:11]);
  BUFF I63 (o_0r0[12:12], i_0r0[12:12]);
  BUFF I64 (o_0r0[13:13], i_0r0[13:13]);
  BUFF I65 (o_0r0[14:14], i_0r0[14:14]);
  BUFF I66 (o_0r0[15:15], i_0r0[15:15]);
  BUFF I67 (o_0r0[16:16], i_0r0[16:16]);
  BUFF I68 (o_0r0[17:17], i_0r0[17:17]);
  BUFF I69 (o_0r0[18:18], i_0r0[18:18]);
  BUFF I70 (o_0r0[19:19], i_0r0[19:19]);
  BUFF I71 (o_0r0[20:20], i_0r0[20:20]);
  BUFF I72 (o_0r0[21:21], i_0r0[21:21]);
  BUFF I73 (o_0r0[22:22], i_0r0[22:22]);
  BUFF I74 (o_0r0[23:23], i_0r0[23:23]);
  BUFF I75 (o_0r0[24:24], i_0r0[24:24]);
  BUFF I76 (o_0r0[25:25], i_0r0[25:25]);
  BUFF I77 (o_0r0[26:26], i_0r0[26:26]);
  BUFF I78 (o_0r0[27:27], i_0r0[27:27]);
  BUFF I79 (o_0r0[28:28], i_0r0[28:28]);
  BUFF I80 (o_0r0[29:29], i_0r0[29:29]);
  BUFF I81 (o_0r0[30:30], termf_1[0:0]);
  BUFF I82 (o_0r0[31:31], termf_1[1:1]);
  BUFF I83 (o_0r1[0:0], i_0r1[0:0]);
  BUFF I84 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I85 (o_0r1[2:2], i_0r1[2:2]);
  BUFF I86 (o_0r1[3:3], i_0r1[3:3]);
  BUFF I87 (o_0r1[4:4], i_0r1[4:4]);
  BUFF I88 (o_0r1[5:5], i_0r1[5:5]);
  BUFF I89 (o_0r1[6:6], i_0r1[6:6]);
  BUFF I90 (o_0r1[7:7], i_0r1[7:7]);
  BUFF I91 (o_0r1[8:8], i_0r1[8:8]);
  BUFF I92 (o_0r1[9:9], i_0r1[9:9]);
  BUFF I93 (o_0r1[10:10], i_0r1[10:10]);
  BUFF I94 (o_0r1[11:11], i_0r1[11:11]);
  BUFF I95 (o_0r1[12:12], i_0r1[12:12]);
  BUFF I96 (o_0r1[13:13], i_0r1[13:13]);
  BUFF I97 (o_0r1[14:14], i_0r1[14:14]);
  BUFF I98 (o_0r1[15:15], i_0r1[15:15]);
  BUFF I99 (o_0r1[16:16], i_0r1[16:16]);
  BUFF I100 (o_0r1[17:17], i_0r1[17:17]);
  BUFF I101 (o_0r1[18:18], i_0r1[18:18]);
  BUFF I102 (o_0r1[19:19], i_0r1[19:19]);
  BUFF I103 (o_0r1[20:20], i_0r1[20:20]);
  BUFF I104 (o_0r1[21:21], i_0r1[21:21]);
  BUFF I105 (o_0r1[22:22], i_0r1[22:22]);
  BUFF I106 (o_0r1[23:23], i_0r1[23:23]);
  BUFF I107 (o_0r1[24:24], i_0r1[24:24]);
  BUFF I108 (o_0r1[25:25], i_0r1[25:25]);
  BUFF I109 (o_0r1[26:26], i_0r1[26:26]);
  BUFF I110 (o_0r1[27:27], i_0r1[27:27]);
  BUFF I111 (o_0r1[28:28], i_0r1[28:28]);
  BUFF I112 (o_0r1[29:29], i_0r1[29:29]);
  BUFF I113 (o_0r1[30:30], termt_1[0:0]);
  BUFF I114 (o_0r1[31:31], termt_1[1:1]);
  BUFF I115 (i_0a, o_0a);
endmodule

// tkvi32_wo0w32_ro0w32o0w30o2w30o2w30 TeakV "i" 32 [] [0] [0,0,2,2] [Many [32],Many [0],Many [0,0,0,0]
//   ,Many [32,30,30,30]]
module tkvi32_wo0w32_ro0w32o0w30o2w30o2w30 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [29:0] rd_1r0;
  output [29:0] rd_1r1;
  input rd_1a;
  output [29:0] rd_2r0;
  output [29:0] rd_2r1;
  input rd_2a;
  output [29:0] rd_3r0;
  output [29:0] rd_3r1;
  input rd_3a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [2:0] simp6521_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_2r0[0:0], df_0[2:2], rg_2r);
  AND2 I487 (rd_2r0[1:1], df_0[3:3], rg_2r);
  AND2 I488 (rd_2r0[2:2], df_0[4:4], rg_2r);
  AND2 I489 (rd_2r0[3:3], df_0[5:5], rg_2r);
  AND2 I490 (rd_2r0[4:4], df_0[6:6], rg_2r);
  AND2 I491 (rd_2r0[5:5], df_0[7:7], rg_2r);
  AND2 I492 (rd_2r0[6:6], df_0[8:8], rg_2r);
  AND2 I493 (rd_2r0[7:7], df_0[9:9], rg_2r);
  AND2 I494 (rd_2r0[8:8], df_0[10:10], rg_2r);
  AND2 I495 (rd_2r0[9:9], df_0[11:11], rg_2r);
  AND2 I496 (rd_2r0[10:10], df_0[12:12], rg_2r);
  AND2 I497 (rd_2r0[11:11], df_0[13:13], rg_2r);
  AND2 I498 (rd_2r0[12:12], df_0[14:14], rg_2r);
  AND2 I499 (rd_2r0[13:13], df_0[15:15], rg_2r);
  AND2 I500 (rd_2r0[14:14], df_0[16:16], rg_2r);
  AND2 I501 (rd_2r0[15:15], df_0[17:17], rg_2r);
  AND2 I502 (rd_2r0[16:16], df_0[18:18], rg_2r);
  AND2 I503 (rd_2r0[17:17], df_0[19:19], rg_2r);
  AND2 I504 (rd_2r0[18:18], df_0[20:20], rg_2r);
  AND2 I505 (rd_2r0[19:19], df_0[21:21], rg_2r);
  AND2 I506 (rd_2r0[20:20], df_0[22:22], rg_2r);
  AND2 I507 (rd_2r0[21:21], df_0[23:23], rg_2r);
  AND2 I508 (rd_2r0[22:22], df_0[24:24], rg_2r);
  AND2 I509 (rd_2r0[23:23], df_0[25:25], rg_2r);
  AND2 I510 (rd_2r0[24:24], df_0[26:26], rg_2r);
  AND2 I511 (rd_2r0[25:25], df_0[27:27], rg_2r);
  AND2 I512 (rd_2r0[26:26], df_0[28:28], rg_2r);
  AND2 I513 (rd_2r0[27:27], df_0[29:29], rg_2r);
  AND2 I514 (rd_2r0[28:28], df_0[30:30], rg_2r);
  AND2 I515 (rd_2r0[29:29], df_0[31:31], rg_2r);
  AND2 I516 (rd_3r0[0:0], df_0[2:2], rg_3r);
  AND2 I517 (rd_3r0[1:1], df_0[3:3], rg_3r);
  AND2 I518 (rd_3r0[2:2], df_0[4:4], rg_3r);
  AND2 I519 (rd_3r0[3:3], df_0[5:5], rg_3r);
  AND2 I520 (rd_3r0[4:4], df_0[6:6], rg_3r);
  AND2 I521 (rd_3r0[5:5], df_0[7:7], rg_3r);
  AND2 I522 (rd_3r0[6:6], df_0[8:8], rg_3r);
  AND2 I523 (rd_3r0[7:7], df_0[9:9], rg_3r);
  AND2 I524 (rd_3r0[8:8], df_0[10:10], rg_3r);
  AND2 I525 (rd_3r0[9:9], df_0[11:11], rg_3r);
  AND2 I526 (rd_3r0[10:10], df_0[12:12], rg_3r);
  AND2 I527 (rd_3r0[11:11], df_0[13:13], rg_3r);
  AND2 I528 (rd_3r0[12:12], df_0[14:14], rg_3r);
  AND2 I529 (rd_3r0[13:13], df_0[15:15], rg_3r);
  AND2 I530 (rd_3r0[14:14], df_0[16:16], rg_3r);
  AND2 I531 (rd_3r0[15:15], df_0[17:17], rg_3r);
  AND2 I532 (rd_3r0[16:16], df_0[18:18], rg_3r);
  AND2 I533 (rd_3r0[17:17], df_0[19:19], rg_3r);
  AND2 I534 (rd_3r0[18:18], df_0[20:20], rg_3r);
  AND2 I535 (rd_3r0[19:19], df_0[21:21], rg_3r);
  AND2 I536 (rd_3r0[20:20], df_0[22:22], rg_3r);
  AND2 I537 (rd_3r0[21:21], df_0[23:23], rg_3r);
  AND2 I538 (rd_3r0[22:22], df_0[24:24], rg_3r);
  AND2 I539 (rd_3r0[23:23], df_0[25:25], rg_3r);
  AND2 I540 (rd_3r0[24:24], df_0[26:26], rg_3r);
  AND2 I541 (rd_3r0[25:25], df_0[27:27], rg_3r);
  AND2 I542 (rd_3r0[26:26], df_0[28:28], rg_3r);
  AND2 I543 (rd_3r0[27:27], df_0[29:29], rg_3r);
  AND2 I544 (rd_3r0[28:28], df_0[30:30], rg_3r);
  AND2 I545 (rd_3r0[29:29], df_0[31:31], rg_3r);
  AND2 I546 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I547 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I548 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I549 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I550 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I551 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I552 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I553 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I554 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I555 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I556 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I557 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I558 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I559 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I560 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I561 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I562 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I563 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I564 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I565 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I566 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I567 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I568 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I569 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I570 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I571 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I572 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I573 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I574 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I575 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I576 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I577 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I578 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I579 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I580 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I581 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I582 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I583 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I584 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I585 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I586 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I587 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I588 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I589 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I590 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I591 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I592 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I593 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I594 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I595 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I596 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I597 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I598 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I599 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I600 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I601 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I602 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I603 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I604 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I605 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I606 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I607 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I608 (rd_2r1[0:0], dt_0[2:2], rg_2r);
  AND2 I609 (rd_2r1[1:1], dt_0[3:3], rg_2r);
  AND2 I610 (rd_2r1[2:2], dt_0[4:4], rg_2r);
  AND2 I611 (rd_2r1[3:3], dt_0[5:5], rg_2r);
  AND2 I612 (rd_2r1[4:4], dt_0[6:6], rg_2r);
  AND2 I613 (rd_2r1[5:5], dt_0[7:7], rg_2r);
  AND2 I614 (rd_2r1[6:6], dt_0[8:8], rg_2r);
  AND2 I615 (rd_2r1[7:7], dt_0[9:9], rg_2r);
  AND2 I616 (rd_2r1[8:8], dt_0[10:10], rg_2r);
  AND2 I617 (rd_2r1[9:9], dt_0[11:11], rg_2r);
  AND2 I618 (rd_2r1[10:10], dt_0[12:12], rg_2r);
  AND2 I619 (rd_2r1[11:11], dt_0[13:13], rg_2r);
  AND2 I620 (rd_2r1[12:12], dt_0[14:14], rg_2r);
  AND2 I621 (rd_2r1[13:13], dt_0[15:15], rg_2r);
  AND2 I622 (rd_2r1[14:14], dt_0[16:16], rg_2r);
  AND2 I623 (rd_2r1[15:15], dt_0[17:17], rg_2r);
  AND2 I624 (rd_2r1[16:16], dt_0[18:18], rg_2r);
  AND2 I625 (rd_2r1[17:17], dt_0[19:19], rg_2r);
  AND2 I626 (rd_2r1[18:18], dt_0[20:20], rg_2r);
  AND2 I627 (rd_2r1[19:19], dt_0[21:21], rg_2r);
  AND2 I628 (rd_2r1[20:20], dt_0[22:22], rg_2r);
  AND2 I629 (rd_2r1[21:21], dt_0[23:23], rg_2r);
  AND2 I630 (rd_2r1[22:22], dt_0[24:24], rg_2r);
  AND2 I631 (rd_2r1[23:23], dt_0[25:25], rg_2r);
  AND2 I632 (rd_2r1[24:24], dt_0[26:26], rg_2r);
  AND2 I633 (rd_2r1[25:25], dt_0[27:27], rg_2r);
  AND2 I634 (rd_2r1[26:26], dt_0[28:28], rg_2r);
  AND2 I635 (rd_2r1[27:27], dt_0[29:29], rg_2r);
  AND2 I636 (rd_2r1[28:28], dt_0[30:30], rg_2r);
  AND2 I637 (rd_2r1[29:29], dt_0[31:31], rg_2r);
  AND2 I638 (rd_3r1[0:0], dt_0[2:2], rg_3r);
  AND2 I639 (rd_3r1[1:1], dt_0[3:3], rg_3r);
  AND2 I640 (rd_3r1[2:2], dt_0[4:4], rg_3r);
  AND2 I641 (rd_3r1[3:3], dt_0[5:5], rg_3r);
  AND2 I642 (rd_3r1[4:4], dt_0[6:6], rg_3r);
  AND2 I643 (rd_3r1[5:5], dt_0[7:7], rg_3r);
  AND2 I644 (rd_3r1[6:6], dt_0[8:8], rg_3r);
  AND2 I645 (rd_3r1[7:7], dt_0[9:9], rg_3r);
  AND2 I646 (rd_3r1[8:8], dt_0[10:10], rg_3r);
  AND2 I647 (rd_3r1[9:9], dt_0[11:11], rg_3r);
  AND2 I648 (rd_3r1[10:10], dt_0[12:12], rg_3r);
  AND2 I649 (rd_3r1[11:11], dt_0[13:13], rg_3r);
  AND2 I650 (rd_3r1[12:12], dt_0[14:14], rg_3r);
  AND2 I651 (rd_3r1[13:13], dt_0[15:15], rg_3r);
  AND2 I652 (rd_3r1[14:14], dt_0[16:16], rg_3r);
  AND2 I653 (rd_3r1[15:15], dt_0[17:17], rg_3r);
  AND2 I654 (rd_3r1[16:16], dt_0[18:18], rg_3r);
  AND2 I655 (rd_3r1[17:17], dt_0[19:19], rg_3r);
  AND2 I656 (rd_3r1[18:18], dt_0[20:20], rg_3r);
  AND2 I657 (rd_3r1[19:19], dt_0[21:21], rg_3r);
  AND2 I658 (rd_3r1[20:20], dt_0[22:22], rg_3r);
  AND2 I659 (rd_3r1[21:21], dt_0[23:23], rg_3r);
  AND2 I660 (rd_3r1[22:22], dt_0[24:24], rg_3r);
  AND2 I661 (rd_3r1[23:23], dt_0[25:25], rg_3r);
  AND2 I662 (rd_3r1[24:24], dt_0[26:26], rg_3r);
  AND2 I663 (rd_3r1[25:25], dt_0[27:27], rg_3r);
  AND2 I664 (rd_3r1[26:26], dt_0[28:28], rg_3r);
  AND2 I665 (rd_3r1[27:27], dt_0[29:29], rg_3r);
  AND2 I666 (rd_3r1[28:28], dt_0[30:30], rg_3r);
  AND2 I667 (rd_3r1[29:29], dt_0[31:31], rg_3r);
  NOR3 I668 (simp6521_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I669 (simp6521_0[1:1], rg_3r, rg_0a, rg_1a);
  NOR2 I670 (simp6521_0[2:2], rg_2a, rg_3a);
  NAND3 I671 (anyread_0, simp6521_0[0:0], simp6521_0[1:1], simp6521_0[2:2]);
  BUFF I672 (wg_0a, wd_0a);
  BUFF I673 (rg_0a, rd_0a);
  BUFF I674 (rg_1a, rd_1a);
  BUFF I675 (rg_2a, rd_2a);
  BUFF I676 (rg_3a, rd_3a);
endmodule

// tkj0m0_0_0 TeakJ [Many [0,0,0],One 0]
module tkj0m0_0_0 (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  output o_0r;
  input o_0a;
  input reset;
  C3 I0 (o_0r, i_0r, i_1r, i_2r);
  BUFF I1 (i_0a, o_0a);
  BUFF I2 (i_1a, o_0a);
  BUFF I3 (i_2a, o_0a);
endmodule

// tkm4x32b TeakM [Many [32,32,32,32],One 32]
module tkm4x32b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  input [31:0] i_2r0;
  input [31:0] i_2r1;
  output i_2a;
  input [31:0] i_3r0;
  input [31:0] i_3r1;
  output i_3a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire [31:0] gfint_0;
  wire [31:0] gfint_1;
  wire [31:0] gfint_2;
  wire [31:0] gfint_3;
  wire [31:0] gtint_0;
  wire [31:0] gtint_1;
  wire [31:0] gtint_2;
  wire [31:0] gtint_3;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire icomp_3;
  wire nchosen_0;
  wire [1:0] simp181_0;
  wire [1:0] simp191_0;
  wire [1:0] simp201_0;
  wire [1:0] simp211_0;
  wire [1:0] simp221_0;
  wire [1:0] simp231_0;
  wire [1:0] simp241_0;
  wire [1:0] simp251_0;
  wire [1:0] simp261_0;
  wire [1:0] simp271_0;
  wire [1:0] simp281_0;
  wire [1:0] simp291_0;
  wire [1:0] simp301_0;
  wire [1:0] simp311_0;
  wire [1:0] simp321_0;
  wire [1:0] simp331_0;
  wire [1:0] simp341_0;
  wire [1:0] simp351_0;
  wire [1:0] simp361_0;
  wire [1:0] simp371_0;
  wire [1:0] simp381_0;
  wire [1:0] simp391_0;
  wire [1:0] simp401_0;
  wire [1:0] simp411_0;
  wire [1:0] simp421_0;
  wire [1:0] simp431_0;
  wire [1:0] simp441_0;
  wire [1:0] simp451_0;
  wire [1:0] simp461_0;
  wire [1:0] simp471_0;
  wire [1:0] simp481_0;
  wire [1:0] simp491_0;
  wire [1:0] simp501_0;
  wire [1:0] simp511_0;
  wire [1:0] simp521_0;
  wire [1:0] simp531_0;
  wire [1:0] simp541_0;
  wire [1:0] simp551_0;
  wire [1:0] simp561_0;
  wire [1:0] simp571_0;
  wire [1:0] simp581_0;
  wire [1:0] simp591_0;
  wire [1:0] simp601_0;
  wire [1:0] simp611_0;
  wire [1:0] simp621_0;
  wire [1:0] simp631_0;
  wire [1:0] simp641_0;
  wire [1:0] simp651_0;
  wire [1:0] simp661_0;
  wire [1:0] simp671_0;
  wire [1:0] simp681_0;
  wire [1:0] simp691_0;
  wire [1:0] simp701_0;
  wire [1:0] simp711_0;
  wire [1:0] simp721_0;
  wire [1:0] simp731_0;
  wire [1:0] simp741_0;
  wire [1:0] simp751_0;
  wire [1:0] simp761_0;
  wire [1:0] simp771_0;
  wire [1:0] simp781_0;
  wire [1:0] simp791_0;
  wire [1:0] simp801_0;
  wire [1:0] simp811_0;
  wire [31:0] comp0_0;
  wire [10:0] simp3711_0;
  wire [3:0] simp3712_0;
  wire [1:0] simp3713_0;
  wire [31:0] comp1_0;
  wire [10:0] simp4051_0;
  wire [3:0] simp4052_0;
  wire [1:0] simp4053_0;
  wire [31:0] comp2_0;
  wire [10:0] simp4391_0;
  wire [3:0] simp4392_0;
  wire [1:0] simp4393_0;
  wire [31:0] comp3_0;
  wire [10:0] simp4731_0;
  wire [3:0] simp4732_0;
  wire [1:0] simp4733_0;
  wire [1:0] simp4781_0;
  NOR3 I0 (simp181_0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  INV I1 (simp181_0[1:1], gfint_3[0:0]);
  NAND2 I2 (o_0r0[0:0], simp181_0[0:0], simp181_0[1:1]);
  NOR3 I3 (simp191_0[0:0], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  INV I4 (simp191_0[1:1], gfint_3[1:1]);
  NAND2 I5 (o_0r0[1:1], simp191_0[0:0], simp191_0[1:1]);
  NOR3 I6 (simp201_0[0:0], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  INV I7 (simp201_0[1:1], gfint_3[2:2]);
  NAND2 I8 (o_0r0[2:2], simp201_0[0:0], simp201_0[1:1]);
  NOR3 I9 (simp211_0[0:0], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  INV I10 (simp211_0[1:1], gfint_3[3:3]);
  NAND2 I11 (o_0r0[3:3], simp211_0[0:0], simp211_0[1:1]);
  NOR3 I12 (simp221_0[0:0], gfint_0[4:4], gfint_1[4:4], gfint_2[4:4]);
  INV I13 (simp221_0[1:1], gfint_3[4:4]);
  NAND2 I14 (o_0r0[4:4], simp221_0[0:0], simp221_0[1:1]);
  NOR3 I15 (simp231_0[0:0], gfint_0[5:5], gfint_1[5:5], gfint_2[5:5]);
  INV I16 (simp231_0[1:1], gfint_3[5:5]);
  NAND2 I17 (o_0r0[5:5], simp231_0[0:0], simp231_0[1:1]);
  NOR3 I18 (simp241_0[0:0], gfint_0[6:6], gfint_1[6:6], gfint_2[6:6]);
  INV I19 (simp241_0[1:1], gfint_3[6:6]);
  NAND2 I20 (o_0r0[6:6], simp241_0[0:0], simp241_0[1:1]);
  NOR3 I21 (simp251_0[0:0], gfint_0[7:7], gfint_1[7:7], gfint_2[7:7]);
  INV I22 (simp251_0[1:1], gfint_3[7:7]);
  NAND2 I23 (o_0r0[7:7], simp251_0[0:0], simp251_0[1:1]);
  NOR3 I24 (simp261_0[0:0], gfint_0[8:8], gfint_1[8:8], gfint_2[8:8]);
  INV I25 (simp261_0[1:1], gfint_3[8:8]);
  NAND2 I26 (o_0r0[8:8], simp261_0[0:0], simp261_0[1:1]);
  NOR3 I27 (simp271_0[0:0], gfint_0[9:9], gfint_1[9:9], gfint_2[9:9]);
  INV I28 (simp271_0[1:1], gfint_3[9:9]);
  NAND2 I29 (o_0r0[9:9], simp271_0[0:0], simp271_0[1:1]);
  NOR3 I30 (simp281_0[0:0], gfint_0[10:10], gfint_1[10:10], gfint_2[10:10]);
  INV I31 (simp281_0[1:1], gfint_3[10:10]);
  NAND2 I32 (o_0r0[10:10], simp281_0[0:0], simp281_0[1:1]);
  NOR3 I33 (simp291_0[0:0], gfint_0[11:11], gfint_1[11:11], gfint_2[11:11]);
  INV I34 (simp291_0[1:1], gfint_3[11:11]);
  NAND2 I35 (o_0r0[11:11], simp291_0[0:0], simp291_0[1:1]);
  NOR3 I36 (simp301_0[0:0], gfint_0[12:12], gfint_1[12:12], gfint_2[12:12]);
  INV I37 (simp301_0[1:1], gfint_3[12:12]);
  NAND2 I38 (o_0r0[12:12], simp301_0[0:0], simp301_0[1:1]);
  NOR3 I39 (simp311_0[0:0], gfint_0[13:13], gfint_1[13:13], gfint_2[13:13]);
  INV I40 (simp311_0[1:1], gfint_3[13:13]);
  NAND2 I41 (o_0r0[13:13], simp311_0[0:0], simp311_0[1:1]);
  NOR3 I42 (simp321_0[0:0], gfint_0[14:14], gfint_1[14:14], gfint_2[14:14]);
  INV I43 (simp321_0[1:1], gfint_3[14:14]);
  NAND2 I44 (o_0r0[14:14], simp321_0[0:0], simp321_0[1:1]);
  NOR3 I45 (simp331_0[0:0], gfint_0[15:15], gfint_1[15:15], gfint_2[15:15]);
  INV I46 (simp331_0[1:1], gfint_3[15:15]);
  NAND2 I47 (o_0r0[15:15], simp331_0[0:0], simp331_0[1:1]);
  NOR3 I48 (simp341_0[0:0], gfint_0[16:16], gfint_1[16:16], gfint_2[16:16]);
  INV I49 (simp341_0[1:1], gfint_3[16:16]);
  NAND2 I50 (o_0r0[16:16], simp341_0[0:0], simp341_0[1:1]);
  NOR3 I51 (simp351_0[0:0], gfint_0[17:17], gfint_1[17:17], gfint_2[17:17]);
  INV I52 (simp351_0[1:1], gfint_3[17:17]);
  NAND2 I53 (o_0r0[17:17], simp351_0[0:0], simp351_0[1:1]);
  NOR3 I54 (simp361_0[0:0], gfint_0[18:18], gfint_1[18:18], gfint_2[18:18]);
  INV I55 (simp361_0[1:1], gfint_3[18:18]);
  NAND2 I56 (o_0r0[18:18], simp361_0[0:0], simp361_0[1:1]);
  NOR3 I57 (simp371_0[0:0], gfint_0[19:19], gfint_1[19:19], gfint_2[19:19]);
  INV I58 (simp371_0[1:1], gfint_3[19:19]);
  NAND2 I59 (o_0r0[19:19], simp371_0[0:0], simp371_0[1:1]);
  NOR3 I60 (simp381_0[0:0], gfint_0[20:20], gfint_1[20:20], gfint_2[20:20]);
  INV I61 (simp381_0[1:1], gfint_3[20:20]);
  NAND2 I62 (o_0r0[20:20], simp381_0[0:0], simp381_0[1:1]);
  NOR3 I63 (simp391_0[0:0], gfint_0[21:21], gfint_1[21:21], gfint_2[21:21]);
  INV I64 (simp391_0[1:1], gfint_3[21:21]);
  NAND2 I65 (o_0r0[21:21], simp391_0[0:0], simp391_0[1:1]);
  NOR3 I66 (simp401_0[0:0], gfint_0[22:22], gfint_1[22:22], gfint_2[22:22]);
  INV I67 (simp401_0[1:1], gfint_3[22:22]);
  NAND2 I68 (o_0r0[22:22], simp401_0[0:0], simp401_0[1:1]);
  NOR3 I69 (simp411_0[0:0], gfint_0[23:23], gfint_1[23:23], gfint_2[23:23]);
  INV I70 (simp411_0[1:1], gfint_3[23:23]);
  NAND2 I71 (o_0r0[23:23], simp411_0[0:0], simp411_0[1:1]);
  NOR3 I72 (simp421_0[0:0], gfint_0[24:24], gfint_1[24:24], gfint_2[24:24]);
  INV I73 (simp421_0[1:1], gfint_3[24:24]);
  NAND2 I74 (o_0r0[24:24], simp421_0[0:0], simp421_0[1:1]);
  NOR3 I75 (simp431_0[0:0], gfint_0[25:25], gfint_1[25:25], gfint_2[25:25]);
  INV I76 (simp431_0[1:1], gfint_3[25:25]);
  NAND2 I77 (o_0r0[25:25], simp431_0[0:0], simp431_0[1:1]);
  NOR3 I78 (simp441_0[0:0], gfint_0[26:26], gfint_1[26:26], gfint_2[26:26]);
  INV I79 (simp441_0[1:1], gfint_3[26:26]);
  NAND2 I80 (o_0r0[26:26], simp441_0[0:0], simp441_0[1:1]);
  NOR3 I81 (simp451_0[0:0], gfint_0[27:27], gfint_1[27:27], gfint_2[27:27]);
  INV I82 (simp451_0[1:1], gfint_3[27:27]);
  NAND2 I83 (o_0r0[27:27], simp451_0[0:0], simp451_0[1:1]);
  NOR3 I84 (simp461_0[0:0], gfint_0[28:28], gfint_1[28:28], gfint_2[28:28]);
  INV I85 (simp461_0[1:1], gfint_3[28:28]);
  NAND2 I86 (o_0r0[28:28], simp461_0[0:0], simp461_0[1:1]);
  NOR3 I87 (simp471_0[0:0], gfint_0[29:29], gfint_1[29:29], gfint_2[29:29]);
  INV I88 (simp471_0[1:1], gfint_3[29:29]);
  NAND2 I89 (o_0r0[29:29], simp471_0[0:0], simp471_0[1:1]);
  NOR3 I90 (simp481_0[0:0], gfint_0[30:30], gfint_1[30:30], gfint_2[30:30]);
  INV I91 (simp481_0[1:1], gfint_3[30:30]);
  NAND2 I92 (o_0r0[30:30], simp481_0[0:0], simp481_0[1:1]);
  NOR3 I93 (simp491_0[0:0], gfint_0[31:31], gfint_1[31:31], gfint_2[31:31]);
  INV I94 (simp491_0[1:1], gfint_3[31:31]);
  NAND2 I95 (o_0r0[31:31], simp491_0[0:0], simp491_0[1:1]);
  NOR3 I96 (simp501_0[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  INV I97 (simp501_0[1:1], gtint_3[0:0]);
  NAND2 I98 (o_0r1[0:0], simp501_0[0:0], simp501_0[1:1]);
  NOR3 I99 (simp511_0[0:0], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  INV I100 (simp511_0[1:1], gtint_3[1:1]);
  NAND2 I101 (o_0r1[1:1], simp511_0[0:0], simp511_0[1:1]);
  NOR3 I102 (simp521_0[0:0], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  INV I103 (simp521_0[1:1], gtint_3[2:2]);
  NAND2 I104 (o_0r1[2:2], simp521_0[0:0], simp521_0[1:1]);
  NOR3 I105 (simp531_0[0:0], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  INV I106 (simp531_0[1:1], gtint_3[3:3]);
  NAND2 I107 (o_0r1[3:3], simp531_0[0:0], simp531_0[1:1]);
  NOR3 I108 (simp541_0[0:0], gtint_0[4:4], gtint_1[4:4], gtint_2[4:4]);
  INV I109 (simp541_0[1:1], gtint_3[4:4]);
  NAND2 I110 (o_0r1[4:4], simp541_0[0:0], simp541_0[1:1]);
  NOR3 I111 (simp551_0[0:0], gtint_0[5:5], gtint_1[5:5], gtint_2[5:5]);
  INV I112 (simp551_0[1:1], gtint_3[5:5]);
  NAND2 I113 (o_0r1[5:5], simp551_0[0:0], simp551_0[1:1]);
  NOR3 I114 (simp561_0[0:0], gtint_0[6:6], gtint_1[6:6], gtint_2[6:6]);
  INV I115 (simp561_0[1:1], gtint_3[6:6]);
  NAND2 I116 (o_0r1[6:6], simp561_0[0:0], simp561_0[1:1]);
  NOR3 I117 (simp571_0[0:0], gtint_0[7:7], gtint_1[7:7], gtint_2[7:7]);
  INV I118 (simp571_0[1:1], gtint_3[7:7]);
  NAND2 I119 (o_0r1[7:7], simp571_0[0:0], simp571_0[1:1]);
  NOR3 I120 (simp581_0[0:0], gtint_0[8:8], gtint_1[8:8], gtint_2[8:8]);
  INV I121 (simp581_0[1:1], gtint_3[8:8]);
  NAND2 I122 (o_0r1[8:8], simp581_0[0:0], simp581_0[1:1]);
  NOR3 I123 (simp591_0[0:0], gtint_0[9:9], gtint_1[9:9], gtint_2[9:9]);
  INV I124 (simp591_0[1:1], gtint_3[9:9]);
  NAND2 I125 (o_0r1[9:9], simp591_0[0:0], simp591_0[1:1]);
  NOR3 I126 (simp601_0[0:0], gtint_0[10:10], gtint_1[10:10], gtint_2[10:10]);
  INV I127 (simp601_0[1:1], gtint_3[10:10]);
  NAND2 I128 (o_0r1[10:10], simp601_0[0:0], simp601_0[1:1]);
  NOR3 I129 (simp611_0[0:0], gtint_0[11:11], gtint_1[11:11], gtint_2[11:11]);
  INV I130 (simp611_0[1:1], gtint_3[11:11]);
  NAND2 I131 (o_0r1[11:11], simp611_0[0:0], simp611_0[1:1]);
  NOR3 I132 (simp621_0[0:0], gtint_0[12:12], gtint_1[12:12], gtint_2[12:12]);
  INV I133 (simp621_0[1:1], gtint_3[12:12]);
  NAND2 I134 (o_0r1[12:12], simp621_0[0:0], simp621_0[1:1]);
  NOR3 I135 (simp631_0[0:0], gtint_0[13:13], gtint_1[13:13], gtint_2[13:13]);
  INV I136 (simp631_0[1:1], gtint_3[13:13]);
  NAND2 I137 (o_0r1[13:13], simp631_0[0:0], simp631_0[1:1]);
  NOR3 I138 (simp641_0[0:0], gtint_0[14:14], gtint_1[14:14], gtint_2[14:14]);
  INV I139 (simp641_0[1:1], gtint_3[14:14]);
  NAND2 I140 (o_0r1[14:14], simp641_0[0:0], simp641_0[1:1]);
  NOR3 I141 (simp651_0[0:0], gtint_0[15:15], gtint_1[15:15], gtint_2[15:15]);
  INV I142 (simp651_0[1:1], gtint_3[15:15]);
  NAND2 I143 (o_0r1[15:15], simp651_0[0:0], simp651_0[1:1]);
  NOR3 I144 (simp661_0[0:0], gtint_0[16:16], gtint_1[16:16], gtint_2[16:16]);
  INV I145 (simp661_0[1:1], gtint_3[16:16]);
  NAND2 I146 (o_0r1[16:16], simp661_0[0:0], simp661_0[1:1]);
  NOR3 I147 (simp671_0[0:0], gtint_0[17:17], gtint_1[17:17], gtint_2[17:17]);
  INV I148 (simp671_0[1:1], gtint_3[17:17]);
  NAND2 I149 (o_0r1[17:17], simp671_0[0:0], simp671_0[1:1]);
  NOR3 I150 (simp681_0[0:0], gtint_0[18:18], gtint_1[18:18], gtint_2[18:18]);
  INV I151 (simp681_0[1:1], gtint_3[18:18]);
  NAND2 I152 (o_0r1[18:18], simp681_0[0:0], simp681_0[1:1]);
  NOR3 I153 (simp691_0[0:0], gtint_0[19:19], gtint_1[19:19], gtint_2[19:19]);
  INV I154 (simp691_0[1:1], gtint_3[19:19]);
  NAND2 I155 (o_0r1[19:19], simp691_0[0:0], simp691_0[1:1]);
  NOR3 I156 (simp701_0[0:0], gtint_0[20:20], gtint_1[20:20], gtint_2[20:20]);
  INV I157 (simp701_0[1:1], gtint_3[20:20]);
  NAND2 I158 (o_0r1[20:20], simp701_0[0:0], simp701_0[1:1]);
  NOR3 I159 (simp711_0[0:0], gtint_0[21:21], gtint_1[21:21], gtint_2[21:21]);
  INV I160 (simp711_0[1:1], gtint_3[21:21]);
  NAND2 I161 (o_0r1[21:21], simp711_0[0:0], simp711_0[1:1]);
  NOR3 I162 (simp721_0[0:0], gtint_0[22:22], gtint_1[22:22], gtint_2[22:22]);
  INV I163 (simp721_0[1:1], gtint_3[22:22]);
  NAND2 I164 (o_0r1[22:22], simp721_0[0:0], simp721_0[1:1]);
  NOR3 I165 (simp731_0[0:0], gtint_0[23:23], gtint_1[23:23], gtint_2[23:23]);
  INV I166 (simp731_0[1:1], gtint_3[23:23]);
  NAND2 I167 (o_0r1[23:23], simp731_0[0:0], simp731_0[1:1]);
  NOR3 I168 (simp741_0[0:0], gtint_0[24:24], gtint_1[24:24], gtint_2[24:24]);
  INV I169 (simp741_0[1:1], gtint_3[24:24]);
  NAND2 I170 (o_0r1[24:24], simp741_0[0:0], simp741_0[1:1]);
  NOR3 I171 (simp751_0[0:0], gtint_0[25:25], gtint_1[25:25], gtint_2[25:25]);
  INV I172 (simp751_0[1:1], gtint_3[25:25]);
  NAND2 I173 (o_0r1[25:25], simp751_0[0:0], simp751_0[1:1]);
  NOR3 I174 (simp761_0[0:0], gtint_0[26:26], gtint_1[26:26], gtint_2[26:26]);
  INV I175 (simp761_0[1:1], gtint_3[26:26]);
  NAND2 I176 (o_0r1[26:26], simp761_0[0:0], simp761_0[1:1]);
  NOR3 I177 (simp771_0[0:0], gtint_0[27:27], gtint_1[27:27], gtint_2[27:27]);
  INV I178 (simp771_0[1:1], gtint_3[27:27]);
  NAND2 I179 (o_0r1[27:27], simp771_0[0:0], simp771_0[1:1]);
  NOR3 I180 (simp781_0[0:0], gtint_0[28:28], gtint_1[28:28], gtint_2[28:28]);
  INV I181 (simp781_0[1:1], gtint_3[28:28]);
  NAND2 I182 (o_0r1[28:28], simp781_0[0:0], simp781_0[1:1]);
  NOR3 I183 (simp791_0[0:0], gtint_0[29:29], gtint_1[29:29], gtint_2[29:29]);
  INV I184 (simp791_0[1:1], gtint_3[29:29]);
  NAND2 I185 (o_0r1[29:29], simp791_0[0:0], simp791_0[1:1]);
  NOR3 I186 (simp801_0[0:0], gtint_0[30:30], gtint_1[30:30], gtint_2[30:30]);
  INV I187 (simp801_0[1:1], gtint_3[30:30]);
  NAND2 I188 (o_0r1[30:30], simp801_0[0:0], simp801_0[1:1]);
  NOR3 I189 (simp811_0[0:0], gtint_0[31:31], gtint_1[31:31], gtint_2[31:31]);
  INV I190 (simp811_0[1:1], gtint_3[31:31]);
  NAND2 I191 (o_0r1[31:31], simp811_0[0:0], simp811_0[1:1]);
  AND2 I192 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I193 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I194 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I195 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I196 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I197 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I198 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I199 (gtint_0[7:7], choice_0, i_0r1[7:7]);
  AND2 I200 (gtint_0[8:8], choice_0, i_0r1[8:8]);
  AND2 I201 (gtint_0[9:9], choice_0, i_0r1[9:9]);
  AND2 I202 (gtint_0[10:10], choice_0, i_0r1[10:10]);
  AND2 I203 (gtint_0[11:11], choice_0, i_0r1[11:11]);
  AND2 I204 (gtint_0[12:12], choice_0, i_0r1[12:12]);
  AND2 I205 (gtint_0[13:13], choice_0, i_0r1[13:13]);
  AND2 I206 (gtint_0[14:14], choice_0, i_0r1[14:14]);
  AND2 I207 (gtint_0[15:15], choice_0, i_0r1[15:15]);
  AND2 I208 (gtint_0[16:16], choice_0, i_0r1[16:16]);
  AND2 I209 (gtint_0[17:17], choice_0, i_0r1[17:17]);
  AND2 I210 (gtint_0[18:18], choice_0, i_0r1[18:18]);
  AND2 I211 (gtint_0[19:19], choice_0, i_0r1[19:19]);
  AND2 I212 (gtint_0[20:20], choice_0, i_0r1[20:20]);
  AND2 I213 (gtint_0[21:21], choice_0, i_0r1[21:21]);
  AND2 I214 (gtint_0[22:22], choice_0, i_0r1[22:22]);
  AND2 I215 (gtint_0[23:23], choice_0, i_0r1[23:23]);
  AND2 I216 (gtint_0[24:24], choice_0, i_0r1[24:24]);
  AND2 I217 (gtint_0[25:25], choice_0, i_0r1[25:25]);
  AND2 I218 (gtint_0[26:26], choice_0, i_0r1[26:26]);
  AND2 I219 (gtint_0[27:27], choice_0, i_0r1[27:27]);
  AND2 I220 (gtint_0[28:28], choice_0, i_0r1[28:28]);
  AND2 I221 (gtint_0[29:29], choice_0, i_0r1[29:29]);
  AND2 I222 (gtint_0[30:30], choice_0, i_0r1[30:30]);
  AND2 I223 (gtint_0[31:31], choice_0, i_0r1[31:31]);
  AND2 I224 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I225 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I226 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I227 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I228 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I229 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I230 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I231 (gtint_1[7:7], choice_1, i_1r1[7:7]);
  AND2 I232 (gtint_1[8:8], choice_1, i_1r1[8:8]);
  AND2 I233 (gtint_1[9:9], choice_1, i_1r1[9:9]);
  AND2 I234 (gtint_1[10:10], choice_1, i_1r1[10:10]);
  AND2 I235 (gtint_1[11:11], choice_1, i_1r1[11:11]);
  AND2 I236 (gtint_1[12:12], choice_1, i_1r1[12:12]);
  AND2 I237 (gtint_1[13:13], choice_1, i_1r1[13:13]);
  AND2 I238 (gtint_1[14:14], choice_1, i_1r1[14:14]);
  AND2 I239 (gtint_1[15:15], choice_1, i_1r1[15:15]);
  AND2 I240 (gtint_1[16:16], choice_1, i_1r1[16:16]);
  AND2 I241 (gtint_1[17:17], choice_1, i_1r1[17:17]);
  AND2 I242 (gtint_1[18:18], choice_1, i_1r1[18:18]);
  AND2 I243 (gtint_1[19:19], choice_1, i_1r1[19:19]);
  AND2 I244 (gtint_1[20:20], choice_1, i_1r1[20:20]);
  AND2 I245 (gtint_1[21:21], choice_1, i_1r1[21:21]);
  AND2 I246 (gtint_1[22:22], choice_1, i_1r1[22:22]);
  AND2 I247 (gtint_1[23:23], choice_1, i_1r1[23:23]);
  AND2 I248 (gtint_1[24:24], choice_1, i_1r1[24:24]);
  AND2 I249 (gtint_1[25:25], choice_1, i_1r1[25:25]);
  AND2 I250 (gtint_1[26:26], choice_1, i_1r1[26:26]);
  AND2 I251 (gtint_1[27:27], choice_1, i_1r1[27:27]);
  AND2 I252 (gtint_1[28:28], choice_1, i_1r1[28:28]);
  AND2 I253 (gtint_1[29:29], choice_1, i_1r1[29:29]);
  AND2 I254 (gtint_1[30:30], choice_1, i_1r1[30:30]);
  AND2 I255 (gtint_1[31:31], choice_1, i_1r1[31:31]);
  AND2 I256 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I257 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I258 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I259 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AND2 I260 (gtint_2[4:4], choice_2, i_2r1[4:4]);
  AND2 I261 (gtint_2[5:5], choice_2, i_2r1[5:5]);
  AND2 I262 (gtint_2[6:6], choice_2, i_2r1[6:6]);
  AND2 I263 (gtint_2[7:7], choice_2, i_2r1[7:7]);
  AND2 I264 (gtint_2[8:8], choice_2, i_2r1[8:8]);
  AND2 I265 (gtint_2[9:9], choice_2, i_2r1[9:9]);
  AND2 I266 (gtint_2[10:10], choice_2, i_2r1[10:10]);
  AND2 I267 (gtint_2[11:11], choice_2, i_2r1[11:11]);
  AND2 I268 (gtint_2[12:12], choice_2, i_2r1[12:12]);
  AND2 I269 (gtint_2[13:13], choice_2, i_2r1[13:13]);
  AND2 I270 (gtint_2[14:14], choice_2, i_2r1[14:14]);
  AND2 I271 (gtint_2[15:15], choice_2, i_2r1[15:15]);
  AND2 I272 (gtint_2[16:16], choice_2, i_2r1[16:16]);
  AND2 I273 (gtint_2[17:17], choice_2, i_2r1[17:17]);
  AND2 I274 (gtint_2[18:18], choice_2, i_2r1[18:18]);
  AND2 I275 (gtint_2[19:19], choice_2, i_2r1[19:19]);
  AND2 I276 (gtint_2[20:20], choice_2, i_2r1[20:20]);
  AND2 I277 (gtint_2[21:21], choice_2, i_2r1[21:21]);
  AND2 I278 (gtint_2[22:22], choice_2, i_2r1[22:22]);
  AND2 I279 (gtint_2[23:23], choice_2, i_2r1[23:23]);
  AND2 I280 (gtint_2[24:24], choice_2, i_2r1[24:24]);
  AND2 I281 (gtint_2[25:25], choice_2, i_2r1[25:25]);
  AND2 I282 (gtint_2[26:26], choice_2, i_2r1[26:26]);
  AND2 I283 (gtint_2[27:27], choice_2, i_2r1[27:27]);
  AND2 I284 (gtint_2[28:28], choice_2, i_2r1[28:28]);
  AND2 I285 (gtint_2[29:29], choice_2, i_2r1[29:29]);
  AND2 I286 (gtint_2[30:30], choice_2, i_2r1[30:30]);
  AND2 I287 (gtint_2[31:31], choice_2, i_2r1[31:31]);
  AND2 I288 (gtint_3[0:0], choice_3, i_3r1[0:0]);
  AND2 I289 (gtint_3[1:1], choice_3, i_3r1[1:1]);
  AND2 I290 (gtint_3[2:2], choice_3, i_3r1[2:2]);
  AND2 I291 (gtint_3[3:3], choice_3, i_3r1[3:3]);
  AND2 I292 (gtint_3[4:4], choice_3, i_3r1[4:4]);
  AND2 I293 (gtint_3[5:5], choice_3, i_3r1[5:5]);
  AND2 I294 (gtint_3[6:6], choice_3, i_3r1[6:6]);
  AND2 I295 (gtint_3[7:7], choice_3, i_3r1[7:7]);
  AND2 I296 (gtint_3[8:8], choice_3, i_3r1[8:8]);
  AND2 I297 (gtint_3[9:9], choice_3, i_3r1[9:9]);
  AND2 I298 (gtint_3[10:10], choice_3, i_3r1[10:10]);
  AND2 I299 (gtint_3[11:11], choice_3, i_3r1[11:11]);
  AND2 I300 (gtint_3[12:12], choice_3, i_3r1[12:12]);
  AND2 I301 (gtint_3[13:13], choice_3, i_3r1[13:13]);
  AND2 I302 (gtint_3[14:14], choice_3, i_3r1[14:14]);
  AND2 I303 (gtint_3[15:15], choice_3, i_3r1[15:15]);
  AND2 I304 (gtint_3[16:16], choice_3, i_3r1[16:16]);
  AND2 I305 (gtint_3[17:17], choice_3, i_3r1[17:17]);
  AND2 I306 (gtint_3[18:18], choice_3, i_3r1[18:18]);
  AND2 I307 (gtint_3[19:19], choice_3, i_3r1[19:19]);
  AND2 I308 (gtint_3[20:20], choice_3, i_3r1[20:20]);
  AND2 I309 (gtint_3[21:21], choice_3, i_3r1[21:21]);
  AND2 I310 (gtint_3[22:22], choice_3, i_3r1[22:22]);
  AND2 I311 (gtint_3[23:23], choice_3, i_3r1[23:23]);
  AND2 I312 (gtint_3[24:24], choice_3, i_3r1[24:24]);
  AND2 I313 (gtint_3[25:25], choice_3, i_3r1[25:25]);
  AND2 I314 (gtint_3[26:26], choice_3, i_3r1[26:26]);
  AND2 I315 (gtint_3[27:27], choice_3, i_3r1[27:27]);
  AND2 I316 (gtint_3[28:28], choice_3, i_3r1[28:28]);
  AND2 I317 (gtint_3[29:29], choice_3, i_3r1[29:29]);
  AND2 I318 (gtint_3[30:30], choice_3, i_3r1[30:30]);
  AND2 I319 (gtint_3[31:31], choice_3, i_3r1[31:31]);
  AND2 I320 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I321 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I322 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I323 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I324 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I325 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I326 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I327 (gfint_0[7:7], choice_0, i_0r0[7:7]);
  AND2 I328 (gfint_0[8:8], choice_0, i_0r0[8:8]);
  AND2 I329 (gfint_0[9:9], choice_0, i_0r0[9:9]);
  AND2 I330 (gfint_0[10:10], choice_0, i_0r0[10:10]);
  AND2 I331 (gfint_0[11:11], choice_0, i_0r0[11:11]);
  AND2 I332 (gfint_0[12:12], choice_0, i_0r0[12:12]);
  AND2 I333 (gfint_0[13:13], choice_0, i_0r0[13:13]);
  AND2 I334 (gfint_0[14:14], choice_0, i_0r0[14:14]);
  AND2 I335 (gfint_0[15:15], choice_0, i_0r0[15:15]);
  AND2 I336 (gfint_0[16:16], choice_0, i_0r0[16:16]);
  AND2 I337 (gfint_0[17:17], choice_0, i_0r0[17:17]);
  AND2 I338 (gfint_0[18:18], choice_0, i_0r0[18:18]);
  AND2 I339 (gfint_0[19:19], choice_0, i_0r0[19:19]);
  AND2 I340 (gfint_0[20:20], choice_0, i_0r0[20:20]);
  AND2 I341 (gfint_0[21:21], choice_0, i_0r0[21:21]);
  AND2 I342 (gfint_0[22:22], choice_0, i_0r0[22:22]);
  AND2 I343 (gfint_0[23:23], choice_0, i_0r0[23:23]);
  AND2 I344 (gfint_0[24:24], choice_0, i_0r0[24:24]);
  AND2 I345 (gfint_0[25:25], choice_0, i_0r0[25:25]);
  AND2 I346 (gfint_0[26:26], choice_0, i_0r0[26:26]);
  AND2 I347 (gfint_0[27:27], choice_0, i_0r0[27:27]);
  AND2 I348 (gfint_0[28:28], choice_0, i_0r0[28:28]);
  AND2 I349 (gfint_0[29:29], choice_0, i_0r0[29:29]);
  AND2 I350 (gfint_0[30:30], choice_0, i_0r0[30:30]);
  AND2 I351 (gfint_0[31:31], choice_0, i_0r0[31:31]);
  AND2 I352 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I353 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I354 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I355 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I356 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I357 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I358 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I359 (gfint_1[7:7], choice_1, i_1r0[7:7]);
  AND2 I360 (gfint_1[8:8], choice_1, i_1r0[8:8]);
  AND2 I361 (gfint_1[9:9], choice_1, i_1r0[9:9]);
  AND2 I362 (gfint_1[10:10], choice_1, i_1r0[10:10]);
  AND2 I363 (gfint_1[11:11], choice_1, i_1r0[11:11]);
  AND2 I364 (gfint_1[12:12], choice_1, i_1r0[12:12]);
  AND2 I365 (gfint_1[13:13], choice_1, i_1r0[13:13]);
  AND2 I366 (gfint_1[14:14], choice_1, i_1r0[14:14]);
  AND2 I367 (gfint_1[15:15], choice_1, i_1r0[15:15]);
  AND2 I368 (gfint_1[16:16], choice_1, i_1r0[16:16]);
  AND2 I369 (gfint_1[17:17], choice_1, i_1r0[17:17]);
  AND2 I370 (gfint_1[18:18], choice_1, i_1r0[18:18]);
  AND2 I371 (gfint_1[19:19], choice_1, i_1r0[19:19]);
  AND2 I372 (gfint_1[20:20], choice_1, i_1r0[20:20]);
  AND2 I373 (gfint_1[21:21], choice_1, i_1r0[21:21]);
  AND2 I374 (gfint_1[22:22], choice_1, i_1r0[22:22]);
  AND2 I375 (gfint_1[23:23], choice_1, i_1r0[23:23]);
  AND2 I376 (gfint_1[24:24], choice_1, i_1r0[24:24]);
  AND2 I377 (gfint_1[25:25], choice_1, i_1r0[25:25]);
  AND2 I378 (gfint_1[26:26], choice_1, i_1r0[26:26]);
  AND2 I379 (gfint_1[27:27], choice_1, i_1r0[27:27]);
  AND2 I380 (gfint_1[28:28], choice_1, i_1r0[28:28]);
  AND2 I381 (gfint_1[29:29], choice_1, i_1r0[29:29]);
  AND2 I382 (gfint_1[30:30], choice_1, i_1r0[30:30]);
  AND2 I383 (gfint_1[31:31], choice_1, i_1r0[31:31]);
  AND2 I384 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I385 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I386 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I387 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AND2 I388 (gfint_2[4:4], choice_2, i_2r0[4:4]);
  AND2 I389 (gfint_2[5:5], choice_2, i_2r0[5:5]);
  AND2 I390 (gfint_2[6:6], choice_2, i_2r0[6:6]);
  AND2 I391 (gfint_2[7:7], choice_2, i_2r0[7:7]);
  AND2 I392 (gfint_2[8:8], choice_2, i_2r0[8:8]);
  AND2 I393 (gfint_2[9:9], choice_2, i_2r0[9:9]);
  AND2 I394 (gfint_2[10:10], choice_2, i_2r0[10:10]);
  AND2 I395 (gfint_2[11:11], choice_2, i_2r0[11:11]);
  AND2 I396 (gfint_2[12:12], choice_2, i_2r0[12:12]);
  AND2 I397 (gfint_2[13:13], choice_2, i_2r0[13:13]);
  AND2 I398 (gfint_2[14:14], choice_2, i_2r0[14:14]);
  AND2 I399 (gfint_2[15:15], choice_2, i_2r0[15:15]);
  AND2 I400 (gfint_2[16:16], choice_2, i_2r0[16:16]);
  AND2 I401 (gfint_2[17:17], choice_2, i_2r0[17:17]);
  AND2 I402 (gfint_2[18:18], choice_2, i_2r0[18:18]);
  AND2 I403 (gfint_2[19:19], choice_2, i_2r0[19:19]);
  AND2 I404 (gfint_2[20:20], choice_2, i_2r0[20:20]);
  AND2 I405 (gfint_2[21:21], choice_2, i_2r0[21:21]);
  AND2 I406 (gfint_2[22:22], choice_2, i_2r0[22:22]);
  AND2 I407 (gfint_2[23:23], choice_2, i_2r0[23:23]);
  AND2 I408 (gfint_2[24:24], choice_2, i_2r0[24:24]);
  AND2 I409 (gfint_2[25:25], choice_2, i_2r0[25:25]);
  AND2 I410 (gfint_2[26:26], choice_2, i_2r0[26:26]);
  AND2 I411 (gfint_2[27:27], choice_2, i_2r0[27:27]);
  AND2 I412 (gfint_2[28:28], choice_2, i_2r0[28:28]);
  AND2 I413 (gfint_2[29:29], choice_2, i_2r0[29:29]);
  AND2 I414 (gfint_2[30:30], choice_2, i_2r0[30:30]);
  AND2 I415 (gfint_2[31:31], choice_2, i_2r0[31:31]);
  AND2 I416 (gfint_3[0:0], choice_3, i_3r0[0:0]);
  AND2 I417 (gfint_3[1:1], choice_3, i_3r0[1:1]);
  AND2 I418 (gfint_3[2:2], choice_3, i_3r0[2:2]);
  AND2 I419 (gfint_3[3:3], choice_3, i_3r0[3:3]);
  AND2 I420 (gfint_3[4:4], choice_3, i_3r0[4:4]);
  AND2 I421 (gfint_3[5:5], choice_3, i_3r0[5:5]);
  AND2 I422 (gfint_3[6:6], choice_3, i_3r0[6:6]);
  AND2 I423 (gfint_3[7:7], choice_3, i_3r0[7:7]);
  AND2 I424 (gfint_3[8:8], choice_3, i_3r0[8:8]);
  AND2 I425 (gfint_3[9:9], choice_3, i_3r0[9:9]);
  AND2 I426 (gfint_3[10:10], choice_3, i_3r0[10:10]);
  AND2 I427 (gfint_3[11:11], choice_3, i_3r0[11:11]);
  AND2 I428 (gfint_3[12:12], choice_3, i_3r0[12:12]);
  AND2 I429 (gfint_3[13:13], choice_3, i_3r0[13:13]);
  AND2 I430 (gfint_3[14:14], choice_3, i_3r0[14:14]);
  AND2 I431 (gfint_3[15:15], choice_3, i_3r0[15:15]);
  AND2 I432 (gfint_3[16:16], choice_3, i_3r0[16:16]);
  AND2 I433 (gfint_3[17:17], choice_3, i_3r0[17:17]);
  AND2 I434 (gfint_3[18:18], choice_3, i_3r0[18:18]);
  AND2 I435 (gfint_3[19:19], choice_3, i_3r0[19:19]);
  AND2 I436 (gfint_3[20:20], choice_3, i_3r0[20:20]);
  AND2 I437 (gfint_3[21:21], choice_3, i_3r0[21:21]);
  AND2 I438 (gfint_3[22:22], choice_3, i_3r0[22:22]);
  AND2 I439 (gfint_3[23:23], choice_3, i_3r0[23:23]);
  AND2 I440 (gfint_3[24:24], choice_3, i_3r0[24:24]);
  AND2 I441 (gfint_3[25:25], choice_3, i_3r0[25:25]);
  AND2 I442 (gfint_3[26:26], choice_3, i_3r0[26:26]);
  AND2 I443 (gfint_3[27:27], choice_3, i_3r0[27:27]);
  AND2 I444 (gfint_3[28:28], choice_3, i_3r0[28:28]);
  AND2 I445 (gfint_3[29:29], choice_3, i_3r0[29:29]);
  AND2 I446 (gfint_3[30:30], choice_3, i_3r0[30:30]);
  AND2 I447 (gfint_3[31:31], choice_3, i_3r0[31:31]);
  OR2 I448 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I449 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I450 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I451 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I452 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I453 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I454 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I455 (comp0_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I456 (comp0_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I457 (comp0_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I458 (comp0_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I459 (comp0_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I460 (comp0_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I461 (comp0_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I462 (comp0_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I463 (comp0_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I464 (comp0_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I465 (comp0_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I466 (comp0_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I467 (comp0_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I468 (comp0_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I469 (comp0_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I470 (comp0_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I471 (comp0_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I472 (comp0_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I473 (comp0_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I474 (comp0_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I475 (comp0_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I476 (comp0_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I477 (comp0_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I478 (comp0_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I479 (comp0_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  C3 I480 (simp3711_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I481 (simp3711_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I482 (simp3711_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I483 (simp3711_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I484 (simp3711_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I485 (simp3711_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I486 (simp3711_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I487 (simp3711_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I488 (simp3711_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I489 (simp3711_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I490 (simp3711_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I491 (simp3712_0[0:0], simp3711_0[0:0], simp3711_0[1:1], simp3711_0[2:2]);
  C3 I492 (simp3712_0[1:1], simp3711_0[3:3], simp3711_0[4:4], simp3711_0[5:5]);
  C3 I493 (simp3712_0[2:2], simp3711_0[6:6], simp3711_0[7:7], simp3711_0[8:8]);
  C2 I494 (simp3712_0[3:3], simp3711_0[9:9], simp3711_0[10:10]);
  C3 I495 (simp3713_0[0:0], simp3712_0[0:0], simp3712_0[1:1], simp3712_0[2:2]);
  BUFF I496 (simp3713_0[1:1], simp3712_0[3:3]);
  C2 I497 (icomp_0, simp3713_0[0:0], simp3713_0[1:1]);
  OR2 I498 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I499 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I500 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I501 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I502 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I503 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I504 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  OR2 I505 (comp1_0[7:7], i_1r0[7:7], i_1r1[7:7]);
  OR2 I506 (comp1_0[8:8], i_1r0[8:8], i_1r1[8:8]);
  OR2 I507 (comp1_0[9:9], i_1r0[9:9], i_1r1[9:9]);
  OR2 I508 (comp1_0[10:10], i_1r0[10:10], i_1r1[10:10]);
  OR2 I509 (comp1_0[11:11], i_1r0[11:11], i_1r1[11:11]);
  OR2 I510 (comp1_0[12:12], i_1r0[12:12], i_1r1[12:12]);
  OR2 I511 (comp1_0[13:13], i_1r0[13:13], i_1r1[13:13]);
  OR2 I512 (comp1_0[14:14], i_1r0[14:14], i_1r1[14:14]);
  OR2 I513 (comp1_0[15:15], i_1r0[15:15], i_1r1[15:15]);
  OR2 I514 (comp1_0[16:16], i_1r0[16:16], i_1r1[16:16]);
  OR2 I515 (comp1_0[17:17], i_1r0[17:17], i_1r1[17:17]);
  OR2 I516 (comp1_0[18:18], i_1r0[18:18], i_1r1[18:18]);
  OR2 I517 (comp1_0[19:19], i_1r0[19:19], i_1r1[19:19]);
  OR2 I518 (comp1_0[20:20], i_1r0[20:20], i_1r1[20:20]);
  OR2 I519 (comp1_0[21:21], i_1r0[21:21], i_1r1[21:21]);
  OR2 I520 (comp1_0[22:22], i_1r0[22:22], i_1r1[22:22]);
  OR2 I521 (comp1_0[23:23], i_1r0[23:23], i_1r1[23:23]);
  OR2 I522 (comp1_0[24:24], i_1r0[24:24], i_1r1[24:24]);
  OR2 I523 (comp1_0[25:25], i_1r0[25:25], i_1r1[25:25]);
  OR2 I524 (comp1_0[26:26], i_1r0[26:26], i_1r1[26:26]);
  OR2 I525 (comp1_0[27:27], i_1r0[27:27], i_1r1[27:27]);
  OR2 I526 (comp1_0[28:28], i_1r0[28:28], i_1r1[28:28]);
  OR2 I527 (comp1_0[29:29], i_1r0[29:29], i_1r1[29:29]);
  OR2 I528 (comp1_0[30:30], i_1r0[30:30], i_1r1[30:30]);
  OR2 I529 (comp1_0[31:31], i_1r0[31:31], i_1r1[31:31]);
  C3 I530 (simp4051_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I531 (simp4051_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  C3 I532 (simp4051_0[2:2], comp1_0[6:6], comp1_0[7:7], comp1_0[8:8]);
  C3 I533 (simp4051_0[3:3], comp1_0[9:9], comp1_0[10:10], comp1_0[11:11]);
  C3 I534 (simp4051_0[4:4], comp1_0[12:12], comp1_0[13:13], comp1_0[14:14]);
  C3 I535 (simp4051_0[5:5], comp1_0[15:15], comp1_0[16:16], comp1_0[17:17]);
  C3 I536 (simp4051_0[6:6], comp1_0[18:18], comp1_0[19:19], comp1_0[20:20]);
  C3 I537 (simp4051_0[7:7], comp1_0[21:21], comp1_0[22:22], comp1_0[23:23]);
  C3 I538 (simp4051_0[8:8], comp1_0[24:24], comp1_0[25:25], comp1_0[26:26]);
  C3 I539 (simp4051_0[9:9], comp1_0[27:27], comp1_0[28:28], comp1_0[29:29]);
  C2 I540 (simp4051_0[10:10], comp1_0[30:30], comp1_0[31:31]);
  C3 I541 (simp4052_0[0:0], simp4051_0[0:0], simp4051_0[1:1], simp4051_0[2:2]);
  C3 I542 (simp4052_0[1:1], simp4051_0[3:3], simp4051_0[4:4], simp4051_0[5:5]);
  C3 I543 (simp4052_0[2:2], simp4051_0[6:6], simp4051_0[7:7], simp4051_0[8:8]);
  C2 I544 (simp4052_0[3:3], simp4051_0[9:9], simp4051_0[10:10]);
  C3 I545 (simp4053_0[0:0], simp4052_0[0:0], simp4052_0[1:1], simp4052_0[2:2]);
  BUFF I546 (simp4053_0[1:1], simp4052_0[3:3]);
  C2 I547 (icomp_1, simp4053_0[0:0], simp4053_0[1:1]);
  OR2 I548 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I549 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I550 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2 I551 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  OR2 I552 (comp2_0[4:4], i_2r0[4:4], i_2r1[4:4]);
  OR2 I553 (comp2_0[5:5], i_2r0[5:5], i_2r1[5:5]);
  OR2 I554 (comp2_0[6:6], i_2r0[6:6], i_2r1[6:6]);
  OR2 I555 (comp2_0[7:7], i_2r0[7:7], i_2r1[7:7]);
  OR2 I556 (comp2_0[8:8], i_2r0[8:8], i_2r1[8:8]);
  OR2 I557 (comp2_0[9:9], i_2r0[9:9], i_2r1[9:9]);
  OR2 I558 (comp2_0[10:10], i_2r0[10:10], i_2r1[10:10]);
  OR2 I559 (comp2_0[11:11], i_2r0[11:11], i_2r1[11:11]);
  OR2 I560 (comp2_0[12:12], i_2r0[12:12], i_2r1[12:12]);
  OR2 I561 (comp2_0[13:13], i_2r0[13:13], i_2r1[13:13]);
  OR2 I562 (comp2_0[14:14], i_2r0[14:14], i_2r1[14:14]);
  OR2 I563 (comp2_0[15:15], i_2r0[15:15], i_2r1[15:15]);
  OR2 I564 (comp2_0[16:16], i_2r0[16:16], i_2r1[16:16]);
  OR2 I565 (comp2_0[17:17], i_2r0[17:17], i_2r1[17:17]);
  OR2 I566 (comp2_0[18:18], i_2r0[18:18], i_2r1[18:18]);
  OR2 I567 (comp2_0[19:19], i_2r0[19:19], i_2r1[19:19]);
  OR2 I568 (comp2_0[20:20], i_2r0[20:20], i_2r1[20:20]);
  OR2 I569 (comp2_0[21:21], i_2r0[21:21], i_2r1[21:21]);
  OR2 I570 (comp2_0[22:22], i_2r0[22:22], i_2r1[22:22]);
  OR2 I571 (comp2_0[23:23], i_2r0[23:23], i_2r1[23:23]);
  OR2 I572 (comp2_0[24:24], i_2r0[24:24], i_2r1[24:24]);
  OR2 I573 (comp2_0[25:25], i_2r0[25:25], i_2r1[25:25]);
  OR2 I574 (comp2_0[26:26], i_2r0[26:26], i_2r1[26:26]);
  OR2 I575 (comp2_0[27:27], i_2r0[27:27], i_2r1[27:27]);
  OR2 I576 (comp2_0[28:28], i_2r0[28:28], i_2r1[28:28]);
  OR2 I577 (comp2_0[29:29], i_2r0[29:29], i_2r1[29:29]);
  OR2 I578 (comp2_0[30:30], i_2r0[30:30], i_2r1[30:30]);
  OR2 I579 (comp2_0[31:31], i_2r0[31:31], i_2r1[31:31]);
  C3 I580 (simp4391_0[0:0], comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C3 I581 (simp4391_0[1:1], comp2_0[3:3], comp2_0[4:4], comp2_0[5:5]);
  C3 I582 (simp4391_0[2:2], comp2_0[6:6], comp2_0[7:7], comp2_0[8:8]);
  C3 I583 (simp4391_0[3:3], comp2_0[9:9], comp2_0[10:10], comp2_0[11:11]);
  C3 I584 (simp4391_0[4:4], comp2_0[12:12], comp2_0[13:13], comp2_0[14:14]);
  C3 I585 (simp4391_0[5:5], comp2_0[15:15], comp2_0[16:16], comp2_0[17:17]);
  C3 I586 (simp4391_0[6:6], comp2_0[18:18], comp2_0[19:19], comp2_0[20:20]);
  C3 I587 (simp4391_0[7:7], comp2_0[21:21], comp2_0[22:22], comp2_0[23:23]);
  C3 I588 (simp4391_0[8:8], comp2_0[24:24], comp2_0[25:25], comp2_0[26:26]);
  C3 I589 (simp4391_0[9:9], comp2_0[27:27], comp2_0[28:28], comp2_0[29:29]);
  C2 I590 (simp4391_0[10:10], comp2_0[30:30], comp2_0[31:31]);
  C3 I591 (simp4392_0[0:0], simp4391_0[0:0], simp4391_0[1:1], simp4391_0[2:2]);
  C3 I592 (simp4392_0[1:1], simp4391_0[3:3], simp4391_0[4:4], simp4391_0[5:5]);
  C3 I593 (simp4392_0[2:2], simp4391_0[6:6], simp4391_0[7:7], simp4391_0[8:8]);
  C2 I594 (simp4392_0[3:3], simp4391_0[9:9], simp4391_0[10:10]);
  C3 I595 (simp4393_0[0:0], simp4392_0[0:0], simp4392_0[1:1], simp4392_0[2:2]);
  BUFF I596 (simp4393_0[1:1], simp4392_0[3:3]);
  C2 I597 (icomp_2, simp4393_0[0:0], simp4393_0[1:1]);
  OR2 I598 (comp3_0[0:0], i_3r0[0:0], i_3r1[0:0]);
  OR2 I599 (comp3_0[1:1], i_3r0[1:1], i_3r1[1:1]);
  OR2 I600 (comp3_0[2:2], i_3r0[2:2], i_3r1[2:2]);
  OR2 I601 (comp3_0[3:3], i_3r0[3:3], i_3r1[3:3]);
  OR2 I602 (comp3_0[4:4], i_3r0[4:4], i_3r1[4:4]);
  OR2 I603 (comp3_0[5:5], i_3r0[5:5], i_3r1[5:5]);
  OR2 I604 (comp3_0[6:6], i_3r0[6:6], i_3r1[6:6]);
  OR2 I605 (comp3_0[7:7], i_3r0[7:7], i_3r1[7:7]);
  OR2 I606 (comp3_0[8:8], i_3r0[8:8], i_3r1[8:8]);
  OR2 I607 (comp3_0[9:9], i_3r0[9:9], i_3r1[9:9]);
  OR2 I608 (comp3_0[10:10], i_3r0[10:10], i_3r1[10:10]);
  OR2 I609 (comp3_0[11:11], i_3r0[11:11], i_3r1[11:11]);
  OR2 I610 (comp3_0[12:12], i_3r0[12:12], i_3r1[12:12]);
  OR2 I611 (comp3_0[13:13], i_3r0[13:13], i_3r1[13:13]);
  OR2 I612 (comp3_0[14:14], i_3r0[14:14], i_3r1[14:14]);
  OR2 I613 (comp3_0[15:15], i_3r0[15:15], i_3r1[15:15]);
  OR2 I614 (comp3_0[16:16], i_3r0[16:16], i_3r1[16:16]);
  OR2 I615 (comp3_0[17:17], i_3r0[17:17], i_3r1[17:17]);
  OR2 I616 (comp3_0[18:18], i_3r0[18:18], i_3r1[18:18]);
  OR2 I617 (comp3_0[19:19], i_3r0[19:19], i_3r1[19:19]);
  OR2 I618 (comp3_0[20:20], i_3r0[20:20], i_3r1[20:20]);
  OR2 I619 (comp3_0[21:21], i_3r0[21:21], i_3r1[21:21]);
  OR2 I620 (comp3_0[22:22], i_3r0[22:22], i_3r1[22:22]);
  OR2 I621 (comp3_0[23:23], i_3r0[23:23], i_3r1[23:23]);
  OR2 I622 (comp3_0[24:24], i_3r0[24:24], i_3r1[24:24]);
  OR2 I623 (comp3_0[25:25], i_3r0[25:25], i_3r1[25:25]);
  OR2 I624 (comp3_0[26:26], i_3r0[26:26], i_3r1[26:26]);
  OR2 I625 (comp3_0[27:27], i_3r0[27:27], i_3r1[27:27]);
  OR2 I626 (comp3_0[28:28], i_3r0[28:28], i_3r1[28:28]);
  OR2 I627 (comp3_0[29:29], i_3r0[29:29], i_3r1[29:29]);
  OR2 I628 (comp3_0[30:30], i_3r0[30:30], i_3r1[30:30]);
  OR2 I629 (comp3_0[31:31], i_3r0[31:31], i_3r1[31:31]);
  C3 I630 (simp4731_0[0:0], comp3_0[0:0], comp3_0[1:1], comp3_0[2:2]);
  C3 I631 (simp4731_0[1:1], comp3_0[3:3], comp3_0[4:4], comp3_0[5:5]);
  C3 I632 (simp4731_0[2:2], comp3_0[6:6], comp3_0[7:7], comp3_0[8:8]);
  C3 I633 (simp4731_0[3:3], comp3_0[9:9], comp3_0[10:10], comp3_0[11:11]);
  C3 I634 (simp4731_0[4:4], comp3_0[12:12], comp3_0[13:13], comp3_0[14:14]);
  C3 I635 (simp4731_0[5:5], comp3_0[15:15], comp3_0[16:16], comp3_0[17:17]);
  C3 I636 (simp4731_0[6:6], comp3_0[18:18], comp3_0[19:19], comp3_0[20:20]);
  C3 I637 (simp4731_0[7:7], comp3_0[21:21], comp3_0[22:22], comp3_0[23:23]);
  C3 I638 (simp4731_0[8:8], comp3_0[24:24], comp3_0[25:25], comp3_0[26:26]);
  C3 I639 (simp4731_0[9:9], comp3_0[27:27], comp3_0[28:28], comp3_0[29:29]);
  C2 I640 (simp4731_0[10:10], comp3_0[30:30], comp3_0[31:31]);
  C3 I641 (simp4732_0[0:0], simp4731_0[0:0], simp4731_0[1:1], simp4731_0[2:2]);
  C3 I642 (simp4732_0[1:1], simp4731_0[3:3], simp4731_0[4:4], simp4731_0[5:5]);
  C3 I643 (simp4732_0[2:2], simp4731_0[6:6], simp4731_0[7:7], simp4731_0[8:8]);
  C2 I644 (simp4732_0[3:3], simp4731_0[9:9], simp4731_0[10:10]);
  C3 I645 (simp4733_0[0:0], simp4732_0[0:0], simp4732_0[1:1], simp4732_0[2:2]);
  BUFF I646 (simp4733_0[1:1], simp4732_0[3:3]);
  C2 I647 (icomp_3, simp4733_0[0:0], simp4733_0[1:1]);
  C2R I648 (choice_0, icomp_0, nchosen_0, reset);
  C2R I649 (choice_1, icomp_1, nchosen_0, reset);
  C2R I650 (choice_2, icomp_2, nchosen_0, reset);
  C2R I651 (choice_3, icomp_3, nchosen_0, reset);
  NOR3 I652 (simp4781_0[0:0], choice_0, choice_1, choice_2);
  INV I653 (simp4781_0[1:1], choice_3);
  NAND2 I654 (anychoice_0, simp4781_0[0:0], simp4781_0[1:1]);
  NOR2 I655 (nchosen_0, anychoice_0, o_0a);
  C2R I656 (i_0a, choice_0, o_0a, reset);
  C2R I657 (i_1a, choice_1, o_0a, reset);
  C2R I658 (i_2a, choice_2, o_0a, reset);
  C2R I659 (i_3a, choice_3, o_0a, reset);
endmodule

// tkj32m32_0 TeakJ [Many [32,0],One 32]
module tkj32m32_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [31:0] joinf_0;
  wire [31:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joint_0[0:0], i_0r1[0:0]);
  BUFF I33 (joint_0[1:1], i_0r1[1:1]);
  BUFF I34 (joint_0[2:2], i_0r1[2:2]);
  BUFF I35 (joint_0[3:3], i_0r1[3:3]);
  BUFF I36 (joint_0[4:4], i_0r1[4:4]);
  BUFF I37 (joint_0[5:5], i_0r1[5:5]);
  BUFF I38 (joint_0[6:6], i_0r1[6:6]);
  BUFF I39 (joint_0[7:7], i_0r1[7:7]);
  BUFF I40 (joint_0[8:8], i_0r1[8:8]);
  BUFF I41 (joint_0[9:9], i_0r1[9:9]);
  BUFF I42 (joint_0[10:10], i_0r1[10:10]);
  BUFF I43 (joint_0[11:11], i_0r1[11:11]);
  BUFF I44 (joint_0[12:12], i_0r1[12:12]);
  BUFF I45 (joint_0[13:13], i_0r1[13:13]);
  BUFF I46 (joint_0[14:14], i_0r1[14:14]);
  BUFF I47 (joint_0[15:15], i_0r1[15:15]);
  BUFF I48 (joint_0[16:16], i_0r1[16:16]);
  BUFF I49 (joint_0[17:17], i_0r1[17:17]);
  BUFF I50 (joint_0[18:18], i_0r1[18:18]);
  BUFF I51 (joint_0[19:19], i_0r1[19:19]);
  BUFF I52 (joint_0[20:20], i_0r1[20:20]);
  BUFF I53 (joint_0[21:21], i_0r1[21:21]);
  BUFF I54 (joint_0[22:22], i_0r1[22:22]);
  BUFF I55 (joint_0[23:23], i_0r1[23:23]);
  BUFF I56 (joint_0[24:24], i_0r1[24:24]);
  BUFF I57 (joint_0[25:25], i_0r1[25:25]);
  BUFF I58 (joint_0[26:26], i_0r1[26:26]);
  BUFF I59 (joint_0[27:27], i_0r1[27:27]);
  BUFF I60 (joint_0[28:28], i_0r1[28:28]);
  BUFF I61 (joint_0[29:29], i_0r1[29:29]);
  BUFF I62 (joint_0[30:30], i_0r1[30:30]);
  BUFF I63 (joint_0[31:31], i_0r1[31:31]);
  BUFF I64 (icomplete_0, i_1r);
  C2 I65 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I66 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I67 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I68 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I69 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I70 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I71 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I72 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I73 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I74 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I75 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I76 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I77 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I78 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I79 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I80 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I81 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I82 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I83 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I84 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I85 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I86 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I87 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I88 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I89 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I90 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I91 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I92 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I93 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I94 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I95 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I96 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I97 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I98 (o_0r1[1:1], joint_0[1:1]);
  BUFF I99 (o_0r1[2:2], joint_0[2:2]);
  BUFF I100 (o_0r1[3:3], joint_0[3:3]);
  BUFF I101 (o_0r1[4:4], joint_0[4:4]);
  BUFF I102 (o_0r1[5:5], joint_0[5:5]);
  BUFF I103 (o_0r1[6:6], joint_0[6:6]);
  BUFF I104 (o_0r1[7:7], joint_0[7:7]);
  BUFF I105 (o_0r1[8:8], joint_0[8:8]);
  BUFF I106 (o_0r1[9:9], joint_0[9:9]);
  BUFF I107 (o_0r1[10:10], joint_0[10:10]);
  BUFF I108 (o_0r1[11:11], joint_0[11:11]);
  BUFF I109 (o_0r1[12:12], joint_0[12:12]);
  BUFF I110 (o_0r1[13:13], joint_0[13:13]);
  BUFF I111 (o_0r1[14:14], joint_0[14:14]);
  BUFF I112 (o_0r1[15:15], joint_0[15:15]);
  BUFF I113 (o_0r1[16:16], joint_0[16:16]);
  BUFF I114 (o_0r1[17:17], joint_0[17:17]);
  BUFF I115 (o_0r1[18:18], joint_0[18:18]);
  BUFF I116 (o_0r1[19:19], joint_0[19:19]);
  BUFF I117 (o_0r1[20:20], joint_0[20:20]);
  BUFF I118 (o_0r1[21:21], joint_0[21:21]);
  BUFF I119 (o_0r1[22:22], joint_0[22:22]);
  BUFF I120 (o_0r1[23:23], joint_0[23:23]);
  BUFF I121 (o_0r1[24:24], joint_0[24:24]);
  BUFF I122 (o_0r1[25:25], joint_0[25:25]);
  BUFF I123 (o_0r1[26:26], joint_0[26:26]);
  BUFF I124 (o_0r1[27:27], joint_0[27:27]);
  BUFF I125 (o_0r1[28:28], joint_0[28:28]);
  BUFF I126 (o_0r1[29:29], joint_0[29:29]);
  BUFF I127 (o_0r1[30:30], joint_0[30:30]);
  BUFF I128 (o_0r1[31:31], joint_0[31:31]);
  BUFF I129 (i_0a, o_0a);
  BUFF I130 (i_1a, o_0a);
endmodule

// tkf32mo0w0_o0w32 TeakF [0,0] [One 32,Many [0,32]]
module tkf32mo0w0_o0w32 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [31:0] o_1r0;
  output [31:0] o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_1r0[0:0], i_0r0[0:0]);
  BUFF I3 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I4 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I5 (o_1r0[3:3], i_0r0[3:3]);
  BUFF I6 (o_1r0[4:4], i_0r0[4:4]);
  BUFF I7 (o_1r0[5:5], i_0r0[5:5]);
  BUFF I8 (o_1r0[6:6], i_0r0[6:6]);
  BUFF I9 (o_1r0[7:7], i_0r0[7:7]);
  BUFF I10 (o_1r0[8:8], i_0r0[8:8]);
  BUFF I11 (o_1r0[9:9], i_0r0[9:9]);
  BUFF I12 (o_1r0[10:10], i_0r0[10:10]);
  BUFF I13 (o_1r0[11:11], i_0r0[11:11]);
  BUFF I14 (o_1r0[12:12], i_0r0[12:12]);
  BUFF I15 (o_1r0[13:13], i_0r0[13:13]);
  BUFF I16 (o_1r0[14:14], i_0r0[14:14]);
  BUFF I17 (o_1r0[15:15], i_0r0[15:15]);
  BUFF I18 (o_1r0[16:16], i_0r0[16:16]);
  BUFF I19 (o_1r0[17:17], i_0r0[17:17]);
  BUFF I20 (o_1r0[18:18], i_0r0[18:18]);
  BUFF I21 (o_1r0[19:19], i_0r0[19:19]);
  BUFF I22 (o_1r0[20:20], i_0r0[20:20]);
  BUFF I23 (o_1r0[21:21], i_0r0[21:21]);
  BUFF I24 (o_1r0[22:22], i_0r0[22:22]);
  BUFF I25 (o_1r0[23:23], i_0r0[23:23]);
  BUFF I26 (o_1r0[24:24], i_0r0[24:24]);
  BUFF I27 (o_1r0[25:25], i_0r0[25:25]);
  BUFF I28 (o_1r0[26:26], i_0r0[26:26]);
  BUFF I29 (o_1r0[27:27], i_0r0[27:27]);
  BUFF I30 (o_1r0[28:28], i_0r0[28:28]);
  BUFF I31 (o_1r0[29:29], i_0r0[29:29]);
  BUFF I32 (o_1r0[30:30], i_0r0[30:30]);
  BUFF I33 (o_1r0[31:31], i_0r0[31:31]);
  BUFF I34 (o_1r1[0:0], i_0r1[0:0]);
  BUFF I35 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I36 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I37 (o_1r1[3:3], i_0r1[3:3]);
  BUFF I38 (o_1r1[4:4], i_0r1[4:4]);
  BUFF I39 (o_1r1[5:5], i_0r1[5:5]);
  BUFF I40 (o_1r1[6:6], i_0r1[6:6]);
  BUFF I41 (o_1r1[7:7], i_0r1[7:7]);
  BUFF I42 (o_1r1[8:8], i_0r1[8:8]);
  BUFF I43 (o_1r1[9:9], i_0r1[9:9]);
  BUFF I44 (o_1r1[10:10], i_0r1[10:10]);
  BUFF I45 (o_1r1[11:11], i_0r1[11:11]);
  BUFF I46 (o_1r1[12:12], i_0r1[12:12]);
  BUFF I47 (o_1r1[13:13], i_0r1[13:13]);
  BUFF I48 (o_1r1[14:14], i_0r1[14:14]);
  BUFF I49 (o_1r1[15:15], i_0r1[15:15]);
  BUFF I50 (o_1r1[16:16], i_0r1[16:16]);
  BUFF I51 (o_1r1[17:17], i_0r1[17:17]);
  BUFF I52 (o_1r1[18:18], i_0r1[18:18]);
  BUFF I53 (o_1r1[19:19], i_0r1[19:19]);
  BUFF I54 (o_1r1[20:20], i_0r1[20:20]);
  BUFF I55 (o_1r1[21:21], i_0r1[21:21]);
  BUFF I56 (o_1r1[22:22], i_0r1[22:22]);
  BUFF I57 (o_1r1[23:23], i_0r1[23:23]);
  BUFF I58 (o_1r1[24:24], i_0r1[24:24]);
  BUFF I59 (o_1r1[25:25], i_0r1[25:25]);
  BUFF I60 (o_1r1[26:26], i_0r1[26:26]);
  BUFF I61 (o_1r1[27:27], i_0r1[27:27]);
  BUFF I62 (o_1r1[28:28], i_0r1[28:28]);
  BUFF I63 (o_1r1[29:29], i_0r1[29:29]);
  BUFF I64 (o_1r1[30:30], i_0r1[30:30]);
  BUFF I65 (o_1r1[31:31], i_0r1[31:31]);
  BUFF I66 (o_0r, icomplete_0);
  C3 I67 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tkj7m5_2_0 TeakJ [Many [5,2,0],One 7]
module tkj7m5_2_0 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r, i_2a, o_0r0, o_0r1, o_0a, reset);
  input [4:0] i_0r0;
  input [4:0] i_0r1;
  output i_0a;
  input [1:0] i_1r0;
  input [1:0] i_1r1;
  output i_1a;
  input i_2r;
  output i_2a;
  output [6:0] o_0r0;
  output [6:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [6:0] joinf_0;
  wire [6:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_1r0[0:0]);
  BUFF I6 (joinf_0[6:6], i_1r0[1:1]);
  BUFF I7 (joint_0[0:0], i_0r1[0:0]);
  BUFF I8 (joint_0[1:1], i_0r1[1:1]);
  BUFF I9 (joint_0[2:2], i_0r1[2:2]);
  BUFF I10 (joint_0[3:3], i_0r1[3:3]);
  BUFF I11 (joint_0[4:4], i_0r1[4:4]);
  BUFF I12 (joint_0[5:5], i_1r1[0:0]);
  BUFF I13 (joint_0[6:6], i_1r1[1:1]);
  OR2 I14 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  C2 I15 (icomplete_0, i_2r, dcomplete_0);
  C2 I16 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I17 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I18 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I19 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I20 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I21 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I22 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I23 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I24 (o_0r1[1:1], joint_0[1:1]);
  BUFF I25 (o_0r1[2:2], joint_0[2:2]);
  BUFF I26 (o_0r1[3:3], joint_0[3:3]);
  BUFF I27 (o_0r1[4:4], joint_0[4:4]);
  BUFF I28 (o_0r1[5:5], joint_0[5:5]);
  BUFF I29 (o_0r1[6:6], joint_0[6:6]);
  BUFF I30 (i_0a, o_0a);
  BUFF I31 (i_1a, o_0a);
  BUFF I32 (i_2a, o_0a);
endmodule

// tkvdistanceIshift7_wo0w7_ro5w2o5w2 TeakV "distanceI-shift" 7 [] [0] [5,5] [Many [7],Many [0],Many [0
//   ,0],Many [2,2]]
module tkvdistanceIshift7_wo0w7_ro5w2o5w2 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, reset);
  input [6:0] wg_0r0;
  input [6:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [1:0] rd_0r0;
  output [1:0] rd_0r1;
  input rd_0a;
  output [1:0] rd_1r0;
  output [1:0] rd_1r1;
  input rd_1a;
  input reset;
  wire [6:0] wf_0;
  wire [6:0] wt_0;
  wire [6:0] df_0;
  wire [6:0] dt_0;
  wire wc_0;
  wire [6:0] wacks_0;
  wire [6:0] wenr_0;
  wire [6:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [6:0] drlgf_0;
  wire [6:0] drlgt_0;
  wire [6:0] comp0_0;
  wire [2:0] simp631_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [6:0] conwgit_0;
  wire [6:0] conwgif_0;
  wire conwig_0;
  wire [2:0] simp1071_0;
  wire [1:0] simp1161_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I9 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I10 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I11 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I12 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I13 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I14 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I15 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I16 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I17 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I18 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I19 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I20 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I21 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  NOR2 I22 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I23 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I24 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I25 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I26 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I27 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I28 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR3 I29 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I30 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I31 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I32 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I33 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I34 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I35 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  AO22 I36 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I37 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I38 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I39 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I40 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I41 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I42 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  OR2 I43 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I44 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I45 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I46 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I47 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I48 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I49 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  C3 I50 (simp631_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I51 (simp631_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  BUFF I52 (simp631_0[2:2], comp0_0[6:6]);
  C3 I53 (wc_0, simp631_0[0:0], simp631_0[1:1], simp631_0[2:2]);
  AND2 I54 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I55 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I56 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I57 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I58 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I59 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I60 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I61 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I62 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I63 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I64 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I65 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I66 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I67 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  BUFF I68 (conwigc_0, wc_0);
  AO22 I69 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I70 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I71 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I72 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I73 (wenr_0[0:0], wc_0);
  BUFF I74 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I75 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I76 (wenr_0[1:1], wc_0);
  BUFF I77 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I78 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I79 (wenr_0[2:2], wc_0);
  BUFF I80 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I81 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I82 (wenr_0[3:3], wc_0);
  BUFF I83 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I84 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I85 (wenr_0[4:4], wc_0);
  BUFF I86 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I87 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I88 (wenr_0[5:5], wc_0);
  BUFF I89 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I90 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I91 (wenr_0[6:6], wc_0);
  C3 I92 (simp1071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I93 (simp1071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C2 I94 (simp1071_0[2:2], wacks_0[5:5], wacks_0[6:6]);
  C3 I95 (wd_0r, simp1071_0[0:0], simp1071_0[1:1], simp1071_0[2:2]);
  AND2 I96 (rd_0r0[0:0], df_0[5:5], rg_0r);
  AND2 I97 (rd_0r0[1:1], df_0[6:6], rg_0r);
  AND2 I98 (rd_1r0[0:0], df_0[5:5], rg_1r);
  AND2 I99 (rd_1r0[1:1], df_0[6:6], rg_1r);
  AND2 I100 (rd_0r1[0:0], dt_0[5:5], rg_0r);
  AND2 I101 (rd_0r1[1:1], dt_0[6:6], rg_0r);
  AND2 I102 (rd_1r1[0:0], dt_0[5:5], rg_1r);
  AND2 I103 (rd_1r1[1:1], dt_0[6:6], rg_1r);
  NOR3 I104 (simp1161_0[0:0], rg_0r, rg_1r, rg_0a);
  INV I105 (simp1161_0[1:1], rg_1a);
  NAND2 I106 (anyread_0, simp1161_0[0:0], simp1161_0[1:1]);
  BUFF I107 (wg_0a, wd_0a);
  BUFF I108 (rg_0a, rd_0a);
  BUFF I109 (rg_1a, rd_1a);
endmodule

// tkf7mo0w7_o2w1_o1w1 TeakF [0,2,1] [One 7,Many [7,1,1]]
module tkf7mo0w7_o2w1_o1w1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r0, o_1r1, o_1a, o_2r0, o_2r1, o_2a, reset);
  input [6:0] i_0r0;
  input [6:0] i_0r1;
  output i_0a;
  output [6:0] o_0r0;
  output [6:0] o_0r1;
  input o_0a;
  output o_1r0;
  output o_1r1;
  input o_1a;
  output o_2r0;
  output o_2r1;
  input o_2a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  wire [1:0] simp231_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_0r0[0:0], i_0r0[0:0]);
  BUFF I3 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I4 (o_0r0[2:2], i_0r0[2:2]);
  BUFF I5 (o_0r0[3:3], i_0r0[3:3]);
  BUFF I6 (o_0r0[4:4], i_0r0[4:4]);
  BUFF I7 (o_0r0[5:5], i_0r0[5:5]);
  BUFF I8 (o_0r0[6:6], i_0r0[6:6]);
  C2 I9 (o_1r0, i_0r0[2:2], icomplete_0);
  C2 I10 (o_2r0, i_0r0[1:1], icomplete_0);
  BUFF I11 (o_0r1[0:0], i_0r1[0:0]);
  BUFF I12 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I13 (o_0r1[2:2], i_0r1[2:2]);
  BUFF I14 (o_0r1[3:3], i_0r1[3:3]);
  BUFF I15 (o_0r1[4:4], i_0r1[4:4]);
  BUFF I16 (o_0r1[5:5], i_0r1[5:5]);
  BUFF I17 (o_0r1[6:6], i_0r1[6:6]);
  C2 I18 (o_1r1, i_0r1[2:2], icomplete_0);
  C2 I19 (o_2r1, i_0r1[1:1], icomplete_0);
  C3 I20 (simp231_0[0:0], acomplete_0, o_0a, o_1a);
  BUFF I21 (simp231_0[1:1], o_2a);
  C2 I22 (i_0a, simp231_0[0:0], simp231_0[1:1]);
endmodule

// tkj1m1_0 TeakJ [Many [1,0],One 1]
module tkj1m1_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire joinf_0;
  wire joint_0;
  BUFF I0 (joinf_0, i_0r0);
  BUFF I1 (joint_0, i_0r1);
  BUFF I2 (icomplete_0, i_1r);
  C2 I3 (o_0r0, joinf_0, icomplete_0);
  C2 I4 (o_0r1, joint_0, icomplete_0);
  BUFF I5 (i_0a, o_0a);
  BUFF I6 (i_1a, o_0a);
endmodule

// tkf0mo0w0_o0w0 TeakF [0,0] [One 0,Many [0,0]]
module tkf0mo0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  C2 I2 (i_0a, o_0a, o_1a);
endmodule

// tks2_o0w2_3o0w0_0c2o0w0_1o0w0 TeakS (0+:2) [([Imp 3 0],0),([Imp 0 2],0),([Imp 1 0],0)] [One 2,Many [
//   0,0,0]]
module tks2_o0w2_3o0w0_0c2o0w0_1o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire match2_0;
  wire [1:0] comp_0;
  BUFF I0 (sel_0, match0_0);
  C2 I1 (match0_0, i_0r1[0:0], i_0r1[1:1]);
  BUFF I2 (sel_1, match1_0);
  BUFF I3 (match1_0, i_0r0[0:0]);
  BUFF I4 (sel_2, match2_0);
  C2 I5 (match2_0, i_0r1[0:0], i_0r0[1:1]);
  C2 I6 (gsel_0, sel_0, icomplete_0);
  C2 I7 (gsel_1, sel_1, icomplete_0);
  C2 I8 (gsel_2, sel_2, icomplete_0);
  OR2 I9 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I10 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  C2 I11 (icomplete_0, comp_0[0:0], comp_0[1:1]);
  BUFF I12 (o_0r, gsel_0);
  BUFF I13 (o_1r, gsel_1);
  BUFF I14 (o_2r, gsel_2);
  OR3 I15 (oack_0, o_0a, o_1a, o_2a);
  C2 I16 (i_0a, oack_0, icomplete_0);
endmodule

// tkf1mo0w1_o0w0 TeakF [0,0] [One 1,Many [1,0]]
module tkf1mo0w1_o0w0 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r, o_1a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0, i_0r1);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_0r0, i_0r0);
  BUFF I3 (o_0r1, i_0r1);
  BUFF I4 (o_1r, icomplete_0);
  C3 I5 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tks1_o0w1_0o0w0_1o0w0 TeakS (0+:1) [([Imp 0 0],0),([Imp 1 0],0)] [One 1,Many [0,0]]
module tks1_o0w1_0o0w0_1o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire comp_0;
  BUFF I0 (sel_0, match0_0);
  BUFF I1 (match0_0, i_0r0);
  BUFF I2 (sel_1, match1_0);
  BUFF I3 (match1_0, i_0r1);
  C2 I4 (gsel_0, sel_0, icomplete_0);
  C2 I5 (gsel_1, sel_1, icomplete_0);
  OR2 I6 (comp_0, i_0r0, i_0r1);
  BUFF I7 (icomplete_0, comp_0);
  BUFF I8 (o_0r, gsel_0);
  BUFF I9 (o_1r, gsel_1);
  OR2 I10 (oack_0, o_0a, o_1a);
  C2 I11 (i_0a, oack_0, icomplete_0);
endmodule

// tki TeakI [One 0,One 0]
module tki (i_0r, i_0a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  input reset;
  wire nreset_0;
  wire firsthsa_0;
  wire nfirsthsa_0;
  wire firsthsd_0;
  wire noa_0;
  INV I0 (nreset_0, reset);
  INV I1 (nfirsthsa_0, firsthsa_0);
  INV I2 (noa_0, o_0a);
  AO22 I3 (o_0r, nreset_0, nfirsthsa_0, i_0r, firsthsd_0);
  AO22 I4 (firsthsa_0, nreset_0, o_0a, nreset_0, firsthsa_0);
  AO22 I5 (firsthsd_0, firsthsa_0, noa_0, firsthsa_0, firsthsd_0);
  AND2 I6 (i_0a, o_0a, firsthsd_0);
endmodule

// latch tkl0x1 width = 0, depth = 1
module tkl0x1 (i_0r, i_0a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  input reset;
  wire b_0;
  C2R I0 (o_0r, i_0r, b_0, reset);
  INV I1 (b_0, o_0a);
  BUFF I2 (i_0a, o_0r);
endmodule

// latch tkl32x1 width = 32, depth = 1
module tkl32x1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire bna_0;
  wire [31:0] bcomp_0;
  wire [10:0] simp991_0;
  wire [3:0] simp992_0;
  wire [1:0] simp993_0;
  C2R I0 (o_0r0[0:0], i_0r0[0:0], bna_0, reset);
  C2R I1 (o_0r0[1:1], i_0r0[1:1], bna_0, reset);
  C2R I2 (o_0r0[2:2], i_0r0[2:2], bna_0, reset);
  C2R I3 (o_0r0[3:3], i_0r0[3:3], bna_0, reset);
  C2R I4 (o_0r0[4:4], i_0r0[4:4], bna_0, reset);
  C2R I5 (o_0r0[5:5], i_0r0[5:5], bna_0, reset);
  C2R I6 (o_0r0[6:6], i_0r0[6:6], bna_0, reset);
  C2R I7 (o_0r0[7:7], i_0r0[7:7], bna_0, reset);
  C2R I8 (o_0r0[8:8], i_0r0[8:8], bna_0, reset);
  C2R I9 (o_0r0[9:9], i_0r0[9:9], bna_0, reset);
  C2R I10 (o_0r0[10:10], i_0r0[10:10], bna_0, reset);
  C2R I11 (o_0r0[11:11], i_0r0[11:11], bna_0, reset);
  C2R I12 (o_0r0[12:12], i_0r0[12:12], bna_0, reset);
  C2R I13 (o_0r0[13:13], i_0r0[13:13], bna_0, reset);
  C2R I14 (o_0r0[14:14], i_0r0[14:14], bna_0, reset);
  C2R I15 (o_0r0[15:15], i_0r0[15:15], bna_0, reset);
  C2R I16 (o_0r0[16:16], i_0r0[16:16], bna_0, reset);
  C2R I17 (o_0r0[17:17], i_0r0[17:17], bna_0, reset);
  C2R I18 (o_0r0[18:18], i_0r0[18:18], bna_0, reset);
  C2R I19 (o_0r0[19:19], i_0r0[19:19], bna_0, reset);
  C2R I20 (o_0r0[20:20], i_0r0[20:20], bna_0, reset);
  C2R I21 (o_0r0[21:21], i_0r0[21:21], bna_0, reset);
  C2R I22 (o_0r0[22:22], i_0r0[22:22], bna_0, reset);
  C2R I23 (o_0r0[23:23], i_0r0[23:23], bna_0, reset);
  C2R I24 (o_0r0[24:24], i_0r0[24:24], bna_0, reset);
  C2R I25 (o_0r0[25:25], i_0r0[25:25], bna_0, reset);
  C2R I26 (o_0r0[26:26], i_0r0[26:26], bna_0, reset);
  C2R I27 (o_0r0[27:27], i_0r0[27:27], bna_0, reset);
  C2R I28 (o_0r0[28:28], i_0r0[28:28], bna_0, reset);
  C2R I29 (o_0r0[29:29], i_0r0[29:29], bna_0, reset);
  C2R I30 (o_0r0[30:30], i_0r0[30:30], bna_0, reset);
  C2R I31 (o_0r0[31:31], i_0r0[31:31], bna_0, reset);
  C2R I32 (o_0r1[0:0], i_0r1[0:0], bna_0, reset);
  C2R I33 (o_0r1[1:1], i_0r1[1:1], bna_0, reset);
  C2R I34 (o_0r1[2:2], i_0r1[2:2], bna_0, reset);
  C2R I35 (o_0r1[3:3], i_0r1[3:3], bna_0, reset);
  C2R I36 (o_0r1[4:4], i_0r1[4:4], bna_0, reset);
  C2R I37 (o_0r1[5:5], i_0r1[5:5], bna_0, reset);
  C2R I38 (o_0r1[6:6], i_0r1[6:6], bna_0, reset);
  C2R I39 (o_0r1[7:7], i_0r1[7:7], bna_0, reset);
  C2R I40 (o_0r1[8:8], i_0r1[8:8], bna_0, reset);
  C2R I41 (o_0r1[9:9], i_0r1[9:9], bna_0, reset);
  C2R I42 (o_0r1[10:10], i_0r1[10:10], bna_0, reset);
  C2R I43 (o_0r1[11:11], i_0r1[11:11], bna_0, reset);
  C2R I44 (o_0r1[12:12], i_0r1[12:12], bna_0, reset);
  C2R I45 (o_0r1[13:13], i_0r1[13:13], bna_0, reset);
  C2R I46 (o_0r1[14:14], i_0r1[14:14], bna_0, reset);
  C2R I47 (o_0r1[15:15], i_0r1[15:15], bna_0, reset);
  C2R I48 (o_0r1[16:16], i_0r1[16:16], bna_0, reset);
  C2R I49 (o_0r1[17:17], i_0r1[17:17], bna_0, reset);
  C2R I50 (o_0r1[18:18], i_0r1[18:18], bna_0, reset);
  C2R I51 (o_0r1[19:19], i_0r1[19:19], bna_0, reset);
  C2R I52 (o_0r1[20:20], i_0r1[20:20], bna_0, reset);
  C2R I53 (o_0r1[21:21], i_0r1[21:21], bna_0, reset);
  C2R I54 (o_0r1[22:22], i_0r1[22:22], bna_0, reset);
  C2R I55 (o_0r1[23:23], i_0r1[23:23], bna_0, reset);
  C2R I56 (o_0r1[24:24], i_0r1[24:24], bna_0, reset);
  C2R I57 (o_0r1[25:25], i_0r1[25:25], bna_0, reset);
  C2R I58 (o_0r1[26:26], i_0r1[26:26], bna_0, reset);
  C2R I59 (o_0r1[27:27], i_0r1[27:27], bna_0, reset);
  C2R I60 (o_0r1[28:28], i_0r1[28:28], bna_0, reset);
  C2R I61 (o_0r1[29:29], i_0r1[29:29], bna_0, reset);
  C2R I62 (o_0r1[30:30], i_0r1[30:30], bna_0, reset);
  C2R I63 (o_0r1[31:31], i_0r1[31:31], bna_0, reset);
  INV I64 (bna_0, o_0a);
  OR2 I65 (bcomp_0[0:0], o_0r0[0:0], o_0r1[0:0]);
  OR2 I66 (bcomp_0[1:1], o_0r0[1:1], o_0r1[1:1]);
  OR2 I67 (bcomp_0[2:2], o_0r0[2:2], o_0r1[2:2]);
  OR2 I68 (bcomp_0[3:3], o_0r0[3:3], o_0r1[3:3]);
  OR2 I69 (bcomp_0[4:4], o_0r0[4:4], o_0r1[4:4]);
  OR2 I70 (bcomp_0[5:5], o_0r0[5:5], o_0r1[5:5]);
  OR2 I71 (bcomp_0[6:6], o_0r0[6:6], o_0r1[6:6]);
  OR2 I72 (bcomp_0[7:7], o_0r0[7:7], o_0r1[7:7]);
  OR2 I73 (bcomp_0[8:8], o_0r0[8:8], o_0r1[8:8]);
  OR2 I74 (bcomp_0[9:9], o_0r0[9:9], o_0r1[9:9]);
  OR2 I75 (bcomp_0[10:10], o_0r0[10:10], o_0r1[10:10]);
  OR2 I76 (bcomp_0[11:11], o_0r0[11:11], o_0r1[11:11]);
  OR2 I77 (bcomp_0[12:12], o_0r0[12:12], o_0r1[12:12]);
  OR2 I78 (bcomp_0[13:13], o_0r0[13:13], o_0r1[13:13]);
  OR2 I79 (bcomp_0[14:14], o_0r0[14:14], o_0r1[14:14]);
  OR2 I80 (bcomp_0[15:15], o_0r0[15:15], o_0r1[15:15]);
  OR2 I81 (bcomp_0[16:16], o_0r0[16:16], o_0r1[16:16]);
  OR2 I82 (bcomp_0[17:17], o_0r0[17:17], o_0r1[17:17]);
  OR2 I83 (bcomp_0[18:18], o_0r0[18:18], o_0r1[18:18]);
  OR2 I84 (bcomp_0[19:19], o_0r0[19:19], o_0r1[19:19]);
  OR2 I85 (bcomp_0[20:20], o_0r0[20:20], o_0r1[20:20]);
  OR2 I86 (bcomp_0[21:21], o_0r0[21:21], o_0r1[21:21]);
  OR2 I87 (bcomp_0[22:22], o_0r0[22:22], o_0r1[22:22]);
  OR2 I88 (bcomp_0[23:23], o_0r0[23:23], o_0r1[23:23]);
  OR2 I89 (bcomp_0[24:24], o_0r0[24:24], o_0r1[24:24]);
  OR2 I90 (bcomp_0[25:25], o_0r0[25:25], o_0r1[25:25]);
  OR2 I91 (bcomp_0[26:26], o_0r0[26:26], o_0r1[26:26]);
  OR2 I92 (bcomp_0[27:27], o_0r0[27:27], o_0r1[27:27]);
  OR2 I93 (bcomp_0[28:28], o_0r0[28:28], o_0r1[28:28]);
  OR2 I94 (bcomp_0[29:29], o_0r0[29:29], o_0r1[29:29]);
  OR2 I95 (bcomp_0[30:30], o_0r0[30:30], o_0r1[30:30]);
  OR2 I96 (bcomp_0[31:31], o_0r0[31:31], o_0r1[31:31]);
  C3 I97 (simp991_0[0:0], bcomp_0[0:0], bcomp_0[1:1], bcomp_0[2:2]);
  C3 I98 (simp991_0[1:1], bcomp_0[3:3], bcomp_0[4:4], bcomp_0[5:5]);
  C3 I99 (simp991_0[2:2], bcomp_0[6:6], bcomp_0[7:7], bcomp_0[8:8]);
  C3 I100 (simp991_0[3:3], bcomp_0[9:9], bcomp_0[10:10], bcomp_0[11:11]);
  C3 I101 (simp991_0[4:4], bcomp_0[12:12], bcomp_0[13:13], bcomp_0[14:14]);
  C3 I102 (simp991_0[5:5], bcomp_0[15:15], bcomp_0[16:16], bcomp_0[17:17]);
  C3 I103 (simp991_0[6:6], bcomp_0[18:18], bcomp_0[19:19], bcomp_0[20:20]);
  C3 I104 (simp991_0[7:7], bcomp_0[21:21], bcomp_0[22:22], bcomp_0[23:23]);
  C3 I105 (simp991_0[8:8], bcomp_0[24:24], bcomp_0[25:25], bcomp_0[26:26]);
  C3 I106 (simp991_0[9:9], bcomp_0[27:27], bcomp_0[28:28], bcomp_0[29:29]);
  C2 I107 (simp991_0[10:10], bcomp_0[30:30], bcomp_0[31:31]);
  C3 I108 (simp992_0[0:0], simp991_0[0:0], simp991_0[1:1], simp991_0[2:2]);
  C3 I109 (simp992_0[1:1], simp991_0[3:3], simp991_0[4:4], simp991_0[5:5]);
  C3 I110 (simp992_0[2:2], simp991_0[6:6], simp991_0[7:7], simp991_0[8:8]);
  C2 I111 (simp992_0[3:3], simp991_0[9:9], simp991_0[10:10]);
  C3 I112 (simp993_0[0:0], simp992_0[0:0], simp992_0[1:1], simp992_0[2:2]);
  BUFF I113 (simp993_0[1:1], simp992_0[3:3]);
  C2 I114 (i_0a, simp993_0[0:0], simp993_0[1:1]);
endmodule

// latch tkl1x3 width = 1, depth = 3
module tkl1x3 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire bf_0;
  wire bt_0;
  wire ba_0;
  wire bbna_0;
  wire bbcomp_0;
  wire bof_0;
  wire bot_0;
  wire boa_0;
  wire bobna_0;
  wire bobcomp_0;
  wire boona_0;
  wire boocomp_0;
  C2R I0 (bf_0, i_0r0, bbna_0, reset);
  C2R I1 (bt_0, i_0r1, bbna_0, reset);
  INV I2 (bbna_0, ba_0);
  OR2 I3 (bbcomp_0, bf_0, bt_0);
  BUFF I4 (i_0a, bbcomp_0);
  C2R I5 (bof_0, bf_0, bobna_0, reset);
  C2R I6 (bot_0, bt_0, bobna_0, reset);
  INV I7 (bobna_0, boa_0);
  OR2 I8 (bobcomp_0, bof_0, bot_0);
  BUFF I9 (ba_0, bobcomp_0);
  C2R I10 (o_0r0, bof_0, boona_0, reset);
  C2R I11 (o_0r1, bot_0, boona_0, reset);
  INV I12 (boona_0, o_0a);
  OR2 I13 (boocomp_0, o_0r0, o_0r1);
  BUFF I14 (boa_0, boocomp_0);
endmodule

// latch tkl1x2 width = 1, depth = 2
module tkl1x2 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire bf_0;
  wire bt_0;
  wire ba_0;
  wire bbna_0;
  wire bbcomp_0;
  wire bona_0;
  wire bocomp_0;
  C2R I0 (bf_0, i_0r0, bbna_0, reset);
  C2R I1 (bt_0, i_0r1, bbna_0, reset);
  INV I2 (bbna_0, ba_0);
  OR2 I3 (bbcomp_0, bf_0, bt_0);
  BUFF I4 (i_0a, bbcomp_0);
  C2R I5 (o_0r0, bf_0, bona_0, reset);
  C2R I6 (o_0r1, bt_0, bona_0, reset);
  INV I7 (bona_0, o_0a);
  OR2 I8 (bocomp_0, o_0r0, o_0r1);
  BUFF I9 (ba_0, bocomp_0);
endmodule

module teak_Shifter (shift_0r0, shift_0r1, shift_0a, distanceI_0r0, distanceI_0r1, distanceI_0a, result_0r0, result_0r1, result_0a, arg_0r0, arg_0r1, arg_0a, reset);
  input [1:0] shift_0r0;
  input [1:0] shift_0r1;
  output shift_0a;
  input [4:0] distanceI_0r0;
  input [4:0] distanceI_0r1;
  output distanceI_0a;
  output [31:0] result_0r0;
  output [31:0] result_0r1;
  input result_0a;
  input [31:0] arg_0r0;
  input [31:0] arg_0r1;
  output arg_0a;
  input reset;
  wire L1_0r;
  wire L1_0a;
  wire [31:0] L35_0r0;
  wire [31:0] L35_0r1;
  wire L35_0a;
  wire L37P_0r;
  wire L37P_0a;
  wire L37A_0r;
  wire L37A_0a;
  wire L38_0r;
  wire L38_0a;
  wire [31:0] L72_0r0;
  wire [31:0] L72_0r1;
  wire L72_0a;
  wire L74_0r;
  wire L74_0a;
  wire L76_0r;
  wire L76_0a;
  wire [31:0] L78_0r0;
  wire [31:0] L78_0r1;
  wire L78_0a;
  wire [31:0] L80_0r0;
  wire [31:0] L80_0r1;
  wire L80_0a;
  wire [31:0] L82_0r0;
  wire [31:0] L82_0r1;
  wire L82_0a;
  wire [31:0] L84_0r0;
  wire [31:0] L84_0r1;
  wire L84_0a;
  wire [31:0] L87_0r0;
  wire [31:0] L87_0r1;
  wire L87_0a;
  wire L100_0r;
  wire L100_0a;
  wire [31:0] L106_0r0;
  wire [31:0] L106_0r1;
  wire L106_0a;
  wire [31:0] L108_0r0;
  wire [31:0] L108_0r1;
  wire L108_0a;
  wire [31:0] L110_0r0;
  wire [31:0] L110_0r1;
  wire L110_0a;
  wire [31:0] L112_0r0;
  wire [31:0] L112_0r1;
  wire L112_0a;
  wire [31:0] L113_0r0;
  wire [31:0] L113_0r1;
  wire L113_0a;
  wire L114_0r;
  wire L114_0a;
  wire [31:0] L122_0r0;
  wire [31:0] L122_0r1;
  wire L122_0a;
  wire [6:0] L129_0r0;
  wire [6:0] L129_0r1;
  wire L129_0a;
  wire [30:0] L137_0r0;
  wire [30:0] L137_0r1;
  wire L137_0a;
  wire [30:0] L138_0r0;
  wire [30:0] L138_0r1;
  wire L138_0a;
  wire [30:0] L139_0r0;
  wire [30:0] L139_0r1;
  wire L139_0a;
  wire [29:0] L140_0r0;
  wire [29:0] L140_0r1;
  wire L140_0a;
  wire [29:0] L141_0r0;
  wire [29:0] L141_0r1;
  wire L141_0a;
  wire [29:0] L142_0r0;
  wire [29:0] L142_0r1;
  wire L142_0a;
  wire L143_0r;
  wire L143_0a;
  wire L144_0r;
  wire L144_0a;
  wire L148P_0r0;
  wire L148P_0r1;
  wire L148P_0a;
  wire L148A_0r0;
  wire L148A_0r1;
  wire L148A_0a;
  wire L149_0r;
  wire L149_0a;
  wire [6:0] L151_0r0;
  wire [6:0] L151_0r1;
  wire L151_0a;
  wire L152P_0r0;
  wire L152P_0r1;
  wire L152P_0a;
  wire L152A_0r0;
  wire L152A_0r1;
  wire L152A_0a;
  wire L154P_0r;
  wire L154P_0a;
  wire L154A_0r;
  wire L154A_0a;
  wire L156_0r;
  wire L156_0a;
  wire L157_0r;
  wire L157_0a;
  wire L158_0r;
  wire L158_0a;
  wire L159_0r;
  wire L159_0a;
  wire L160_0r;
  wire L160_0a;
  wire L161_0r;
  wire L161_0a;
  wire L162_0r;
  wire L162_0a;
  wire [1:0] L175_0r0;
  wire [1:0] L175_0r1;
  wire L175_0a;
  wire [1:0] L181_0r0;
  wire [1:0] L181_0r1;
  wire L181_0a;
  wire L183_0r;
  wire L183_0a;
  wire L184_0r;
  wire L184_0a;
  wire L185_0r0;
  wire L185_0r1;
  wire L185_0a;
  wire L186_0r0;
  wire L186_0r1;
  wire L186_0a;
  wire L188_0r0;
  wire L188_0r1;
  wire L188_0a;
  wire L189_0r0;
  wire L189_0r1;
  wire L189_0a;
  tko31m32_1nm1b0_2apt1o0w1bi0w31b I0 (L137_0r0[30:0], L137_0r1[30:0], L137_0a, L108_0r0[31:0], L108_0r1[31:0], L108_0a, reset);
  tko31m32_1nm1b0_2api0w31bt1o0w1b I1 (L138_0r0[30:0], L138_0r1[30:0], L138_0a, L110_0r0[31:0], L110_0r1[31:0], L110_0a, reset);
  tko31m32_1nm1b1_2api0w31bt1o0w1b I2 (L139_0r0[30:0], L139_0r1[30:0], L139_0a, L112_0r0[31:0], L112_0r1[31:0], L112_0a, reset);
  tkvi32_wo0w32_ro0w32o0w31o1w31o1w31 I3 (L35_0r0[31:0], L35_0r1[31:0], L35_0a, L1_0r, L1_0a, L144_0r, L144_0a, L160_0r, L160_0a, L161_0r, L161_0a, L162_0r, L162_0a, L106_0r0[31:0], L106_0r1[31:0], L106_0a, L137_0r0[30:0], L137_0r1[30:0], L137_0a, L138_0r0[30:0], L138_0r1[30:0], L138_0a, L139_0r0[30:0], L139_0r1[30:0], L139_0a, reset);
  tko30m32_1nm2b0_2apt1o0w2bi0w30b I4 (L140_0r0[29:0], L140_0r1[29:0], L140_0a, L80_0r0[31:0], L80_0r1[31:0], L80_0a, reset);
  tko30m32_1nm2b0_2api0w30bt1o0w2b I5 (L141_0r0[29:0], L141_0r1[29:0], L141_0a, L82_0r0[31:0], L82_0r1[31:0], L82_0a, reset);
  tko30m32_1nm2b3_2api0w30bt1o0w2b I6 (L142_0r0[29:0], L142_0r1[29:0], L142_0a, L84_0r0[31:0], L84_0r1[31:0], L84_0a, reset);
  tkvi32_wo0w32_ro0w32o0w30o2w30o2w30 I7 (L72_0r0[31:0], L72_0r1[31:0], L72_0a, L38_0r, L38_0a, L143_0r, L143_0a, L157_0r, L157_0a, L158_0r, L158_0a, L159_0r, L159_0a, L78_0r0[31:0], L78_0r1[31:0], L78_0a, L140_0r0[29:0], L140_0r1[29:0], L140_0a, L141_0r0[29:0], L141_0r1[29:0], L141_0a, L142_0r0[29:0], L142_0r1[29:0], L142_0a, reset);
  tkj0m0_0_0 I8 (L114_0r, L114_0a, L156_0r, L156_0a, L154P_0r, L154P_0a, L76_0r, L76_0a, reset);
  tkm4x32b I9 (L78_0r0[31:0], L78_0r1[31:0], L78_0a, L80_0r0[31:0], L80_0r1[31:0], L80_0a, L82_0r0[31:0], L82_0r1[31:0], L82_0a, L84_0r0[31:0], L84_0r1[31:0], L84_0a, L87_0r0[31:0], L87_0r1[31:0], L87_0a, reset);
  tkj32m32_0 I10 (L87_0r0[31:0], L87_0r1[31:0], L87_0a, L37P_0r, L37P_0a, L35_0r0[31:0], L35_0r1[31:0], L35_0a, reset);
  tkm4x32b I11 (L106_0r0[31:0], L106_0r1[31:0], L106_0a, L108_0r0[31:0], L108_0r1[31:0], L108_0a, L110_0r0[31:0], L110_0r1[31:0], L110_0a, L112_0r0[31:0], L112_0r1[31:0], L112_0a, L113_0r0[31:0], L113_0r1[31:0], L113_0a, reset);
  tkf32mo0w0_o0w32 I12 (L113_0r0[31:0], L113_0r1[31:0], L113_0a, L114_0r, L114_0a, result_0r0[31:0], result_0r1[31:0], result_0a, reset);
  tkj32m32_0 I13 (L122_0r0[31:0], L122_0r1[31:0], L122_0a, L74_0r, L74_0a, L72_0r0[31:0], L72_0r1[31:0], L72_0a, reset);
  tkj7m5_2_0 I14 (distanceI_0r0[4:0], distanceI_0r1[4:0], distanceI_0a, shift_0r0[1:0], shift_0r1[1:0], shift_0a, L100_0r, L100_0a, L129_0r0[6:0], L129_0r1[6:0], L129_0a, reset);
  tkvdistanceIshift7_wo0w7_ro5w2o5w2 I15 (L151_0r0[6:0], L151_0r1[6:0], L151_0a, L149_0r, L149_0a, L183_0r, L183_0a, L184_0r, L184_0a, L175_0r0[1:0], L175_0r1[1:0], L175_0a, L181_0r0[1:0], L181_0r1[1:0], L181_0a, reset);
  tkf7mo0w7_o2w1_o1w1 I16 (L129_0r0[6:0], L129_0r1[6:0], L129_0a, L151_0r0[6:0], L151_0r1[6:0], L151_0a, L152A_0r0, L152A_0r1, L152A_0a, L148A_0r0, L148A_0r1, L148A_0a, reset);
  tkj1m1_0 I17 (L148P_0r0, L148P_0r1, L148P_0a, L1_0r, L1_0a, L185_0r0, L185_0r1, L185_0a, reset);
  tkj1m1_0 I18 (L152P_0r0, L152P_0r1, L152P_0a, L38_0r, L38_0a, L188_0r0, L188_0r1, L188_0a, reset);
  tkf0mo0w0_o0w0 I19 (L149_0r, L149_0a, L74_0r, L74_0a, L37A_0r, L37A_0a, reset);
  tks2_o0w2_3o0w0_0c2o0w0_1o0w0 I20 (L175_0r0[1:0], L175_0r1[1:0], L175_0a, L162_0r, L162_0a, L160_0r, L160_0a, L161_0r, L161_0a, reset);
  tks2_o0w2_3o0w0_0c2o0w0_1o0w0 I21 (L181_0r0[1:0], L181_0r1[1:0], L181_0a, L159_0r, L159_0a, L157_0r, L157_0a, L158_0r, L158_0a, reset);
  tkf1mo0w1_o0w0 I22 (L185_0r0, L185_0r1, L185_0a, L186_0r0, L186_0r1, L186_0a, L156_0r, L156_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I23 (L186_0r0, L186_0r1, L186_0a, L144_0r, L144_0a, L183_0r, L183_0a, reset);
  tkf1mo0w1_o0w0 I24 (L188_0r0, L188_0r1, L188_0a, L189_0r0, L189_0r1, L189_0a, L154A_0r, L154A_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I25 (L189_0r0, L189_0r1, L189_0a, L143_0r, L143_0a, L184_0r, L184_0a, reset);
  tki I26 (L76_0r, L76_0a, L100_0r, L100_0a, reset);
  tkl0x1 I27 (L37A_0r, L37A_0a, L37P_0r, L37P_0a, reset);
  tkl32x1 I28 (arg_0r0[31:0], arg_0r1[31:0], arg_0a, L122_0r0[31:0], L122_0r1[31:0], L122_0a, reset);
  tkl1x3 I29 (L148A_0r0, L148A_0r1, L148A_0a, L148P_0r0, L148P_0r1, L148P_0a, reset);
  tkl1x2 I30 (L152A_0r0, L152A_0r1, L152A_0a, L152P_0r0, L152P_0r1, L152P_0a, reset);
  tkl0x1 I31 (L154A_0r, L154A_0a, L154P_0r, L154P_0a, reset);
  tkr_ra_monitor #("Shifter.L1.L") I32 (L1_0r, L1_0a);
  tkr_dr_monitor #("Shifter.L35.L", 32) I33 (L35_0r0[31:0], L35_0r1[31:0], L35_0a);
  tkr_ra_monitor #("Shifter.L37.P") I34 (L37P_0r, L37P_0a);
  tkr_ra_monitor #("Shifter.L37.A") I35 (L37A_0r, L37A_0a);
  tkr_ra_monitor #("Shifter.L38.L") I36 (L38_0r, L38_0a);
  tkr_dr_monitor #("Shifter.L72.L", 32) I37 (L72_0r0[31:0], L72_0r1[31:0], L72_0a);
  tkr_ra_monitor #("Shifter.L74.L") I38 (L74_0r, L74_0a);
  tkr_ra_monitor #("Shifter.L76.L") I39 (L76_0r, L76_0a);
  tkr_dr_monitor #("Shifter.L78.L", 32) I40 (L78_0r0[31:0], L78_0r1[31:0], L78_0a);
  tkr_dr_monitor #("Shifter.L80.L", 32) I41 (L80_0r0[31:0], L80_0r1[31:0], L80_0a);
  tkr_dr_monitor #("Shifter.L82.L", 32) I42 (L82_0r0[31:0], L82_0r1[31:0], L82_0a);
  tkr_dr_monitor #("Shifter.L84.L", 32) I43 (L84_0r0[31:0], L84_0r1[31:0], L84_0a);
  tkr_dr_monitor #("Shifter.L87.L", 32) I44 (L87_0r0[31:0], L87_0r1[31:0], L87_0a);
  tkr_ra_monitor #("Shifter.L100.L") I45 (L100_0r, L100_0a);
  tkr_dr_monitor #("Shifter.L103.L", 2) I46 (shift_0r0[1:0], shift_0r1[1:0], shift_0a);
  tkr_dr_monitor #("Shifter.L104.L", 5) I47 (distanceI_0r0[4:0], distanceI_0r1[4:0], distanceI_0a);
  tkr_dr_monitor #("Shifter.L106.L", 32) I48 (L106_0r0[31:0], L106_0r1[31:0], L106_0a);
  tkr_dr_monitor #("Shifter.L108.L", 32) I49 (L108_0r0[31:0], L108_0r1[31:0], L108_0a);
  tkr_dr_monitor #("Shifter.L110.L", 32) I50 (L110_0r0[31:0], L110_0r1[31:0], L110_0a);
  tkr_dr_monitor #("Shifter.L112.L", 32) I51 (L112_0r0[31:0], L112_0r1[31:0], L112_0a);
  tkr_dr_monitor #("Shifter.L113.L", 32) I52 (L113_0r0[31:0], L113_0r1[31:0], L113_0a);
  tkr_ra_monitor #("Shifter.L114.L") I53 (L114_0r, L114_0a);
  tkr_dr_monitor #("Shifter.L115.L", 32) I54 (result_0r0[31:0], result_0r1[31:0], result_0a);
  tkr_dr_monitor #("Shifter.L122.P", 32) I55 (L122_0r0[31:0], L122_0r1[31:0], L122_0a);
  tkr_dr_monitor #("Shifter.L122.A", 32) I56 (arg_0r0[31:0], arg_0r1[31:0], arg_0a);
  tkr_dr_monitor #("Shifter.L129.L", 7) I57 (L129_0r0[6:0], L129_0r1[6:0], L129_0a);
  tkr_dr_monitor #("Shifter.L137.L", 31) I58 (L137_0r0[30:0], L137_0r1[30:0], L137_0a);
  tkr_dr_monitor #("Shifter.L138.L", 31) I59 (L138_0r0[30:0], L138_0r1[30:0], L138_0a);
  tkr_dr_monitor #("Shifter.L139.L", 31) I60 (L139_0r0[30:0], L139_0r1[30:0], L139_0a);
  tkr_dr_monitor #("Shifter.L140.L", 30) I61 (L140_0r0[29:0], L140_0r1[29:0], L140_0a);
  tkr_dr_monitor #("Shifter.L141.L", 30) I62 (L141_0r0[29:0], L141_0r1[29:0], L141_0a);
  tkr_dr_monitor #("Shifter.L142.L", 30) I63 (L142_0r0[29:0], L142_0r1[29:0], L142_0a);
  tkr_ra_monitor #("Shifter.L143.L") I64 (L143_0r, L143_0a);
  tkr_ra_monitor #("Shifter.L144.L") I65 (L144_0r, L144_0a);
  tkr_dr_monitor #("Shifter.L148.P", 1) I66 (L148P_0r0, L148P_0r1, L148P_0a);
  tkr_dr_monitor #("Shifter.L148.A", 1) I67 (L148A_0r0, L148A_0r1, L148A_0a);
  tkr_ra_monitor #("Shifter.L149.L") I68 (L149_0r, L149_0a);
  tkr_dr_monitor #("Shifter.L151.L", 7) I69 (L151_0r0[6:0], L151_0r1[6:0], L151_0a);
  tkr_dr_monitor #("Shifter.L152.P", 1) I70 (L152P_0r0, L152P_0r1, L152P_0a);
  tkr_dr_monitor #("Shifter.L152.A", 1) I71 (L152A_0r0, L152A_0r1, L152A_0a);
  tkr_ra_monitor #("Shifter.L154.P") I72 (L154P_0r, L154P_0a);
  tkr_ra_monitor #("Shifter.L154.A") I73 (L154A_0r, L154A_0a);
  tkr_ra_monitor #("Shifter.L156.L") I74 (L156_0r, L156_0a);
  tkr_ra_monitor #("Shifter.L157.L") I75 (L157_0r, L157_0a);
  tkr_ra_monitor #("Shifter.L158.L") I76 (L158_0r, L158_0a);
  tkr_ra_monitor #("Shifter.L159.L") I77 (L159_0r, L159_0a);
  tkr_ra_monitor #("Shifter.L160.L") I78 (L160_0r, L160_0a);
  tkr_ra_monitor #("Shifter.L161.L") I79 (L161_0r, L161_0a);
  tkr_ra_monitor #("Shifter.L162.L") I80 (L162_0r, L162_0a);
  tkr_dr_monitor #("Shifter.L175.L", 2) I81 (L175_0r0[1:0], L175_0r1[1:0], L175_0a);
  tkr_dr_monitor #("Shifter.L181.L", 2) I82 (L181_0r0[1:0], L181_0r1[1:0], L181_0a);
  tkr_ra_monitor #("Shifter.L183.L") I83 (L183_0r, L183_0a);
  tkr_ra_monitor #("Shifter.L184.L") I84 (L184_0r, L184_0a);
  tkr_dr_monitor #("Shifter.L185.L", 1) I85 (L185_0r0, L185_0r1, L185_0a);
  tkr_dr_monitor #("Shifter.L186.L", 1) I86 (L186_0r0, L186_0r1, L186_0a);
  tkr_dr_monitor #("Shifter.L188.L", 1) I87 (L188_0r0, L188_0r1, L188_0a);
  tkr_dr_monitor #("Shifter.L189.L", 1) I88 (L189_0r0, L189_0r1, L189_0a);
endmodule

// Netlist costs:
// teak_Shifter: AND2*1370 AO22*77 BUFF*1081 C2*84 C2R*92 C3*279 GND*9 INV*145 NAND2*131 NAND3*2 NOR2*78 NOR3*206 OR2*560 OR3*2
// tkf0mo0w0_o0w0: BUFF*2 C2*1
// tkf1mo0w1_o0w0: BUFF*4 C3*1 OR2*1
// tkf32mo0w0_o0w32: BUFF*66 C3*1 OR2*1
// tkf7mo0w7_o2w1_o1w1: BUFF*16 C2*5 C3*1 OR2*1
// tki: AND2*1 AO22*3 INV*3
// tkj0m0_0_0: BUFF*3 C3*1
// tkj1m1_0: BUFF*5 C2*2
// tkj32m32_0: BUFF*129 C2*2
// tkj7m5_2_0: BUFF*29 C2*3 OR2*1
// tkl0x1: BUFF*1 C2R*1 INV*1
// tkl1x2: BUFF*2 C2R*4 INV*2 OR2*2
// tkl1x3: BUFF*3 C2R*6 INV*3 OR2*3
// tkl32x1: BUFF*1 C2*3 C2R*64 C3*14 INV*1 OR2*32
// tkm4x32b: AND2*256 BUFF*4 C2*12 C2R*8 C3*56 INV*65 NAND2*65 NOR2*1 NOR3*65 OR2*128
// tko30m32_1nm2b0_2api0w30bt1o0w2b: BUFF*69 C2*1 C3*14 GND*2 OR2*30
// tko30m32_1nm2b0_2apt1o0w2bi0w30b: BUFF*69 C2*1 C3*14 GND*2 OR2*30
// tko30m32_1nm2b3_2api0w30bt1o0w2b: BUFF*69 C2*1 C3*14 GND*2 OR2*30
// tko31m32_1nm1b0_2api0w31bt1o0w1b: BUFF*68 C2*2 C3*14 GND*1 OR2*31
// tko31m32_1nm1b0_2apt1o0w1bi0w31b: BUFF*68 C2*2 C3*14 GND*1 OR2*31
// tko31m32_1nm1b1_2api0w31bt1o0w1b: BUFF*68 C2*2 C3*14 GND*1 OR2*31
// tks1_o0w1_0o0w0_1o0w0: BUFF*7 C2*3 OR2*2
// tks2_o0w2_3o0w0_0c2o0w0_1o0w0: BUFF*7 C2*7 OR2*2 OR3*1
// tkvdistanceIshift7_wo0w7_ro5w2o5w2: AND2*43 AO22*8 BUFF*26 C2*1 C3*6 INV*2 NAND2*1 NOR2*8 NOR3*8 OR2*7
// tkvi32_wo0w32_ro0w32o0w30o2w30o2w30: AND2*404 AO22*33 BUFF*104 C2*5 C3*29 INV*1 NAND3*1 NOR2*34 NOR3*34 OR2*32
// tkvi32_wo0w32_ro0w32o0w31o1w31o1w31: AND2*410 AO22*33 BUFF*104 C2*5 C3*29 INV*1 NAND3*1 NOR2*34 NOR3*34 OR2*32
