//
// by teak gui
//
// Generated on: Thu Feb  7 11:25:01 GMT 2013
//


`timescale 1ns/1ps

// tko0m1_1nm1b0 TeakO [
//     (1,TeakOConstant 1 0)] [One 0,One 1]
module tko0m1_1nm1b0 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0, i_0r);
  GND I1 (o_0r1);
  BUFF I2 (i_0a, o_0a);
endmodule

// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0 TeakF [0,0,0,0,0,0] [One 0,Many [0,0,0,0,0,0]]
module tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, o_5r, o_5a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  input reset;
  wire [1:0] simp11_0;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  BUFF I2 (o_2r, i_0r);
  BUFF I3 (o_3r, i_0r);
  BUFF I4 (o_4r, i_0r);
  BUFF I5 (o_5r, i_0r);
  C3 I6 (simp11_0[0:0], o_0a, o_1a, o_2a);
  C3 I7 (simp11_0[1:1], o_3a, o_4a, o_5a);
  C2 I8 (i_0a, simp11_0[0:0], simp11_0[1:1]);
endmodule

// tkj0m0_0_0 TeakJ [Many [0,0,0],One 0]
module tkj0m0_0_0 (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  output o_0r;
  input o_0a;
  input reset;
  C3 I0 (o_0r, i_0r, i_1r, i_2r);
  BUFF I1 (i_0a, o_0a);
  BUFF I2 (i_1a, o_0a);
  BUFF I3 (i_2a, o_0a);
endmodule

// tko1m1_1noti0w1b TeakO [
//     (1,TeakOp TeakOpNot [(0,0+:1)])] [One 1,One 1]
module tko1m1_1noti0w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1, i_0r0);
  BUFF I1 (o_0r0, i_0r1);
  BUFF I2 (i_0a, o_0a);
endmodule

// tko0m5_1nm5b1 TeakO [
//     (1,TeakOConstant 5 1)] [One 0,One 5]
module tko0m5_1nm5b1 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [4:0] o_0r0;
  output [4:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  GND I1 (o_0r0[0:0]);
  BUFF I2 (o_0r0[1:1], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  GND I6 (o_0r1[1:1]);
  GND I7 (o_0r1[2:2]);
  GND I8 (o_0r1[3:3]);
  GND I9 (o_0r1[4:4]);
  BUFF I10 (i_0a, o_0a);
endmodule

// tko0m1_1nm1b1 TeakO [
//     (1,TeakOConstant 1 1)] [One 0,One 1]
module tko0m1_1nm1b1 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1, i_0r);
  GND I1 (o_0r0);
  BUFF I2 (i_0a, o_0a);
endmodule

// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0 TeakF [0,0,0,0,0] [One 0,Many [0,0,0,0,0]]
module tkf0mo0w0_o0w0_o0w0_o0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  input reset;
  wire [1:0] simp11_0;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  BUFF I2 (o_2r, i_0r);
  BUFF I3 (o_3r, i_0r);
  BUFF I4 (o_4r, i_0r);
  C3 I5 (simp11_0[0:0], o_0a, o_1a, o_2a);
  C2 I6 (simp11_0[1:1], o_3a, o_4a);
  C2 I7 (i_0a, simp11_0[0:0], simp11_0[1:1]);
endmodule

// tks1_o0w1_0o0w0_1o0w0 TeakS (0+:1) [([Imp 0 0],0),([Imp 1 0],0)] [One 1,Many [0,0]]
module tks1_o0w1_0o0w0_1o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire comp_0;
  BUFF I0 (sel_0, match0_0);
  BUFF I1 (match0_0, i_0r0);
  BUFF I2 (sel_1, match1_0);
  BUFF I3 (match1_0, i_0r1);
  C2 I4 (gsel_0, sel_0, icomplete_0);
  C2 I5 (gsel_1, sel_1, icomplete_0);
  OR2 I6 (comp_0, i_0r0, i_0r1);
  BUFF I7 (icomplete_0, comp_0);
  BUFF I8 (o_0r, gsel_0);
  BUFF I9 (o_1r, gsel_1);
  OR2 I10 (oack_0, o_0a, o_1a);
  C2 I11 (i_0a, oack_0, icomplete_0);
endmodule

// tks3_o0w3_2o0w0_3o0w0_4c1o0w0_6o0w0_7o0w0_0m1o0w3 TeakS (0+:3) [([Imp 2 0],0),([Imp 3 0],0),([Imp 4 
//   1],0),([Imp 6 0],0),([Imp 7 0],0),([Imp 0 0,Imp 1 0],0)] [One 3,Many [0,0,0,0,0,3]]
module tks3_o0w3_2o0w0_3o0w0_4c1o0w0_6o0w0_7o0w0_0m1o0w3 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, o_5r0, o_5r1, o_5a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output [2:0] o_5r0;
  output [2:0] o_5r1;
  input o_5a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire sel_4;
  wire sel_5;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire gsel_4;
  wire gsel_5;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire match2_0;
  wire match3_0;
  wire match4_0;
  wire [1:0] match5_0;
  wire [2:0] comp_0;
  wire [1:0] simp551_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (match0_0, i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I2 (sel_1, match1_0);
  C3 I3 (match1_0, i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I4 (sel_2, match2_0);
  C2 I5 (match2_0, i_0r0[1:1], i_0r1[2:2]);
  BUFF I6 (sel_3, match3_0);
  C3 I7 (match3_0, i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I8 (sel_4, match4_0);
  C3 I9 (match4_0, i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  OR2 I10 (sel_5, match5_0[0:0], match5_0[1:1]);
  C3 I11 (match5_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I12 (match5_0[1:1], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C2 I13 (gsel_0, sel_0, icomplete_0);
  C2 I14 (gsel_1, sel_1, icomplete_0);
  C2 I15 (gsel_2, sel_2, icomplete_0);
  C2 I16 (gsel_3, sel_3, icomplete_0);
  C2 I17 (gsel_4, sel_4, icomplete_0);
  C2 I18 (gsel_5, sel_5, icomplete_0);
  OR2 I19 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I20 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I21 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I22 (icomplete_0, comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C2 I23 (o_5r0[0:0], i_0r0[0:0], gsel_5);
  C2 I24 (o_5r0[1:1], i_0r0[1:1], gsel_5);
  C2 I25 (o_5r0[2:2], i_0r0[2:2], gsel_5);
  C2 I26 (o_5r1[0:0], i_0r1[0:0], gsel_5);
  C2 I27 (o_5r1[1:1], i_0r1[1:1], gsel_5);
  C2 I28 (o_5r1[2:2], i_0r1[2:2], gsel_5);
  BUFF I29 (o_0r, gsel_0);
  BUFF I30 (o_1r, gsel_1);
  BUFF I31 (o_2r, gsel_2);
  BUFF I32 (o_3r, gsel_3);
  BUFF I33 (o_4r, gsel_4);
  NOR3 I34 (simp551_0[0:0], o_0a, o_1a, o_2a);
  NOR3 I35 (simp551_0[1:1], o_3a, o_4a, o_5a);
  NAND2 I36 (oack_0, simp551_0[0:0], simp551_0[1:1]);
  C2 I37 (i_0a, oack_0, icomplete_0);
endmodule

// tkm6x0b TeakM [Many [0,0,0,0,0,0],One 0]
module tkm6x0b (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, i_3r, i_3a, i_4r, i_4a, i_5r, i_5a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  input i_4r;
  output i_4a;
  input i_5r;
  output i_5a;
  output o_0r;
  input o_0a;
  input reset;
  wire nchosen_0;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire choice_4;
  wire choice_5;
  wire [1:0] simp141_0;
  C2R I0 (choice_0, i_0r, nchosen_0, reset);
  C2R I1 (choice_1, i_1r, nchosen_0, reset);
  C2R I2 (choice_2, i_2r, nchosen_0, reset);
  C2R I3 (choice_3, i_3r, nchosen_0, reset);
  C2R I4 (choice_4, i_4r, nchosen_0, reset);
  C2R I5 (choice_5, i_5r, nchosen_0, reset);
  NOR2 I6 (nchosen_0, o_0r, o_0a);
  NOR3 I7 (simp141_0[0:0], choice_0, choice_1, choice_2);
  NOR3 I8 (simp141_0[1:1], choice_3, choice_4, choice_5);
  NAND2 I9 (o_0r, simp141_0[0:0], simp141_0[1:1]);
  C2R I10 (i_0a, choice_0, o_0a, reset);
  C2R I11 (i_1a, choice_1, o_0a, reset);
  C2R I12 (i_2a, choice_2, o_0a, reset);
  C2R I13 (i_3a, choice_3, o_0a, reset);
  C2R I14 (i_4a, choice_4, o_0a, reset);
  C2R I15 (i_5a, choice_5, o_0a, reset);
endmodule

// tkm2x0b TeakM [Many [0,0],One 0]
module tkm2x0b (i_0r, i_0a, i_1r, i_1a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  output o_0r;
  input o_0a;
  input reset;
  wire nchosen_0;
  wire choice_0;
  wire choice_1;
  C2R I0 (choice_0, i_0r, nchosen_0, reset);
  C2R I1 (choice_1, i_1r, nchosen_0, reset);
  NOR2 I2 (nchosen_0, o_0r, o_0a);
  OR2 I3 (o_0r, choice_0, choice_1);
  C2R I4 (i_0a, choice_0, o_0a, reset);
  C2R I5 (i_1a, choice_1, o_0a, reset);
endmodule

// tkj0m0_0 TeakJ [Many [0,0],One 0]
module tkj0m0_0 (i_0r, i_0a, i_1r, i_1a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  output o_0r;
  input o_0a;
  input reset;
  C2 I0 (o_0r, i_0r, i_1r);
  BUFF I1 (i_0a, o_0a);
  BUFF I2 (i_1a, o_0a);
endmodule

// tkj10m5_5 TeakJ [Many [5,5],One 10]
module tkj10m5_5 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [4:0] i_0r0;
  input [4:0] i_0r1;
  output i_0a;
  input [4:0] i_1r0;
  input [4:0] i_1r1;
  output i_1a;
  output [9:0] o_0r0;
  output [9:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [9:0] joinf_0;
  wire [9:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_1r0[0:0]);
  BUFF I6 (joinf_0[6:6], i_1r0[1:1]);
  BUFF I7 (joinf_0[7:7], i_1r0[2:2]);
  BUFF I8 (joinf_0[8:8], i_1r0[3:3]);
  BUFF I9 (joinf_0[9:9], i_1r0[4:4]);
  BUFF I10 (joint_0[0:0], i_0r1[0:0]);
  BUFF I11 (joint_0[1:1], i_0r1[1:1]);
  BUFF I12 (joint_0[2:2], i_0r1[2:2]);
  BUFF I13 (joint_0[3:3], i_0r1[3:3]);
  BUFF I14 (joint_0[4:4], i_0r1[4:4]);
  BUFF I15 (joint_0[5:5], i_1r1[0:0]);
  BUFF I16 (joint_0[6:6], i_1r1[1:1]);
  BUFF I17 (joint_0[7:7], i_1r1[2:2]);
  BUFF I18 (joint_0[8:8], i_1r1[3:3]);
  BUFF I19 (joint_0[9:9], i_1r1[4:4]);
  OR2 I20 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I21 (icomplete_0, dcomplete_0);
  C2 I22 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I23 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I24 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I25 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I26 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I27 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I28 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I29 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I30 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I31 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I32 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I33 (o_0r1[1:1], joint_0[1:1]);
  BUFF I34 (o_0r1[2:2], joint_0[2:2]);
  BUFF I35 (o_0r1[3:3], joint_0[3:3]);
  BUFF I36 (o_0r1[4:4], joint_0[4:4]);
  BUFF I37 (o_0r1[5:5], joint_0[5:5]);
  BUFF I38 (o_0r1[6:6], joint_0[6:6]);
  BUFF I39 (o_0r1[7:7], joint_0[7:7]);
  BUFF I40 (o_0r1[8:8], joint_0[8:8]);
  BUFF I41 (o_0r1[9:9], joint_0[9:9]);
  BUFF I42 (i_0a, o_0a);
  BUFF I43 (i_1a, o_0a);
endmodule

// tko10m6_1nm1b0_2api0w5bt1o0w1b_3nm1b0_4api5w5bt3o0w1b_5addt2o0w6bt4o0w6b TeakO [
//     (1,TeakOConstant 1 0),
//     (2,TeakOAppend 1 [(0,0+:5),(1,0+:1)]),
//     (3,TeakOConstant 1 0),
//     (4,TeakOAppend 1 [(0,5+:5),(3,0+:1)]),
//     (5,TeakOp TeakOpAdd [(2,0+:6),(4,0+:6)])] [One 10,One 6]
module tko10m6_1nm1b0_2api0w5bt1o0w1b_3nm1b0_4api5w5bt3o0w1b_5addt2o0w6bt4o0w6b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [9:0] i_0r0;
  input [9:0] i_0r1;
  output i_0a;
  output [5:0] o_0r0;
  output [5:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [9:0] gocomp_0;
  wire [3:0] simp121_0;
  wire [1:0] simp122_0;
  wire termf_1;
  wire [5:0] termf_2;
  wire termf_3;
  wire [5:0] termf_4;
  wire termt_1;
  wire [5:0] termt_2;
  wire termt_3;
  wire [5:0] termt_4;
  wire [5:0] cf5__0;
  wire [5:0] ct5__0;
  wire [3:0] ha5__0;
  wire [7:0] fa5_1min_0;
  wire [1:0] simp711_0;
  wire [1:0] simp721_0;
  wire [7:0] fa5_2min_0;
  wire [1:0] simp841_0;
  wire [1:0] simp851_0;
  wire [7:0] fa5_3min_0;
  wire [1:0] simp971_0;
  wire [1:0] simp981_0;
  wire [7:0] fa5_4min_0;
  wire [1:0] simp1101_0;
  wire [1:0] simp1111_0;
  wire [7:0] fa5_5min_0;
  wire [1:0] simp1231_0;
  wire [1:0] simp1241_0;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  C3 I10 (simp121_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  C3 I11 (simp121_0[1:1], gocomp_0[3:3], gocomp_0[4:4], gocomp_0[5:5]);
  C3 I12 (simp121_0[2:2], gocomp_0[6:6], gocomp_0[7:7], gocomp_0[8:8]);
  BUFF I13 (simp121_0[3:3], gocomp_0[9:9]);
  C3 I14 (simp122_0[0:0], simp121_0[0:0], simp121_0[1:1], simp121_0[2:2]);
  BUFF I15 (simp122_0[1:1], simp121_0[3:3]);
  C2 I16 (go_0, simp122_0[0:0], simp122_0[1:1]);
  BUFF I17 (termf_1, go_0);
  GND I18 (termt_1);
  BUFF I19 (termf_2[0:0], i_0r0[0:0]);
  BUFF I20 (termf_2[1:1], i_0r0[1:1]);
  BUFF I21 (termf_2[2:2], i_0r0[2:2]);
  BUFF I22 (termf_2[3:3], i_0r0[3:3]);
  BUFF I23 (termf_2[4:4], i_0r0[4:4]);
  BUFF I24 (termf_2[5:5], termf_1);
  BUFF I25 (termt_2[0:0], i_0r1[0:0]);
  BUFF I26 (termt_2[1:1], i_0r1[1:1]);
  BUFF I27 (termt_2[2:2], i_0r1[2:2]);
  BUFF I28 (termt_2[3:3], i_0r1[3:3]);
  BUFF I29 (termt_2[4:4], i_0r1[4:4]);
  BUFF I30 (termt_2[5:5], termt_1);
  BUFF I31 (termf_3, go_0);
  GND I32 (termt_3);
  BUFF I33 (termf_4[0:0], i_0r0[5:5]);
  BUFF I34 (termf_4[1:1], i_0r0[6:6]);
  BUFF I35 (termf_4[2:2], i_0r0[7:7]);
  BUFF I36 (termf_4[3:3], i_0r0[8:8]);
  BUFF I37 (termf_4[4:4], i_0r0[9:9]);
  BUFF I38 (termf_4[5:5], termf_3);
  BUFF I39 (termt_4[0:0], i_0r1[5:5]);
  BUFF I40 (termt_4[1:1], i_0r1[6:6]);
  BUFF I41 (termt_4[2:2], i_0r1[7:7]);
  BUFF I42 (termt_4[3:3], i_0r1[8:8]);
  BUFF I43 (termt_4[4:4], i_0r1[9:9]);
  BUFF I44 (termt_4[5:5], termt_3);
  C2 I45 (ha5__0[0:0], termf_4[0:0], termf_2[0:0]);
  C2 I46 (ha5__0[1:1], termf_4[0:0], termt_2[0:0]);
  C2 I47 (ha5__0[2:2], termt_4[0:0], termf_2[0:0]);
  C2 I48 (ha5__0[3:3], termt_4[0:0], termt_2[0:0]);
  OR3 I49 (cf5__0[0:0], ha5__0[0:0], ha5__0[1:1], ha5__0[2:2]);
  BUFF I50 (ct5__0[0:0], ha5__0[3:3]);
  OR2 I51 (o_0r0[0:0], ha5__0[0:0], ha5__0[3:3]);
  OR2 I52 (o_0r1[0:0], ha5__0[1:1], ha5__0[2:2]);
  C3 I53 (fa5_1min_0[0:0], cf5__0[0:0], termf_4[1:1], termf_2[1:1]);
  C3 I54 (fa5_1min_0[1:1], cf5__0[0:0], termf_4[1:1], termt_2[1:1]);
  C3 I55 (fa5_1min_0[2:2], cf5__0[0:0], termt_4[1:1], termf_2[1:1]);
  C3 I56 (fa5_1min_0[3:3], cf5__0[0:0], termt_4[1:1], termt_2[1:1]);
  C3 I57 (fa5_1min_0[4:4], ct5__0[0:0], termf_4[1:1], termf_2[1:1]);
  C3 I58 (fa5_1min_0[5:5], ct5__0[0:0], termf_4[1:1], termt_2[1:1]);
  C3 I59 (fa5_1min_0[6:6], ct5__0[0:0], termt_4[1:1], termf_2[1:1]);
  C3 I60 (fa5_1min_0[7:7], ct5__0[0:0], termt_4[1:1], termt_2[1:1]);
  NOR3 I61 (simp711_0[0:0], fa5_1min_0[0:0], fa5_1min_0[3:3], fa5_1min_0[5:5]);
  INV I62 (simp711_0[1:1], fa5_1min_0[6:6]);
  NAND2 I63 (o_0r0[1:1], simp711_0[0:0], simp711_0[1:1]);
  NOR3 I64 (simp721_0[0:0], fa5_1min_0[1:1], fa5_1min_0[2:2], fa5_1min_0[4:4]);
  INV I65 (simp721_0[1:1], fa5_1min_0[7:7]);
  NAND2 I66 (o_0r1[1:1], simp721_0[0:0], simp721_0[1:1]);
  AO222 I67 (ct5__0[1:1], termt_2[1:1], termt_4[1:1], termt_2[1:1], ct5__0[0:0], termt_4[1:1], ct5__0[0:0]);
  AO222 I68 (cf5__0[1:1], termf_2[1:1], termf_4[1:1], termf_2[1:1], cf5__0[0:0], termf_4[1:1], cf5__0[0:0]);
  C3 I69 (fa5_2min_0[0:0], cf5__0[1:1], termf_4[2:2], termf_2[2:2]);
  C3 I70 (fa5_2min_0[1:1], cf5__0[1:1], termf_4[2:2], termt_2[2:2]);
  C3 I71 (fa5_2min_0[2:2], cf5__0[1:1], termt_4[2:2], termf_2[2:2]);
  C3 I72 (fa5_2min_0[3:3], cf5__0[1:1], termt_4[2:2], termt_2[2:2]);
  C3 I73 (fa5_2min_0[4:4], ct5__0[1:1], termf_4[2:2], termf_2[2:2]);
  C3 I74 (fa5_2min_0[5:5], ct5__0[1:1], termf_4[2:2], termt_2[2:2]);
  C3 I75 (fa5_2min_0[6:6], ct5__0[1:1], termt_4[2:2], termf_2[2:2]);
  C3 I76 (fa5_2min_0[7:7], ct5__0[1:1], termt_4[2:2], termt_2[2:2]);
  NOR3 I77 (simp841_0[0:0], fa5_2min_0[0:0], fa5_2min_0[3:3], fa5_2min_0[5:5]);
  INV I78 (simp841_0[1:1], fa5_2min_0[6:6]);
  NAND2 I79 (o_0r0[2:2], simp841_0[0:0], simp841_0[1:1]);
  NOR3 I80 (simp851_0[0:0], fa5_2min_0[1:1], fa5_2min_0[2:2], fa5_2min_0[4:4]);
  INV I81 (simp851_0[1:1], fa5_2min_0[7:7]);
  NAND2 I82 (o_0r1[2:2], simp851_0[0:0], simp851_0[1:1]);
  AO222 I83 (ct5__0[2:2], termt_2[2:2], termt_4[2:2], termt_2[2:2], ct5__0[1:1], termt_4[2:2], ct5__0[1:1]);
  AO222 I84 (cf5__0[2:2], termf_2[2:2], termf_4[2:2], termf_2[2:2], cf5__0[1:1], termf_4[2:2], cf5__0[1:1]);
  C3 I85 (fa5_3min_0[0:0], cf5__0[2:2], termf_4[3:3], termf_2[3:3]);
  C3 I86 (fa5_3min_0[1:1], cf5__0[2:2], termf_4[3:3], termt_2[3:3]);
  C3 I87 (fa5_3min_0[2:2], cf5__0[2:2], termt_4[3:3], termf_2[3:3]);
  C3 I88 (fa5_3min_0[3:3], cf5__0[2:2], termt_4[3:3], termt_2[3:3]);
  C3 I89 (fa5_3min_0[4:4], ct5__0[2:2], termf_4[3:3], termf_2[3:3]);
  C3 I90 (fa5_3min_0[5:5], ct5__0[2:2], termf_4[3:3], termt_2[3:3]);
  C3 I91 (fa5_3min_0[6:6], ct5__0[2:2], termt_4[3:3], termf_2[3:3]);
  C3 I92 (fa5_3min_0[7:7], ct5__0[2:2], termt_4[3:3], termt_2[3:3]);
  NOR3 I93 (simp971_0[0:0], fa5_3min_0[0:0], fa5_3min_0[3:3], fa5_3min_0[5:5]);
  INV I94 (simp971_0[1:1], fa5_3min_0[6:6]);
  NAND2 I95 (o_0r0[3:3], simp971_0[0:0], simp971_0[1:1]);
  NOR3 I96 (simp981_0[0:0], fa5_3min_0[1:1], fa5_3min_0[2:2], fa5_3min_0[4:4]);
  INV I97 (simp981_0[1:1], fa5_3min_0[7:7]);
  NAND2 I98 (o_0r1[3:3], simp981_0[0:0], simp981_0[1:1]);
  AO222 I99 (ct5__0[3:3], termt_2[3:3], termt_4[3:3], termt_2[3:3], ct5__0[2:2], termt_4[3:3], ct5__0[2:2]);
  AO222 I100 (cf5__0[3:3], termf_2[3:3], termf_4[3:3], termf_2[3:3], cf5__0[2:2], termf_4[3:3], cf5__0[2:2]);
  C3 I101 (fa5_4min_0[0:0], cf5__0[3:3], termf_4[4:4], termf_2[4:4]);
  C3 I102 (fa5_4min_0[1:1], cf5__0[3:3], termf_4[4:4], termt_2[4:4]);
  C3 I103 (fa5_4min_0[2:2], cf5__0[3:3], termt_4[4:4], termf_2[4:4]);
  C3 I104 (fa5_4min_0[3:3], cf5__0[3:3], termt_4[4:4], termt_2[4:4]);
  C3 I105 (fa5_4min_0[4:4], ct5__0[3:3], termf_4[4:4], termf_2[4:4]);
  C3 I106 (fa5_4min_0[5:5], ct5__0[3:3], termf_4[4:4], termt_2[4:4]);
  C3 I107 (fa5_4min_0[6:6], ct5__0[3:3], termt_4[4:4], termf_2[4:4]);
  C3 I108 (fa5_4min_0[7:7], ct5__0[3:3], termt_4[4:4], termt_2[4:4]);
  NOR3 I109 (simp1101_0[0:0], fa5_4min_0[0:0], fa5_4min_0[3:3], fa5_4min_0[5:5]);
  INV I110 (simp1101_0[1:1], fa5_4min_0[6:6]);
  NAND2 I111 (o_0r0[4:4], simp1101_0[0:0], simp1101_0[1:1]);
  NOR3 I112 (simp1111_0[0:0], fa5_4min_0[1:1], fa5_4min_0[2:2], fa5_4min_0[4:4]);
  INV I113 (simp1111_0[1:1], fa5_4min_0[7:7]);
  NAND2 I114 (o_0r1[4:4], simp1111_0[0:0], simp1111_0[1:1]);
  AO222 I115 (ct5__0[4:4], termt_2[4:4], termt_4[4:4], termt_2[4:4], ct5__0[3:3], termt_4[4:4], ct5__0[3:3]);
  AO222 I116 (cf5__0[4:4], termf_2[4:4], termf_4[4:4], termf_2[4:4], cf5__0[3:3], termf_4[4:4], cf5__0[3:3]);
  C3 I117 (fa5_5min_0[0:0], cf5__0[4:4], termf_4[5:5], termf_2[5:5]);
  C3 I118 (fa5_5min_0[1:1], cf5__0[4:4], termf_4[5:5], termt_2[5:5]);
  C3 I119 (fa5_5min_0[2:2], cf5__0[4:4], termt_4[5:5], termf_2[5:5]);
  C3 I120 (fa5_5min_0[3:3], cf5__0[4:4], termt_4[5:5], termt_2[5:5]);
  C3 I121 (fa5_5min_0[4:4], ct5__0[4:4], termf_4[5:5], termf_2[5:5]);
  C3 I122 (fa5_5min_0[5:5], ct5__0[4:4], termf_4[5:5], termt_2[5:5]);
  C3 I123 (fa5_5min_0[6:6], ct5__0[4:4], termt_4[5:5], termf_2[5:5]);
  C3 I124 (fa5_5min_0[7:7], ct5__0[4:4], termt_4[5:5], termt_2[5:5]);
  NOR3 I125 (simp1231_0[0:0], fa5_5min_0[0:0], fa5_5min_0[3:3], fa5_5min_0[5:5]);
  INV I126 (simp1231_0[1:1], fa5_5min_0[6:6]);
  NAND2 I127 (o_0r0[5:5], simp1231_0[0:0], simp1231_0[1:1]);
  NOR3 I128 (simp1241_0[0:0], fa5_5min_0[1:1], fa5_5min_0[2:2], fa5_5min_0[4:4]);
  INV I129 (simp1241_0[1:1], fa5_5min_0[7:7]);
  NAND2 I130 (o_0r1[5:5], simp1241_0[0:0], simp1241_0[1:1]);
  AO222 I131 (ct5__0[5:5], termt_2[5:5], termt_4[5:5], termt_2[5:5], ct5__0[4:4], termt_4[5:5], ct5__0[4:4]);
  AO222 I132 (cf5__0[5:5], termf_2[5:5], termf_4[5:5], termf_2[5:5], cf5__0[4:4], termf_4[5:5], cf5__0[4:4]);
  BUFF I133 (i_0a, o_0a);
endmodule

// tkf6mo0w0_o0w5 TeakF [0,0] [One 6,Many [0,5]]
module tkf6mo0w0_o0w5 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [5:0] i_0r0;
  input [5:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [4:0] o_1r0;
  output [4:0] o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  wire ucomplete_0;
  wire comp_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (comp_0, i_0r0[5:5], i_0r1[5:5]);
  BUFF I2 (ucomplete_0, comp_0);
  C2 I3 (acomplete_0, ucomplete_0, icomplete_0);
  C2 I4 (o_1r0[0:0], i_0r0[0:0], icomplete_0);
  BUFF I5 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I6 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I7 (o_1r0[3:3], i_0r0[3:3]);
  BUFF I8 (o_1r0[4:4], i_0r0[4:4]);
  C2 I9 (o_1r1[0:0], i_0r1[0:0], icomplete_0);
  BUFF I10 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I11 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I12 (o_1r1[3:3], i_0r1[3:3]);
  BUFF I13 (o_1r1[4:4], i_0r1[4:4]);
  BUFF I14 (o_0r, icomplete_0);
  C3 I15 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tkf0mo0w0_o0w0 TeakF [0,0] [One 0,Many [0,0]]
module tkf0mo0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  C2 I2 (i_0a, o_0a, o_1a);
endmodule

// tko0m3_1nm3b2 TeakO [
//     (1,TeakOConstant 3 2)] [One 0,One 3]
module tko0m3_1nm3b2 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[1:1], i_0r);
  GND I1 (o_0r0[1:1]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  GND I4 (o_0r1[0:0]);
  GND I5 (o_0r1[2:2]);
  BUFF I6 (i_0a, o_0a);
endmodule

// tkm2x3b TeakM [Many [3,3],One 3]
module tkm2x3b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  input [2:0] i_1r0;
  input [2:0] i_1r1;
  output i_1a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire [2:0] gfint_0;
  wire [2:0] gfint_1;
  wire [2:0] gtint_0;
  wire [2:0] gtint_1;
  wire choice_0;
  wire choice_1;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire nchosen_0;
  wire [2:0] comp0_0;
  wire [2:0] comp1_0;
  OR2 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0]);
  OR2 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1]);
  OR2 I2 (o_0r0[2:2], gfint_0[2:2], gfint_1[2:2]);
  OR2 I3 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0]);
  OR2 I4 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1]);
  OR2 I5 (o_0r1[2:2], gtint_0[2:2], gtint_1[2:2]);
  AND2 I6 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I7 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I8 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I9 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I10 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I11 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I12 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I13 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I14 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I15 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I16 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I17 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  OR2 I18 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I19 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I20 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I21 (icomp_0, comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  OR2 I22 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I23 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I24 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  C3 I25 (icomp_1, comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C2R I26 (choice_0, icomp_0, nchosen_0, reset);
  C2R I27 (choice_1, icomp_1, nchosen_0, reset);
  OR2 I28 (anychoice_0, choice_0, choice_1);
  NOR2 I29 (nchosen_0, anychoice_0, o_0a);
  C2R I30 (i_0a, choice_0, o_0a, reset);
  C2R I31 (i_1a, choice_1, o_0a, reset);
endmodule

// tkj3m0_3 TeakJ [Many [0,3],One 3]
module tkj3m0_3 (i_0r, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  input [2:0] i_1r0;
  input [2:0] i_1r1;
  output i_1a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [2:0] joinf_0;
  wire [2:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_1r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_1r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_1r0[2:2]);
  BUFF I3 (joint_0[0:0], i_1r1[0:0]);
  BUFF I4 (joint_0[1:1], i_1r1[1:1]);
  BUFF I5 (joint_0[2:2], i_1r1[2:2]);
  BUFF I6 (icomplete_0, i_0r);
  C2 I7 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I8 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I9 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I10 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I11 (o_0r1[1:1], joint_0[1:1]);
  BUFF I12 (o_0r1[2:2], joint_0[2:2]);
  BUFF I13 (i_0a, o_0a);
  BUFF I14 (i_1a, o_0a);
endmodule

// tks3_o0w3_1o0w0_2o0w0_4o0w0 TeakS (0+:3) [([Imp 1 0],0),([Imp 2 0],0),([Imp 4 0],0)] [One 3,Many [0,
//   0,0]]
module tks3_o0w3_1o0w0_2o0w0_4o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire match2_0;
  wire [2:0] comp_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (match0_0, i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I2 (sel_1, match1_0);
  C3 I3 (match1_0, i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I4 (sel_2, match2_0);
  C3 I5 (match2_0, i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C2 I6 (gsel_0, sel_0, icomplete_0);
  C2 I7 (gsel_1, sel_1, icomplete_0);
  C2 I8 (gsel_2, sel_2, icomplete_0);
  OR2 I9 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I10 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I11 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I12 (icomplete_0, comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  BUFF I13 (o_0r, gsel_0);
  BUFF I14 (o_1r, gsel_1);
  BUFF I15 (o_2r, gsel_2);
  OR3 I16 (oack_0, o_0a, o_1a, o_2a);
  C2 I17 (i_0a, oack_0, icomplete_0);
endmodule

// tkj64m32_32 TeakJ [Many [32,32],One 64]
module tkj64m32_32 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  output [63:0] o_0r0;
  output [63:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [63:0] joinf_0;
  wire [63:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joinf_0[32:32], i_1r0[0:0]);
  BUFF I33 (joinf_0[33:33], i_1r0[1:1]);
  BUFF I34 (joinf_0[34:34], i_1r0[2:2]);
  BUFF I35 (joinf_0[35:35], i_1r0[3:3]);
  BUFF I36 (joinf_0[36:36], i_1r0[4:4]);
  BUFF I37 (joinf_0[37:37], i_1r0[5:5]);
  BUFF I38 (joinf_0[38:38], i_1r0[6:6]);
  BUFF I39 (joinf_0[39:39], i_1r0[7:7]);
  BUFF I40 (joinf_0[40:40], i_1r0[8:8]);
  BUFF I41 (joinf_0[41:41], i_1r0[9:9]);
  BUFF I42 (joinf_0[42:42], i_1r0[10:10]);
  BUFF I43 (joinf_0[43:43], i_1r0[11:11]);
  BUFF I44 (joinf_0[44:44], i_1r0[12:12]);
  BUFF I45 (joinf_0[45:45], i_1r0[13:13]);
  BUFF I46 (joinf_0[46:46], i_1r0[14:14]);
  BUFF I47 (joinf_0[47:47], i_1r0[15:15]);
  BUFF I48 (joinf_0[48:48], i_1r0[16:16]);
  BUFF I49 (joinf_0[49:49], i_1r0[17:17]);
  BUFF I50 (joinf_0[50:50], i_1r0[18:18]);
  BUFF I51 (joinf_0[51:51], i_1r0[19:19]);
  BUFF I52 (joinf_0[52:52], i_1r0[20:20]);
  BUFF I53 (joinf_0[53:53], i_1r0[21:21]);
  BUFF I54 (joinf_0[54:54], i_1r0[22:22]);
  BUFF I55 (joinf_0[55:55], i_1r0[23:23]);
  BUFF I56 (joinf_0[56:56], i_1r0[24:24]);
  BUFF I57 (joinf_0[57:57], i_1r0[25:25]);
  BUFF I58 (joinf_0[58:58], i_1r0[26:26]);
  BUFF I59 (joinf_0[59:59], i_1r0[27:27]);
  BUFF I60 (joinf_0[60:60], i_1r0[28:28]);
  BUFF I61 (joinf_0[61:61], i_1r0[29:29]);
  BUFF I62 (joinf_0[62:62], i_1r0[30:30]);
  BUFF I63 (joinf_0[63:63], i_1r0[31:31]);
  BUFF I64 (joint_0[0:0], i_0r1[0:0]);
  BUFF I65 (joint_0[1:1], i_0r1[1:1]);
  BUFF I66 (joint_0[2:2], i_0r1[2:2]);
  BUFF I67 (joint_0[3:3], i_0r1[3:3]);
  BUFF I68 (joint_0[4:4], i_0r1[4:4]);
  BUFF I69 (joint_0[5:5], i_0r1[5:5]);
  BUFF I70 (joint_0[6:6], i_0r1[6:6]);
  BUFF I71 (joint_0[7:7], i_0r1[7:7]);
  BUFF I72 (joint_0[8:8], i_0r1[8:8]);
  BUFF I73 (joint_0[9:9], i_0r1[9:9]);
  BUFF I74 (joint_0[10:10], i_0r1[10:10]);
  BUFF I75 (joint_0[11:11], i_0r1[11:11]);
  BUFF I76 (joint_0[12:12], i_0r1[12:12]);
  BUFF I77 (joint_0[13:13], i_0r1[13:13]);
  BUFF I78 (joint_0[14:14], i_0r1[14:14]);
  BUFF I79 (joint_0[15:15], i_0r1[15:15]);
  BUFF I80 (joint_0[16:16], i_0r1[16:16]);
  BUFF I81 (joint_0[17:17], i_0r1[17:17]);
  BUFF I82 (joint_0[18:18], i_0r1[18:18]);
  BUFF I83 (joint_0[19:19], i_0r1[19:19]);
  BUFF I84 (joint_0[20:20], i_0r1[20:20]);
  BUFF I85 (joint_0[21:21], i_0r1[21:21]);
  BUFF I86 (joint_0[22:22], i_0r1[22:22]);
  BUFF I87 (joint_0[23:23], i_0r1[23:23]);
  BUFF I88 (joint_0[24:24], i_0r1[24:24]);
  BUFF I89 (joint_0[25:25], i_0r1[25:25]);
  BUFF I90 (joint_0[26:26], i_0r1[26:26]);
  BUFF I91 (joint_0[27:27], i_0r1[27:27]);
  BUFF I92 (joint_0[28:28], i_0r1[28:28]);
  BUFF I93 (joint_0[29:29], i_0r1[29:29]);
  BUFF I94 (joint_0[30:30], i_0r1[30:30]);
  BUFF I95 (joint_0[31:31], i_0r1[31:31]);
  BUFF I96 (joint_0[32:32], i_1r1[0:0]);
  BUFF I97 (joint_0[33:33], i_1r1[1:1]);
  BUFF I98 (joint_0[34:34], i_1r1[2:2]);
  BUFF I99 (joint_0[35:35], i_1r1[3:3]);
  BUFF I100 (joint_0[36:36], i_1r1[4:4]);
  BUFF I101 (joint_0[37:37], i_1r1[5:5]);
  BUFF I102 (joint_0[38:38], i_1r1[6:6]);
  BUFF I103 (joint_0[39:39], i_1r1[7:7]);
  BUFF I104 (joint_0[40:40], i_1r1[8:8]);
  BUFF I105 (joint_0[41:41], i_1r1[9:9]);
  BUFF I106 (joint_0[42:42], i_1r1[10:10]);
  BUFF I107 (joint_0[43:43], i_1r1[11:11]);
  BUFF I108 (joint_0[44:44], i_1r1[12:12]);
  BUFF I109 (joint_0[45:45], i_1r1[13:13]);
  BUFF I110 (joint_0[46:46], i_1r1[14:14]);
  BUFF I111 (joint_0[47:47], i_1r1[15:15]);
  BUFF I112 (joint_0[48:48], i_1r1[16:16]);
  BUFF I113 (joint_0[49:49], i_1r1[17:17]);
  BUFF I114 (joint_0[50:50], i_1r1[18:18]);
  BUFF I115 (joint_0[51:51], i_1r1[19:19]);
  BUFF I116 (joint_0[52:52], i_1r1[20:20]);
  BUFF I117 (joint_0[53:53], i_1r1[21:21]);
  BUFF I118 (joint_0[54:54], i_1r1[22:22]);
  BUFF I119 (joint_0[55:55], i_1r1[23:23]);
  BUFF I120 (joint_0[56:56], i_1r1[24:24]);
  BUFF I121 (joint_0[57:57], i_1r1[25:25]);
  BUFF I122 (joint_0[58:58], i_1r1[26:26]);
  BUFF I123 (joint_0[59:59], i_1r1[27:27]);
  BUFF I124 (joint_0[60:60], i_1r1[28:28]);
  BUFF I125 (joint_0[61:61], i_1r1[29:29]);
  BUFF I126 (joint_0[62:62], i_1r1[30:30]);
  BUFF I127 (joint_0[63:63], i_1r1[31:31]);
  OR2 I128 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I129 (icomplete_0, dcomplete_0);
  C2 I130 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I131 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I132 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I133 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I134 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I135 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I136 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I137 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I138 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I139 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I140 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I141 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I142 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I143 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I144 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I145 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I146 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I147 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I148 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I149 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I150 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I151 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I152 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I153 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I154 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I155 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I156 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I157 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I158 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I159 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I160 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I161 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I162 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I163 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I164 (o_0r0[33:33], joinf_0[33:33]);
  BUFF I165 (o_0r0[34:34], joinf_0[34:34]);
  BUFF I166 (o_0r0[35:35], joinf_0[35:35]);
  BUFF I167 (o_0r0[36:36], joinf_0[36:36]);
  BUFF I168 (o_0r0[37:37], joinf_0[37:37]);
  BUFF I169 (o_0r0[38:38], joinf_0[38:38]);
  BUFF I170 (o_0r0[39:39], joinf_0[39:39]);
  BUFF I171 (o_0r0[40:40], joinf_0[40:40]);
  BUFF I172 (o_0r0[41:41], joinf_0[41:41]);
  BUFF I173 (o_0r0[42:42], joinf_0[42:42]);
  BUFF I174 (o_0r0[43:43], joinf_0[43:43]);
  BUFF I175 (o_0r0[44:44], joinf_0[44:44]);
  BUFF I176 (o_0r0[45:45], joinf_0[45:45]);
  BUFF I177 (o_0r0[46:46], joinf_0[46:46]);
  BUFF I178 (o_0r0[47:47], joinf_0[47:47]);
  BUFF I179 (o_0r0[48:48], joinf_0[48:48]);
  BUFF I180 (o_0r0[49:49], joinf_0[49:49]);
  BUFF I181 (o_0r0[50:50], joinf_0[50:50]);
  BUFF I182 (o_0r0[51:51], joinf_0[51:51]);
  BUFF I183 (o_0r0[52:52], joinf_0[52:52]);
  BUFF I184 (o_0r0[53:53], joinf_0[53:53]);
  BUFF I185 (o_0r0[54:54], joinf_0[54:54]);
  BUFF I186 (o_0r0[55:55], joinf_0[55:55]);
  BUFF I187 (o_0r0[56:56], joinf_0[56:56]);
  BUFF I188 (o_0r0[57:57], joinf_0[57:57]);
  BUFF I189 (o_0r0[58:58], joinf_0[58:58]);
  BUFF I190 (o_0r0[59:59], joinf_0[59:59]);
  BUFF I191 (o_0r0[60:60], joinf_0[60:60]);
  BUFF I192 (o_0r0[61:61], joinf_0[61:61]);
  BUFF I193 (o_0r0[62:62], joinf_0[62:62]);
  BUFF I194 (o_0r0[63:63], joinf_0[63:63]);
  BUFF I195 (o_0r1[1:1], joint_0[1:1]);
  BUFF I196 (o_0r1[2:2], joint_0[2:2]);
  BUFF I197 (o_0r1[3:3], joint_0[3:3]);
  BUFF I198 (o_0r1[4:4], joint_0[4:4]);
  BUFF I199 (o_0r1[5:5], joint_0[5:5]);
  BUFF I200 (o_0r1[6:6], joint_0[6:6]);
  BUFF I201 (o_0r1[7:7], joint_0[7:7]);
  BUFF I202 (o_0r1[8:8], joint_0[8:8]);
  BUFF I203 (o_0r1[9:9], joint_0[9:9]);
  BUFF I204 (o_0r1[10:10], joint_0[10:10]);
  BUFF I205 (o_0r1[11:11], joint_0[11:11]);
  BUFF I206 (o_0r1[12:12], joint_0[12:12]);
  BUFF I207 (o_0r1[13:13], joint_0[13:13]);
  BUFF I208 (o_0r1[14:14], joint_0[14:14]);
  BUFF I209 (o_0r1[15:15], joint_0[15:15]);
  BUFF I210 (o_0r1[16:16], joint_0[16:16]);
  BUFF I211 (o_0r1[17:17], joint_0[17:17]);
  BUFF I212 (o_0r1[18:18], joint_0[18:18]);
  BUFF I213 (o_0r1[19:19], joint_0[19:19]);
  BUFF I214 (o_0r1[20:20], joint_0[20:20]);
  BUFF I215 (o_0r1[21:21], joint_0[21:21]);
  BUFF I216 (o_0r1[22:22], joint_0[22:22]);
  BUFF I217 (o_0r1[23:23], joint_0[23:23]);
  BUFF I218 (o_0r1[24:24], joint_0[24:24]);
  BUFF I219 (o_0r1[25:25], joint_0[25:25]);
  BUFF I220 (o_0r1[26:26], joint_0[26:26]);
  BUFF I221 (o_0r1[27:27], joint_0[27:27]);
  BUFF I222 (o_0r1[28:28], joint_0[28:28]);
  BUFF I223 (o_0r1[29:29], joint_0[29:29]);
  BUFF I224 (o_0r1[30:30], joint_0[30:30]);
  BUFF I225 (o_0r1[31:31], joint_0[31:31]);
  BUFF I226 (o_0r1[32:32], joint_0[32:32]);
  BUFF I227 (o_0r1[33:33], joint_0[33:33]);
  BUFF I228 (o_0r1[34:34], joint_0[34:34]);
  BUFF I229 (o_0r1[35:35], joint_0[35:35]);
  BUFF I230 (o_0r1[36:36], joint_0[36:36]);
  BUFF I231 (o_0r1[37:37], joint_0[37:37]);
  BUFF I232 (o_0r1[38:38], joint_0[38:38]);
  BUFF I233 (o_0r1[39:39], joint_0[39:39]);
  BUFF I234 (o_0r1[40:40], joint_0[40:40]);
  BUFF I235 (o_0r1[41:41], joint_0[41:41]);
  BUFF I236 (o_0r1[42:42], joint_0[42:42]);
  BUFF I237 (o_0r1[43:43], joint_0[43:43]);
  BUFF I238 (o_0r1[44:44], joint_0[44:44]);
  BUFF I239 (o_0r1[45:45], joint_0[45:45]);
  BUFF I240 (o_0r1[46:46], joint_0[46:46]);
  BUFF I241 (o_0r1[47:47], joint_0[47:47]);
  BUFF I242 (o_0r1[48:48], joint_0[48:48]);
  BUFF I243 (o_0r1[49:49], joint_0[49:49]);
  BUFF I244 (o_0r1[50:50], joint_0[50:50]);
  BUFF I245 (o_0r1[51:51], joint_0[51:51]);
  BUFF I246 (o_0r1[52:52], joint_0[52:52]);
  BUFF I247 (o_0r1[53:53], joint_0[53:53]);
  BUFF I248 (o_0r1[54:54], joint_0[54:54]);
  BUFF I249 (o_0r1[55:55], joint_0[55:55]);
  BUFF I250 (o_0r1[56:56], joint_0[56:56]);
  BUFF I251 (o_0r1[57:57], joint_0[57:57]);
  BUFF I252 (o_0r1[58:58], joint_0[58:58]);
  BUFF I253 (o_0r1[59:59], joint_0[59:59]);
  BUFF I254 (o_0r1[60:60], joint_0[60:60]);
  BUFF I255 (o_0r1[61:61], joint_0[61:61]);
  BUFF I256 (o_0r1[62:62], joint_0[62:62]);
  BUFF I257 (o_0r1[63:63], joint_0[63:63]);
  BUFF I258 (i_0a, o_0a);
  BUFF I259 (i_1a, o_0a);
endmodule

// tko0m5_1nm5b0 TeakO [
//     (1,TeakOConstant 5 0)] [One 0,One 5]
module tko0m5_1nm5b0 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [4:0] o_0r0;
  output [4:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r);
  BUFF I1 (o_0r0[1:1], i_0r);
  BUFF I2 (o_0r0[2:2], i_0r);
  BUFF I3 (o_0r0[3:3], i_0r);
  BUFF I4 (o_0r0[4:4], i_0r);
  GND I5 (o_0r1[0:0]);
  GND I6 (o_0r1[1:1]);
  GND I7 (o_0r1[2:2]);
  GND I8 (o_0r1[3:3]);
  GND I9 (o_0r1[4:4]);
  BUFF I10 (i_0a, o_0a);
endmodule

// tko0m2_1nm2b1 TeakO [
//     (1,TeakOConstant 2 1)] [One 0,One 2]
module tko0m2_1nm2b1 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  GND I1 (o_0r0[0:0]);
  BUFF I2 (o_0r0[1:1], i_0r);
  GND I3 (o_0r1[1:1]);
  BUFF I4 (i_0a, o_0a);
endmodule

// tko0m2_1nm2b2 TeakO [
//     (1,TeakOConstant 2 2)] [One 0,One 2]
module tko0m2_1nm2b2 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[1:1], i_0r);
  GND I1 (o_0r0[1:1]);
  BUFF I2 (o_0r0[0:0], i_0r);
  GND I3 (o_0r1[0:0]);
  BUFF I4 (i_0a, o_0a);
endmodule

// tkm2x2b TeakM [Many [2,2],One 2]
module tkm2x2b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  input [1:0] i_1r0;
  input [1:0] i_1r1;
  output i_1a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  wire [1:0] gfint_0;
  wire [1:0] gfint_1;
  wire [1:0] gtint_0;
  wire [1:0] gtint_1;
  wire choice_0;
  wire choice_1;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire nchosen_0;
  wire [1:0] comp0_0;
  wire [1:0] comp1_0;
  OR2 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0]);
  OR2 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1]);
  OR2 I2 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0]);
  OR2 I3 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1]);
  AND2 I4 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I5 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I6 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I7 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I8 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I9 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I10 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I11 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  OR2 I12 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I13 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  C2 I14 (icomp_0, comp0_0[0:0], comp0_0[1:1]);
  OR2 I15 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I16 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  C2 I17 (icomp_1, comp1_0[0:0], comp1_0[1:1]);
  C2R I18 (choice_0, icomp_0, nchosen_0, reset);
  C2R I19 (choice_1, icomp_1, nchosen_0, reset);
  OR2 I20 (anychoice_0, choice_0, choice_1);
  NOR2 I21 (nchosen_0, anychoice_0, o_0a);
  C2R I22 (i_0a, choice_0, o_0a, reset);
  C2R I23 (i_1a, choice_1, o_0a, reset);
endmodule

// tkj2m0_2 TeakJ [Many [0,2],One 2]
module tkj2m0_2 (i_0r, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  input [1:0] i_1r0;
  input [1:0] i_1r1;
  output i_1a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [1:0] joinf_0;
  wire [1:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_1r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_1r0[1:1]);
  BUFF I2 (joint_0[0:0], i_1r1[0:0]);
  BUFF I3 (joint_0[1:1], i_1r1[1:1]);
  BUFF I4 (icomplete_0, i_0r);
  C2 I5 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I6 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I7 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I8 (o_0r1[1:1], joint_0[1:1]);
  BUFF I9 (i_0a, o_0a);
  BUFF I10 (i_1a, o_0a);
endmodule

// tks2_o0w2_1o0w0_2o0w0 TeakS (0+:2) [([Imp 1 0],0),([Imp 2 0],0)] [One 2,Many [0,0]]
module tks2_o0w2_1o0w0_2o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire [1:0] comp_0;
  BUFF I0 (sel_0, match0_0);
  C2 I1 (match0_0, i_0r1[0:0], i_0r0[1:1]);
  BUFF I2 (sel_1, match1_0);
  C2 I3 (match1_0, i_0r0[0:0], i_0r1[1:1]);
  C2 I4 (gsel_0, sel_0, icomplete_0);
  C2 I5 (gsel_1, sel_1, icomplete_0);
  OR2 I6 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I7 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  C2 I8 (icomplete_0, comp_0[0:0], comp_0[1:1]);
  BUFF I9 (o_0r, gsel_0);
  BUFF I10 (o_1r, gsel_1);
  OR2 I11 (oack_0, o_0a, o_1a);
  C2 I12 (i_0a, oack_0, icomplete_0);
endmodule

// tko0m32_1nm32b0 TeakO [
//     (1,TeakOConstant 32 0)] [One 0,One 32]
module tko0m32_1nm32b0 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r);
  BUFF I1 (o_0r0[1:1], i_0r);
  BUFF I2 (o_0r0[2:2], i_0r);
  BUFF I3 (o_0r0[3:3], i_0r);
  BUFF I4 (o_0r0[4:4], i_0r);
  BUFF I5 (o_0r0[5:5], i_0r);
  BUFF I6 (o_0r0[6:6], i_0r);
  BUFF I7 (o_0r0[7:7], i_0r);
  BUFF I8 (o_0r0[8:8], i_0r);
  BUFF I9 (o_0r0[9:9], i_0r);
  BUFF I10 (o_0r0[10:10], i_0r);
  BUFF I11 (o_0r0[11:11], i_0r);
  BUFF I12 (o_0r0[12:12], i_0r);
  BUFF I13 (o_0r0[13:13], i_0r);
  BUFF I14 (o_0r0[14:14], i_0r);
  BUFF I15 (o_0r0[15:15], i_0r);
  BUFF I16 (o_0r0[16:16], i_0r);
  BUFF I17 (o_0r0[17:17], i_0r);
  BUFF I18 (o_0r0[18:18], i_0r);
  BUFF I19 (o_0r0[19:19], i_0r);
  BUFF I20 (o_0r0[20:20], i_0r);
  BUFF I21 (o_0r0[21:21], i_0r);
  BUFF I22 (o_0r0[22:22], i_0r);
  BUFF I23 (o_0r0[23:23], i_0r);
  BUFF I24 (o_0r0[24:24], i_0r);
  BUFF I25 (o_0r0[25:25], i_0r);
  BUFF I26 (o_0r0[26:26], i_0r);
  BUFF I27 (o_0r0[27:27], i_0r);
  BUFF I28 (o_0r0[28:28], i_0r);
  BUFF I29 (o_0r0[29:29], i_0r);
  BUFF I30 (o_0r0[30:30], i_0r);
  BUFF I31 (o_0r0[31:31], i_0r);
  GND I32 (o_0r1[0:0]);
  GND I33 (o_0r1[1:1]);
  GND I34 (o_0r1[2:2]);
  GND I35 (o_0r1[3:3]);
  GND I36 (o_0r1[4:4]);
  GND I37 (o_0r1[5:5]);
  GND I38 (o_0r1[6:6]);
  GND I39 (o_0r1[7:7]);
  GND I40 (o_0r1[8:8]);
  GND I41 (o_0r1[9:9]);
  GND I42 (o_0r1[10:10]);
  GND I43 (o_0r1[11:11]);
  GND I44 (o_0r1[12:12]);
  GND I45 (o_0r1[13:13]);
  GND I46 (o_0r1[14:14]);
  GND I47 (o_0r1[15:15]);
  GND I48 (o_0r1[16:16]);
  GND I49 (o_0r1[17:17]);
  GND I50 (o_0r1[18:18]);
  GND I51 (o_0r1[19:19]);
  GND I52 (o_0r1[20:20]);
  GND I53 (o_0r1[21:21]);
  GND I54 (o_0r1[22:22]);
  GND I55 (o_0r1[23:23]);
  GND I56 (o_0r1[24:24]);
  GND I57 (o_0r1[25:25]);
  GND I58 (o_0r1[26:26]);
  GND I59 (o_0r1[27:27]);
  GND I60 (o_0r1[28:28]);
  GND I61 (o_0r1[29:29]);
  GND I62 (o_0r1[30:30]);
  GND I63 (o_0r1[31:31]);
  BUFF I64 (i_0a, o_0a);
endmodule

// tko0m3_1nm3b4 TeakO [
//     (1,TeakOConstant 3 4)] [One 0,One 3]
module tko0m3_1nm3b4 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[2:2], i_0r);
  GND I1 (o_0r0[2:2]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  GND I4 (o_0r1[0:0]);
  GND I5 (o_0r1[1:1]);
  BUFF I6 (i_0a, o_0a);
endmodule

// tkj3m0_0_0_3 TeakJ [Many [0,0,0,3],One 3]
module tkj3m0_0_0_3 (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, i_3r0, i_3r1, i_3a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input [2:0] i_3r0;
  input [2:0] i_3r1;
  output i_3a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [2:0] joinf_0;
  wire [2:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_3r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_3r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_3r0[2:2]);
  BUFF I3 (joint_0[0:0], i_3r1[0:0]);
  BUFF I4 (joint_0[1:1], i_3r1[1:1]);
  BUFF I5 (joint_0[2:2], i_3r1[2:2]);
  C3 I6 (icomplete_0, i_0r, i_1r, i_2r);
  C2 I7 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I8 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I9 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I10 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I11 (o_0r1[1:1], joint_0[1:1]);
  BUFF I12 (o_0r1[2:2], joint_0[2:2]);
  BUFF I13 (i_0a, o_0a);
  BUFF I14 (i_1a, o_0a);
  BUFF I15 (i_2a, o_0a);
  BUFF I16 (i_3a, o_0a);
endmodule

// tkm2x1b TeakM [Many [1,1],One 1]
module tkm2x1b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input i_1r0;
  input i_1r1;
  output i_1a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire gfint_0;
  wire gfint_1;
  wire gtint_0;
  wire gtint_1;
  wire choice_0;
  wire choice_1;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire nchosen_0;
  wire comp0_0;
  wire comp1_0;
  OR2 I0 (o_0r0, gfint_0, gfint_1);
  OR2 I1 (o_0r1, gtint_0, gtint_1);
  AND2 I2 (gtint_0, choice_0, i_0r1);
  AND2 I3 (gtint_1, choice_1, i_1r1);
  AND2 I4 (gfint_0, choice_0, i_0r0);
  AND2 I5 (gfint_1, choice_1, i_1r0);
  OR2 I6 (comp0_0, i_0r0, i_0r1);
  BUFF I7 (icomp_0, comp0_0);
  OR2 I8 (comp1_0, i_1r0, i_1r1);
  BUFF I9 (icomp_1, comp1_0);
  C2R I10 (choice_0, icomp_0, nchosen_0, reset);
  C2R I11 (choice_1, icomp_1, nchosen_0, reset);
  OR2 I12 (anychoice_0, choice_0, choice_1);
  NOR2 I13 (nchosen_0, anychoice_0, o_0a);
  C2R I14 (i_0a, choice_0, o_0a, reset);
  C2R I15 (i_1a, choice_1, o_0a, reset);
endmodule

// tkvStopped1_wo0w1_ro0w1 TeakV "Stopped" 1 [] [0] [0] [Many [1],Many [0],Many [0],Many [1]]
module tkvStopped1_wo0w1_ro0w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input wg_0r0;
  input wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  input reset;
  wire wf_0;
  wire wt_0;
  wire df_0;
  wire dt_0;
  wire wc_0;
  wire wacks_0;
  wire wenr_0;
  wire wen_0;
  wire anyread_0;
  wire nreset_0;
  wire drlgf_0;
  wire drlgt_0;
  wire comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire conwgit_0;
  wire conwgif_0;
  wire conwig_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0, wenr_0, nreset_0);
  AND2 I2 (drlgf_0, wf_0, wen_0);
  AND2 I3 (drlgt_0, wt_0, wen_0);
  NOR2 I4 (df_0, dt_0, drlgt_0);
  NOR3 I5 (dt_0, df_0, drlgf_0, reset);
  AO22 I6 (wacks_0, drlgf_0, df_0, drlgt_0, dt_0);
  OR2 I7 (comp0_0, wg_0r0, wg_0r1);
  BUFF I8 (wc_0, comp0_0);
  AND2 I9 (conwgif_0, wg_0r0, conwig_0);
  AND2 I10 (conwgit_0, wg_0r1, conwig_0);
  BUFF I11 (conwigc_0, wc_0);
  AO22 I12 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I13 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I14 (wf_0, conwgif_0);
  BUFF I15 (wt_0, conwgit_0);
  BUFF I16 (wenr_0, wc_0);
  C2 I17 (wd_0r, conwig_0, wacks_0);
  AND2 I18 (rd_0r0, df_0, rg_0r);
  AND2 I19 (rd_0r1, dt_0, rg_0r);
  OR2 I20 (anyread_0, rg_0r, rg_0a);
  BUFF I21 (wg_0a, wd_0a);
  BUFF I22 (rg_0a, rd_0a);
endmodule

// tkvMDR32_wo0w32_ro0w32o0w5 TeakV "MDR" 32 [] [0] [0,0] [Many [32],Many [0],Many [0,0],Many [32,5]]
module tkvMDR32_wo0w32_ro0w32o0w5 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [4:0] rd_1r0;
  output [4:0] rd_1r1;
  input rd_1a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp4821_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I462 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I463 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I464 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I465 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I466 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I467 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I468 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I469 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I470 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I471 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I472 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I473 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I474 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I475 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I476 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I477 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I478 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I479 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I480 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I481 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I482 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I483 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I484 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I485 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I486 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I487 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I488 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I489 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I490 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I491 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I492 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I493 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I494 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I495 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I496 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I497 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  NOR3 I498 (simp4821_0[0:0], rg_0r, rg_1r, rg_0a);
  INV I499 (simp4821_0[1:1], rg_1a);
  NAND2 I500 (anyread_0, simp4821_0[0:0], simp4821_0[1:1]);
  BUFF I501 (wg_0a, wd_0a);
  BUFF I502 (rg_0a, rd_0a);
  BUFF I503 (rg_1a, rd_1a);
endmodule

// tkm2x5b TeakM [Many [5,5],One 5]
module tkm2x5b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [4:0] i_0r0;
  input [4:0] i_0r1;
  output i_0a;
  input [4:0] i_1r0;
  input [4:0] i_1r1;
  output i_1a;
  output [4:0] o_0r0;
  output [4:0] o_0r1;
  input o_0a;
  input reset;
  wire [4:0] gfint_0;
  wire [4:0] gfint_1;
  wire [4:0] gtint_0;
  wire [4:0] gtint_1;
  wire choice_0;
  wire choice_1;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire nchosen_0;
  wire [4:0] comp0_0;
  wire [1:0] simp461_0;
  wire [4:0] comp1_0;
  wire [1:0] simp531_0;
  OR2 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0]);
  OR2 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1]);
  OR2 I2 (o_0r0[2:2], gfint_0[2:2], gfint_1[2:2]);
  OR2 I3 (o_0r0[3:3], gfint_0[3:3], gfint_1[3:3]);
  OR2 I4 (o_0r0[4:4], gfint_0[4:4], gfint_1[4:4]);
  OR2 I5 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0]);
  OR2 I6 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1]);
  OR2 I7 (o_0r1[2:2], gtint_0[2:2], gtint_1[2:2]);
  OR2 I8 (o_0r1[3:3], gtint_0[3:3], gtint_1[3:3]);
  OR2 I9 (o_0r1[4:4], gtint_0[4:4], gtint_1[4:4]);
  AND2 I10 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I11 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I12 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I13 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I14 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I15 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I16 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I17 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I18 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I19 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I20 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I21 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I22 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I23 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I24 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I25 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I26 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I27 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I28 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I29 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  OR2 I30 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I31 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I32 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I33 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I34 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  C3 I35 (simp461_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C2 I36 (simp461_0[1:1], comp0_0[3:3], comp0_0[4:4]);
  C2 I37 (icomp_0, simp461_0[0:0], simp461_0[1:1]);
  OR2 I38 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I39 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I40 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I41 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I42 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  C3 I43 (simp531_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C2 I44 (simp531_0[1:1], comp1_0[3:3], comp1_0[4:4]);
  C2 I45 (icomp_1, simp531_0[0:0], simp531_0[1:1]);
  C2R I46 (choice_0, icomp_0, nchosen_0, reset);
  C2R I47 (choice_1, icomp_1, nchosen_0, reset);
  OR2 I48 (anychoice_0, choice_0, choice_1);
  NOR2 I49 (nchosen_0, anychoice_0, o_0a);
  C2R I50 (i_0a, choice_0, o_0a, reset);
  C2R I51 (i_1a, choice_1, o_0a, reset);
endmodule

// tkvPCstep5_wo0w5_ro0w5 TeakV "PC_step" 5 [] [0] [0] [Many [5],Many [0],Many [0],Many [5]]
module tkvPCstep5_wo0w5_ro0w5 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [4:0] wg_0r0;
  input [4:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [4:0] rd_0r0;
  output [4:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [4:0] wf_0;
  wire [4:0] wt_0;
  wire [4:0] df_0;
  wire [4:0] dt_0;
  wire wc_0;
  wire [4:0] wacks_0;
  wire [4:0] wenr_0;
  wire [4:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [4:0] drlgf_0;
  wire [4:0] drlgt_0;
  wire [4:0] comp0_0;
  wire [1:0] simp491_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [4:0] conwgit_0;
  wire [4:0] conwgif_0;
  wire conwig_0;
  wire [1:0] simp831_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I7 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I8 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I9 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I10 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I11 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I12 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I13 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I14 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I15 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  NOR2 I16 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I17 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I18 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I19 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I20 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR3 I21 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I22 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I23 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I24 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I25 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  AO22 I26 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I27 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I28 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I29 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I30 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  OR2 I31 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I32 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I33 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I34 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I35 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  C3 I36 (simp491_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C2 I37 (simp491_0[1:1], comp0_0[3:3], comp0_0[4:4]);
  C2 I38 (wc_0, simp491_0[0:0], simp491_0[1:1]);
  AND2 I39 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I40 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I41 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I42 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I43 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I44 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I45 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I46 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I47 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I48 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  BUFF I49 (conwigc_0, wc_0);
  AO22 I50 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I51 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I52 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I53 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I54 (wenr_0[0:0], wc_0);
  BUFF I55 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I56 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I57 (wenr_0[1:1], wc_0);
  BUFF I58 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I59 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I60 (wenr_0[2:2], wc_0);
  BUFF I61 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I62 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I63 (wenr_0[3:3], wc_0);
  BUFF I64 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I65 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I66 (wenr_0[4:4], wc_0);
  C3 I67 (simp831_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I68 (simp831_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C2 I69 (wd_0r, simp831_0[0:0], simp831_0[1:1]);
  AND2 I70 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I71 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I72 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I73 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I74 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I75 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I76 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I77 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I78 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I79 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  OR2 I80 (anyread_0, rg_0r, rg_0a);
  BUFF I81 (wg_0a, wd_0a);
  BUFF I82 (rg_0a, rd_0a);
endmodule

// tkvPC5_wo0w5_ro0w5o0w5 TeakV "PC" 5 [] [0] [0,0] [Many [5],Many [0],Many [0,0],Many [5,5]]
module tkvPC5_wo0w5_ro0w5o0w5 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, reset);
  input [4:0] wg_0r0;
  input [4:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [4:0] rd_0r0;
  output [4:0] rd_0r1;
  input rd_0a;
  output [4:0] rd_1r0;
  output [4:0] rd_1r1;
  input rd_1a;
  input reset;
  wire [4:0] wf_0;
  wire [4:0] wt_0;
  wire [4:0] df_0;
  wire [4:0] dt_0;
  wire wc_0;
  wire [4:0] wacks_0;
  wire [4:0] wenr_0;
  wire [4:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [4:0] drlgf_0;
  wire [4:0] drlgt_0;
  wire [4:0] comp0_0;
  wire [1:0] simp491_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [4:0] conwgit_0;
  wire [4:0] conwgif_0;
  wire conwig_0;
  wire [1:0] simp831_0;
  wire [1:0] simp1041_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I7 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I8 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I9 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I10 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I11 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I12 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I13 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I14 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I15 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  NOR2 I16 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I17 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I18 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I19 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I20 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR3 I21 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I22 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I23 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I24 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I25 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  AO22 I26 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I27 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I28 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I29 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I30 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  OR2 I31 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I32 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I33 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I34 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I35 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  C3 I36 (simp491_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C2 I37 (simp491_0[1:1], comp0_0[3:3], comp0_0[4:4]);
  C2 I38 (wc_0, simp491_0[0:0], simp491_0[1:1]);
  AND2 I39 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I40 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I41 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I42 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I43 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I44 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I45 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I46 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I47 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I48 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  BUFF I49 (conwigc_0, wc_0);
  AO22 I50 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I51 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I52 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I53 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I54 (wenr_0[0:0], wc_0);
  BUFF I55 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I56 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I57 (wenr_0[1:1], wc_0);
  BUFF I58 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I59 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I60 (wenr_0[2:2], wc_0);
  BUFF I61 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I62 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I63 (wenr_0[3:3], wc_0);
  BUFF I64 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I65 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I66 (wenr_0[4:4], wc_0);
  C3 I67 (simp831_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I68 (simp831_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C2 I69 (wd_0r, simp831_0[0:0], simp831_0[1:1]);
  AND2 I70 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I71 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I72 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I73 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I74 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I75 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I76 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I77 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I78 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I79 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I80 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I81 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I82 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I83 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I84 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I85 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I86 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I87 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I88 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I89 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  NOR3 I90 (simp1041_0[0:0], rg_0r, rg_1r, rg_0a);
  INV I91 (simp1041_0[1:1], rg_1a);
  NAND2 I92 (anyread_0, simp1041_0[0:0], simp1041_0[1:1]);
  BUFF I93 (wg_0a, wd_0a);
  BUFF I94 (rg_0a, rd_0a);
  BUFF I95 (rg_1a, rd_1a);
endmodule

// tkvIR32_wo0w32_ro0w5 TeakV "IR" 32 [] [0] [0] [Many [32],Many [0],Many [0],Many [5]]
module tkvIR32_wo0w32_ro0w5 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [4:0] rd_0r0;
  output [4:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I430 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I431 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I432 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I433 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  OR2 I434 (anyread_0, rg_0r, rg_0a);
  BUFF I435 (wg_0a, wd_0a);
  BUFF I436 (rg_0a, rd_0a);
endmodule

// tkvACCslave32_wo0w32_ro0w32o0w32 TeakV "ACC_slave" 32 [] [0] [0,0] [Many [32],Many [0],Many [0,0],Ma
//   ny [32,32]]
module tkvACCslave32_wo0w32_ro0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp5361_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I489 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I490 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I491 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I492 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I493 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I494 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I495 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I496 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I497 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I498 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I499 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I500 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I501 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I502 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I503 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I504 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I505 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I506 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I507 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I508 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I509 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I510 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I511 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I512 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I513 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I514 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I515 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I516 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I517 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I518 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I519 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I520 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I521 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I522 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I523 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I524 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I525 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I526 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I527 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I528 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I529 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I530 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I531 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I532 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I533 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I534 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I535 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I536 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I537 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I538 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I539 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I540 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I541 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I542 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I543 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I544 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I545 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I546 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I547 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I548 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I549 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I550 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I551 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  NOR3 I552 (simp5361_0[0:0], rg_0r, rg_1r, rg_0a);
  INV I553 (simp5361_0[1:1], rg_1a);
  NAND2 I554 (anyread_0, simp5361_0[0:0], simp5361_0[1:1]);
  BUFF I555 (wg_0a, wd_0a);
  BUFF I556 (rg_0a, rd_0a);
  BUFF I557 (rg_1a, rd_1a);
endmodule

// tkm2x32b TeakM [Many [32,32],One 32]
module tkm2x32b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire [31:0] gfint_0;
  wire [31:0] gfint_1;
  wire [31:0] gtint_0;
  wire [31:0] gtint_1;
  wire choice_0;
  wire choice_1;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire nchosen_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2351_0;
  wire [3:0] simp2352_0;
  wire [1:0] simp2353_0;
  wire [31:0] comp1_0;
  wire [10:0] simp2691_0;
  wire [3:0] simp2692_0;
  wire [1:0] simp2693_0;
  OR2 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0]);
  OR2 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1]);
  OR2 I2 (o_0r0[2:2], gfint_0[2:2], gfint_1[2:2]);
  OR2 I3 (o_0r0[3:3], gfint_0[3:3], gfint_1[3:3]);
  OR2 I4 (o_0r0[4:4], gfint_0[4:4], gfint_1[4:4]);
  OR2 I5 (o_0r0[5:5], gfint_0[5:5], gfint_1[5:5]);
  OR2 I6 (o_0r0[6:6], gfint_0[6:6], gfint_1[6:6]);
  OR2 I7 (o_0r0[7:7], gfint_0[7:7], gfint_1[7:7]);
  OR2 I8 (o_0r0[8:8], gfint_0[8:8], gfint_1[8:8]);
  OR2 I9 (o_0r0[9:9], gfint_0[9:9], gfint_1[9:9]);
  OR2 I10 (o_0r0[10:10], gfint_0[10:10], gfint_1[10:10]);
  OR2 I11 (o_0r0[11:11], gfint_0[11:11], gfint_1[11:11]);
  OR2 I12 (o_0r0[12:12], gfint_0[12:12], gfint_1[12:12]);
  OR2 I13 (o_0r0[13:13], gfint_0[13:13], gfint_1[13:13]);
  OR2 I14 (o_0r0[14:14], gfint_0[14:14], gfint_1[14:14]);
  OR2 I15 (o_0r0[15:15], gfint_0[15:15], gfint_1[15:15]);
  OR2 I16 (o_0r0[16:16], gfint_0[16:16], gfint_1[16:16]);
  OR2 I17 (o_0r0[17:17], gfint_0[17:17], gfint_1[17:17]);
  OR2 I18 (o_0r0[18:18], gfint_0[18:18], gfint_1[18:18]);
  OR2 I19 (o_0r0[19:19], gfint_0[19:19], gfint_1[19:19]);
  OR2 I20 (o_0r0[20:20], gfint_0[20:20], gfint_1[20:20]);
  OR2 I21 (o_0r0[21:21], gfint_0[21:21], gfint_1[21:21]);
  OR2 I22 (o_0r0[22:22], gfint_0[22:22], gfint_1[22:22]);
  OR2 I23 (o_0r0[23:23], gfint_0[23:23], gfint_1[23:23]);
  OR2 I24 (o_0r0[24:24], gfint_0[24:24], gfint_1[24:24]);
  OR2 I25 (o_0r0[25:25], gfint_0[25:25], gfint_1[25:25]);
  OR2 I26 (o_0r0[26:26], gfint_0[26:26], gfint_1[26:26]);
  OR2 I27 (o_0r0[27:27], gfint_0[27:27], gfint_1[27:27]);
  OR2 I28 (o_0r0[28:28], gfint_0[28:28], gfint_1[28:28]);
  OR2 I29 (o_0r0[29:29], gfint_0[29:29], gfint_1[29:29]);
  OR2 I30 (o_0r0[30:30], gfint_0[30:30], gfint_1[30:30]);
  OR2 I31 (o_0r0[31:31], gfint_0[31:31], gfint_1[31:31]);
  OR2 I32 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0]);
  OR2 I33 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1]);
  OR2 I34 (o_0r1[2:2], gtint_0[2:2], gtint_1[2:2]);
  OR2 I35 (o_0r1[3:3], gtint_0[3:3], gtint_1[3:3]);
  OR2 I36 (o_0r1[4:4], gtint_0[4:4], gtint_1[4:4]);
  OR2 I37 (o_0r1[5:5], gtint_0[5:5], gtint_1[5:5]);
  OR2 I38 (o_0r1[6:6], gtint_0[6:6], gtint_1[6:6]);
  OR2 I39 (o_0r1[7:7], gtint_0[7:7], gtint_1[7:7]);
  OR2 I40 (o_0r1[8:8], gtint_0[8:8], gtint_1[8:8]);
  OR2 I41 (o_0r1[9:9], gtint_0[9:9], gtint_1[9:9]);
  OR2 I42 (o_0r1[10:10], gtint_0[10:10], gtint_1[10:10]);
  OR2 I43 (o_0r1[11:11], gtint_0[11:11], gtint_1[11:11]);
  OR2 I44 (o_0r1[12:12], gtint_0[12:12], gtint_1[12:12]);
  OR2 I45 (o_0r1[13:13], gtint_0[13:13], gtint_1[13:13]);
  OR2 I46 (o_0r1[14:14], gtint_0[14:14], gtint_1[14:14]);
  OR2 I47 (o_0r1[15:15], gtint_0[15:15], gtint_1[15:15]);
  OR2 I48 (o_0r1[16:16], gtint_0[16:16], gtint_1[16:16]);
  OR2 I49 (o_0r1[17:17], gtint_0[17:17], gtint_1[17:17]);
  OR2 I50 (o_0r1[18:18], gtint_0[18:18], gtint_1[18:18]);
  OR2 I51 (o_0r1[19:19], gtint_0[19:19], gtint_1[19:19]);
  OR2 I52 (o_0r1[20:20], gtint_0[20:20], gtint_1[20:20]);
  OR2 I53 (o_0r1[21:21], gtint_0[21:21], gtint_1[21:21]);
  OR2 I54 (o_0r1[22:22], gtint_0[22:22], gtint_1[22:22]);
  OR2 I55 (o_0r1[23:23], gtint_0[23:23], gtint_1[23:23]);
  OR2 I56 (o_0r1[24:24], gtint_0[24:24], gtint_1[24:24]);
  OR2 I57 (o_0r1[25:25], gtint_0[25:25], gtint_1[25:25]);
  OR2 I58 (o_0r1[26:26], gtint_0[26:26], gtint_1[26:26]);
  OR2 I59 (o_0r1[27:27], gtint_0[27:27], gtint_1[27:27]);
  OR2 I60 (o_0r1[28:28], gtint_0[28:28], gtint_1[28:28]);
  OR2 I61 (o_0r1[29:29], gtint_0[29:29], gtint_1[29:29]);
  OR2 I62 (o_0r1[30:30], gtint_0[30:30], gtint_1[30:30]);
  OR2 I63 (o_0r1[31:31], gtint_0[31:31], gtint_1[31:31]);
  AND2 I64 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I65 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I66 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I67 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I68 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I69 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I70 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I71 (gtint_0[7:7], choice_0, i_0r1[7:7]);
  AND2 I72 (gtint_0[8:8], choice_0, i_0r1[8:8]);
  AND2 I73 (gtint_0[9:9], choice_0, i_0r1[9:9]);
  AND2 I74 (gtint_0[10:10], choice_0, i_0r1[10:10]);
  AND2 I75 (gtint_0[11:11], choice_0, i_0r1[11:11]);
  AND2 I76 (gtint_0[12:12], choice_0, i_0r1[12:12]);
  AND2 I77 (gtint_0[13:13], choice_0, i_0r1[13:13]);
  AND2 I78 (gtint_0[14:14], choice_0, i_0r1[14:14]);
  AND2 I79 (gtint_0[15:15], choice_0, i_0r1[15:15]);
  AND2 I80 (gtint_0[16:16], choice_0, i_0r1[16:16]);
  AND2 I81 (gtint_0[17:17], choice_0, i_0r1[17:17]);
  AND2 I82 (gtint_0[18:18], choice_0, i_0r1[18:18]);
  AND2 I83 (gtint_0[19:19], choice_0, i_0r1[19:19]);
  AND2 I84 (gtint_0[20:20], choice_0, i_0r1[20:20]);
  AND2 I85 (gtint_0[21:21], choice_0, i_0r1[21:21]);
  AND2 I86 (gtint_0[22:22], choice_0, i_0r1[22:22]);
  AND2 I87 (gtint_0[23:23], choice_0, i_0r1[23:23]);
  AND2 I88 (gtint_0[24:24], choice_0, i_0r1[24:24]);
  AND2 I89 (gtint_0[25:25], choice_0, i_0r1[25:25]);
  AND2 I90 (gtint_0[26:26], choice_0, i_0r1[26:26]);
  AND2 I91 (gtint_0[27:27], choice_0, i_0r1[27:27]);
  AND2 I92 (gtint_0[28:28], choice_0, i_0r1[28:28]);
  AND2 I93 (gtint_0[29:29], choice_0, i_0r1[29:29]);
  AND2 I94 (gtint_0[30:30], choice_0, i_0r1[30:30]);
  AND2 I95 (gtint_0[31:31], choice_0, i_0r1[31:31]);
  AND2 I96 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I97 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I98 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I99 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I100 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I101 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I102 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I103 (gtint_1[7:7], choice_1, i_1r1[7:7]);
  AND2 I104 (gtint_1[8:8], choice_1, i_1r1[8:8]);
  AND2 I105 (gtint_1[9:9], choice_1, i_1r1[9:9]);
  AND2 I106 (gtint_1[10:10], choice_1, i_1r1[10:10]);
  AND2 I107 (gtint_1[11:11], choice_1, i_1r1[11:11]);
  AND2 I108 (gtint_1[12:12], choice_1, i_1r1[12:12]);
  AND2 I109 (gtint_1[13:13], choice_1, i_1r1[13:13]);
  AND2 I110 (gtint_1[14:14], choice_1, i_1r1[14:14]);
  AND2 I111 (gtint_1[15:15], choice_1, i_1r1[15:15]);
  AND2 I112 (gtint_1[16:16], choice_1, i_1r1[16:16]);
  AND2 I113 (gtint_1[17:17], choice_1, i_1r1[17:17]);
  AND2 I114 (gtint_1[18:18], choice_1, i_1r1[18:18]);
  AND2 I115 (gtint_1[19:19], choice_1, i_1r1[19:19]);
  AND2 I116 (gtint_1[20:20], choice_1, i_1r1[20:20]);
  AND2 I117 (gtint_1[21:21], choice_1, i_1r1[21:21]);
  AND2 I118 (gtint_1[22:22], choice_1, i_1r1[22:22]);
  AND2 I119 (gtint_1[23:23], choice_1, i_1r1[23:23]);
  AND2 I120 (gtint_1[24:24], choice_1, i_1r1[24:24]);
  AND2 I121 (gtint_1[25:25], choice_1, i_1r1[25:25]);
  AND2 I122 (gtint_1[26:26], choice_1, i_1r1[26:26]);
  AND2 I123 (gtint_1[27:27], choice_1, i_1r1[27:27]);
  AND2 I124 (gtint_1[28:28], choice_1, i_1r1[28:28]);
  AND2 I125 (gtint_1[29:29], choice_1, i_1r1[29:29]);
  AND2 I126 (gtint_1[30:30], choice_1, i_1r1[30:30]);
  AND2 I127 (gtint_1[31:31], choice_1, i_1r1[31:31]);
  AND2 I128 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I129 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I130 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I131 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I132 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I133 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I134 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I135 (gfint_0[7:7], choice_0, i_0r0[7:7]);
  AND2 I136 (gfint_0[8:8], choice_0, i_0r0[8:8]);
  AND2 I137 (gfint_0[9:9], choice_0, i_0r0[9:9]);
  AND2 I138 (gfint_0[10:10], choice_0, i_0r0[10:10]);
  AND2 I139 (gfint_0[11:11], choice_0, i_0r0[11:11]);
  AND2 I140 (gfint_0[12:12], choice_0, i_0r0[12:12]);
  AND2 I141 (gfint_0[13:13], choice_0, i_0r0[13:13]);
  AND2 I142 (gfint_0[14:14], choice_0, i_0r0[14:14]);
  AND2 I143 (gfint_0[15:15], choice_0, i_0r0[15:15]);
  AND2 I144 (gfint_0[16:16], choice_0, i_0r0[16:16]);
  AND2 I145 (gfint_0[17:17], choice_0, i_0r0[17:17]);
  AND2 I146 (gfint_0[18:18], choice_0, i_0r0[18:18]);
  AND2 I147 (gfint_0[19:19], choice_0, i_0r0[19:19]);
  AND2 I148 (gfint_0[20:20], choice_0, i_0r0[20:20]);
  AND2 I149 (gfint_0[21:21], choice_0, i_0r0[21:21]);
  AND2 I150 (gfint_0[22:22], choice_0, i_0r0[22:22]);
  AND2 I151 (gfint_0[23:23], choice_0, i_0r0[23:23]);
  AND2 I152 (gfint_0[24:24], choice_0, i_0r0[24:24]);
  AND2 I153 (gfint_0[25:25], choice_0, i_0r0[25:25]);
  AND2 I154 (gfint_0[26:26], choice_0, i_0r0[26:26]);
  AND2 I155 (gfint_0[27:27], choice_0, i_0r0[27:27]);
  AND2 I156 (gfint_0[28:28], choice_0, i_0r0[28:28]);
  AND2 I157 (gfint_0[29:29], choice_0, i_0r0[29:29]);
  AND2 I158 (gfint_0[30:30], choice_0, i_0r0[30:30]);
  AND2 I159 (gfint_0[31:31], choice_0, i_0r0[31:31]);
  AND2 I160 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I161 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I162 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I163 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I164 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I165 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I166 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I167 (gfint_1[7:7], choice_1, i_1r0[7:7]);
  AND2 I168 (gfint_1[8:8], choice_1, i_1r0[8:8]);
  AND2 I169 (gfint_1[9:9], choice_1, i_1r0[9:9]);
  AND2 I170 (gfint_1[10:10], choice_1, i_1r0[10:10]);
  AND2 I171 (gfint_1[11:11], choice_1, i_1r0[11:11]);
  AND2 I172 (gfint_1[12:12], choice_1, i_1r0[12:12]);
  AND2 I173 (gfint_1[13:13], choice_1, i_1r0[13:13]);
  AND2 I174 (gfint_1[14:14], choice_1, i_1r0[14:14]);
  AND2 I175 (gfint_1[15:15], choice_1, i_1r0[15:15]);
  AND2 I176 (gfint_1[16:16], choice_1, i_1r0[16:16]);
  AND2 I177 (gfint_1[17:17], choice_1, i_1r0[17:17]);
  AND2 I178 (gfint_1[18:18], choice_1, i_1r0[18:18]);
  AND2 I179 (gfint_1[19:19], choice_1, i_1r0[19:19]);
  AND2 I180 (gfint_1[20:20], choice_1, i_1r0[20:20]);
  AND2 I181 (gfint_1[21:21], choice_1, i_1r0[21:21]);
  AND2 I182 (gfint_1[22:22], choice_1, i_1r0[22:22]);
  AND2 I183 (gfint_1[23:23], choice_1, i_1r0[23:23]);
  AND2 I184 (gfint_1[24:24], choice_1, i_1r0[24:24]);
  AND2 I185 (gfint_1[25:25], choice_1, i_1r0[25:25]);
  AND2 I186 (gfint_1[26:26], choice_1, i_1r0[26:26]);
  AND2 I187 (gfint_1[27:27], choice_1, i_1r0[27:27]);
  AND2 I188 (gfint_1[28:28], choice_1, i_1r0[28:28]);
  AND2 I189 (gfint_1[29:29], choice_1, i_1r0[29:29]);
  AND2 I190 (gfint_1[30:30], choice_1, i_1r0[30:30]);
  AND2 I191 (gfint_1[31:31], choice_1, i_1r0[31:31]);
  OR2 I192 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I193 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I194 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I195 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I196 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I197 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I198 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I199 (comp0_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I200 (comp0_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I201 (comp0_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I202 (comp0_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I203 (comp0_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I204 (comp0_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I205 (comp0_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I206 (comp0_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I207 (comp0_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I208 (comp0_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I209 (comp0_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I210 (comp0_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I211 (comp0_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I212 (comp0_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I213 (comp0_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I214 (comp0_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I215 (comp0_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I216 (comp0_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I217 (comp0_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I218 (comp0_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I219 (comp0_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I220 (comp0_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I221 (comp0_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I222 (comp0_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I223 (comp0_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  C3 I224 (simp2351_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I225 (simp2351_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I226 (simp2351_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I227 (simp2351_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I228 (simp2351_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I229 (simp2351_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I230 (simp2351_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I231 (simp2351_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I232 (simp2351_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I233 (simp2351_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I234 (simp2351_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I235 (simp2352_0[0:0], simp2351_0[0:0], simp2351_0[1:1], simp2351_0[2:2]);
  C3 I236 (simp2352_0[1:1], simp2351_0[3:3], simp2351_0[4:4], simp2351_0[5:5]);
  C3 I237 (simp2352_0[2:2], simp2351_0[6:6], simp2351_0[7:7], simp2351_0[8:8]);
  C2 I238 (simp2352_0[3:3], simp2351_0[9:9], simp2351_0[10:10]);
  C3 I239 (simp2353_0[0:0], simp2352_0[0:0], simp2352_0[1:1], simp2352_0[2:2]);
  BUFF I240 (simp2353_0[1:1], simp2352_0[3:3]);
  C2 I241 (icomp_0, simp2353_0[0:0], simp2353_0[1:1]);
  OR2 I242 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I243 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I244 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I245 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I246 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I247 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I248 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  OR2 I249 (comp1_0[7:7], i_1r0[7:7], i_1r1[7:7]);
  OR2 I250 (comp1_0[8:8], i_1r0[8:8], i_1r1[8:8]);
  OR2 I251 (comp1_0[9:9], i_1r0[9:9], i_1r1[9:9]);
  OR2 I252 (comp1_0[10:10], i_1r0[10:10], i_1r1[10:10]);
  OR2 I253 (comp1_0[11:11], i_1r0[11:11], i_1r1[11:11]);
  OR2 I254 (comp1_0[12:12], i_1r0[12:12], i_1r1[12:12]);
  OR2 I255 (comp1_0[13:13], i_1r0[13:13], i_1r1[13:13]);
  OR2 I256 (comp1_0[14:14], i_1r0[14:14], i_1r1[14:14]);
  OR2 I257 (comp1_0[15:15], i_1r0[15:15], i_1r1[15:15]);
  OR2 I258 (comp1_0[16:16], i_1r0[16:16], i_1r1[16:16]);
  OR2 I259 (comp1_0[17:17], i_1r0[17:17], i_1r1[17:17]);
  OR2 I260 (comp1_0[18:18], i_1r0[18:18], i_1r1[18:18]);
  OR2 I261 (comp1_0[19:19], i_1r0[19:19], i_1r1[19:19]);
  OR2 I262 (comp1_0[20:20], i_1r0[20:20], i_1r1[20:20]);
  OR2 I263 (comp1_0[21:21], i_1r0[21:21], i_1r1[21:21]);
  OR2 I264 (comp1_0[22:22], i_1r0[22:22], i_1r1[22:22]);
  OR2 I265 (comp1_0[23:23], i_1r0[23:23], i_1r1[23:23]);
  OR2 I266 (comp1_0[24:24], i_1r0[24:24], i_1r1[24:24]);
  OR2 I267 (comp1_0[25:25], i_1r0[25:25], i_1r1[25:25]);
  OR2 I268 (comp1_0[26:26], i_1r0[26:26], i_1r1[26:26]);
  OR2 I269 (comp1_0[27:27], i_1r0[27:27], i_1r1[27:27]);
  OR2 I270 (comp1_0[28:28], i_1r0[28:28], i_1r1[28:28]);
  OR2 I271 (comp1_0[29:29], i_1r0[29:29], i_1r1[29:29]);
  OR2 I272 (comp1_0[30:30], i_1r0[30:30], i_1r1[30:30]);
  OR2 I273 (comp1_0[31:31], i_1r0[31:31], i_1r1[31:31]);
  C3 I274 (simp2691_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I275 (simp2691_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  C3 I276 (simp2691_0[2:2], comp1_0[6:6], comp1_0[7:7], comp1_0[8:8]);
  C3 I277 (simp2691_0[3:3], comp1_0[9:9], comp1_0[10:10], comp1_0[11:11]);
  C3 I278 (simp2691_0[4:4], comp1_0[12:12], comp1_0[13:13], comp1_0[14:14]);
  C3 I279 (simp2691_0[5:5], comp1_0[15:15], comp1_0[16:16], comp1_0[17:17]);
  C3 I280 (simp2691_0[6:6], comp1_0[18:18], comp1_0[19:19], comp1_0[20:20]);
  C3 I281 (simp2691_0[7:7], comp1_0[21:21], comp1_0[22:22], comp1_0[23:23]);
  C3 I282 (simp2691_0[8:8], comp1_0[24:24], comp1_0[25:25], comp1_0[26:26]);
  C3 I283 (simp2691_0[9:9], comp1_0[27:27], comp1_0[28:28], comp1_0[29:29]);
  C2 I284 (simp2691_0[10:10], comp1_0[30:30], comp1_0[31:31]);
  C3 I285 (simp2692_0[0:0], simp2691_0[0:0], simp2691_0[1:1], simp2691_0[2:2]);
  C3 I286 (simp2692_0[1:1], simp2691_0[3:3], simp2691_0[4:4], simp2691_0[5:5]);
  C3 I287 (simp2692_0[2:2], simp2691_0[6:6], simp2691_0[7:7], simp2691_0[8:8]);
  C2 I288 (simp2692_0[3:3], simp2691_0[9:9], simp2691_0[10:10]);
  C3 I289 (simp2693_0[0:0], simp2692_0[0:0], simp2692_0[1:1], simp2692_0[2:2]);
  BUFF I290 (simp2693_0[1:1], simp2692_0[3:3]);
  C2 I291 (icomp_1, simp2693_0[0:0], simp2693_0[1:1]);
  C2R I292 (choice_0, icomp_0, nchosen_0, reset);
  C2R I293 (choice_1, icomp_1, nchosen_0, reset);
  OR2 I294 (anychoice_0, choice_0, choice_1);
  NOR2 I295 (nchosen_0, anychoice_0, o_0a);
  C2R I296 (i_0a, choice_0, o_0a, reset);
  C2R I297 (i_1a, choice_1, o_0a, reset);
endmodule

// tkvACC32_wo0w32_ro0w32o31w1 TeakV "ACC" 32 [] [0] [0,31] [Many [32],Many [0],Many [0,0],Many [32,1]]
module tkvACC32_wo0w32_ro0w32o31w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output rd_1r0;
  output rd_1r1;
  input rd_1a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp4741_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0, df_0[31:31], rg_1r);
  AND2 I457 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I458 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I459 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I460 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I461 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I462 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I463 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I464 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I465 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I466 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I467 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I468 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I469 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I470 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I471 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I472 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I473 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I474 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I475 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I476 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I477 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I478 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I479 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I480 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I481 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I482 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I483 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I484 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I485 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I486 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I487 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I488 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I489 (rd_1r1, dt_0[31:31], rg_1r);
  NOR3 I490 (simp4741_0[0:0], rg_0r, rg_1r, rg_0a);
  INV I491 (simp4741_0[1:1], rg_1a);
  NAND2 I492 (anyread_0, simp4741_0[0:0], simp4741_0[1:1]);
  BUFF I493 (wg_0a, wd_0a);
  BUFF I494 (rg_0a, rd_0a);
  BUFF I495 (rg_1a, rd_1a);
endmodule

// tkf5mo0w0_o0w5 TeakF [0,0] [One 5,Many [0,5]]
module tkf5mo0w0_o0w5 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [4:0] i_0r0;
  input [4:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [4:0] o_1r0;
  output [4:0] o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_1r0[0:0], i_0r0[0:0]);
  BUFF I3 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I4 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I5 (o_1r0[3:3], i_0r0[3:3]);
  BUFF I6 (o_1r0[4:4], i_0r0[4:4]);
  BUFF I7 (o_1r1[0:0], i_0r1[0:0]);
  BUFF I8 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I9 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I10 (o_1r1[3:3], i_0r1[3:3]);
  BUFF I11 (o_1r1[4:4], i_0r1[4:4]);
  BUFF I12 (o_0r, icomplete_0);
  C3 I13 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tkm3x1b TeakM [Many [1,1,1],One 1]
module tkm3x1b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input i_1r0;
  input i_1r1;
  output i_1a;
  input i_2r0;
  input i_2r1;
  output i_2a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire gfint_0;
  wire gfint_1;
  wire gfint_2;
  wire gtint_0;
  wire gtint_1;
  wire gtint_2;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire nchosen_0;
  wire comp0_0;
  wire comp1_0;
  wire comp2_0;
  OR3 I0 (o_0r0, gfint_0, gfint_1, gfint_2);
  OR3 I1 (o_0r1, gtint_0, gtint_1, gtint_2);
  AND2 I2 (gtint_0, choice_0, i_0r1);
  AND2 I3 (gtint_1, choice_1, i_1r1);
  AND2 I4 (gtint_2, choice_2, i_2r1);
  AND2 I5 (gfint_0, choice_0, i_0r0);
  AND2 I6 (gfint_1, choice_1, i_1r0);
  AND2 I7 (gfint_2, choice_2, i_2r0);
  OR2 I8 (comp0_0, i_0r0, i_0r1);
  BUFF I9 (icomp_0, comp0_0);
  OR2 I10 (comp1_0, i_1r0, i_1r1);
  BUFF I11 (icomp_1, comp1_0);
  OR2 I12 (comp2_0, i_2r0, i_2r1);
  BUFF I13 (icomp_2, comp2_0);
  C2R I14 (choice_0, icomp_0, nchosen_0, reset);
  C2R I15 (choice_1, icomp_1, nchosen_0, reset);
  C2R I16 (choice_2, icomp_2, nchosen_0, reset);
  OR3 I17 (anychoice_0, choice_0, choice_1, choice_2);
  NOR2 I18 (nchosen_0, anychoice_0, o_0a);
  C2R I19 (i_0a, choice_0, o_0a, reset);
  C2R I20 (i_1a, choice_1, o_0a, reset);
  C2R I21 (i_2a, choice_2, o_0a, reset);
endmodule

// tkf1mo0w0_o0w1 TeakF [0,0] [One 1,Many [0,1]]
module tkf1mo0w0_o0w1 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r0;
  output o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0, i_0r1);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_1r0, i_0r0);
  BUFF I3 (o_1r1, i_0r1);
  BUFF I4 (o_0r, icomplete_0);
  C3 I5 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tko0m3_1nm3b1 TeakO [
//     (1,TeakOConstant 3 1)] [One 0,One 3]
module tko0m3_1nm3b1 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  GND I1 (o_0r0[0:0]);
  BUFF I2 (o_0r0[1:1], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  GND I4 (o_0r1[1:1]);
  GND I5 (o_0r1[2:2]);
  BUFF I6 (i_0a, o_0a);
endmodule

// tkm3x3b TeakM [Many [3,3,3],One 3]
module tkm3x3b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, o_0r0, o_0r1, o_0a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  input [2:0] i_1r0;
  input [2:0] i_1r1;
  output i_1a;
  input [2:0] i_2r0;
  input [2:0] i_2r1;
  output i_2a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire [2:0] gfint_0;
  wire [2:0] gfint_1;
  wire [2:0] gfint_2;
  wire [2:0] gtint_0;
  wire [2:0] gtint_1;
  wire [2:0] gtint_2;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire nchosen_0;
  wire [2:0] comp0_0;
  wire [2:0] comp1_0;
  wire [2:0] comp2_0;
  OR3 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  OR3 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  OR3 I2 (o_0r0[2:2], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  OR3 I3 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  OR3 I4 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  OR3 I5 (o_0r1[2:2], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  AND2 I6 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I7 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I8 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I9 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I10 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I11 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I12 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I13 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I14 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I15 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I16 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I17 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I18 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I19 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I20 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I21 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I22 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I23 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  OR2 I24 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I25 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I26 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I27 (icomp_0, comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  OR2 I28 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I29 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I30 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  C3 I31 (icomp_1, comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  OR2 I32 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I33 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I34 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  C3 I35 (icomp_2, comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C2R I36 (choice_0, icomp_0, nchosen_0, reset);
  C2R I37 (choice_1, icomp_1, nchosen_0, reset);
  C2R I38 (choice_2, icomp_2, nchosen_0, reset);
  OR3 I39 (anychoice_0, choice_0, choice_1, choice_2);
  NOR2 I40 (nchosen_0, anychoice_0, o_0a);
  C2R I41 (i_0a, choice_0, o_0a, reset);
  C2R I42 (i_1a, choice_1, o_0a, reset);
  C2R I43 (i_2a, choice_2, o_0a, reset);
endmodule

// tkj34m32_2 TeakJ [Many [32,2],One 34]
module tkj34m32_2 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [1:0] i_1r0;
  input [1:0] i_1r1;
  output i_1a;
  output [33:0] o_0r0;
  output [33:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [33:0] joinf_0;
  wire [33:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joinf_0[32:32], i_1r0[0:0]);
  BUFF I33 (joinf_0[33:33], i_1r0[1:1]);
  BUFF I34 (joint_0[0:0], i_0r1[0:0]);
  BUFF I35 (joint_0[1:1], i_0r1[1:1]);
  BUFF I36 (joint_0[2:2], i_0r1[2:2]);
  BUFF I37 (joint_0[3:3], i_0r1[3:3]);
  BUFF I38 (joint_0[4:4], i_0r1[4:4]);
  BUFF I39 (joint_0[5:5], i_0r1[5:5]);
  BUFF I40 (joint_0[6:6], i_0r1[6:6]);
  BUFF I41 (joint_0[7:7], i_0r1[7:7]);
  BUFF I42 (joint_0[8:8], i_0r1[8:8]);
  BUFF I43 (joint_0[9:9], i_0r1[9:9]);
  BUFF I44 (joint_0[10:10], i_0r1[10:10]);
  BUFF I45 (joint_0[11:11], i_0r1[11:11]);
  BUFF I46 (joint_0[12:12], i_0r1[12:12]);
  BUFF I47 (joint_0[13:13], i_0r1[13:13]);
  BUFF I48 (joint_0[14:14], i_0r1[14:14]);
  BUFF I49 (joint_0[15:15], i_0r1[15:15]);
  BUFF I50 (joint_0[16:16], i_0r1[16:16]);
  BUFF I51 (joint_0[17:17], i_0r1[17:17]);
  BUFF I52 (joint_0[18:18], i_0r1[18:18]);
  BUFF I53 (joint_0[19:19], i_0r1[19:19]);
  BUFF I54 (joint_0[20:20], i_0r1[20:20]);
  BUFF I55 (joint_0[21:21], i_0r1[21:21]);
  BUFF I56 (joint_0[22:22], i_0r1[22:22]);
  BUFF I57 (joint_0[23:23], i_0r1[23:23]);
  BUFF I58 (joint_0[24:24], i_0r1[24:24]);
  BUFF I59 (joint_0[25:25], i_0r1[25:25]);
  BUFF I60 (joint_0[26:26], i_0r1[26:26]);
  BUFF I61 (joint_0[27:27], i_0r1[27:27]);
  BUFF I62 (joint_0[28:28], i_0r1[28:28]);
  BUFF I63 (joint_0[29:29], i_0r1[29:29]);
  BUFF I64 (joint_0[30:30], i_0r1[30:30]);
  BUFF I65 (joint_0[31:31], i_0r1[31:31]);
  BUFF I66 (joint_0[32:32], i_1r1[0:0]);
  BUFF I67 (joint_0[33:33], i_1r1[1:1]);
  OR2 I68 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I69 (icomplete_0, dcomplete_0);
  C2 I70 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I71 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I72 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I73 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I74 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I75 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I76 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I77 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I78 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I79 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I80 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I81 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I82 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I83 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I84 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I85 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I86 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I87 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I88 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I89 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I90 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I91 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I92 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I93 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I94 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I95 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I96 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I97 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I98 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I99 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I100 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I101 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I102 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I103 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I104 (o_0r0[33:33], joinf_0[33:33]);
  BUFF I105 (o_0r1[1:1], joint_0[1:1]);
  BUFF I106 (o_0r1[2:2], joint_0[2:2]);
  BUFF I107 (o_0r1[3:3], joint_0[3:3]);
  BUFF I108 (o_0r1[4:4], joint_0[4:4]);
  BUFF I109 (o_0r1[5:5], joint_0[5:5]);
  BUFF I110 (o_0r1[6:6], joint_0[6:6]);
  BUFF I111 (o_0r1[7:7], joint_0[7:7]);
  BUFF I112 (o_0r1[8:8], joint_0[8:8]);
  BUFF I113 (o_0r1[9:9], joint_0[9:9]);
  BUFF I114 (o_0r1[10:10], joint_0[10:10]);
  BUFF I115 (o_0r1[11:11], joint_0[11:11]);
  BUFF I116 (o_0r1[12:12], joint_0[12:12]);
  BUFF I117 (o_0r1[13:13], joint_0[13:13]);
  BUFF I118 (o_0r1[14:14], joint_0[14:14]);
  BUFF I119 (o_0r1[15:15], joint_0[15:15]);
  BUFF I120 (o_0r1[16:16], joint_0[16:16]);
  BUFF I121 (o_0r1[17:17], joint_0[17:17]);
  BUFF I122 (o_0r1[18:18], joint_0[18:18]);
  BUFF I123 (o_0r1[19:19], joint_0[19:19]);
  BUFF I124 (o_0r1[20:20], joint_0[20:20]);
  BUFF I125 (o_0r1[21:21], joint_0[21:21]);
  BUFF I126 (o_0r1[22:22], joint_0[22:22]);
  BUFF I127 (o_0r1[23:23], joint_0[23:23]);
  BUFF I128 (o_0r1[24:24], joint_0[24:24]);
  BUFF I129 (o_0r1[25:25], joint_0[25:25]);
  BUFF I130 (o_0r1[26:26], joint_0[26:26]);
  BUFF I131 (o_0r1[27:27], joint_0[27:27]);
  BUFF I132 (o_0r1[28:28], joint_0[28:28]);
  BUFF I133 (o_0r1[29:29], joint_0[29:29]);
  BUFF I134 (o_0r1[30:30], joint_0[30:30]);
  BUFF I135 (o_0r1[31:31], joint_0[31:31]);
  BUFF I136 (o_0r1[32:32], joint_0[32:32]);
  BUFF I137 (o_0r1[33:33], joint_0[33:33]);
  BUFF I138 (i_0a, o_0a);
  BUFF I139 (i_1a, o_0a);
endmodule

// tks34_o32w2_1o0w32_2o0w32 TeakS (32+:2) [([Imp 1 0],0),([Imp 2 0],0)] [One 34,Many [32,32]]
module tks34_o32w2_1o0w32_2o0w32 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [33:0] i_0r0;
  input [33:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  output [31:0] o_1r0;
  output [31:0] o_1r1;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire [33:0] comp_0;
  wire [11:0] simp491_0;
  wire [3:0] simp492_0;
  wire [1:0] simp493_0;
  BUFF I0 (sel_0, match0_0);
  C2 I1 (match0_0, i_0r1[32:32], i_0r0[33:33]);
  BUFF I2 (sel_1, match1_0);
  C2 I3 (match1_0, i_0r0[32:32], i_0r1[33:33]);
  C2 I4 (gsel_0, sel_0, icomplete_0);
  C2 I5 (gsel_1, sel_1, icomplete_0);
  OR2 I6 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I7 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I8 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I9 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I10 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I11 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I12 (comp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I13 (comp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I14 (comp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I15 (comp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I16 (comp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I17 (comp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I18 (comp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I19 (comp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I20 (comp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I21 (comp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I22 (comp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I23 (comp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I24 (comp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I25 (comp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I26 (comp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I27 (comp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I28 (comp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I29 (comp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I30 (comp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I31 (comp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I32 (comp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I33 (comp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I34 (comp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I35 (comp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I36 (comp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I37 (comp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I38 (comp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  OR2 I39 (comp_0[33:33], i_0r0[33:33], i_0r1[33:33]);
  C3 I40 (simp491_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I41 (simp491_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C3 I42 (simp491_0[2:2], comp_0[6:6], comp_0[7:7], comp_0[8:8]);
  C3 I43 (simp491_0[3:3], comp_0[9:9], comp_0[10:10], comp_0[11:11]);
  C3 I44 (simp491_0[4:4], comp_0[12:12], comp_0[13:13], comp_0[14:14]);
  C3 I45 (simp491_0[5:5], comp_0[15:15], comp_0[16:16], comp_0[17:17]);
  C3 I46 (simp491_0[6:6], comp_0[18:18], comp_0[19:19], comp_0[20:20]);
  C3 I47 (simp491_0[7:7], comp_0[21:21], comp_0[22:22], comp_0[23:23]);
  C3 I48 (simp491_0[8:8], comp_0[24:24], comp_0[25:25], comp_0[26:26]);
  C3 I49 (simp491_0[9:9], comp_0[27:27], comp_0[28:28], comp_0[29:29]);
  C3 I50 (simp491_0[10:10], comp_0[30:30], comp_0[31:31], comp_0[32:32]);
  BUFF I51 (simp491_0[11:11], comp_0[33:33]);
  C3 I52 (simp492_0[0:0], simp491_0[0:0], simp491_0[1:1], simp491_0[2:2]);
  C3 I53 (simp492_0[1:1], simp491_0[3:3], simp491_0[4:4], simp491_0[5:5]);
  C3 I54 (simp492_0[2:2], simp491_0[6:6], simp491_0[7:7], simp491_0[8:8]);
  C3 I55 (simp492_0[3:3], simp491_0[9:9], simp491_0[10:10], simp491_0[11:11]);
  C3 I56 (simp493_0[0:0], simp492_0[0:0], simp492_0[1:1], simp492_0[2:2]);
  BUFF I57 (simp493_0[1:1], simp492_0[3:3]);
  C2 I58 (icomplete_0, simp493_0[0:0], simp493_0[1:1]);
  C2 I59 (o_0r0[0:0], i_0r0[0:0], gsel_0);
  C2 I60 (o_0r0[1:1], i_0r0[1:1], gsel_0);
  C2 I61 (o_0r0[2:2], i_0r0[2:2], gsel_0);
  C2 I62 (o_0r0[3:3], i_0r0[3:3], gsel_0);
  C2 I63 (o_0r0[4:4], i_0r0[4:4], gsel_0);
  C2 I64 (o_0r0[5:5], i_0r0[5:5], gsel_0);
  C2 I65 (o_0r0[6:6], i_0r0[6:6], gsel_0);
  C2 I66 (o_0r0[7:7], i_0r0[7:7], gsel_0);
  C2 I67 (o_0r0[8:8], i_0r0[8:8], gsel_0);
  C2 I68 (o_0r0[9:9], i_0r0[9:9], gsel_0);
  C2 I69 (o_0r0[10:10], i_0r0[10:10], gsel_0);
  C2 I70 (o_0r0[11:11], i_0r0[11:11], gsel_0);
  C2 I71 (o_0r0[12:12], i_0r0[12:12], gsel_0);
  C2 I72 (o_0r0[13:13], i_0r0[13:13], gsel_0);
  C2 I73 (o_0r0[14:14], i_0r0[14:14], gsel_0);
  C2 I74 (o_0r0[15:15], i_0r0[15:15], gsel_0);
  C2 I75 (o_0r0[16:16], i_0r0[16:16], gsel_0);
  C2 I76 (o_0r0[17:17], i_0r0[17:17], gsel_0);
  C2 I77 (o_0r0[18:18], i_0r0[18:18], gsel_0);
  C2 I78 (o_0r0[19:19], i_0r0[19:19], gsel_0);
  C2 I79 (o_0r0[20:20], i_0r0[20:20], gsel_0);
  C2 I80 (o_0r0[21:21], i_0r0[21:21], gsel_0);
  C2 I81 (o_0r0[22:22], i_0r0[22:22], gsel_0);
  C2 I82 (o_0r0[23:23], i_0r0[23:23], gsel_0);
  C2 I83 (o_0r0[24:24], i_0r0[24:24], gsel_0);
  C2 I84 (o_0r0[25:25], i_0r0[25:25], gsel_0);
  C2 I85 (o_0r0[26:26], i_0r0[26:26], gsel_0);
  C2 I86 (o_0r0[27:27], i_0r0[27:27], gsel_0);
  C2 I87 (o_0r0[28:28], i_0r0[28:28], gsel_0);
  C2 I88 (o_0r0[29:29], i_0r0[29:29], gsel_0);
  C2 I89 (o_0r0[30:30], i_0r0[30:30], gsel_0);
  C2 I90 (o_0r0[31:31], i_0r0[31:31], gsel_0);
  C2 I91 (o_1r0[0:0], i_0r0[0:0], gsel_1);
  C2 I92 (o_1r0[1:1], i_0r0[1:1], gsel_1);
  C2 I93 (o_1r0[2:2], i_0r0[2:2], gsel_1);
  C2 I94 (o_1r0[3:3], i_0r0[3:3], gsel_1);
  C2 I95 (o_1r0[4:4], i_0r0[4:4], gsel_1);
  C2 I96 (o_1r0[5:5], i_0r0[5:5], gsel_1);
  C2 I97 (o_1r0[6:6], i_0r0[6:6], gsel_1);
  C2 I98 (o_1r0[7:7], i_0r0[7:7], gsel_1);
  C2 I99 (o_1r0[8:8], i_0r0[8:8], gsel_1);
  C2 I100 (o_1r0[9:9], i_0r0[9:9], gsel_1);
  C2 I101 (o_1r0[10:10], i_0r0[10:10], gsel_1);
  C2 I102 (o_1r0[11:11], i_0r0[11:11], gsel_1);
  C2 I103 (o_1r0[12:12], i_0r0[12:12], gsel_1);
  C2 I104 (o_1r0[13:13], i_0r0[13:13], gsel_1);
  C2 I105 (o_1r0[14:14], i_0r0[14:14], gsel_1);
  C2 I106 (o_1r0[15:15], i_0r0[15:15], gsel_1);
  C2 I107 (o_1r0[16:16], i_0r0[16:16], gsel_1);
  C2 I108 (o_1r0[17:17], i_0r0[17:17], gsel_1);
  C2 I109 (o_1r0[18:18], i_0r0[18:18], gsel_1);
  C2 I110 (o_1r0[19:19], i_0r0[19:19], gsel_1);
  C2 I111 (o_1r0[20:20], i_0r0[20:20], gsel_1);
  C2 I112 (o_1r0[21:21], i_0r0[21:21], gsel_1);
  C2 I113 (o_1r0[22:22], i_0r0[22:22], gsel_1);
  C2 I114 (o_1r0[23:23], i_0r0[23:23], gsel_1);
  C2 I115 (o_1r0[24:24], i_0r0[24:24], gsel_1);
  C2 I116 (o_1r0[25:25], i_0r0[25:25], gsel_1);
  C2 I117 (o_1r0[26:26], i_0r0[26:26], gsel_1);
  C2 I118 (o_1r0[27:27], i_0r0[27:27], gsel_1);
  C2 I119 (o_1r0[28:28], i_0r0[28:28], gsel_1);
  C2 I120 (o_1r0[29:29], i_0r0[29:29], gsel_1);
  C2 I121 (o_1r0[30:30], i_0r0[30:30], gsel_1);
  C2 I122 (o_1r0[31:31], i_0r0[31:31], gsel_1);
  C2 I123 (o_0r1[0:0], i_0r1[0:0], gsel_0);
  C2 I124 (o_0r1[1:1], i_0r1[1:1], gsel_0);
  C2 I125 (o_0r1[2:2], i_0r1[2:2], gsel_0);
  C2 I126 (o_0r1[3:3], i_0r1[3:3], gsel_0);
  C2 I127 (o_0r1[4:4], i_0r1[4:4], gsel_0);
  C2 I128 (o_0r1[5:5], i_0r1[5:5], gsel_0);
  C2 I129 (o_0r1[6:6], i_0r1[6:6], gsel_0);
  C2 I130 (o_0r1[7:7], i_0r1[7:7], gsel_0);
  C2 I131 (o_0r1[8:8], i_0r1[8:8], gsel_0);
  C2 I132 (o_0r1[9:9], i_0r1[9:9], gsel_0);
  C2 I133 (o_0r1[10:10], i_0r1[10:10], gsel_0);
  C2 I134 (o_0r1[11:11], i_0r1[11:11], gsel_0);
  C2 I135 (o_0r1[12:12], i_0r1[12:12], gsel_0);
  C2 I136 (o_0r1[13:13], i_0r1[13:13], gsel_0);
  C2 I137 (o_0r1[14:14], i_0r1[14:14], gsel_0);
  C2 I138 (o_0r1[15:15], i_0r1[15:15], gsel_0);
  C2 I139 (o_0r1[16:16], i_0r1[16:16], gsel_0);
  C2 I140 (o_0r1[17:17], i_0r1[17:17], gsel_0);
  C2 I141 (o_0r1[18:18], i_0r1[18:18], gsel_0);
  C2 I142 (o_0r1[19:19], i_0r1[19:19], gsel_0);
  C2 I143 (o_0r1[20:20], i_0r1[20:20], gsel_0);
  C2 I144 (o_0r1[21:21], i_0r1[21:21], gsel_0);
  C2 I145 (o_0r1[22:22], i_0r1[22:22], gsel_0);
  C2 I146 (o_0r1[23:23], i_0r1[23:23], gsel_0);
  C2 I147 (o_0r1[24:24], i_0r1[24:24], gsel_0);
  C2 I148 (o_0r1[25:25], i_0r1[25:25], gsel_0);
  C2 I149 (o_0r1[26:26], i_0r1[26:26], gsel_0);
  C2 I150 (o_0r1[27:27], i_0r1[27:27], gsel_0);
  C2 I151 (o_0r1[28:28], i_0r1[28:28], gsel_0);
  C2 I152 (o_0r1[29:29], i_0r1[29:29], gsel_0);
  C2 I153 (o_0r1[30:30], i_0r1[30:30], gsel_0);
  C2 I154 (o_0r1[31:31], i_0r1[31:31], gsel_0);
  C2 I155 (o_1r1[0:0], i_0r1[0:0], gsel_1);
  C2 I156 (o_1r1[1:1], i_0r1[1:1], gsel_1);
  C2 I157 (o_1r1[2:2], i_0r1[2:2], gsel_1);
  C2 I158 (o_1r1[3:3], i_0r1[3:3], gsel_1);
  C2 I159 (o_1r1[4:4], i_0r1[4:4], gsel_1);
  C2 I160 (o_1r1[5:5], i_0r1[5:5], gsel_1);
  C2 I161 (o_1r1[6:6], i_0r1[6:6], gsel_1);
  C2 I162 (o_1r1[7:7], i_0r1[7:7], gsel_1);
  C2 I163 (o_1r1[8:8], i_0r1[8:8], gsel_1);
  C2 I164 (o_1r1[9:9], i_0r1[9:9], gsel_1);
  C2 I165 (o_1r1[10:10], i_0r1[10:10], gsel_1);
  C2 I166 (o_1r1[11:11], i_0r1[11:11], gsel_1);
  C2 I167 (o_1r1[12:12], i_0r1[12:12], gsel_1);
  C2 I168 (o_1r1[13:13], i_0r1[13:13], gsel_1);
  C2 I169 (o_1r1[14:14], i_0r1[14:14], gsel_1);
  C2 I170 (o_1r1[15:15], i_0r1[15:15], gsel_1);
  C2 I171 (o_1r1[16:16], i_0r1[16:16], gsel_1);
  C2 I172 (o_1r1[17:17], i_0r1[17:17], gsel_1);
  C2 I173 (o_1r1[18:18], i_0r1[18:18], gsel_1);
  C2 I174 (o_1r1[19:19], i_0r1[19:19], gsel_1);
  C2 I175 (o_1r1[20:20], i_0r1[20:20], gsel_1);
  C2 I176 (o_1r1[21:21], i_0r1[21:21], gsel_1);
  C2 I177 (o_1r1[22:22], i_0r1[22:22], gsel_1);
  C2 I178 (o_1r1[23:23], i_0r1[23:23], gsel_1);
  C2 I179 (o_1r1[24:24], i_0r1[24:24], gsel_1);
  C2 I180 (o_1r1[25:25], i_0r1[25:25], gsel_1);
  C2 I181 (o_1r1[26:26], i_0r1[26:26], gsel_1);
  C2 I182 (o_1r1[27:27], i_0r1[27:27], gsel_1);
  C2 I183 (o_1r1[28:28], i_0r1[28:28], gsel_1);
  C2 I184 (o_1r1[29:29], i_0r1[29:29], gsel_1);
  C2 I185 (o_1r1[30:30], i_0r1[30:30], gsel_1);
  C2 I186 (o_1r1[31:31], i_0r1[31:31], gsel_1);
  OR2 I187 (oack_0, o_0a, o_1a);
  C2 I188 (i_0a, oack_0, icomplete_0);
endmodule

// tkf32mo0w32_o13w3 TeakF [0,13] [One 32,Many [32,3]]
module tkf32mo0w32_o13w3 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  output [2:0] o_1r0;
  output [2:0] o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_0r0[0:0], i_0r0[0:0]);
  BUFF I3 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I4 (o_0r0[2:2], i_0r0[2:2]);
  BUFF I5 (o_0r0[3:3], i_0r0[3:3]);
  BUFF I6 (o_0r0[4:4], i_0r0[4:4]);
  BUFF I7 (o_0r0[5:5], i_0r0[5:5]);
  BUFF I8 (o_0r0[6:6], i_0r0[6:6]);
  BUFF I9 (o_0r0[7:7], i_0r0[7:7]);
  BUFF I10 (o_0r0[8:8], i_0r0[8:8]);
  BUFF I11 (o_0r0[9:9], i_0r0[9:9]);
  BUFF I12 (o_0r0[10:10], i_0r0[10:10]);
  BUFF I13 (o_0r0[11:11], i_0r0[11:11]);
  BUFF I14 (o_0r0[12:12], i_0r0[12:12]);
  BUFF I15 (o_0r0[13:13], i_0r0[13:13]);
  BUFF I16 (o_0r0[14:14], i_0r0[14:14]);
  BUFF I17 (o_0r0[15:15], i_0r0[15:15]);
  BUFF I18 (o_0r0[16:16], i_0r0[16:16]);
  BUFF I19 (o_0r0[17:17], i_0r0[17:17]);
  BUFF I20 (o_0r0[18:18], i_0r0[18:18]);
  BUFF I21 (o_0r0[19:19], i_0r0[19:19]);
  BUFF I22 (o_0r0[20:20], i_0r0[20:20]);
  BUFF I23 (o_0r0[21:21], i_0r0[21:21]);
  BUFF I24 (o_0r0[22:22], i_0r0[22:22]);
  BUFF I25 (o_0r0[23:23], i_0r0[23:23]);
  BUFF I26 (o_0r0[24:24], i_0r0[24:24]);
  BUFF I27 (o_0r0[25:25], i_0r0[25:25]);
  BUFF I28 (o_0r0[26:26], i_0r0[26:26]);
  BUFF I29 (o_0r0[27:27], i_0r0[27:27]);
  BUFF I30 (o_0r0[28:28], i_0r0[28:28]);
  BUFF I31 (o_0r0[29:29], i_0r0[29:29]);
  BUFF I32 (o_0r0[30:30], i_0r0[30:30]);
  BUFF I33 (o_0r0[31:31], i_0r0[31:31]);
  C2 I34 (o_1r0[0:0], i_0r0[13:13], icomplete_0);
  BUFF I35 (o_1r0[1:1], i_0r0[14:14]);
  BUFF I36 (o_1r0[2:2], i_0r0[15:15]);
  BUFF I37 (o_0r1[0:0], i_0r1[0:0]);
  BUFF I38 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I39 (o_0r1[2:2], i_0r1[2:2]);
  BUFF I40 (o_0r1[3:3], i_0r1[3:3]);
  BUFF I41 (o_0r1[4:4], i_0r1[4:4]);
  BUFF I42 (o_0r1[5:5], i_0r1[5:5]);
  BUFF I43 (o_0r1[6:6], i_0r1[6:6]);
  BUFF I44 (o_0r1[7:7], i_0r1[7:7]);
  BUFF I45 (o_0r1[8:8], i_0r1[8:8]);
  BUFF I46 (o_0r1[9:9], i_0r1[9:9]);
  BUFF I47 (o_0r1[10:10], i_0r1[10:10]);
  BUFF I48 (o_0r1[11:11], i_0r1[11:11]);
  BUFF I49 (o_0r1[12:12], i_0r1[12:12]);
  BUFF I50 (o_0r1[13:13], i_0r1[13:13]);
  BUFF I51 (o_0r1[14:14], i_0r1[14:14]);
  BUFF I52 (o_0r1[15:15], i_0r1[15:15]);
  BUFF I53 (o_0r1[16:16], i_0r1[16:16]);
  BUFF I54 (o_0r1[17:17], i_0r1[17:17]);
  BUFF I55 (o_0r1[18:18], i_0r1[18:18]);
  BUFF I56 (o_0r1[19:19], i_0r1[19:19]);
  BUFF I57 (o_0r1[20:20], i_0r1[20:20]);
  BUFF I58 (o_0r1[21:21], i_0r1[21:21]);
  BUFF I59 (o_0r1[22:22], i_0r1[22:22]);
  BUFF I60 (o_0r1[23:23], i_0r1[23:23]);
  BUFF I61 (o_0r1[24:24], i_0r1[24:24]);
  BUFF I62 (o_0r1[25:25], i_0r1[25:25]);
  BUFF I63 (o_0r1[26:26], i_0r1[26:26]);
  BUFF I64 (o_0r1[27:27], i_0r1[27:27]);
  BUFF I65 (o_0r1[28:28], i_0r1[28:28]);
  BUFF I66 (o_0r1[29:29], i_0r1[29:29]);
  BUFF I67 (o_0r1[30:30], i_0r1[30:30]);
  BUFF I68 (o_0r1[31:31], i_0r1[31:31]);
  C2 I69 (o_1r1[0:0], i_0r1[13:13], icomplete_0);
  BUFF I70 (o_1r1[1:1], i_0r1[14:14]);
  BUFF I71 (o_1r1[2:2], i_0r1[15:15]);
  C3 I72 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tkj3m3_0_0_0 TeakJ [Many [3,0,0,0],One 3]
module tkj3m3_0_0_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, i_2r, i_2a, i_3r, i_3a, o_0r0, o_0r1, o_0a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [2:0] joinf_0;
  wire [2:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joint_0[0:0], i_0r1[0:0]);
  BUFF I4 (joint_0[1:1], i_0r1[1:1]);
  BUFF I5 (joint_0[2:2], i_0r1[2:2]);
  C3 I6 (icomplete_0, i_1r, i_2r, i_3r);
  C2 I7 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I8 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I9 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I10 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I11 (o_0r1[1:1], joint_0[1:1]);
  BUFF I12 (o_0r1[2:2], joint_0[2:2]);
  BUFF I13 (i_0a, o_0a);
  BUFF I14 (i_1a, o_0a);
  BUFF I15 (i_2a, o_0a);
  BUFF I16 (i_3a, o_0a);
endmodule

// tkf3mo0w3_o0w0 TeakF [0,0] [One 3,Many [3,0]]
module tkf3mo0w3_o0w0 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r, o_1a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_0r0[0:0], i_0r0[0:0]);
  BUFF I3 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I4 (o_0r0[2:2], i_0r0[2:2]);
  BUFF I5 (o_0r1[0:0], i_0r1[0:0]);
  BUFF I6 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I7 (o_0r1[2:2], i_0r1[2:2]);
  BUFF I8 (o_1r, icomplete_0);
  C3 I9 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tkf2mo0w2_o0w0 TeakF [0,0] [One 2,Many [2,0]]
module tkf2mo0w2_o0w0 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r, o_1a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_0r0[0:0], i_0r0[0:0]);
  BUFF I3 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I4 (o_0r1[0:0], i_0r1[0:0]);
  BUFF I5 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I6 (o_1r, icomplete_0);
  C3 I7 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tko64m32_1nm2b0_2api0w32bt1o0w2b_3nm2b0_4api32w32bt3o0w2b_5subt2o0w34bt4o0w34b_6apt5o0w32b TeakO [
//     (1,TeakOConstant 2 0),
//     (2,TeakOAppend 1 [(0,0+:32),(1,0+:2)]),
//     (3,TeakOConstant 2 0),
//     (4,TeakOAppend 1 [(0,32+:32),(3,0+:2)]),
//     (5,TeakOp TeakOpSub [(2,0+:34),(4,0+:34)]),
//     (6,TeakOAppend 1 [(5,0+:32)])] [One 64,One 32]
module tko64m32_1nm2b0_2api0w32bt1o0w2b_3nm2b0_4api32w32bt3o0w2b_5subt2o0w34bt4o0w34b_6apt5o0w32b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [63:0] i_0r0;
  input [63:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [63:0] gocomp_0;
  wire [21:0] simp661_0;
  wire [7:0] simp662_0;
  wire [2:0] simp663_0;
  wire [1:0] termf_1;
  wire [33:0] termf_2;
  wire [1:0] termf_3;
  wire [33:0] termf_4;
  wire [33:0] termf_5;
  wire [1:0] termt_1;
  wire [33:0] termt_2;
  wire [1:0] termt_3;
  wire [33:0] termt_4;
  wire [33:0] termt_5;
  wire [33:0] cf5__0;
  wire [33:0] ct5__0;
  wire [3:0] ha5__0;
  wire [7:0] fa5_1min_0;
  wire [1:0] simp2391_0;
  wire [1:0] simp2401_0;
  wire [7:0] fa5_2min_0;
  wire [1:0] simp2521_0;
  wire [1:0] simp2531_0;
  wire [7:0] fa5_3min_0;
  wire [1:0] simp2651_0;
  wire [1:0] simp2661_0;
  wire [7:0] fa5_4min_0;
  wire [1:0] simp2781_0;
  wire [1:0] simp2791_0;
  wire [7:0] fa5_5min_0;
  wire [1:0] simp2911_0;
  wire [1:0] simp2921_0;
  wire [7:0] fa5_6min_0;
  wire [1:0] simp3041_0;
  wire [1:0] simp3051_0;
  wire [7:0] fa5_7min_0;
  wire [1:0] simp3171_0;
  wire [1:0] simp3181_0;
  wire [7:0] fa5_8min_0;
  wire [1:0] simp3301_0;
  wire [1:0] simp3311_0;
  wire [7:0] fa5_9min_0;
  wire [1:0] simp3431_0;
  wire [1:0] simp3441_0;
  wire [7:0] fa5_10min_0;
  wire [1:0] simp3561_0;
  wire [1:0] simp3571_0;
  wire [7:0] fa5_11min_0;
  wire [1:0] simp3691_0;
  wire [1:0] simp3701_0;
  wire [7:0] fa5_12min_0;
  wire [1:0] simp3821_0;
  wire [1:0] simp3831_0;
  wire [7:0] fa5_13min_0;
  wire [1:0] simp3951_0;
  wire [1:0] simp3961_0;
  wire [7:0] fa5_14min_0;
  wire [1:0] simp4081_0;
  wire [1:0] simp4091_0;
  wire [7:0] fa5_15min_0;
  wire [1:0] simp4211_0;
  wire [1:0] simp4221_0;
  wire [7:0] fa5_16min_0;
  wire [1:0] simp4341_0;
  wire [1:0] simp4351_0;
  wire [7:0] fa5_17min_0;
  wire [1:0] simp4471_0;
  wire [1:0] simp4481_0;
  wire [7:0] fa5_18min_0;
  wire [1:0] simp4601_0;
  wire [1:0] simp4611_0;
  wire [7:0] fa5_19min_0;
  wire [1:0] simp4731_0;
  wire [1:0] simp4741_0;
  wire [7:0] fa5_20min_0;
  wire [1:0] simp4861_0;
  wire [1:0] simp4871_0;
  wire [7:0] fa5_21min_0;
  wire [1:0] simp4991_0;
  wire [1:0] simp5001_0;
  wire [7:0] fa5_22min_0;
  wire [1:0] simp5121_0;
  wire [1:0] simp5131_0;
  wire [7:0] fa5_23min_0;
  wire [1:0] simp5251_0;
  wire [1:0] simp5261_0;
  wire [7:0] fa5_24min_0;
  wire [1:0] simp5381_0;
  wire [1:0] simp5391_0;
  wire [7:0] fa5_25min_0;
  wire [1:0] simp5511_0;
  wire [1:0] simp5521_0;
  wire [7:0] fa5_26min_0;
  wire [1:0] simp5641_0;
  wire [1:0] simp5651_0;
  wire [7:0] fa5_27min_0;
  wire [1:0] simp5771_0;
  wire [1:0] simp5781_0;
  wire [7:0] fa5_28min_0;
  wire [1:0] simp5901_0;
  wire [1:0] simp5911_0;
  wire [7:0] fa5_29min_0;
  wire [1:0] simp6031_0;
  wire [1:0] simp6041_0;
  wire [7:0] fa5_30min_0;
  wire [1:0] simp6161_0;
  wire [1:0] simp6171_0;
  wire [7:0] fa5_31min_0;
  wire [1:0] simp6291_0;
  wire [1:0] simp6301_0;
  wire [7:0] fa5_32min_0;
  wire [1:0] simp6421_0;
  wire [1:0] simp6431_0;
  wire [7:0] fa5_33min_0;
  wire [1:0] simp6551_0;
  wire [1:0] simp6561_0;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I30 (gocomp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I31 (gocomp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I32 (gocomp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  OR2 I33 (gocomp_0[33:33], i_0r0[33:33], i_0r1[33:33]);
  OR2 I34 (gocomp_0[34:34], i_0r0[34:34], i_0r1[34:34]);
  OR2 I35 (gocomp_0[35:35], i_0r0[35:35], i_0r1[35:35]);
  OR2 I36 (gocomp_0[36:36], i_0r0[36:36], i_0r1[36:36]);
  OR2 I37 (gocomp_0[37:37], i_0r0[37:37], i_0r1[37:37]);
  OR2 I38 (gocomp_0[38:38], i_0r0[38:38], i_0r1[38:38]);
  OR2 I39 (gocomp_0[39:39], i_0r0[39:39], i_0r1[39:39]);
  OR2 I40 (gocomp_0[40:40], i_0r0[40:40], i_0r1[40:40]);
  OR2 I41 (gocomp_0[41:41], i_0r0[41:41], i_0r1[41:41]);
  OR2 I42 (gocomp_0[42:42], i_0r0[42:42], i_0r1[42:42]);
  OR2 I43 (gocomp_0[43:43], i_0r0[43:43], i_0r1[43:43]);
  OR2 I44 (gocomp_0[44:44], i_0r0[44:44], i_0r1[44:44]);
  OR2 I45 (gocomp_0[45:45], i_0r0[45:45], i_0r1[45:45]);
  OR2 I46 (gocomp_0[46:46], i_0r0[46:46], i_0r1[46:46]);
  OR2 I47 (gocomp_0[47:47], i_0r0[47:47], i_0r1[47:47]);
  OR2 I48 (gocomp_0[48:48], i_0r0[48:48], i_0r1[48:48]);
  OR2 I49 (gocomp_0[49:49], i_0r0[49:49], i_0r1[49:49]);
  OR2 I50 (gocomp_0[50:50], i_0r0[50:50], i_0r1[50:50]);
  OR2 I51 (gocomp_0[51:51], i_0r0[51:51], i_0r1[51:51]);
  OR2 I52 (gocomp_0[52:52], i_0r0[52:52], i_0r1[52:52]);
  OR2 I53 (gocomp_0[53:53], i_0r0[53:53], i_0r1[53:53]);
  OR2 I54 (gocomp_0[54:54], i_0r0[54:54], i_0r1[54:54]);
  OR2 I55 (gocomp_0[55:55], i_0r0[55:55], i_0r1[55:55]);
  OR2 I56 (gocomp_0[56:56], i_0r0[56:56], i_0r1[56:56]);
  OR2 I57 (gocomp_0[57:57], i_0r0[57:57], i_0r1[57:57]);
  OR2 I58 (gocomp_0[58:58], i_0r0[58:58], i_0r1[58:58]);
  OR2 I59 (gocomp_0[59:59], i_0r0[59:59], i_0r1[59:59]);
  OR2 I60 (gocomp_0[60:60], i_0r0[60:60], i_0r1[60:60]);
  OR2 I61 (gocomp_0[61:61], i_0r0[61:61], i_0r1[61:61]);
  OR2 I62 (gocomp_0[62:62], i_0r0[62:62], i_0r1[62:62]);
  OR2 I63 (gocomp_0[63:63], i_0r0[63:63], i_0r1[63:63]);
  C3 I64 (simp661_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  C3 I65 (simp661_0[1:1], gocomp_0[3:3], gocomp_0[4:4], gocomp_0[5:5]);
  C3 I66 (simp661_0[2:2], gocomp_0[6:6], gocomp_0[7:7], gocomp_0[8:8]);
  C3 I67 (simp661_0[3:3], gocomp_0[9:9], gocomp_0[10:10], gocomp_0[11:11]);
  C3 I68 (simp661_0[4:4], gocomp_0[12:12], gocomp_0[13:13], gocomp_0[14:14]);
  C3 I69 (simp661_0[5:5], gocomp_0[15:15], gocomp_0[16:16], gocomp_0[17:17]);
  C3 I70 (simp661_0[6:6], gocomp_0[18:18], gocomp_0[19:19], gocomp_0[20:20]);
  C3 I71 (simp661_0[7:7], gocomp_0[21:21], gocomp_0[22:22], gocomp_0[23:23]);
  C3 I72 (simp661_0[8:8], gocomp_0[24:24], gocomp_0[25:25], gocomp_0[26:26]);
  C3 I73 (simp661_0[9:9], gocomp_0[27:27], gocomp_0[28:28], gocomp_0[29:29]);
  C3 I74 (simp661_0[10:10], gocomp_0[30:30], gocomp_0[31:31], gocomp_0[32:32]);
  C3 I75 (simp661_0[11:11], gocomp_0[33:33], gocomp_0[34:34], gocomp_0[35:35]);
  C3 I76 (simp661_0[12:12], gocomp_0[36:36], gocomp_0[37:37], gocomp_0[38:38]);
  C3 I77 (simp661_0[13:13], gocomp_0[39:39], gocomp_0[40:40], gocomp_0[41:41]);
  C3 I78 (simp661_0[14:14], gocomp_0[42:42], gocomp_0[43:43], gocomp_0[44:44]);
  C3 I79 (simp661_0[15:15], gocomp_0[45:45], gocomp_0[46:46], gocomp_0[47:47]);
  C3 I80 (simp661_0[16:16], gocomp_0[48:48], gocomp_0[49:49], gocomp_0[50:50]);
  C3 I81 (simp661_0[17:17], gocomp_0[51:51], gocomp_0[52:52], gocomp_0[53:53]);
  C3 I82 (simp661_0[18:18], gocomp_0[54:54], gocomp_0[55:55], gocomp_0[56:56]);
  C3 I83 (simp661_0[19:19], gocomp_0[57:57], gocomp_0[58:58], gocomp_0[59:59]);
  C3 I84 (simp661_0[20:20], gocomp_0[60:60], gocomp_0[61:61], gocomp_0[62:62]);
  BUFF I85 (simp661_0[21:21], gocomp_0[63:63]);
  C3 I86 (simp662_0[0:0], simp661_0[0:0], simp661_0[1:1], simp661_0[2:2]);
  C3 I87 (simp662_0[1:1], simp661_0[3:3], simp661_0[4:4], simp661_0[5:5]);
  C3 I88 (simp662_0[2:2], simp661_0[6:6], simp661_0[7:7], simp661_0[8:8]);
  C3 I89 (simp662_0[3:3], simp661_0[9:9], simp661_0[10:10], simp661_0[11:11]);
  C3 I90 (simp662_0[4:4], simp661_0[12:12], simp661_0[13:13], simp661_0[14:14]);
  C3 I91 (simp662_0[5:5], simp661_0[15:15], simp661_0[16:16], simp661_0[17:17]);
  C3 I92 (simp662_0[6:6], simp661_0[18:18], simp661_0[19:19], simp661_0[20:20]);
  BUFF I93 (simp662_0[7:7], simp661_0[21:21]);
  C3 I94 (simp663_0[0:0], simp662_0[0:0], simp662_0[1:1], simp662_0[2:2]);
  C3 I95 (simp663_0[1:1], simp662_0[3:3], simp662_0[4:4], simp662_0[5:5]);
  C2 I96 (simp663_0[2:2], simp662_0[6:6], simp662_0[7:7]);
  C3 I97 (go_0, simp663_0[0:0], simp663_0[1:1], simp663_0[2:2]);
  BUFF I98 (termf_1[0:0], go_0);
  BUFF I99 (termf_1[1:1], go_0);
  GND I100 (termt_1[0:0]);
  GND I101 (termt_1[1:1]);
  BUFF I102 (termf_2[0:0], i_0r0[0:0]);
  BUFF I103 (termf_2[1:1], i_0r0[1:1]);
  BUFF I104 (termf_2[2:2], i_0r0[2:2]);
  BUFF I105 (termf_2[3:3], i_0r0[3:3]);
  BUFF I106 (termf_2[4:4], i_0r0[4:4]);
  BUFF I107 (termf_2[5:5], i_0r0[5:5]);
  BUFF I108 (termf_2[6:6], i_0r0[6:6]);
  BUFF I109 (termf_2[7:7], i_0r0[7:7]);
  BUFF I110 (termf_2[8:8], i_0r0[8:8]);
  BUFF I111 (termf_2[9:9], i_0r0[9:9]);
  BUFF I112 (termf_2[10:10], i_0r0[10:10]);
  BUFF I113 (termf_2[11:11], i_0r0[11:11]);
  BUFF I114 (termf_2[12:12], i_0r0[12:12]);
  BUFF I115 (termf_2[13:13], i_0r0[13:13]);
  BUFF I116 (termf_2[14:14], i_0r0[14:14]);
  BUFF I117 (termf_2[15:15], i_0r0[15:15]);
  BUFF I118 (termf_2[16:16], i_0r0[16:16]);
  BUFF I119 (termf_2[17:17], i_0r0[17:17]);
  BUFF I120 (termf_2[18:18], i_0r0[18:18]);
  BUFF I121 (termf_2[19:19], i_0r0[19:19]);
  BUFF I122 (termf_2[20:20], i_0r0[20:20]);
  BUFF I123 (termf_2[21:21], i_0r0[21:21]);
  BUFF I124 (termf_2[22:22], i_0r0[22:22]);
  BUFF I125 (termf_2[23:23], i_0r0[23:23]);
  BUFF I126 (termf_2[24:24], i_0r0[24:24]);
  BUFF I127 (termf_2[25:25], i_0r0[25:25]);
  BUFF I128 (termf_2[26:26], i_0r0[26:26]);
  BUFF I129 (termf_2[27:27], i_0r0[27:27]);
  BUFF I130 (termf_2[28:28], i_0r0[28:28]);
  BUFF I131 (termf_2[29:29], i_0r0[29:29]);
  BUFF I132 (termf_2[30:30], i_0r0[30:30]);
  BUFF I133 (termf_2[31:31], i_0r0[31:31]);
  BUFF I134 (termf_2[32:32], termf_1[0:0]);
  BUFF I135 (termf_2[33:33], termf_1[1:1]);
  BUFF I136 (termt_2[0:0], i_0r1[0:0]);
  BUFF I137 (termt_2[1:1], i_0r1[1:1]);
  BUFF I138 (termt_2[2:2], i_0r1[2:2]);
  BUFF I139 (termt_2[3:3], i_0r1[3:3]);
  BUFF I140 (termt_2[4:4], i_0r1[4:4]);
  BUFF I141 (termt_2[5:5], i_0r1[5:5]);
  BUFF I142 (termt_2[6:6], i_0r1[6:6]);
  BUFF I143 (termt_2[7:7], i_0r1[7:7]);
  BUFF I144 (termt_2[8:8], i_0r1[8:8]);
  BUFF I145 (termt_2[9:9], i_0r1[9:9]);
  BUFF I146 (termt_2[10:10], i_0r1[10:10]);
  BUFF I147 (termt_2[11:11], i_0r1[11:11]);
  BUFF I148 (termt_2[12:12], i_0r1[12:12]);
  BUFF I149 (termt_2[13:13], i_0r1[13:13]);
  BUFF I150 (termt_2[14:14], i_0r1[14:14]);
  BUFF I151 (termt_2[15:15], i_0r1[15:15]);
  BUFF I152 (termt_2[16:16], i_0r1[16:16]);
  BUFF I153 (termt_2[17:17], i_0r1[17:17]);
  BUFF I154 (termt_2[18:18], i_0r1[18:18]);
  BUFF I155 (termt_2[19:19], i_0r1[19:19]);
  BUFF I156 (termt_2[20:20], i_0r1[20:20]);
  BUFF I157 (termt_2[21:21], i_0r1[21:21]);
  BUFF I158 (termt_2[22:22], i_0r1[22:22]);
  BUFF I159 (termt_2[23:23], i_0r1[23:23]);
  BUFF I160 (termt_2[24:24], i_0r1[24:24]);
  BUFF I161 (termt_2[25:25], i_0r1[25:25]);
  BUFF I162 (termt_2[26:26], i_0r1[26:26]);
  BUFF I163 (termt_2[27:27], i_0r1[27:27]);
  BUFF I164 (termt_2[28:28], i_0r1[28:28]);
  BUFF I165 (termt_2[29:29], i_0r1[29:29]);
  BUFF I166 (termt_2[30:30], i_0r1[30:30]);
  BUFF I167 (termt_2[31:31], i_0r1[31:31]);
  BUFF I168 (termt_2[32:32], termt_1[0:0]);
  BUFF I169 (termt_2[33:33], termt_1[1:1]);
  BUFF I170 (termf_3[0:0], go_0);
  BUFF I171 (termf_3[1:1], go_0);
  GND I172 (termt_3[0:0]);
  GND I173 (termt_3[1:1]);
  BUFF I174 (termf_4[0:0], i_0r0[32:32]);
  BUFF I175 (termf_4[1:1], i_0r0[33:33]);
  BUFF I176 (termf_4[2:2], i_0r0[34:34]);
  BUFF I177 (termf_4[3:3], i_0r0[35:35]);
  BUFF I178 (termf_4[4:4], i_0r0[36:36]);
  BUFF I179 (termf_4[5:5], i_0r0[37:37]);
  BUFF I180 (termf_4[6:6], i_0r0[38:38]);
  BUFF I181 (termf_4[7:7], i_0r0[39:39]);
  BUFF I182 (termf_4[8:8], i_0r0[40:40]);
  BUFF I183 (termf_4[9:9], i_0r0[41:41]);
  BUFF I184 (termf_4[10:10], i_0r0[42:42]);
  BUFF I185 (termf_4[11:11], i_0r0[43:43]);
  BUFF I186 (termf_4[12:12], i_0r0[44:44]);
  BUFF I187 (termf_4[13:13], i_0r0[45:45]);
  BUFF I188 (termf_4[14:14], i_0r0[46:46]);
  BUFF I189 (termf_4[15:15], i_0r0[47:47]);
  BUFF I190 (termf_4[16:16], i_0r0[48:48]);
  BUFF I191 (termf_4[17:17], i_0r0[49:49]);
  BUFF I192 (termf_4[18:18], i_0r0[50:50]);
  BUFF I193 (termf_4[19:19], i_0r0[51:51]);
  BUFF I194 (termf_4[20:20], i_0r0[52:52]);
  BUFF I195 (termf_4[21:21], i_0r0[53:53]);
  BUFF I196 (termf_4[22:22], i_0r0[54:54]);
  BUFF I197 (termf_4[23:23], i_0r0[55:55]);
  BUFF I198 (termf_4[24:24], i_0r0[56:56]);
  BUFF I199 (termf_4[25:25], i_0r0[57:57]);
  BUFF I200 (termf_4[26:26], i_0r0[58:58]);
  BUFF I201 (termf_4[27:27], i_0r0[59:59]);
  BUFF I202 (termf_4[28:28], i_0r0[60:60]);
  BUFF I203 (termf_4[29:29], i_0r0[61:61]);
  BUFF I204 (termf_4[30:30], i_0r0[62:62]);
  BUFF I205 (termf_4[31:31], i_0r0[63:63]);
  BUFF I206 (termf_4[32:32], termf_3[0:0]);
  BUFF I207 (termf_4[33:33], termf_3[1:1]);
  BUFF I208 (termt_4[0:0], i_0r1[32:32]);
  BUFF I209 (termt_4[1:1], i_0r1[33:33]);
  BUFF I210 (termt_4[2:2], i_0r1[34:34]);
  BUFF I211 (termt_4[3:3], i_0r1[35:35]);
  BUFF I212 (termt_4[4:4], i_0r1[36:36]);
  BUFF I213 (termt_4[5:5], i_0r1[37:37]);
  BUFF I214 (termt_4[6:6], i_0r1[38:38]);
  BUFF I215 (termt_4[7:7], i_0r1[39:39]);
  BUFF I216 (termt_4[8:8], i_0r1[40:40]);
  BUFF I217 (termt_4[9:9], i_0r1[41:41]);
  BUFF I218 (termt_4[10:10], i_0r1[42:42]);
  BUFF I219 (termt_4[11:11], i_0r1[43:43]);
  BUFF I220 (termt_4[12:12], i_0r1[44:44]);
  BUFF I221 (termt_4[13:13], i_0r1[45:45]);
  BUFF I222 (termt_4[14:14], i_0r1[46:46]);
  BUFF I223 (termt_4[15:15], i_0r1[47:47]);
  BUFF I224 (termt_4[16:16], i_0r1[48:48]);
  BUFF I225 (termt_4[17:17], i_0r1[49:49]);
  BUFF I226 (termt_4[18:18], i_0r1[50:50]);
  BUFF I227 (termt_4[19:19], i_0r1[51:51]);
  BUFF I228 (termt_4[20:20], i_0r1[52:52]);
  BUFF I229 (termt_4[21:21], i_0r1[53:53]);
  BUFF I230 (termt_4[22:22], i_0r1[54:54]);
  BUFF I231 (termt_4[23:23], i_0r1[55:55]);
  BUFF I232 (termt_4[24:24], i_0r1[56:56]);
  BUFF I233 (termt_4[25:25], i_0r1[57:57]);
  BUFF I234 (termt_4[26:26], i_0r1[58:58]);
  BUFF I235 (termt_4[27:27], i_0r1[59:59]);
  BUFF I236 (termt_4[28:28], i_0r1[60:60]);
  BUFF I237 (termt_4[29:29], i_0r1[61:61]);
  BUFF I238 (termt_4[30:30], i_0r1[62:62]);
  BUFF I239 (termt_4[31:31], i_0r1[63:63]);
  BUFF I240 (termt_4[32:32], termt_3[0:0]);
  BUFF I241 (termt_4[33:33], termt_3[1:1]);
  C2 I242 (ha5__0[0:0], termt_4[0:0], termf_2[0:0]);
  C2 I243 (ha5__0[1:1], termt_4[0:0], termt_2[0:0]);
  C2 I244 (ha5__0[2:2], termf_4[0:0], termf_2[0:0]);
  C2 I245 (ha5__0[3:3], termf_4[0:0], termt_2[0:0]);
  BUFF I246 (cf5__0[0:0], ha5__0[0:0]);
  OR3 I247 (ct5__0[0:0], ha5__0[1:1], ha5__0[2:2], ha5__0[3:3]);
  OR2 I248 (termf_5[0:0], ha5__0[1:1], ha5__0[2:2]);
  OR2 I249 (termt_5[0:0], ha5__0[0:0], ha5__0[3:3]);
  C3 I250 (fa5_1min_0[0:0], cf5__0[0:0], termt_4[1:1], termf_2[1:1]);
  C3 I251 (fa5_1min_0[1:1], cf5__0[0:0], termt_4[1:1], termt_2[1:1]);
  C3 I252 (fa5_1min_0[2:2], cf5__0[0:0], termf_4[1:1], termf_2[1:1]);
  C3 I253 (fa5_1min_0[3:3], cf5__0[0:0], termf_4[1:1], termt_2[1:1]);
  C3 I254 (fa5_1min_0[4:4], ct5__0[0:0], termt_4[1:1], termf_2[1:1]);
  C3 I255 (fa5_1min_0[5:5], ct5__0[0:0], termt_4[1:1], termt_2[1:1]);
  C3 I256 (fa5_1min_0[6:6], ct5__0[0:0], termf_4[1:1], termf_2[1:1]);
  C3 I257 (fa5_1min_0[7:7], ct5__0[0:0], termf_4[1:1], termt_2[1:1]);
  NOR3 I258 (simp2391_0[0:0], fa5_1min_0[0:0], fa5_1min_0[3:3], fa5_1min_0[5:5]);
  INV I259 (simp2391_0[1:1], fa5_1min_0[6:6]);
  NAND2 I260 (termf_5[1:1], simp2391_0[0:0], simp2391_0[1:1]);
  NOR3 I261 (simp2401_0[0:0], fa5_1min_0[1:1], fa5_1min_0[2:2], fa5_1min_0[4:4]);
  INV I262 (simp2401_0[1:1], fa5_1min_0[7:7]);
  NAND2 I263 (termt_5[1:1], simp2401_0[0:0], simp2401_0[1:1]);
  AO222 I264 (ct5__0[1:1], termt_2[1:1], termf_4[1:1], termt_2[1:1], ct5__0[0:0], termf_4[1:1], ct5__0[0:0]);
  AO222 I265 (cf5__0[1:1], termf_2[1:1], termt_4[1:1], termf_2[1:1], cf5__0[0:0], termt_4[1:1], cf5__0[0:0]);
  C3 I266 (fa5_2min_0[0:0], cf5__0[1:1], termt_4[2:2], termf_2[2:2]);
  C3 I267 (fa5_2min_0[1:1], cf5__0[1:1], termt_4[2:2], termt_2[2:2]);
  C3 I268 (fa5_2min_0[2:2], cf5__0[1:1], termf_4[2:2], termf_2[2:2]);
  C3 I269 (fa5_2min_0[3:3], cf5__0[1:1], termf_4[2:2], termt_2[2:2]);
  C3 I270 (fa5_2min_0[4:4], ct5__0[1:1], termt_4[2:2], termf_2[2:2]);
  C3 I271 (fa5_2min_0[5:5], ct5__0[1:1], termt_4[2:2], termt_2[2:2]);
  C3 I272 (fa5_2min_0[6:6], ct5__0[1:1], termf_4[2:2], termf_2[2:2]);
  C3 I273 (fa5_2min_0[7:7], ct5__0[1:1], termf_4[2:2], termt_2[2:2]);
  NOR3 I274 (simp2521_0[0:0], fa5_2min_0[0:0], fa5_2min_0[3:3], fa5_2min_0[5:5]);
  INV I275 (simp2521_0[1:1], fa5_2min_0[6:6]);
  NAND2 I276 (termf_5[2:2], simp2521_0[0:0], simp2521_0[1:1]);
  NOR3 I277 (simp2531_0[0:0], fa5_2min_0[1:1], fa5_2min_0[2:2], fa5_2min_0[4:4]);
  INV I278 (simp2531_0[1:1], fa5_2min_0[7:7]);
  NAND2 I279 (termt_5[2:2], simp2531_0[0:0], simp2531_0[1:1]);
  AO222 I280 (ct5__0[2:2], termt_2[2:2], termf_4[2:2], termt_2[2:2], ct5__0[1:1], termf_4[2:2], ct5__0[1:1]);
  AO222 I281 (cf5__0[2:2], termf_2[2:2], termt_4[2:2], termf_2[2:2], cf5__0[1:1], termt_4[2:2], cf5__0[1:1]);
  C3 I282 (fa5_3min_0[0:0], cf5__0[2:2], termt_4[3:3], termf_2[3:3]);
  C3 I283 (fa5_3min_0[1:1], cf5__0[2:2], termt_4[3:3], termt_2[3:3]);
  C3 I284 (fa5_3min_0[2:2], cf5__0[2:2], termf_4[3:3], termf_2[3:3]);
  C3 I285 (fa5_3min_0[3:3], cf5__0[2:2], termf_4[3:3], termt_2[3:3]);
  C3 I286 (fa5_3min_0[4:4], ct5__0[2:2], termt_4[3:3], termf_2[3:3]);
  C3 I287 (fa5_3min_0[5:5], ct5__0[2:2], termt_4[3:3], termt_2[3:3]);
  C3 I288 (fa5_3min_0[6:6], ct5__0[2:2], termf_4[3:3], termf_2[3:3]);
  C3 I289 (fa5_3min_0[7:7], ct5__0[2:2], termf_4[3:3], termt_2[3:3]);
  NOR3 I290 (simp2651_0[0:0], fa5_3min_0[0:0], fa5_3min_0[3:3], fa5_3min_0[5:5]);
  INV I291 (simp2651_0[1:1], fa5_3min_0[6:6]);
  NAND2 I292 (termf_5[3:3], simp2651_0[0:0], simp2651_0[1:1]);
  NOR3 I293 (simp2661_0[0:0], fa5_3min_0[1:1], fa5_3min_0[2:2], fa5_3min_0[4:4]);
  INV I294 (simp2661_0[1:1], fa5_3min_0[7:7]);
  NAND2 I295 (termt_5[3:3], simp2661_0[0:0], simp2661_0[1:1]);
  AO222 I296 (ct5__0[3:3], termt_2[3:3], termf_4[3:3], termt_2[3:3], ct5__0[2:2], termf_4[3:3], ct5__0[2:2]);
  AO222 I297 (cf5__0[3:3], termf_2[3:3], termt_4[3:3], termf_2[3:3], cf5__0[2:2], termt_4[3:3], cf5__0[2:2]);
  C3 I298 (fa5_4min_0[0:0], cf5__0[3:3], termt_4[4:4], termf_2[4:4]);
  C3 I299 (fa5_4min_0[1:1], cf5__0[3:3], termt_4[4:4], termt_2[4:4]);
  C3 I300 (fa5_4min_0[2:2], cf5__0[3:3], termf_4[4:4], termf_2[4:4]);
  C3 I301 (fa5_4min_0[3:3], cf5__0[3:3], termf_4[4:4], termt_2[4:4]);
  C3 I302 (fa5_4min_0[4:4], ct5__0[3:3], termt_4[4:4], termf_2[4:4]);
  C3 I303 (fa5_4min_0[5:5], ct5__0[3:3], termt_4[4:4], termt_2[4:4]);
  C3 I304 (fa5_4min_0[6:6], ct5__0[3:3], termf_4[4:4], termf_2[4:4]);
  C3 I305 (fa5_4min_0[7:7], ct5__0[3:3], termf_4[4:4], termt_2[4:4]);
  NOR3 I306 (simp2781_0[0:0], fa5_4min_0[0:0], fa5_4min_0[3:3], fa5_4min_0[5:5]);
  INV I307 (simp2781_0[1:1], fa5_4min_0[6:6]);
  NAND2 I308 (termf_5[4:4], simp2781_0[0:0], simp2781_0[1:1]);
  NOR3 I309 (simp2791_0[0:0], fa5_4min_0[1:1], fa5_4min_0[2:2], fa5_4min_0[4:4]);
  INV I310 (simp2791_0[1:1], fa5_4min_0[7:7]);
  NAND2 I311 (termt_5[4:4], simp2791_0[0:0], simp2791_0[1:1]);
  AO222 I312 (ct5__0[4:4], termt_2[4:4], termf_4[4:4], termt_2[4:4], ct5__0[3:3], termf_4[4:4], ct5__0[3:3]);
  AO222 I313 (cf5__0[4:4], termf_2[4:4], termt_4[4:4], termf_2[4:4], cf5__0[3:3], termt_4[4:4], cf5__0[3:3]);
  C3 I314 (fa5_5min_0[0:0], cf5__0[4:4], termt_4[5:5], termf_2[5:5]);
  C3 I315 (fa5_5min_0[1:1], cf5__0[4:4], termt_4[5:5], termt_2[5:5]);
  C3 I316 (fa5_5min_0[2:2], cf5__0[4:4], termf_4[5:5], termf_2[5:5]);
  C3 I317 (fa5_5min_0[3:3], cf5__0[4:4], termf_4[5:5], termt_2[5:5]);
  C3 I318 (fa5_5min_0[4:4], ct5__0[4:4], termt_4[5:5], termf_2[5:5]);
  C3 I319 (fa5_5min_0[5:5], ct5__0[4:4], termt_4[5:5], termt_2[5:5]);
  C3 I320 (fa5_5min_0[6:6], ct5__0[4:4], termf_4[5:5], termf_2[5:5]);
  C3 I321 (fa5_5min_0[7:7], ct5__0[4:4], termf_4[5:5], termt_2[5:5]);
  NOR3 I322 (simp2911_0[0:0], fa5_5min_0[0:0], fa5_5min_0[3:3], fa5_5min_0[5:5]);
  INV I323 (simp2911_0[1:1], fa5_5min_0[6:6]);
  NAND2 I324 (termf_5[5:5], simp2911_0[0:0], simp2911_0[1:1]);
  NOR3 I325 (simp2921_0[0:0], fa5_5min_0[1:1], fa5_5min_0[2:2], fa5_5min_0[4:4]);
  INV I326 (simp2921_0[1:1], fa5_5min_0[7:7]);
  NAND2 I327 (termt_5[5:5], simp2921_0[0:0], simp2921_0[1:1]);
  AO222 I328 (ct5__0[5:5], termt_2[5:5], termf_4[5:5], termt_2[5:5], ct5__0[4:4], termf_4[5:5], ct5__0[4:4]);
  AO222 I329 (cf5__0[5:5], termf_2[5:5], termt_4[5:5], termf_2[5:5], cf5__0[4:4], termt_4[5:5], cf5__0[4:4]);
  C3 I330 (fa5_6min_0[0:0], cf5__0[5:5], termt_4[6:6], termf_2[6:6]);
  C3 I331 (fa5_6min_0[1:1], cf5__0[5:5], termt_4[6:6], termt_2[6:6]);
  C3 I332 (fa5_6min_0[2:2], cf5__0[5:5], termf_4[6:6], termf_2[6:6]);
  C3 I333 (fa5_6min_0[3:3], cf5__0[5:5], termf_4[6:6], termt_2[6:6]);
  C3 I334 (fa5_6min_0[4:4], ct5__0[5:5], termt_4[6:6], termf_2[6:6]);
  C3 I335 (fa5_6min_0[5:5], ct5__0[5:5], termt_4[6:6], termt_2[6:6]);
  C3 I336 (fa5_6min_0[6:6], ct5__0[5:5], termf_4[6:6], termf_2[6:6]);
  C3 I337 (fa5_6min_0[7:7], ct5__0[5:5], termf_4[6:6], termt_2[6:6]);
  NOR3 I338 (simp3041_0[0:0], fa5_6min_0[0:0], fa5_6min_0[3:3], fa5_6min_0[5:5]);
  INV I339 (simp3041_0[1:1], fa5_6min_0[6:6]);
  NAND2 I340 (termf_5[6:6], simp3041_0[0:0], simp3041_0[1:1]);
  NOR3 I341 (simp3051_0[0:0], fa5_6min_0[1:1], fa5_6min_0[2:2], fa5_6min_0[4:4]);
  INV I342 (simp3051_0[1:1], fa5_6min_0[7:7]);
  NAND2 I343 (termt_5[6:6], simp3051_0[0:0], simp3051_0[1:1]);
  AO222 I344 (ct5__0[6:6], termt_2[6:6], termf_4[6:6], termt_2[6:6], ct5__0[5:5], termf_4[6:6], ct5__0[5:5]);
  AO222 I345 (cf5__0[6:6], termf_2[6:6], termt_4[6:6], termf_2[6:6], cf5__0[5:5], termt_4[6:6], cf5__0[5:5]);
  C3 I346 (fa5_7min_0[0:0], cf5__0[6:6], termt_4[7:7], termf_2[7:7]);
  C3 I347 (fa5_7min_0[1:1], cf5__0[6:6], termt_4[7:7], termt_2[7:7]);
  C3 I348 (fa5_7min_0[2:2], cf5__0[6:6], termf_4[7:7], termf_2[7:7]);
  C3 I349 (fa5_7min_0[3:3], cf5__0[6:6], termf_4[7:7], termt_2[7:7]);
  C3 I350 (fa5_7min_0[4:4], ct5__0[6:6], termt_4[7:7], termf_2[7:7]);
  C3 I351 (fa5_7min_0[5:5], ct5__0[6:6], termt_4[7:7], termt_2[7:7]);
  C3 I352 (fa5_7min_0[6:6], ct5__0[6:6], termf_4[7:7], termf_2[7:7]);
  C3 I353 (fa5_7min_0[7:7], ct5__0[6:6], termf_4[7:7], termt_2[7:7]);
  NOR3 I354 (simp3171_0[0:0], fa5_7min_0[0:0], fa5_7min_0[3:3], fa5_7min_0[5:5]);
  INV I355 (simp3171_0[1:1], fa5_7min_0[6:6]);
  NAND2 I356 (termf_5[7:7], simp3171_0[0:0], simp3171_0[1:1]);
  NOR3 I357 (simp3181_0[0:0], fa5_7min_0[1:1], fa5_7min_0[2:2], fa5_7min_0[4:4]);
  INV I358 (simp3181_0[1:1], fa5_7min_0[7:7]);
  NAND2 I359 (termt_5[7:7], simp3181_0[0:0], simp3181_0[1:1]);
  AO222 I360 (ct5__0[7:7], termt_2[7:7], termf_4[7:7], termt_2[7:7], ct5__0[6:6], termf_4[7:7], ct5__0[6:6]);
  AO222 I361 (cf5__0[7:7], termf_2[7:7], termt_4[7:7], termf_2[7:7], cf5__0[6:6], termt_4[7:7], cf5__0[6:6]);
  C3 I362 (fa5_8min_0[0:0], cf5__0[7:7], termt_4[8:8], termf_2[8:8]);
  C3 I363 (fa5_8min_0[1:1], cf5__0[7:7], termt_4[8:8], termt_2[8:8]);
  C3 I364 (fa5_8min_0[2:2], cf5__0[7:7], termf_4[8:8], termf_2[8:8]);
  C3 I365 (fa5_8min_0[3:3], cf5__0[7:7], termf_4[8:8], termt_2[8:8]);
  C3 I366 (fa5_8min_0[4:4], ct5__0[7:7], termt_4[8:8], termf_2[8:8]);
  C3 I367 (fa5_8min_0[5:5], ct5__0[7:7], termt_4[8:8], termt_2[8:8]);
  C3 I368 (fa5_8min_0[6:6], ct5__0[7:7], termf_4[8:8], termf_2[8:8]);
  C3 I369 (fa5_8min_0[7:7], ct5__0[7:7], termf_4[8:8], termt_2[8:8]);
  NOR3 I370 (simp3301_0[0:0], fa5_8min_0[0:0], fa5_8min_0[3:3], fa5_8min_0[5:5]);
  INV I371 (simp3301_0[1:1], fa5_8min_0[6:6]);
  NAND2 I372 (termf_5[8:8], simp3301_0[0:0], simp3301_0[1:1]);
  NOR3 I373 (simp3311_0[0:0], fa5_8min_0[1:1], fa5_8min_0[2:2], fa5_8min_0[4:4]);
  INV I374 (simp3311_0[1:1], fa5_8min_0[7:7]);
  NAND2 I375 (termt_5[8:8], simp3311_0[0:0], simp3311_0[1:1]);
  AO222 I376 (ct5__0[8:8], termt_2[8:8], termf_4[8:8], termt_2[8:8], ct5__0[7:7], termf_4[8:8], ct5__0[7:7]);
  AO222 I377 (cf5__0[8:8], termf_2[8:8], termt_4[8:8], termf_2[8:8], cf5__0[7:7], termt_4[8:8], cf5__0[7:7]);
  C3 I378 (fa5_9min_0[0:0], cf5__0[8:8], termt_4[9:9], termf_2[9:9]);
  C3 I379 (fa5_9min_0[1:1], cf5__0[8:8], termt_4[9:9], termt_2[9:9]);
  C3 I380 (fa5_9min_0[2:2], cf5__0[8:8], termf_4[9:9], termf_2[9:9]);
  C3 I381 (fa5_9min_0[3:3], cf5__0[8:8], termf_4[9:9], termt_2[9:9]);
  C3 I382 (fa5_9min_0[4:4], ct5__0[8:8], termt_4[9:9], termf_2[9:9]);
  C3 I383 (fa5_9min_0[5:5], ct5__0[8:8], termt_4[9:9], termt_2[9:9]);
  C3 I384 (fa5_9min_0[6:6], ct5__0[8:8], termf_4[9:9], termf_2[9:9]);
  C3 I385 (fa5_9min_0[7:7], ct5__0[8:8], termf_4[9:9], termt_2[9:9]);
  NOR3 I386 (simp3431_0[0:0], fa5_9min_0[0:0], fa5_9min_0[3:3], fa5_9min_0[5:5]);
  INV I387 (simp3431_0[1:1], fa5_9min_0[6:6]);
  NAND2 I388 (termf_5[9:9], simp3431_0[0:0], simp3431_0[1:1]);
  NOR3 I389 (simp3441_0[0:0], fa5_9min_0[1:1], fa5_9min_0[2:2], fa5_9min_0[4:4]);
  INV I390 (simp3441_0[1:1], fa5_9min_0[7:7]);
  NAND2 I391 (termt_5[9:9], simp3441_0[0:0], simp3441_0[1:1]);
  AO222 I392 (ct5__0[9:9], termt_2[9:9], termf_4[9:9], termt_2[9:9], ct5__0[8:8], termf_4[9:9], ct5__0[8:8]);
  AO222 I393 (cf5__0[9:9], termf_2[9:9], termt_4[9:9], termf_2[9:9], cf5__0[8:8], termt_4[9:9], cf5__0[8:8]);
  C3 I394 (fa5_10min_0[0:0], cf5__0[9:9], termt_4[10:10], termf_2[10:10]);
  C3 I395 (fa5_10min_0[1:1], cf5__0[9:9], termt_4[10:10], termt_2[10:10]);
  C3 I396 (fa5_10min_0[2:2], cf5__0[9:9], termf_4[10:10], termf_2[10:10]);
  C3 I397 (fa5_10min_0[3:3], cf5__0[9:9], termf_4[10:10], termt_2[10:10]);
  C3 I398 (fa5_10min_0[4:4], ct5__0[9:9], termt_4[10:10], termf_2[10:10]);
  C3 I399 (fa5_10min_0[5:5], ct5__0[9:9], termt_4[10:10], termt_2[10:10]);
  C3 I400 (fa5_10min_0[6:6], ct5__0[9:9], termf_4[10:10], termf_2[10:10]);
  C3 I401 (fa5_10min_0[7:7], ct5__0[9:9], termf_4[10:10], termt_2[10:10]);
  NOR3 I402 (simp3561_0[0:0], fa5_10min_0[0:0], fa5_10min_0[3:3], fa5_10min_0[5:5]);
  INV I403 (simp3561_0[1:1], fa5_10min_0[6:6]);
  NAND2 I404 (termf_5[10:10], simp3561_0[0:0], simp3561_0[1:1]);
  NOR3 I405 (simp3571_0[0:0], fa5_10min_0[1:1], fa5_10min_0[2:2], fa5_10min_0[4:4]);
  INV I406 (simp3571_0[1:1], fa5_10min_0[7:7]);
  NAND2 I407 (termt_5[10:10], simp3571_0[0:0], simp3571_0[1:1]);
  AO222 I408 (ct5__0[10:10], termt_2[10:10], termf_4[10:10], termt_2[10:10], ct5__0[9:9], termf_4[10:10], ct5__0[9:9]);
  AO222 I409 (cf5__0[10:10], termf_2[10:10], termt_4[10:10], termf_2[10:10], cf5__0[9:9], termt_4[10:10], cf5__0[9:9]);
  C3 I410 (fa5_11min_0[0:0], cf5__0[10:10], termt_4[11:11], termf_2[11:11]);
  C3 I411 (fa5_11min_0[1:1], cf5__0[10:10], termt_4[11:11], termt_2[11:11]);
  C3 I412 (fa5_11min_0[2:2], cf5__0[10:10], termf_4[11:11], termf_2[11:11]);
  C3 I413 (fa5_11min_0[3:3], cf5__0[10:10], termf_4[11:11], termt_2[11:11]);
  C3 I414 (fa5_11min_0[4:4], ct5__0[10:10], termt_4[11:11], termf_2[11:11]);
  C3 I415 (fa5_11min_0[5:5], ct5__0[10:10], termt_4[11:11], termt_2[11:11]);
  C3 I416 (fa5_11min_0[6:6], ct5__0[10:10], termf_4[11:11], termf_2[11:11]);
  C3 I417 (fa5_11min_0[7:7], ct5__0[10:10], termf_4[11:11], termt_2[11:11]);
  NOR3 I418 (simp3691_0[0:0], fa5_11min_0[0:0], fa5_11min_0[3:3], fa5_11min_0[5:5]);
  INV I419 (simp3691_0[1:1], fa5_11min_0[6:6]);
  NAND2 I420 (termf_5[11:11], simp3691_0[0:0], simp3691_0[1:1]);
  NOR3 I421 (simp3701_0[0:0], fa5_11min_0[1:1], fa5_11min_0[2:2], fa5_11min_0[4:4]);
  INV I422 (simp3701_0[1:1], fa5_11min_0[7:7]);
  NAND2 I423 (termt_5[11:11], simp3701_0[0:0], simp3701_0[1:1]);
  AO222 I424 (ct5__0[11:11], termt_2[11:11], termf_4[11:11], termt_2[11:11], ct5__0[10:10], termf_4[11:11], ct5__0[10:10]);
  AO222 I425 (cf5__0[11:11], termf_2[11:11], termt_4[11:11], termf_2[11:11], cf5__0[10:10], termt_4[11:11], cf5__0[10:10]);
  C3 I426 (fa5_12min_0[0:0], cf5__0[11:11], termt_4[12:12], termf_2[12:12]);
  C3 I427 (fa5_12min_0[1:1], cf5__0[11:11], termt_4[12:12], termt_2[12:12]);
  C3 I428 (fa5_12min_0[2:2], cf5__0[11:11], termf_4[12:12], termf_2[12:12]);
  C3 I429 (fa5_12min_0[3:3], cf5__0[11:11], termf_4[12:12], termt_2[12:12]);
  C3 I430 (fa5_12min_0[4:4], ct5__0[11:11], termt_4[12:12], termf_2[12:12]);
  C3 I431 (fa5_12min_0[5:5], ct5__0[11:11], termt_4[12:12], termt_2[12:12]);
  C3 I432 (fa5_12min_0[6:6], ct5__0[11:11], termf_4[12:12], termf_2[12:12]);
  C3 I433 (fa5_12min_0[7:7], ct5__0[11:11], termf_4[12:12], termt_2[12:12]);
  NOR3 I434 (simp3821_0[0:0], fa5_12min_0[0:0], fa5_12min_0[3:3], fa5_12min_0[5:5]);
  INV I435 (simp3821_0[1:1], fa5_12min_0[6:6]);
  NAND2 I436 (termf_5[12:12], simp3821_0[0:0], simp3821_0[1:1]);
  NOR3 I437 (simp3831_0[0:0], fa5_12min_0[1:1], fa5_12min_0[2:2], fa5_12min_0[4:4]);
  INV I438 (simp3831_0[1:1], fa5_12min_0[7:7]);
  NAND2 I439 (termt_5[12:12], simp3831_0[0:0], simp3831_0[1:1]);
  AO222 I440 (ct5__0[12:12], termt_2[12:12], termf_4[12:12], termt_2[12:12], ct5__0[11:11], termf_4[12:12], ct5__0[11:11]);
  AO222 I441 (cf5__0[12:12], termf_2[12:12], termt_4[12:12], termf_2[12:12], cf5__0[11:11], termt_4[12:12], cf5__0[11:11]);
  C3 I442 (fa5_13min_0[0:0], cf5__0[12:12], termt_4[13:13], termf_2[13:13]);
  C3 I443 (fa5_13min_0[1:1], cf5__0[12:12], termt_4[13:13], termt_2[13:13]);
  C3 I444 (fa5_13min_0[2:2], cf5__0[12:12], termf_4[13:13], termf_2[13:13]);
  C3 I445 (fa5_13min_0[3:3], cf5__0[12:12], termf_4[13:13], termt_2[13:13]);
  C3 I446 (fa5_13min_0[4:4], ct5__0[12:12], termt_4[13:13], termf_2[13:13]);
  C3 I447 (fa5_13min_0[5:5], ct5__0[12:12], termt_4[13:13], termt_2[13:13]);
  C3 I448 (fa5_13min_0[6:6], ct5__0[12:12], termf_4[13:13], termf_2[13:13]);
  C3 I449 (fa5_13min_0[7:7], ct5__0[12:12], termf_4[13:13], termt_2[13:13]);
  NOR3 I450 (simp3951_0[0:0], fa5_13min_0[0:0], fa5_13min_0[3:3], fa5_13min_0[5:5]);
  INV I451 (simp3951_0[1:1], fa5_13min_0[6:6]);
  NAND2 I452 (termf_5[13:13], simp3951_0[0:0], simp3951_0[1:1]);
  NOR3 I453 (simp3961_0[0:0], fa5_13min_0[1:1], fa5_13min_0[2:2], fa5_13min_0[4:4]);
  INV I454 (simp3961_0[1:1], fa5_13min_0[7:7]);
  NAND2 I455 (termt_5[13:13], simp3961_0[0:0], simp3961_0[1:1]);
  AO222 I456 (ct5__0[13:13], termt_2[13:13], termf_4[13:13], termt_2[13:13], ct5__0[12:12], termf_4[13:13], ct5__0[12:12]);
  AO222 I457 (cf5__0[13:13], termf_2[13:13], termt_4[13:13], termf_2[13:13], cf5__0[12:12], termt_4[13:13], cf5__0[12:12]);
  C3 I458 (fa5_14min_0[0:0], cf5__0[13:13], termt_4[14:14], termf_2[14:14]);
  C3 I459 (fa5_14min_0[1:1], cf5__0[13:13], termt_4[14:14], termt_2[14:14]);
  C3 I460 (fa5_14min_0[2:2], cf5__0[13:13], termf_4[14:14], termf_2[14:14]);
  C3 I461 (fa5_14min_0[3:3], cf5__0[13:13], termf_4[14:14], termt_2[14:14]);
  C3 I462 (fa5_14min_0[4:4], ct5__0[13:13], termt_4[14:14], termf_2[14:14]);
  C3 I463 (fa5_14min_0[5:5], ct5__0[13:13], termt_4[14:14], termt_2[14:14]);
  C3 I464 (fa5_14min_0[6:6], ct5__0[13:13], termf_4[14:14], termf_2[14:14]);
  C3 I465 (fa5_14min_0[7:7], ct5__0[13:13], termf_4[14:14], termt_2[14:14]);
  NOR3 I466 (simp4081_0[0:0], fa5_14min_0[0:0], fa5_14min_0[3:3], fa5_14min_0[5:5]);
  INV I467 (simp4081_0[1:1], fa5_14min_0[6:6]);
  NAND2 I468 (termf_5[14:14], simp4081_0[0:0], simp4081_0[1:1]);
  NOR3 I469 (simp4091_0[0:0], fa5_14min_0[1:1], fa5_14min_0[2:2], fa5_14min_0[4:4]);
  INV I470 (simp4091_0[1:1], fa5_14min_0[7:7]);
  NAND2 I471 (termt_5[14:14], simp4091_0[0:0], simp4091_0[1:1]);
  AO222 I472 (ct5__0[14:14], termt_2[14:14], termf_4[14:14], termt_2[14:14], ct5__0[13:13], termf_4[14:14], ct5__0[13:13]);
  AO222 I473 (cf5__0[14:14], termf_2[14:14], termt_4[14:14], termf_2[14:14], cf5__0[13:13], termt_4[14:14], cf5__0[13:13]);
  C3 I474 (fa5_15min_0[0:0], cf5__0[14:14], termt_4[15:15], termf_2[15:15]);
  C3 I475 (fa5_15min_0[1:1], cf5__0[14:14], termt_4[15:15], termt_2[15:15]);
  C3 I476 (fa5_15min_0[2:2], cf5__0[14:14], termf_4[15:15], termf_2[15:15]);
  C3 I477 (fa5_15min_0[3:3], cf5__0[14:14], termf_4[15:15], termt_2[15:15]);
  C3 I478 (fa5_15min_0[4:4], ct5__0[14:14], termt_4[15:15], termf_2[15:15]);
  C3 I479 (fa5_15min_0[5:5], ct5__0[14:14], termt_4[15:15], termt_2[15:15]);
  C3 I480 (fa5_15min_0[6:6], ct5__0[14:14], termf_4[15:15], termf_2[15:15]);
  C3 I481 (fa5_15min_0[7:7], ct5__0[14:14], termf_4[15:15], termt_2[15:15]);
  NOR3 I482 (simp4211_0[0:0], fa5_15min_0[0:0], fa5_15min_0[3:3], fa5_15min_0[5:5]);
  INV I483 (simp4211_0[1:1], fa5_15min_0[6:6]);
  NAND2 I484 (termf_5[15:15], simp4211_0[0:0], simp4211_0[1:1]);
  NOR3 I485 (simp4221_0[0:0], fa5_15min_0[1:1], fa5_15min_0[2:2], fa5_15min_0[4:4]);
  INV I486 (simp4221_0[1:1], fa5_15min_0[7:7]);
  NAND2 I487 (termt_5[15:15], simp4221_0[0:0], simp4221_0[1:1]);
  AO222 I488 (ct5__0[15:15], termt_2[15:15], termf_4[15:15], termt_2[15:15], ct5__0[14:14], termf_4[15:15], ct5__0[14:14]);
  AO222 I489 (cf5__0[15:15], termf_2[15:15], termt_4[15:15], termf_2[15:15], cf5__0[14:14], termt_4[15:15], cf5__0[14:14]);
  C3 I490 (fa5_16min_0[0:0], cf5__0[15:15], termt_4[16:16], termf_2[16:16]);
  C3 I491 (fa5_16min_0[1:1], cf5__0[15:15], termt_4[16:16], termt_2[16:16]);
  C3 I492 (fa5_16min_0[2:2], cf5__0[15:15], termf_4[16:16], termf_2[16:16]);
  C3 I493 (fa5_16min_0[3:3], cf5__0[15:15], termf_4[16:16], termt_2[16:16]);
  C3 I494 (fa5_16min_0[4:4], ct5__0[15:15], termt_4[16:16], termf_2[16:16]);
  C3 I495 (fa5_16min_0[5:5], ct5__0[15:15], termt_4[16:16], termt_2[16:16]);
  C3 I496 (fa5_16min_0[6:6], ct5__0[15:15], termf_4[16:16], termf_2[16:16]);
  C3 I497 (fa5_16min_0[7:7], ct5__0[15:15], termf_4[16:16], termt_2[16:16]);
  NOR3 I498 (simp4341_0[0:0], fa5_16min_0[0:0], fa5_16min_0[3:3], fa5_16min_0[5:5]);
  INV I499 (simp4341_0[1:1], fa5_16min_0[6:6]);
  NAND2 I500 (termf_5[16:16], simp4341_0[0:0], simp4341_0[1:1]);
  NOR3 I501 (simp4351_0[0:0], fa5_16min_0[1:1], fa5_16min_0[2:2], fa5_16min_0[4:4]);
  INV I502 (simp4351_0[1:1], fa5_16min_0[7:7]);
  NAND2 I503 (termt_5[16:16], simp4351_0[0:0], simp4351_0[1:1]);
  AO222 I504 (ct5__0[16:16], termt_2[16:16], termf_4[16:16], termt_2[16:16], ct5__0[15:15], termf_4[16:16], ct5__0[15:15]);
  AO222 I505 (cf5__0[16:16], termf_2[16:16], termt_4[16:16], termf_2[16:16], cf5__0[15:15], termt_4[16:16], cf5__0[15:15]);
  C3 I506 (fa5_17min_0[0:0], cf5__0[16:16], termt_4[17:17], termf_2[17:17]);
  C3 I507 (fa5_17min_0[1:1], cf5__0[16:16], termt_4[17:17], termt_2[17:17]);
  C3 I508 (fa5_17min_0[2:2], cf5__0[16:16], termf_4[17:17], termf_2[17:17]);
  C3 I509 (fa5_17min_0[3:3], cf5__0[16:16], termf_4[17:17], termt_2[17:17]);
  C3 I510 (fa5_17min_0[4:4], ct5__0[16:16], termt_4[17:17], termf_2[17:17]);
  C3 I511 (fa5_17min_0[5:5], ct5__0[16:16], termt_4[17:17], termt_2[17:17]);
  C3 I512 (fa5_17min_0[6:6], ct5__0[16:16], termf_4[17:17], termf_2[17:17]);
  C3 I513 (fa5_17min_0[7:7], ct5__0[16:16], termf_4[17:17], termt_2[17:17]);
  NOR3 I514 (simp4471_0[0:0], fa5_17min_0[0:0], fa5_17min_0[3:3], fa5_17min_0[5:5]);
  INV I515 (simp4471_0[1:1], fa5_17min_0[6:6]);
  NAND2 I516 (termf_5[17:17], simp4471_0[0:0], simp4471_0[1:1]);
  NOR3 I517 (simp4481_0[0:0], fa5_17min_0[1:1], fa5_17min_0[2:2], fa5_17min_0[4:4]);
  INV I518 (simp4481_0[1:1], fa5_17min_0[7:7]);
  NAND2 I519 (termt_5[17:17], simp4481_0[0:0], simp4481_0[1:1]);
  AO222 I520 (ct5__0[17:17], termt_2[17:17], termf_4[17:17], termt_2[17:17], ct5__0[16:16], termf_4[17:17], ct5__0[16:16]);
  AO222 I521 (cf5__0[17:17], termf_2[17:17], termt_4[17:17], termf_2[17:17], cf5__0[16:16], termt_4[17:17], cf5__0[16:16]);
  C3 I522 (fa5_18min_0[0:0], cf5__0[17:17], termt_4[18:18], termf_2[18:18]);
  C3 I523 (fa5_18min_0[1:1], cf5__0[17:17], termt_4[18:18], termt_2[18:18]);
  C3 I524 (fa5_18min_0[2:2], cf5__0[17:17], termf_4[18:18], termf_2[18:18]);
  C3 I525 (fa5_18min_0[3:3], cf5__0[17:17], termf_4[18:18], termt_2[18:18]);
  C3 I526 (fa5_18min_0[4:4], ct5__0[17:17], termt_4[18:18], termf_2[18:18]);
  C3 I527 (fa5_18min_0[5:5], ct5__0[17:17], termt_4[18:18], termt_2[18:18]);
  C3 I528 (fa5_18min_0[6:6], ct5__0[17:17], termf_4[18:18], termf_2[18:18]);
  C3 I529 (fa5_18min_0[7:7], ct5__0[17:17], termf_4[18:18], termt_2[18:18]);
  NOR3 I530 (simp4601_0[0:0], fa5_18min_0[0:0], fa5_18min_0[3:3], fa5_18min_0[5:5]);
  INV I531 (simp4601_0[1:1], fa5_18min_0[6:6]);
  NAND2 I532 (termf_5[18:18], simp4601_0[0:0], simp4601_0[1:1]);
  NOR3 I533 (simp4611_0[0:0], fa5_18min_0[1:1], fa5_18min_0[2:2], fa5_18min_0[4:4]);
  INV I534 (simp4611_0[1:1], fa5_18min_0[7:7]);
  NAND2 I535 (termt_5[18:18], simp4611_0[0:0], simp4611_0[1:1]);
  AO222 I536 (ct5__0[18:18], termt_2[18:18], termf_4[18:18], termt_2[18:18], ct5__0[17:17], termf_4[18:18], ct5__0[17:17]);
  AO222 I537 (cf5__0[18:18], termf_2[18:18], termt_4[18:18], termf_2[18:18], cf5__0[17:17], termt_4[18:18], cf5__0[17:17]);
  C3 I538 (fa5_19min_0[0:0], cf5__0[18:18], termt_4[19:19], termf_2[19:19]);
  C3 I539 (fa5_19min_0[1:1], cf5__0[18:18], termt_4[19:19], termt_2[19:19]);
  C3 I540 (fa5_19min_0[2:2], cf5__0[18:18], termf_4[19:19], termf_2[19:19]);
  C3 I541 (fa5_19min_0[3:3], cf5__0[18:18], termf_4[19:19], termt_2[19:19]);
  C3 I542 (fa5_19min_0[4:4], ct5__0[18:18], termt_4[19:19], termf_2[19:19]);
  C3 I543 (fa5_19min_0[5:5], ct5__0[18:18], termt_4[19:19], termt_2[19:19]);
  C3 I544 (fa5_19min_0[6:6], ct5__0[18:18], termf_4[19:19], termf_2[19:19]);
  C3 I545 (fa5_19min_0[7:7], ct5__0[18:18], termf_4[19:19], termt_2[19:19]);
  NOR3 I546 (simp4731_0[0:0], fa5_19min_0[0:0], fa5_19min_0[3:3], fa5_19min_0[5:5]);
  INV I547 (simp4731_0[1:1], fa5_19min_0[6:6]);
  NAND2 I548 (termf_5[19:19], simp4731_0[0:0], simp4731_0[1:1]);
  NOR3 I549 (simp4741_0[0:0], fa5_19min_0[1:1], fa5_19min_0[2:2], fa5_19min_0[4:4]);
  INV I550 (simp4741_0[1:1], fa5_19min_0[7:7]);
  NAND2 I551 (termt_5[19:19], simp4741_0[0:0], simp4741_0[1:1]);
  AO222 I552 (ct5__0[19:19], termt_2[19:19], termf_4[19:19], termt_2[19:19], ct5__0[18:18], termf_4[19:19], ct5__0[18:18]);
  AO222 I553 (cf5__0[19:19], termf_2[19:19], termt_4[19:19], termf_2[19:19], cf5__0[18:18], termt_4[19:19], cf5__0[18:18]);
  C3 I554 (fa5_20min_0[0:0], cf5__0[19:19], termt_4[20:20], termf_2[20:20]);
  C3 I555 (fa5_20min_0[1:1], cf5__0[19:19], termt_4[20:20], termt_2[20:20]);
  C3 I556 (fa5_20min_0[2:2], cf5__0[19:19], termf_4[20:20], termf_2[20:20]);
  C3 I557 (fa5_20min_0[3:3], cf5__0[19:19], termf_4[20:20], termt_2[20:20]);
  C3 I558 (fa5_20min_0[4:4], ct5__0[19:19], termt_4[20:20], termf_2[20:20]);
  C3 I559 (fa5_20min_0[5:5], ct5__0[19:19], termt_4[20:20], termt_2[20:20]);
  C3 I560 (fa5_20min_0[6:6], ct5__0[19:19], termf_4[20:20], termf_2[20:20]);
  C3 I561 (fa5_20min_0[7:7], ct5__0[19:19], termf_4[20:20], termt_2[20:20]);
  NOR3 I562 (simp4861_0[0:0], fa5_20min_0[0:0], fa5_20min_0[3:3], fa5_20min_0[5:5]);
  INV I563 (simp4861_0[1:1], fa5_20min_0[6:6]);
  NAND2 I564 (termf_5[20:20], simp4861_0[0:0], simp4861_0[1:1]);
  NOR3 I565 (simp4871_0[0:0], fa5_20min_0[1:1], fa5_20min_0[2:2], fa5_20min_0[4:4]);
  INV I566 (simp4871_0[1:1], fa5_20min_0[7:7]);
  NAND2 I567 (termt_5[20:20], simp4871_0[0:0], simp4871_0[1:1]);
  AO222 I568 (ct5__0[20:20], termt_2[20:20], termf_4[20:20], termt_2[20:20], ct5__0[19:19], termf_4[20:20], ct5__0[19:19]);
  AO222 I569 (cf5__0[20:20], termf_2[20:20], termt_4[20:20], termf_2[20:20], cf5__0[19:19], termt_4[20:20], cf5__0[19:19]);
  C3 I570 (fa5_21min_0[0:0], cf5__0[20:20], termt_4[21:21], termf_2[21:21]);
  C3 I571 (fa5_21min_0[1:1], cf5__0[20:20], termt_4[21:21], termt_2[21:21]);
  C3 I572 (fa5_21min_0[2:2], cf5__0[20:20], termf_4[21:21], termf_2[21:21]);
  C3 I573 (fa5_21min_0[3:3], cf5__0[20:20], termf_4[21:21], termt_2[21:21]);
  C3 I574 (fa5_21min_0[4:4], ct5__0[20:20], termt_4[21:21], termf_2[21:21]);
  C3 I575 (fa5_21min_0[5:5], ct5__0[20:20], termt_4[21:21], termt_2[21:21]);
  C3 I576 (fa5_21min_0[6:6], ct5__0[20:20], termf_4[21:21], termf_2[21:21]);
  C3 I577 (fa5_21min_0[7:7], ct5__0[20:20], termf_4[21:21], termt_2[21:21]);
  NOR3 I578 (simp4991_0[0:0], fa5_21min_0[0:0], fa5_21min_0[3:3], fa5_21min_0[5:5]);
  INV I579 (simp4991_0[1:1], fa5_21min_0[6:6]);
  NAND2 I580 (termf_5[21:21], simp4991_0[0:0], simp4991_0[1:1]);
  NOR3 I581 (simp5001_0[0:0], fa5_21min_0[1:1], fa5_21min_0[2:2], fa5_21min_0[4:4]);
  INV I582 (simp5001_0[1:1], fa5_21min_0[7:7]);
  NAND2 I583 (termt_5[21:21], simp5001_0[0:0], simp5001_0[1:1]);
  AO222 I584 (ct5__0[21:21], termt_2[21:21], termf_4[21:21], termt_2[21:21], ct5__0[20:20], termf_4[21:21], ct5__0[20:20]);
  AO222 I585 (cf5__0[21:21], termf_2[21:21], termt_4[21:21], termf_2[21:21], cf5__0[20:20], termt_4[21:21], cf5__0[20:20]);
  C3 I586 (fa5_22min_0[0:0], cf5__0[21:21], termt_4[22:22], termf_2[22:22]);
  C3 I587 (fa5_22min_0[1:1], cf5__0[21:21], termt_4[22:22], termt_2[22:22]);
  C3 I588 (fa5_22min_0[2:2], cf5__0[21:21], termf_4[22:22], termf_2[22:22]);
  C3 I589 (fa5_22min_0[3:3], cf5__0[21:21], termf_4[22:22], termt_2[22:22]);
  C3 I590 (fa5_22min_0[4:4], ct5__0[21:21], termt_4[22:22], termf_2[22:22]);
  C3 I591 (fa5_22min_0[5:5], ct5__0[21:21], termt_4[22:22], termt_2[22:22]);
  C3 I592 (fa5_22min_0[6:6], ct5__0[21:21], termf_4[22:22], termf_2[22:22]);
  C3 I593 (fa5_22min_0[7:7], ct5__0[21:21], termf_4[22:22], termt_2[22:22]);
  NOR3 I594 (simp5121_0[0:0], fa5_22min_0[0:0], fa5_22min_0[3:3], fa5_22min_0[5:5]);
  INV I595 (simp5121_0[1:1], fa5_22min_0[6:6]);
  NAND2 I596 (termf_5[22:22], simp5121_0[0:0], simp5121_0[1:1]);
  NOR3 I597 (simp5131_0[0:0], fa5_22min_0[1:1], fa5_22min_0[2:2], fa5_22min_0[4:4]);
  INV I598 (simp5131_0[1:1], fa5_22min_0[7:7]);
  NAND2 I599 (termt_5[22:22], simp5131_0[0:0], simp5131_0[1:1]);
  AO222 I600 (ct5__0[22:22], termt_2[22:22], termf_4[22:22], termt_2[22:22], ct5__0[21:21], termf_4[22:22], ct5__0[21:21]);
  AO222 I601 (cf5__0[22:22], termf_2[22:22], termt_4[22:22], termf_2[22:22], cf5__0[21:21], termt_4[22:22], cf5__0[21:21]);
  C3 I602 (fa5_23min_0[0:0], cf5__0[22:22], termt_4[23:23], termf_2[23:23]);
  C3 I603 (fa5_23min_0[1:1], cf5__0[22:22], termt_4[23:23], termt_2[23:23]);
  C3 I604 (fa5_23min_0[2:2], cf5__0[22:22], termf_4[23:23], termf_2[23:23]);
  C3 I605 (fa5_23min_0[3:3], cf5__0[22:22], termf_4[23:23], termt_2[23:23]);
  C3 I606 (fa5_23min_0[4:4], ct5__0[22:22], termt_4[23:23], termf_2[23:23]);
  C3 I607 (fa5_23min_0[5:5], ct5__0[22:22], termt_4[23:23], termt_2[23:23]);
  C3 I608 (fa5_23min_0[6:6], ct5__0[22:22], termf_4[23:23], termf_2[23:23]);
  C3 I609 (fa5_23min_0[7:7], ct5__0[22:22], termf_4[23:23], termt_2[23:23]);
  NOR3 I610 (simp5251_0[0:0], fa5_23min_0[0:0], fa5_23min_0[3:3], fa5_23min_0[5:5]);
  INV I611 (simp5251_0[1:1], fa5_23min_0[6:6]);
  NAND2 I612 (termf_5[23:23], simp5251_0[0:0], simp5251_0[1:1]);
  NOR3 I613 (simp5261_0[0:0], fa5_23min_0[1:1], fa5_23min_0[2:2], fa5_23min_0[4:4]);
  INV I614 (simp5261_0[1:1], fa5_23min_0[7:7]);
  NAND2 I615 (termt_5[23:23], simp5261_0[0:0], simp5261_0[1:1]);
  AO222 I616 (ct5__0[23:23], termt_2[23:23], termf_4[23:23], termt_2[23:23], ct5__0[22:22], termf_4[23:23], ct5__0[22:22]);
  AO222 I617 (cf5__0[23:23], termf_2[23:23], termt_4[23:23], termf_2[23:23], cf5__0[22:22], termt_4[23:23], cf5__0[22:22]);
  C3 I618 (fa5_24min_0[0:0], cf5__0[23:23], termt_4[24:24], termf_2[24:24]);
  C3 I619 (fa5_24min_0[1:1], cf5__0[23:23], termt_4[24:24], termt_2[24:24]);
  C3 I620 (fa5_24min_0[2:2], cf5__0[23:23], termf_4[24:24], termf_2[24:24]);
  C3 I621 (fa5_24min_0[3:3], cf5__0[23:23], termf_4[24:24], termt_2[24:24]);
  C3 I622 (fa5_24min_0[4:4], ct5__0[23:23], termt_4[24:24], termf_2[24:24]);
  C3 I623 (fa5_24min_0[5:5], ct5__0[23:23], termt_4[24:24], termt_2[24:24]);
  C3 I624 (fa5_24min_0[6:6], ct5__0[23:23], termf_4[24:24], termf_2[24:24]);
  C3 I625 (fa5_24min_0[7:7], ct5__0[23:23], termf_4[24:24], termt_2[24:24]);
  NOR3 I626 (simp5381_0[0:0], fa5_24min_0[0:0], fa5_24min_0[3:3], fa5_24min_0[5:5]);
  INV I627 (simp5381_0[1:1], fa5_24min_0[6:6]);
  NAND2 I628 (termf_5[24:24], simp5381_0[0:0], simp5381_0[1:1]);
  NOR3 I629 (simp5391_0[0:0], fa5_24min_0[1:1], fa5_24min_0[2:2], fa5_24min_0[4:4]);
  INV I630 (simp5391_0[1:1], fa5_24min_0[7:7]);
  NAND2 I631 (termt_5[24:24], simp5391_0[0:0], simp5391_0[1:1]);
  AO222 I632 (ct5__0[24:24], termt_2[24:24], termf_4[24:24], termt_2[24:24], ct5__0[23:23], termf_4[24:24], ct5__0[23:23]);
  AO222 I633 (cf5__0[24:24], termf_2[24:24], termt_4[24:24], termf_2[24:24], cf5__0[23:23], termt_4[24:24], cf5__0[23:23]);
  C3 I634 (fa5_25min_0[0:0], cf5__0[24:24], termt_4[25:25], termf_2[25:25]);
  C3 I635 (fa5_25min_0[1:1], cf5__0[24:24], termt_4[25:25], termt_2[25:25]);
  C3 I636 (fa5_25min_0[2:2], cf5__0[24:24], termf_4[25:25], termf_2[25:25]);
  C3 I637 (fa5_25min_0[3:3], cf5__0[24:24], termf_4[25:25], termt_2[25:25]);
  C3 I638 (fa5_25min_0[4:4], ct5__0[24:24], termt_4[25:25], termf_2[25:25]);
  C3 I639 (fa5_25min_0[5:5], ct5__0[24:24], termt_4[25:25], termt_2[25:25]);
  C3 I640 (fa5_25min_0[6:6], ct5__0[24:24], termf_4[25:25], termf_2[25:25]);
  C3 I641 (fa5_25min_0[7:7], ct5__0[24:24], termf_4[25:25], termt_2[25:25]);
  NOR3 I642 (simp5511_0[0:0], fa5_25min_0[0:0], fa5_25min_0[3:3], fa5_25min_0[5:5]);
  INV I643 (simp5511_0[1:1], fa5_25min_0[6:6]);
  NAND2 I644 (termf_5[25:25], simp5511_0[0:0], simp5511_0[1:1]);
  NOR3 I645 (simp5521_0[0:0], fa5_25min_0[1:1], fa5_25min_0[2:2], fa5_25min_0[4:4]);
  INV I646 (simp5521_0[1:1], fa5_25min_0[7:7]);
  NAND2 I647 (termt_5[25:25], simp5521_0[0:0], simp5521_0[1:1]);
  AO222 I648 (ct5__0[25:25], termt_2[25:25], termf_4[25:25], termt_2[25:25], ct5__0[24:24], termf_4[25:25], ct5__0[24:24]);
  AO222 I649 (cf5__0[25:25], termf_2[25:25], termt_4[25:25], termf_2[25:25], cf5__0[24:24], termt_4[25:25], cf5__0[24:24]);
  C3 I650 (fa5_26min_0[0:0], cf5__0[25:25], termt_4[26:26], termf_2[26:26]);
  C3 I651 (fa5_26min_0[1:1], cf5__0[25:25], termt_4[26:26], termt_2[26:26]);
  C3 I652 (fa5_26min_0[2:2], cf5__0[25:25], termf_4[26:26], termf_2[26:26]);
  C3 I653 (fa5_26min_0[3:3], cf5__0[25:25], termf_4[26:26], termt_2[26:26]);
  C3 I654 (fa5_26min_0[4:4], ct5__0[25:25], termt_4[26:26], termf_2[26:26]);
  C3 I655 (fa5_26min_0[5:5], ct5__0[25:25], termt_4[26:26], termt_2[26:26]);
  C3 I656 (fa5_26min_0[6:6], ct5__0[25:25], termf_4[26:26], termf_2[26:26]);
  C3 I657 (fa5_26min_0[7:7], ct5__0[25:25], termf_4[26:26], termt_2[26:26]);
  NOR3 I658 (simp5641_0[0:0], fa5_26min_0[0:0], fa5_26min_0[3:3], fa5_26min_0[5:5]);
  INV I659 (simp5641_0[1:1], fa5_26min_0[6:6]);
  NAND2 I660 (termf_5[26:26], simp5641_0[0:0], simp5641_0[1:1]);
  NOR3 I661 (simp5651_0[0:0], fa5_26min_0[1:1], fa5_26min_0[2:2], fa5_26min_0[4:4]);
  INV I662 (simp5651_0[1:1], fa5_26min_0[7:7]);
  NAND2 I663 (termt_5[26:26], simp5651_0[0:0], simp5651_0[1:1]);
  AO222 I664 (ct5__0[26:26], termt_2[26:26], termf_4[26:26], termt_2[26:26], ct5__0[25:25], termf_4[26:26], ct5__0[25:25]);
  AO222 I665 (cf5__0[26:26], termf_2[26:26], termt_4[26:26], termf_2[26:26], cf5__0[25:25], termt_4[26:26], cf5__0[25:25]);
  C3 I666 (fa5_27min_0[0:0], cf5__0[26:26], termt_4[27:27], termf_2[27:27]);
  C3 I667 (fa5_27min_0[1:1], cf5__0[26:26], termt_4[27:27], termt_2[27:27]);
  C3 I668 (fa5_27min_0[2:2], cf5__0[26:26], termf_4[27:27], termf_2[27:27]);
  C3 I669 (fa5_27min_0[3:3], cf5__0[26:26], termf_4[27:27], termt_2[27:27]);
  C3 I670 (fa5_27min_0[4:4], ct5__0[26:26], termt_4[27:27], termf_2[27:27]);
  C3 I671 (fa5_27min_0[5:5], ct5__0[26:26], termt_4[27:27], termt_2[27:27]);
  C3 I672 (fa5_27min_0[6:6], ct5__0[26:26], termf_4[27:27], termf_2[27:27]);
  C3 I673 (fa5_27min_0[7:7], ct5__0[26:26], termf_4[27:27], termt_2[27:27]);
  NOR3 I674 (simp5771_0[0:0], fa5_27min_0[0:0], fa5_27min_0[3:3], fa5_27min_0[5:5]);
  INV I675 (simp5771_0[1:1], fa5_27min_0[6:6]);
  NAND2 I676 (termf_5[27:27], simp5771_0[0:0], simp5771_0[1:1]);
  NOR3 I677 (simp5781_0[0:0], fa5_27min_0[1:1], fa5_27min_0[2:2], fa5_27min_0[4:4]);
  INV I678 (simp5781_0[1:1], fa5_27min_0[7:7]);
  NAND2 I679 (termt_5[27:27], simp5781_0[0:0], simp5781_0[1:1]);
  AO222 I680 (ct5__0[27:27], termt_2[27:27], termf_4[27:27], termt_2[27:27], ct5__0[26:26], termf_4[27:27], ct5__0[26:26]);
  AO222 I681 (cf5__0[27:27], termf_2[27:27], termt_4[27:27], termf_2[27:27], cf5__0[26:26], termt_4[27:27], cf5__0[26:26]);
  C3 I682 (fa5_28min_0[0:0], cf5__0[27:27], termt_4[28:28], termf_2[28:28]);
  C3 I683 (fa5_28min_0[1:1], cf5__0[27:27], termt_4[28:28], termt_2[28:28]);
  C3 I684 (fa5_28min_0[2:2], cf5__0[27:27], termf_4[28:28], termf_2[28:28]);
  C3 I685 (fa5_28min_0[3:3], cf5__0[27:27], termf_4[28:28], termt_2[28:28]);
  C3 I686 (fa5_28min_0[4:4], ct5__0[27:27], termt_4[28:28], termf_2[28:28]);
  C3 I687 (fa5_28min_0[5:5], ct5__0[27:27], termt_4[28:28], termt_2[28:28]);
  C3 I688 (fa5_28min_0[6:6], ct5__0[27:27], termf_4[28:28], termf_2[28:28]);
  C3 I689 (fa5_28min_0[7:7], ct5__0[27:27], termf_4[28:28], termt_2[28:28]);
  NOR3 I690 (simp5901_0[0:0], fa5_28min_0[0:0], fa5_28min_0[3:3], fa5_28min_0[5:5]);
  INV I691 (simp5901_0[1:1], fa5_28min_0[6:6]);
  NAND2 I692 (termf_5[28:28], simp5901_0[0:0], simp5901_0[1:1]);
  NOR3 I693 (simp5911_0[0:0], fa5_28min_0[1:1], fa5_28min_0[2:2], fa5_28min_0[4:4]);
  INV I694 (simp5911_0[1:1], fa5_28min_0[7:7]);
  NAND2 I695 (termt_5[28:28], simp5911_0[0:0], simp5911_0[1:1]);
  AO222 I696 (ct5__0[28:28], termt_2[28:28], termf_4[28:28], termt_2[28:28], ct5__0[27:27], termf_4[28:28], ct5__0[27:27]);
  AO222 I697 (cf5__0[28:28], termf_2[28:28], termt_4[28:28], termf_2[28:28], cf5__0[27:27], termt_4[28:28], cf5__0[27:27]);
  C3 I698 (fa5_29min_0[0:0], cf5__0[28:28], termt_4[29:29], termf_2[29:29]);
  C3 I699 (fa5_29min_0[1:1], cf5__0[28:28], termt_4[29:29], termt_2[29:29]);
  C3 I700 (fa5_29min_0[2:2], cf5__0[28:28], termf_4[29:29], termf_2[29:29]);
  C3 I701 (fa5_29min_0[3:3], cf5__0[28:28], termf_4[29:29], termt_2[29:29]);
  C3 I702 (fa5_29min_0[4:4], ct5__0[28:28], termt_4[29:29], termf_2[29:29]);
  C3 I703 (fa5_29min_0[5:5], ct5__0[28:28], termt_4[29:29], termt_2[29:29]);
  C3 I704 (fa5_29min_0[6:6], ct5__0[28:28], termf_4[29:29], termf_2[29:29]);
  C3 I705 (fa5_29min_0[7:7], ct5__0[28:28], termf_4[29:29], termt_2[29:29]);
  NOR3 I706 (simp6031_0[0:0], fa5_29min_0[0:0], fa5_29min_0[3:3], fa5_29min_0[5:5]);
  INV I707 (simp6031_0[1:1], fa5_29min_0[6:6]);
  NAND2 I708 (termf_5[29:29], simp6031_0[0:0], simp6031_0[1:1]);
  NOR3 I709 (simp6041_0[0:0], fa5_29min_0[1:1], fa5_29min_0[2:2], fa5_29min_0[4:4]);
  INV I710 (simp6041_0[1:1], fa5_29min_0[7:7]);
  NAND2 I711 (termt_5[29:29], simp6041_0[0:0], simp6041_0[1:1]);
  AO222 I712 (ct5__0[29:29], termt_2[29:29], termf_4[29:29], termt_2[29:29], ct5__0[28:28], termf_4[29:29], ct5__0[28:28]);
  AO222 I713 (cf5__0[29:29], termf_2[29:29], termt_4[29:29], termf_2[29:29], cf5__0[28:28], termt_4[29:29], cf5__0[28:28]);
  C3 I714 (fa5_30min_0[0:0], cf5__0[29:29], termt_4[30:30], termf_2[30:30]);
  C3 I715 (fa5_30min_0[1:1], cf5__0[29:29], termt_4[30:30], termt_2[30:30]);
  C3 I716 (fa5_30min_0[2:2], cf5__0[29:29], termf_4[30:30], termf_2[30:30]);
  C3 I717 (fa5_30min_0[3:3], cf5__0[29:29], termf_4[30:30], termt_2[30:30]);
  C3 I718 (fa5_30min_0[4:4], ct5__0[29:29], termt_4[30:30], termf_2[30:30]);
  C3 I719 (fa5_30min_0[5:5], ct5__0[29:29], termt_4[30:30], termt_2[30:30]);
  C3 I720 (fa5_30min_0[6:6], ct5__0[29:29], termf_4[30:30], termf_2[30:30]);
  C3 I721 (fa5_30min_0[7:7], ct5__0[29:29], termf_4[30:30], termt_2[30:30]);
  NOR3 I722 (simp6161_0[0:0], fa5_30min_0[0:0], fa5_30min_0[3:3], fa5_30min_0[5:5]);
  INV I723 (simp6161_0[1:1], fa5_30min_0[6:6]);
  NAND2 I724 (termf_5[30:30], simp6161_0[0:0], simp6161_0[1:1]);
  NOR3 I725 (simp6171_0[0:0], fa5_30min_0[1:1], fa5_30min_0[2:2], fa5_30min_0[4:4]);
  INV I726 (simp6171_0[1:1], fa5_30min_0[7:7]);
  NAND2 I727 (termt_5[30:30], simp6171_0[0:0], simp6171_0[1:1]);
  AO222 I728 (ct5__0[30:30], termt_2[30:30], termf_4[30:30], termt_2[30:30], ct5__0[29:29], termf_4[30:30], ct5__0[29:29]);
  AO222 I729 (cf5__0[30:30], termf_2[30:30], termt_4[30:30], termf_2[30:30], cf5__0[29:29], termt_4[30:30], cf5__0[29:29]);
  C3 I730 (fa5_31min_0[0:0], cf5__0[30:30], termt_4[31:31], termf_2[31:31]);
  C3 I731 (fa5_31min_0[1:1], cf5__0[30:30], termt_4[31:31], termt_2[31:31]);
  C3 I732 (fa5_31min_0[2:2], cf5__0[30:30], termf_4[31:31], termf_2[31:31]);
  C3 I733 (fa5_31min_0[3:3], cf5__0[30:30], termf_4[31:31], termt_2[31:31]);
  C3 I734 (fa5_31min_0[4:4], ct5__0[30:30], termt_4[31:31], termf_2[31:31]);
  C3 I735 (fa5_31min_0[5:5], ct5__0[30:30], termt_4[31:31], termt_2[31:31]);
  C3 I736 (fa5_31min_0[6:6], ct5__0[30:30], termf_4[31:31], termf_2[31:31]);
  C3 I737 (fa5_31min_0[7:7], ct5__0[30:30], termf_4[31:31], termt_2[31:31]);
  NOR3 I738 (simp6291_0[0:0], fa5_31min_0[0:0], fa5_31min_0[3:3], fa5_31min_0[5:5]);
  INV I739 (simp6291_0[1:1], fa5_31min_0[6:6]);
  NAND2 I740 (termf_5[31:31], simp6291_0[0:0], simp6291_0[1:1]);
  NOR3 I741 (simp6301_0[0:0], fa5_31min_0[1:1], fa5_31min_0[2:2], fa5_31min_0[4:4]);
  INV I742 (simp6301_0[1:1], fa5_31min_0[7:7]);
  NAND2 I743 (termt_5[31:31], simp6301_0[0:0], simp6301_0[1:1]);
  AO222 I744 (ct5__0[31:31], termt_2[31:31], termf_4[31:31], termt_2[31:31], ct5__0[30:30], termf_4[31:31], ct5__0[30:30]);
  AO222 I745 (cf5__0[31:31], termf_2[31:31], termt_4[31:31], termf_2[31:31], cf5__0[30:30], termt_4[31:31], cf5__0[30:30]);
  C3 I746 (fa5_32min_0[0:0], cf5__0[31:31], termt_4[32:32], termf_2[32:32]);
  C3 I747 (fa5_32min_0[1:1], cf5__0[31:31], termt_4[32:32], termt_2[32:32]);
  C3 I748 (fa5_32min_0[2:2], cf5__0[31:31], termf_4[32:32], termf_2[32:32]);
  C3 I749 (fa5_32min_0[3:3], cf5__0[31:31], termf_4[32:32], termt_2[32:32]);
  C3 I750 (fa5_32min_0[4:4], ct5__0[31:31], termt_4[32:32], termf_2[32:32]);
  C3 I751 (fa5_32min_0[5:5], ct5__0[31:31], termt_4[32:32], termt_2[32:32]);
  C3 I752 (fa5_32min_0[6:6], ct5__0[31:31], termf_4[32:32], termf_2[32:32]);
  C3 I753 (fa5_32min_0[7:7], ct5__0[31:31], termf_4[32:32], termt_2[32:32]);
  NOR3 I754 (simp6421_0[0:0], fa5_32min_0[0:0], fa5_32min_0[3:3], fa5_32min_0[5:5]);
  INV I755 (simp6421_0[1:1], fa5_32min_0[6:6]);
  NAND2 I756 (termf_5[32:32], simp6421_0[0:0], simp6421_0[1:1]);
  NOR3 I757 (simp6431_0[0:0], fa5_32min_0[1:1], fa5_32min_0[2:2], fa5_32min_0[4:4]);
  INV I758 (simp6431_0[1:1], fa5_32min_0[7:7]);
  NAND2 I759 (termt_5[32:32], simp6431_0[0:0], simp6431_0[1:1]);
  AO222 I760 (ct5__0[32:32], termt_2[32:32], termf_4[32:32], termt_2[32:32], ct5__0[31:31], termf_4[32:32], ct5__0[31:31]);
  AO222 I761 (cf5__0[32:32], termf_2[32:32], termt_4[32:32], termf_2[32:32], cf5__0[31:31], termt_4[32:32], cf5__0[31:31]);
  C3 I762 (fa5_33min_0[0:0], cf5__0[32:32], termt_4[33:33], termf_2[33:33]);
  C3 I763 (fa5_33min_0[1:1], cf5__0[32:32], termt_4[33:33], termt_2[33:33]);
  C3 I764 (fa5_33min_0[2:2], cf5__0[32:32], termf_4[33:33], termf_2[33:33]);
  C3 I765 (fa5_33min_0[3:3], cf5__0[32:32], termf_4[33:33], termt_2[33:33]);
  C3 I766 (fa5_33min_0[4:4], ct5__0[32:32], termt_4[33:33], termf_2[33:33]);
  C3 I767 (fa5_33min_0[5:5], ct5__0[32:32], termt_4[33:33], termt_2[33:33]);
  C3 I768 (fa5_33min_0[6:6], ct5__0[32:32], termf_4[33:33], termf_2[33:33]);
  C3 I769 (fa5_33min_0[7:7], ct5__0[32:32], termf_4[33:33], termt_2[33:33]);
  NOR3 I770 (simp6551_0[0:0], fa5_33min_0[0:0], fa5_33min_0[3:3], fa5_33min_0[5:5]);
  INV I771 (simp6551_0[1:1], fa5_33min_0[6:6]);
  NAND2 I772 (termf_5[33:33], simp6551_0[0:0], simp6551_0[1:1]);
  NOR3 I773 (simp6561_0[0:0], fa5_33min_0[1:1], fa5_33min_0[2:2], fa5_33min_0[4:4]);
  INV I774 (simp6561_0[1:1], fa5_33min_0[7:7]);
  NAND2 I775 (termt_5[33:33], simp6561_0[0:0], simp6561_0[1:1]);
  AO222 I776 (ct5__0[33:33], termt_2[33:33], termf_4[33:33], termt_2[33:33], ct5__0[32:32], termf_4[33:33], ct5__0[32:32]);
  AO222 I777 (cf5__0[33:33], termf_2[33:33], termt_4[33:33], termf_2[33:33], cf5__0[32:32], termt_4[33:33], cf5__0[32:32]);
  BUFF I778 (o_0r0[0:0], termf_5[0:0]);
  BUFF I779 (o_0r0[1:1], termf_5[1:1]);
  BUFF I780 (o_0r0[2:2], termf_5[2:2]);
  BUFF I781 (o_0r0[3:3], termf_5[3:3]);
  BUFF I782 (o_0r0[4:4], termf_5[4:4]);
  BUFF I783 (o_0r0[5:5], termf_5[5:5]);
  BUFF I784 (o_0r0[6:6], termf_5[6:6]);
  BUFF I785 (o_0r0[7:7], termf_5[7:7]);
  BUFF I786 (o_0r0[8:8], termf_5[8:8]);
  BUFF I787 (o_0r0[9:9], termf_5[9:9]);
  BUFF I788 (o_0r0[10:10], termf_5[10:10]);
  BUFF I789 (o_0r0[11:11], termf_5[11:11]);
  BUFF I790 (o_0r0[12:12], termf_5[12:12]);
  BUFF I791 (o_0r0[13:13], termf_5[13:13]);
  BUFF I792 (o_0r0[14:14], termf_5[14:14]);
  BUFF I793 (o_0r0[15:15], termf_5[15:15]);
  BUFF I794 (o_0r0[16:16], termf_5[16:16]);
  BUFF I795 (o_0r0[17:17], termf_5[17:17]);
  BUFF I796 (o_0r0[18:18], termf_5[18:18]);
  BUFF I797 (o_0r0[19:19], termf_5[19:19]);
  BUFF I798 (o_0r0[20:20], termf_5[20:20]);
  BUFF I799 (o_0r0[21:21], termf_5[21:21]);
  BUFF I800 (o_0r0[22:22], termf_5[22:22]);
  BUFF I801 (o_0r0[23:23], termf_5[23:23]);
  BUFF I802 (o_0r0[24:24], termf_5[24:24]);
  BUFF I803 (o_0r0[25:25], termf_5[25:25]);
  BUFF I804 (o_0r0[26:26], termf_5[26:26]);
  BUFF I805 (o_0r0[27:27], termf_5[27:27]);
  BUFF I806 (o_0r0[28:28], termf_5[28:28]);
  BUFF I807 (o_0r0[29:29], termf_5[29:29]);
  BUFF I808 (o_0r0[30:30], termf_5[30:30]);
  BUFF I809 (o_0r0[31:31], termf_5[31:31]);
  BUFF I810 (o_0r1[0:0], termt_5[0:0]);
  BUFF I811 (o_0r1[1:1], termt_5[1:1]);
  BUFF I812 (o_0r1[2:2], termt_5[2:2]);
  BUFF I813 (o_0r1[3:3], termt_5[3:3]);
  BUFF I814 (o_0r1[4:4], termt_5[4:4]);
  BUFF I815 (o_0r1[5:5], termt_5[5:5]);
  BUFF I816 (o_0r1[6:6], termt_5[6:6]);
  BUFF I817 (o_0r1[7:7], termt_5[7:7]);
  BUFF I818 (o_0r1[8:8], termt_5[8:8]);
  BUFF I819 (o_0r1[9:9], termt_5[9:9]);
  BUFF I820 (o_0r1[10:10], termt_5[10:10]);
  BUFF I821 (o_0r1[11:11], termt_5[11:11]);
  BUFF I822 (o_0r1[12:12], termt_5[12:12]);
  BUFF I823 (o_0r1[13:13], termt_5[13:13]);
  BUFF I824 (o_0r1[14:14], termt_5[14:14]);
  BUFF I825 (o_0r1[15:15], termt_5[15:15]);
  BUFF I826 (o_0r1[16:16], termt_5[16:16]);
  BUFF I827 (o_0r1[17:17], termt_5[17:17]);
  BUFF I828 (o_0r1[18:18], termt_5[18:18]);
  BUFF I829 (o_0r1[19:19], termt_5[19:19]);
  BUFF I830 (o_0r1[20:20], termt_5[20:20]);
  BUFF I831 (o_0r1[21:21], termt_5[21:21]);
  BUFF I832 (o_0r1[22:22], termt_5[22:22]);
  BUFF I833 (o_0r1[23:23], termt_5[23:23]);
  BUFF I834 (o_0r1[24:24], termt_5[24:24]);
  BUFF I835 (o_0r1[25:25], termt_5[25:25]);
  BUFF I836 (o_0r1[26:26], termt_5[26:26]);
  BUFF I837 (o_0r1[27:27], termt_5[27:27]);
  BUFF I838 (o_0r1[28:28], termt_5[28:28]);
  BUFF I839 (o_0r1[29:29], termt_5[29:29]);
  BUFF I840 (o_0r1[30:30], termt_5[30:30]);
  BUFF I841 (o_0r1[31:31], termt_5[31:31]);
  BUFF I842 (i_0a, o_0a);
endmodule

// tko3m3_1nm3b1_2nm3b2_3mx0_1_i0w3bt1o0w3bt2o0w3b TeakO [
//     (1,TeakOConstant 3 1),
//     (2,TeakOConstant 3 2),
//     (3,TeakOMux [[Imp 0 0],[Imp 1 0]] [(0,0+:3),(1,0+:3),(2,0+:3)])] [One 3,One 3]
module tko3m3_1nm3b1_2nm3b2_3mx0_1_i0w3bt1o0w3bt2o0w3b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [2:0] gocomp_0;
  wire [2:0] termf_1;
  wire [2:0] termf_2;
  wire [2:0] termt_1;
  wire [2:0] termt_2;
  wire [2:0] gfint3_0;
  wire [2:0] gfint3_1;
  wire [2:0] gtint3_0;
  wire [2:0] gtint3_1;
  wire selcomp3_0;
  wire selcomp3_1;
  wire sel3_0;
  wire sel3_1;
  wire selg3_0;
  wire selg3_1;
  wire icomplete3_0;
  wire scomplete3_0;
  wire [2:0] comp30_0;
  wire [2:0] comp31_0;
  wire [2:0] dcomp3_0;
  wire match30_0;
  wire match31_0;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I3 (go_0, gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  BUFF I4 (termt_1[0:0], go_0);
  GND I5 (termf_1[0:0]);
  BUFF I6 (termf_1[1:1], go_0);
  BUFF I7 (termf_1[2:2], go_0);
  GND I8 (termt_1[1:1]);
  GND I9 (termt_1[2:2]);
  BUFF I10 (termt_2[1:1], go_0);
  GND I11 (termf_2[1:1]);
  BUFF I12 (termf_2[0:0], go_0);
  BUFF I13 (termf_2[2:2], go_0);
  GND I14 (termt_2[0:0]);
  GND I15 (termt_2[2:2]);
  OR2 I16 (comp30_0[0:0], termf_1[0:0], termt_1[0:0]);
  OR2 I17 (comp30_0[1:1], termf_1[1:1], termt_1[1:1]);
  OR2 I18 (comp30_0[2:2], termf_1[2:2], termt_1[2:2]);
  C3 I19 (selcomp3_0, comp30_0[0:0], comp30_0[1:1], comp30_0[2:2]);
  OR2 I20 (comp31_0[0:0], termf_2[0:0], termt_2[0:0]);
  OR2 I21 (comp31_0[1:1], termf_2[1:1], termt_2[1:1]);
  OR2 I22 (comp31_0[2:2], termf_2[2:2], termt_2[2:2]);
  C3 I23 (selcomp3_1, comp31_0[0:0], comp31_0[1:1], comp31_0[2:2]);
  OR2 I24 (dcomp3_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I25 (dcomp3_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I26 (dcomp3_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I27 (scomplete3_0, dcomp3_0[0:0], dcomp3_0[1:1], dcomp3_0[2:2]);
  C3 I28 (icomplete3_0, scomplete3_0, selcomp3_0, selcomp3_1);
  OR2 I29 (o_0r0[0:0], gfint3_0[0:0], gfint3_1[0:0]);
  OR2 I30 (o_0r0[1:1], gfint3_0[1:1], gfint3_1[1:1]);
  OR2 I31 (o_0r0[2:2], gfint3_0[2:2], gfint3_1[2:2]);
  OR2 I32 (o_0r1[0:0], gtint3_0[0:0], gtint3_1[0:0]);
  OR2 I33 (o_0r1[1:1], gtint3_0[1:1], gtint3_1[1:1]);
  OR2 I34 (o_0r1[2:2], gtint3_0[2:2], gtint3_1[2:2]);
  C2R I35 (sel3_0, selg3_0, icomplete3_0, reset);
  C2R I36 (sel3_1, selg3_1, icomplete3_0, reset);
  C2R I37 (gfint3_0[0:0], sel3_0, termf_1[0:0], reset);
  C2R I38 (gfint3_0[1:1], sel3_0, termf_1[1:1], reset);
  C2R I39 (gfint3_0[2:2], sel3_0, termf_1[2:2], reset);
  C2R I40 (gfint3_1[0:0], sel3_1, termf_2[0:0], reset);
  C2R I41 (gfint3_1[1:1], sel3_1, termf_2[1:1], reset);
  C2R I42 (gfint3_1[2:2], sel3_1, termf_2[2:2], reset);
  C2R I43 (gtint3_0[0:0], sel3_0, termt_1[0:0], reset);
  C2R I44 (gtint3_0[1:1], sel3_0, termt_1[1:1], reset);
  C2R I45 (gtint3_0[2:2], sel3_0, termt_1[2:2], reset);
  C2R I46 (gtint3_1[0:0], sel3_1, termt_2[0:0], reset);
  C2R I47 (gtint3_1[1:1], sel3_1, termt_2[1:1], reset);
  C2R I48 (gtint3_1[2:2], sel3_1, termt_2[2:2], reset);
  BUFF I49 (selg3_0, match30_0);
  C3 I50 (match30_0, i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I51 (selg3_1, match31_0);
  C3 I52 (match31_0, i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I53 (i_0a, o_0a);
endmodule

// tko2m3_1nm3b4_2nm3b1_3mx1_2_i0w2bt1o0w3bt2o0w3b TeakO [
//     (1,TeakOConstant 3 4),
//     (2,TeakOConstant 3 1),
//     (3,TeakOMux [[Imp 1 0],[Imp 2 0]] [(0,0+:2),(1,0+:3),(2,0+:3)])] [One 2,One 3]
module tko2m3_1nm3b4_2nm3b1_3mx1_2_i0w2bt1o0w3bt2o0w3b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [1:0] gocomp_0;
  wire [2:0] termf_1;
  wire [2:0] termf_2;
  wire [2:0] termt_1;
  wire [2:0] termt_2;
  wire [2:0] gfint3_0;
  wire [2:0] gfint3_1;
  wire [2:0] gtint3_0;
  wire [2:0] gtint3_1;
  wire selcomp3_0;
  wire selcomp3_1;
  wire sel3_0;
  wire sel3_1;
  wire selg3_0;
  wire selg3_1;
  wire icomplete3_0;
  wire scomplete3_0;
  wire [2:0] comp30_0;
  wire [2:0] comp31_0;
  wire [1:0] dcomp3_0;
  wire match30_0;
  wire match31_0;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  C2 I2 (go_0, gocomp_0[0:0], gocomp_0[1:1]);
  BUFF I3 (termt_1[2:2], go_0);
  GND I4 (termf_1[2:2]);
  BUFF I5 (termf_1[0:0], go_0);
  BUFF I6 (termf_1[1:1], go_0);
  GND I7 (termt_1[0:0]);
  GND I8 (termt_1[1:1]);
  BUFF I9 (termt_2[0:0], go_0);
  GND I10 (termf_2[0:0]);
  BUFF I11 (termf_2[1:1], go_0);
  BUFF I12 (termf_2[2:2], go_0);
  GND I13 (termt_2[1:1]);
  GND I14 (termt_2[2:2]);
  OR2 I15 (comp30_0[0:0], termf_1[0:0], termt_1[0:0]);
  OR2 I16 (comp30_0[1:1], termf_1[1:1], termt_1[1:1]);
  OR2 I17 (comp30_0[2:2], termf_1[2:2], termt_1[2:2]);
  C3 I18 (selcomp3_0, comp30_0[0:0], comp30_0[1:1], comp30_0[2:2]);
  OR2 I19 (comp31_0[0:0], termf_2[0:0], termt_2[0:0]);
  OR2 I20 (comp31_0[1:1], termf_2[1:1], termt_2[1:1]);
  OR2 I21 (comp31_0[2:2], termf_2[2:2], termt_2[2:2]);
  C3 I22 (selcomp3_1, comp31_0[0:0], comp31_0[1:1], comp31_0[2:2]);
  OR2 I23 (dcomp3_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I24 (dcomp3_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  C2 I25 (scomplete3_0, dcomp3_0[0:0], dcomp3_0[1:1]);
  C3 I26 (icomplete3_0, scomplete3_0, selcomp3_0, selcomp3_1);
  OR2 I27 (o_0r0[0:0], gfint3_0[0:0], gfint3_1[0:0]);
  OR2 I28 (o_0r0[1:1], gfint3_0[1:1], gfint3_1[1:1]);
  OR2 I29 (o_0r0[2:2], gfint3_0[2:2], gfint3_1[2:2]);
  OR2 I30 (o_0r1[0:0], gtint3_0[0:0], gtint3_1[0:0]);
  OR2 I31 (o_0r1[1:1], gtint3_0[1:1], gtint3_1[1:1]);
  OR2 I32 (o_0r1[2:2], gtint3_0[2:2], gtint3_1[2:2]);
  C2R I33 (sel3_0, selg3_0, icomplete3_0, reset);
  C2R I34 (sel3_1, selg3_1, icomplete3_0, reset);
  C2R I35 (gfint3_0[0:0], sel3_0, termf_1[0:0], reset);
  C2R I36 (gfint3_0[1:1], sel3_0, termf_1[1:1], reset);
  C2R I37 (gfint3_0[2:2], sel3_0, termf_1[2:2], reset);
  C2R I38 (gfint3_1[0:0], sel3_1, termf_2[0:0], reset);
  C2R I39 (gfint3_1[1:1], sel3_1, termf_2[1:1], reset);
  C2R I40 (gfint3_1[2:2], sel3_1, termf_2[2:2], reset);
  C2R I41 (gtint3_0[0:0], sel3_0, termt_1[0:0], reset);
  C2R I42 (gtint3_0[1:1], sel3_0, termt_1[1:1], reset);
  C2R I43 (gtint3_0[2:2], sel3_0, termt_1[2:2], reset);
  C2R I44 (gtint3_1[0:0], sel3_1, termt_2[0:0], reset);
  C2R I45 (gtint3_1[1:1], sel3_1, termt_2[1:1], reset);
  C2R I46 (gtint3_1[2:2], sel3_1, termt_2[2:2], reset);
  BUFF I47 (selg3_0, match30_0);
  C2 I48 (match30_0, i_0r1[0:0], i_0r0[1:1]);
  BUFF I49 (selg3_1, match31_0);
  C2 I50 (match31_0, i_0r0[0:0], i_0r1[1:1]);
  BUFF I51 (i_0a, o_0a);
endmodule

// tkf0mo0w0_o0w0_o0w0 TeakF [0,0,0] [One 0,Many [0,0,0]]
module tkf0mo0w0_o0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  input reset;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  BUFF I2 (o_2r, i_0r);
  C3 I3 (i_0a, o_0a, o_1a, o_2a);
endmodule

// latch tkl0x1 width = 0, depth = 1
module tkl0x1 (i_0r, i_0a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  input reset;
  wire b_0;
  C2R I0 (o_0r, i_0r, b_0, reset);
  INV I1 (b_0, o_0a);
  BUFF I2 (i_0a, o_0r);
endmodule

// latch tkl1x1 width = 1, depth = 1
module tkl1x1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire bna_0;
  wire bcomp_0;
  C2R I0 (o_0r0, i_0r0, bna_0, reset);
  C2R I1 (o_0r1, i_0r1, bna_0, reset);
  INV I2 (bna_0, o_0a);
  OR2 I3 (bcomp_0, o_0r0, o_0r1);
  BUFF I4 (i_0a, bcomp_0);
endmodule

// latch tkl32x1 width = 32, depth = 1
module tkl32x1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire bna_0;
  wire [31:0] bcomp_0;
  wire [10:0] simp991_0;
  wire [3:0] simp992_0;
  wire [1:0] simp993_0;
  C2R I0 (o_0r0[0:0], i_0r0[0:0], bna_0, reset);
  C2R I1 (o_0r0[1:1], i_0r0[1:1], bna_0, reset);
  C2R I2 (o_0r0[2:2], i_0r0[2:2], bna_0, reset);
  C2R I3 (o_0r0[3:3], i_0r0[3:3], bna_0, reset);
  C2R I4 (o_0r0[4:4], i_0r0[4:4], bna_0, reset);
  C2R I5 (o_0r0[5:5], i_0r0[5:5], bna_0, reset);
  C2R I6 (o_0r0[6:6], i_0r0[6:6], bna_0, reset);
  C2R I7 (o_0r0[7:7], i_0r0[7:7], bna_0, reset);
  C2R I8 (o_0r0[8:8], i_0r0[8:8], bna_0, reset);
  C2R I9 (o_0r0[9:9], i_0r0[9:9], bna_0, reset);
  C2R I10 (o_0r0[10:10], i_0r0[10:10], bna_0, reset);
  C2R I11 (o_0r0[11:11], i_0r0[11:11], bna_0, reset);
  C2R I12 (o_0r0[12:12], i_0r0[12:12], bna_0, reset);
  C2R I13 (o_0r0[13:13], i_0r0[13:13], bna_0, reset);
  C2R I14 (o_0r0[14:14], i_0r0[14:14], bna_0, reset);
  C2R I15 (o_0r0[15:15], i_0r0[15:15], bna_0, reset);
  C2R I16 (o_0r0[16:16], i_0r0[16:16], bna_0, reset);
  C2R I17 (o_0r0[17:17], i_0r0[17:17], bna_0, reset);
  C2R I18 (o_0r0[18:18], i_0r0[18:18], bna_0, reset);
  C2R I19 (o_0r0[19:19], i_0r0[19:19], bna_0, reset);
  C2R I20 (o_0r0[20:20], i_0r0[20:20], bna_0, reset);
  C2R I21 (o_0r0[21:21], i_0r0[21:21], bna_0, reset);
  C2R I22 (o_0r0[22:22], i_0r0[22:22], bna_0, reset);
  C2R I23 (o_0r0[23:23], i_0r0[23:23], bna_0, reset);
  C2R I24 (o_0r0[24:24], i_0r0[24:24], bna_0, reset);
  C2R I25 (o_0r0[25:25], i_0r0[25:25], bna_0, reset);
  C2R I26 (o_0r0[26:26], i_0r0[26:26], bna_0, reset);
  C2R I27 (o_0r0[27:27], i_0r0[27:27], bna_0, reset);
  C2R I28 (o_0r0[28:28], i_0r0[28:28], bna_0, reset);
  C2R I29 (o_0r0[29:29], i_0r0[29:29], bna_0, reset);
  C2R I30 (o_0r0[30:30], i_0r0[30:30], bna_0, reset);
  C2R I31 (o_0r0[31:31], i_0r0[31:31], bna_0, reset);
  C2R I32 (o_0r1[0:0], i_0r1[0:0], bna_0, reset);
  C2R I33 (o_0r1[1:1], i_0r1[1:1], bna_0, reset);
  C2R I34 (o_0r1[2:2], i_0r1[2:2], bna_0, reset);
  C2R I35 (o_0r1[3:3], i_0r1[3:3], bna_0, reset);
  C2R I36 (o_0r1[4:4], i_0r1[4:4], bna_0, reset);
  C2R I37 (o_0r1[5:5], i_0r1[5:5], bna_0, reset);
  C2R I38 (o_0r1[6:6], i_0r1[6:6], bna_0, reset);
  C2R I39 (o_0r1[7:7], i_0r1[7:7], bna_0, reset);
  C2R I40 (o_0r1[8:8], i_0r1[8:8], bna_0, reset);
  C2R I41 (o_0r1[9:9], i_0r1[9:9], bna_0, reset);
  C2R I42 (o_0r1[10:10], i_0r1[10:10], bna_0, reset);
  C2R I43 (o_0r1[11:11], i_0r1[11:11], bna_0, reset);
  C2R I44 (o_0r1[12:12], i_0r1[12:12], bna_0, reset);
  C2R I45 (o_0r1[13:13], i_0r1[13:13], bna_0, reset);
  C2R I46 (o_0r1[14:14], i_0r1[14:14], bna_0, reset);
  C2R I47 (o_0r1[15:15], i_0r1[15:15], bna_0, reset);
  C2R I48 (o_0r1[16:16], i_0r1[16:16], bna_0, reset);
  C2R I49 (o_0r1[17:17], i_0r1[17:17], bna_0, reset);
  C2R I50 (o_0r1[18:18], i_0r1[18:18], bna_0, reset);
  C2R I51 (o_0r1[19:19], i_0r1[19:19], bna_0, reset);
  C2R I52 (o_0r1[20:20], i_0r1[20:20], bna_0, reset);
  C2R I53 (o_0r1[21:21], i_0r1[21:21], bna_0, reset);
  C2R I54 (o_0r1[22:22], i_0r1[22:22], bna_0, reset);
  C2R I55 (o_0r1[23:23], i_0r1[23:23], bna_0, reset);
  C2R I56 (o_0r1[24:24], i_0r1[24:24], bna_0, reset);
  C2R I57 (o_0r1[25:25], i_0r1[25:25], bna_0, reset);
  C2R I58 (o_0r1[26:26], i_0r1[26:26], bna_0, reset);
  C2R I59 (o_0r1[27:27], i_0r1[27:27], bna_0, reset);
  C2R I60 (o_0r1[28:28], i_0r1[28:28], bna_0, reset);
  C2R I61 (o_0r1[29:29], i_0r1[29:29], bna_0, reset);
  C2R I62 (o_0r1[30:30], i_0r1[30:30], bna_0, reset);
  C2R I63 (o_0r1[31:31], i_0r1[31:31], bna_0, reset);
  INV I64 (bna_0, o_0a);
  OR2 I65 (bcomp_0[0:0], o_0r0[0:0], o_0r1[0:0]);
  OR2 I66 (bcomp_0[1:1], o_0r0[1:1], o_0r1[1:1]);
  OR2 I67 (bcomp_0[2:2], o_0r0[2:2], o_0r1[2:2]);
  OR2 I68 (bcomp_0[3:3], o_0r0[3:3], o_0r1[3:3]);
  OR2 I69 (bcomp_0[4:4], o_0r0[4:4], o_0r1[4:4]);
  OR2 I70 (bcomp_0[5:5], o_0r0[5:5], o_0r1[5:5]);
  OR2 I71 (bcomp_0[6:6], o_0r0[6:6], o_0r1[6:6]);
  OR2 I72 (bcomp_0[7:7], o_0r0[7:7], o_0r1[7:7]);
  OR2 I73 (bcomp_0[8:8], o_0r0[8:8], o_0r1[8:8]);
  OR2 I74 (bcomp_0[9:9], o_0r0[9:9], o_0r1[9:9]);
  OR2 I75 (bcomp_0[10:10], o_0r0[10:10], o_0r1[10:10]);
  OR2 I76 (bcomp_0[11:11], o_0r0[11:11], o_0r1[11:11]);
  OR2 I77 (bcomp_0[12:12], o_0r0[12:12], o_0r1[12:12]);
  OR2 I78 (bcomp_0[13:13], o_0r0[13:13], o_0r1[13:13]);
  OR2 I79 (bcomp_0[14:14], o_0r0[14:14], o_0r1[14:14]);
  OR2 I80 (bcomp_0[15:15], o_0r0[15:15], o_0r1[15:15]);
  OR2 I81 (bcomp_0[16:16], o_0r0[16:16], o_0r1[16:16]);
  OR2 I82 (bcomp_0[17:17], o_0r0[17:17], o_0r1[17:17]);
  OR2 I83 (bcomp_0[18:18], o_0r0[18:18], o_0r1[18:18]);
  OR2 I84 (bcomp_0[19:19], o_0r0[19:19], o_0r1[19:19]);
  OR2 I85 (bcomp_0[20:20], o_0r0[20:20], o_0r1[20:20]);
  OR2 I86 (bcomp_0[21:21], o_0r0[21:21], o_0r1[21:21]);
  OR2 I87 (bcomp_0[22:22], o_0r0[22:22], o_0r1[22:22]);
  OR2 I88 (bcomp_0[23:23], o_0r0[23:23], o_0r1[23:23]);
  OR2 I89 (bcomp_0[24:24], o_0r0[24:24], o_0r1[24:24]);
  OR2 I90 (bcomp_0[25:25], o_0r0[25:25], o_0r1[25:25]);
  OR2 I91 (bcomp_0[26:26], o_0r0[26:26], o_0r1[26:26]);
  OR2 I92 (bcomp_0[27:27], o_0r0[27:27], o_0r1[27:27]);
  OR2 I93 (bcomp_0[28:28], o_0r0[28:28], o_0r1[28:28]);
  OR2 I94 (bcomp_0[29:29], o_0r0[29:29], o_0r1[29:29]);
  OR2 I95 (bcomp_0[30:30], o_0r0[30:30], o_0r1[30:30]);
  OR2 I96 (bcomp_0[31:31], o_0r0[31:31], o_0r1[31:31]);
  C3 I97 (simp991_0[0:0], bcomp_0[0:0], bcomp_0[1:1], bcomp_0[2:2]);
  C3 I98 (simp991_0[1:1], bcomp_0[3:3], bcomp_0[4:4], bcomp_0[5:5]);
  C3 I99 (simp991_0[2:2], bcomp_0[6:6], bcomp_0[7:7], bcomp_0[8:8]);
  C3 I100 (simp991_0[3:3], bcomp_0[9:9], bcomp_0[10:10], bcomp_0[11:11]);
  C3 I101 (simp991_0[4:4], bcomp_0[12:12], bcomp_0[13:13], bcomp_0[14:14]);
  C3 I102 (simp991_0[5:5], bcomp_0[15:15], bcomp_0[16:16], bcomp_0[17:17]);
  C3 I103 (simp991_0[6:6], bcomp_0[18:18], bcomp_0[19:19], bcomp_0[20:20]);
  C3 I104 (simp991_0[7:7], bcomp_0[21:21], bcomp_0[22:22], bcomp_0[23:23]);
  C3 I105 (simp991_0[8:8], bcomp_0[24:24], bcomp_0[25:25], bcomp_0[26:26]);
  C3 I106 (simp991_0[9:9], bcomp_0[27:27], bcomp_0[28:28], bcomp_0[29:29]);
  C2 I107 (simp991_0[10:10], bcomp_0[30:30], bcomp_0[31:31]);
  C3 I108 (simp992_0[0:0], simp991_0[0:0], simp991_0[1:1], simp991_0[2:2]);
  C3 I109 (simp992_0[1:1], simp991_0[3:3], simp991_0[4:4], simp991_0[5:5]);
  C3 I110 (simp992_0[2:2], simp991_0[6:6], simp991_0[7:7], simp991_0[8:8]);
  C2 I111 (simp992_0[3:3], simp991_0[9:9], simp991_0[10:10]);
  C3 I112 (simp993_0[0:0], simp992_0[0:0], simp992_0[1:1], simp992_0[2:2]);
  BUFF I113 (simp993_0[1:1], simp992_0[3:3]);
  C2 I114 (i_0a, simp993_0[0:0], simp993_0[1:1]);
endmodule

// latch tkl3x1 width = 3, depth = 1
module tkl3x1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire bna_0;
  wire [2:0] bcomp_0;
  C2R I0 (o_0r0[0:0], i_0r0[0:0], bna_0, reset);
  C2R I1 (o_0r0[1:1], i_0r0[1:1], bna_0, reset);
  C2R I2 (o_0r0[2:2], i_0r0[2:2], bna_0, reset);
  C2R I3 (o_0r1[0:0], i_0r1[0:0], bna_0, reset);
  C2R I4 (o_0r1[1:1], i_0r1[1:1], bna_0, reset);
  C2R I5 (o_0r1[2:2], i_0r1[2:2], bna_0, reset);
  INV I6 (bna_0, o_0a);
  OR2 I7 (bcomp_0[0:0], o_0r0[0:0], o_0r1[0:0]);
  OR2 I8 (bcomp_0[1:1], o_0r0[1:1], o_0r1[1:1]);
  OR2 I9 (bcomp_0[2:2], o_0r0[2:2], o_0r1[2:2]);
  C3 I10 (i_0a, bcomp_0[0:0], bcomp_0[1:1], bcomp_0[2:2]);
endmodule

// latch tkl10x1 width = 10, depth = 1
module tkl10x1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [9:0] i_0r0;
  input [9:0] i_0r1;
  output i_0a;
  output [9:0] o_0r0;
  output [9:0] o_0r1;
  input o_0a;
  input reset;
  wire bna_0;
  wire [9:0] bcomp_0;
  wire [3:0] simp331_0;
  wire [1:0] simp332_0;
  C2R I0 (o_0r0[0:0], i_0r0[0:0], bna_0, reset);
  C2R I1 (o_0r0[1:1], i_0r0[1:1], bna_0, reset);
  C2R I2 (o_0r0[2:2], i_0r0[2:2], bna_0, reset);
  C2R I3 (o_0r0[3:3], i_0r0[3:3], bna_0, reset);
  C2R I4 (o_0r0[4:4], i_0r0[4:4], bna_0, reset);
  C2R I5 (o_0r0[5:5], i_0r0[5:5], bna_0, reset);
  C2R I6 (o_0r0[6:6], i_0r0[6:6], bna_0, reset);
  C2R I7 (o_0r0[7:7], i_0r0[7:7], bna_0, reset);
  C2R I8 (o_0r0[8:8], i_0r0[8:8], bna_0, reset);
  C2R I9 (o_0r0[9:9], i_0r0[9:9], bna_0, reset);
  C2R I10 (o_0r1[0:0], i_0r1[0:0], bna_0, reset);
  C2R I11 (o_0r1[1:1], i_0r1[1:1], bna_0, reset);
  C2R I12 (o_0r1[2:2], i_0r1[2:2], bna_0, reset);
  C2R I13 (o_0r1[3:3], i_0r1[3:3], bna_0, reset);
  C2R I14 (o_0r1[4:4], i_0r1[4:4], bna_0, reset);
  C2R I15 (o_0r1[5:5], i_0r1[5:5], bna_0, reset);
  C2R I16 (o_0r1[6:6], i_0r1[6:6], bna_0, reset);
  C2R I17 (o_0r1[7:7], i_0r1[7:7], bna_0, reset);
  C2R I18 (o_0r1[8:8], i_0r1[8:8], bna_0, reset);
  C2R I19 (o_0r1[9:9], i_0r1[9:9], bna_0, reset);
  INV I20 (bna_0, o_0a);
  OR2 I21 (bcomp_0[0:0], o_0r0[0:0], o_0r1[0:0]);
  OR2 I22 (bcomp_0[1:1], o_0r0[1:1], o_0r1[1:1]);
  OR2 I23 (bcomp_0[2:2], o_0r0[2:2], o_0r1[2:2]);
  OR2 I24 (bcomp_0[3:3], o_0r0[3:3], o_0r1[3:3]);
  OR2 I25 (bcomp_0[4:4], o_0r0[4:4], o_0r1[4:4]);
  OR2 I26 (bcomp_0[5:5], o_0r0[5:5], o_0r1[5:5]);
  OR2 I27 (bcomp_0[6:6], o_0r0[6:6], o_0r1[6:6]);
  OR2 I28 (bcomp_0[7:7], o_0r0[7:7], o_0r1[7:7]);
  OR2 I29 (bcomp_0[8:8], o_0r0[8:8], o_0r1[8:8]);
  OR2 I30 (bcomp_0[9:9], o_0r0[9:9], o_0r1[9:9]);
  C3 I31 (simp331_0[0:0], bcomp_0[0:0], bcomp_0[1:1], bcomp_0[2:2]);
  C3 I32 (simp331_0[1:1], bcomp_0[3:3], bcomp_0[4:4], bcomp_0[5:5]);
  C3 I33 (simp331_0[2:2], bcomp_0[6:6], bcomp_0[7:7], bcomp_0[8:8]);
  BUFF I34 (simp331_0[3:3], bcomp_0[9:9]);
  C3 I35 (simp332_0[0:0], simp331_0[0:0], simp331_0[1:1], simp331_0[2:2]);
  BUFF I36 (simp332_0[1:1], simp331_0[3:3]);
  C2 I37 (i_0a, simp332_0[0:0], simp332_0[1:1]);
endmodule

// latch tkl6x1 width = 6, depth = 1
module tkl6x1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [5:0] i_0r0;
  input [5:0] i_0r1;
  output i_0a;
  output [5:0] o_0r0;
  output [5:0] o_0r1;
  input o_0a;
  input reset;
  wire bna_0;
  wire [5:0] bcomp_0;
  wire [1:0] simp211_0;
  C2R I0 (o_0r0[0:0], i_0r0[0:0], bna_0, reset);
  C2R I1 (o_0r0[1:1], i_0r0[1:1], bna_0, reset);
  C2R I2 (o_0r0[2:2], i_0r0[2:2], bna_0, reset);
  C2R I3 (o_0r0[3:3], i_0r0[3:3], bna_0, reset);
  C2R I4 (o_0r0[4:4], i_0r0[4:4], bna_0, reset);
  C2R I5 (o_0r0[5:5], i_0r0[5:5], bna_0, reset);
  C2R I6 (o_0r1[0:0], i_0r1[0:0], bna_0, reset);
  C2R I7 (o_0r1[1:1], i_0r1[1:1], bna_0, reset);
  C2R I8 (o_0r1[2:2], i_0r1[2:2], bna_0, reset);
  C2R I9 (o_0r1[3:3], i_0r1[3:3], bna_0, reset);
  C2R I10 (o_0r1[4:4], i_0r1[4:4], bna_0, reset);
  C2R I11 (o_0r1[5:5], i_0r1[5:5], bna_0, reset);
  INV I12 (bna_0, o_0a);
  OR2 I13 (bcomp_0[0:0], o_0r0[0:0], o_0r1[0:0]);
  OR2 I14 (bcomp_0[1:1], o_0r0[1:1], o_0r1[1:1]);
  OR2 I15 (bcomp_0[2:2], o_0r0[2:2], o_0r1[2:2]);
  OR2 I16 (bcomp_0[3:3], o_0r0[3:3], o_0r1[3:3]);
  OR2 I17 (bcomp_0[4:4], o_0r0[4:4], o_0r1[4:4]);
  OR2 I18 (bcomp_0[5:5], o_0r0[5:5], o_0r1[5:5]);
  C3 I19 (simp211_0[0:0], bcomp_0[0:0], bcomp_0[1:1], bcomp_0[2:2]);
  C3 I20 (simp211_0[1:1], bcomp_0[3:3], bcomp_0[4:4], bcomp_0[5:5]);
  C2 I21 (i_0a, simp211_0[0:0], simp211_0[1:1]);
endmodule

// latch tkl64x1 width = 64, depth = 1
module tkl64x1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [63:0] i_0r0;
  input [63:0] i_0r1;
  output i_0a;
  output [63:0] o_0r0;
  output [63:0] o_0r1;
  input o_0a;
  input reset;
  wire bna_0;
  wire [63:0] bcomp_0;
  wire [21:0] simp1951_0;
  wire [7:0] simp1952_0;
  wire [2:0] simp1953_0;
  C2R I0 (o_0r0[0:0], i_0r0[0:0], bna_0, reset);
  C2R I1 (o_0r0[1:1], i_0r0[1:1], bna_0, reset);
  C2R I2 (o_0r0[2:2], i_0r0[2:2], bna_0, reset);
  C2R I3 (o_0r0[3:3], i_0r0[3:3], bna_0, reset);
  C2R I4 (o_0r0[4:4], i_0r0[4:4], bna_0, reset);
  C2R I5 (o_0r0[5:5], i_0r0[5:5], bna_0, reset);
  C2R I6 (o_0r0[6:6], i_0r0[6:6], bna_0, reset);
  C2R I7 (o_0r0[7:7], i_0r0[7:7], bna_0, reset);
  C2R I8 (o_0r0[8:8], i_0r0[8:8], bna_0, reset);
  C2R I9 (o_0r0[9:9], i_0r0[9:9], bna_0, reset);
  C2R I10 (o_0r0[10:10], i_0r0[10:10], bna_0, reset);
  C2R I11 (o_0r0[11:11], i_0r0[11:11], bna_0, reset);
  C2R I12 (o_0r0[12:12], i_0r0[12:12], bna_0, reset);
  C2R I13 (o_0r0[13:13], i_0r0[13:13], bna_0, reset);
  C2R I14 (o_0r0[14:14], i_0r0[14:14], bna_0, reset);
  C2R I15 (o_0r0[15:15], i_0r0[15:15], bna_0, reset);
  C2R I16 (o_0r0[16:16], i_0r0[16:16], bna_0, reset);
  C2R I17 (o_0r0[17:17], i_0r0[17:17], bna_0, reset);
  C2R I18 (o_0r0[18:18], i_0r0[18:18], bna_0, reset);
  C2R I19 (o_0r0[19:19], i_0r0[19:19], bna_0, reset);
  C2R I20 (o_0r0[20:20], i_0r0[20:20], bna_0, reset);
  C2R I21 (o_0r0[21:21], i_0r0[21:21], bna_0, reset);
  C2R I22 (o_0r0[22:22], i_0r0[22:22], bna_0, reset);
  C2R I23 (o_0r0[23:23], i_0r0[23:23], bna_0, reset);
  C2R I24 (o_0r0[24:24], i_0r0[24:24], bna_0, reset);
  C2R I25 (o_0r0[25:25], i_0r0[25:25], bna_0, reset);
  C2R I26 (o_0r0[26:26], i_0r0[26:26], bna_0, reset);
  C2R I27 (o_0r0[27:27], i_0r0[27:27], bna_0, reset);
  C2R I28 (o_0r0[28:28], i_0r0[28:28], bna_0, reset);
  C2R I29 (o_0r0[29:29], i_0r0[29:29], bna_0, reset);
  C2R I30 (o_0r0[30:30], i_0r0[30:30], bna_0, reset);
  C2R I31 (o_0r0[31:31], i_0r0[31:31], bna_0, reset);
  C2R I32 (o_0r0[32:32], i_0r0[32:32], bna_0, reset);
  C2R I33 (o_0r0[33:33], i_0r0[33:33], bna_0, reset);
  C2R I34 (o_0r0[34:34], i_0r0[34:34], bna_0, reset);
  C2R I35 (o_0r0[35:35], i_0r0[35:35], bna_0, reset);
  C2R I36 (o_0r0[36:36], i_0r0[36:36], bna_0, reset);
  C2R I37 (o_0r0[37:37], i_0r0[37:37], bna_0, reset);
  C2R I38 (o_0r0[38:38], i_0r0[38:38], bna_0, reset);
  C2R I39 (o_0r0[39:39], i_0r0[39:39], bna_0, reset);
  C2R I40 (o_0r0[40:40], i_0r0[40:40], bna_0, reset);
  C2R I41 (o_0r0[41:41], i_0r0[41:41], bna_0, reset);
  C2R I42 (o_0r0[42:42], i_0r0[42:42], bna_0, reset);
  C2R I43 (o_0r0[43:43], i_0r0[43:43], bna_0, reset);
  C2R I44 (o_0r0[44:44], i_0r0[44:44], bna_0, reset);
  C2R I45 (o_0r0[45:45], i_0r0[45:45], bna_0, reset);
  C2R I46 (o_0r0[46:46], i_0r0[46:46], bna_0, reset);
  C2R I47 (o_0r0[47:47], i_0r0[47:47], bna_0, reset);
  C2R I48 (o_0r0[48:48], i_0r0[48:48], bna_0, reset);
  C2R I49 (o_0r0[49:49], i_0r0[49:49], bna_0, reset);
  C2R I50 (o_0r0[50:50], i_0r0[50:50], bna_0, reset);
  C2R I51 (o_0r0[51:51], i_0r0[51:51], bna_0, reset);
  C2R I52 (o_0r0[52:52], i_0r0[52:52], bna_0, reset);
  C2R I53 (o_0r0[53:53], i_0r0[53:53], bna_0, reset);
  C2R I54 (o_0r0[54:54], i_0r0[54:54], bna_0, reset);
  C2R I55 (o_0r0[55:55], i_0r0[55:55], bna_0, reset);
  C2R I56 (o_0r0[56:56], i_0r0[56:56], bna_0, reset);
  C2R I57 (o_0r0[57:57], i_0r0[57:57], bna_0, reset);
  C2R I58 (o_0r0[58:58], i_0r0[58:58], bna_0, reset);
  C2R I59 (o_0r0[59:59], i_0r0[59:59], bna_0, reset);
  C2R I60 (o_0r0[60:60], i_0r0[60:60], bna_0, reset);
  C2R I61 (o_0r0[61:61], i_0r0[61:61], bna_0, reset);
  C2R I62 (o_0r0[62:62], i_0r0[62:62], bna_0, reset);
  C2R I63 (o_0r0[63:63], i_0r0[63:63], bna_0, reset);
  C2R I64 (o_0r1[0:0], i_0r1[0:0], bna_0, reset);
  C2R I65 (o_0r1[1:1], i_0r1[1:1], bna_0, reset);
  C2R I66 (o_0r1[2:2], i_0r1[2:2], bna_0, reset);
  C2R I67 (o_0r1[3:3], i_0r1[3:3], bna_0, reset);
  C2R I68 (o_0r1[4:4], i_0r1[4:4], bna_0, reset);
  C2R I69 (o_0r1[5:5], i_0r1[5:5], bna_0, reset);
  C2R I70 (o_0r1[6:6], i_0r1[6:6], bna_0, reset);
  C2R I71 (o_0r1[7:7], i_0r1[7:7], bna_0, reset);
  C2R I72 (o_0r1[8:8], i_0r1[8:8], bna_0, reset);
  C2R I73 (o_0r1[9:9], i_0r1[9:9], bna_0, reset);
  C2R I74 (o_0r1[10:10], i_0r1[10:10], bna_0, reset);
  C2R I75 (o_0r1[11:11], i_0r1[11:11], bna_0, reset);
  C2R I76 (o_0r1[12:12], i_0r1[12:12], bna_0, reset);
  C2R I77 (o_0r1[13:13], i_0r1[13:13], bna_0, reset);
  C2R I78 (o_0r1[14:14], i_0r1[14:14], bna_0, reset);
  C2R I79 (o_0r1[15:15], i_0r1[15:15], bna_0, reset);
  C2R I80 (o_0r1[16:16], i_0r1[16:16], bna_0, reset);
  C2R I81 (o_0r1[17:17], i_0r1[17:17], bna_0, reset);
  C2R I82 (o_0r1[18:18], i_0r1[18:18], bna_0, reset);
  C2R I83 (o_0r1[19:19], i_0r1[19:19], bna_0, reset);
  C2R I84 (o_0r1[20:20], i_0r1[20:20], bna_0, reset);
  C2R I85 (o_0r1[21:21], i_0r1[21:21], bna_0, reset);
  C2R I86 (o_0r1[22:22], i_0r1[22:22], bna_0, reset);
  C2R I87 (o_0r1[23:23], i_0r1[23:23], bna_0, reset);
  C2R I88 (o_0r1[24:24], i_0r1[24:24], bna_0, reset);
  C2R I89 (o_0r1[25:25], i_0r1[25:25], bna_0, reset);
  C2R I90 (o_0r1[26:26], i_0r1[26:26], bna_0, reset);
  C2R I91 (o_0r1[27:27], i_0r1[27:27], bna_0, reset);
  C2R I92 (o_0r1[28:28], i_0r1[28:28], bna_0, reset);
  C2R I93 (o_0r1[29:29], i_0r1[29:29], bna_0, reset);
  C2R I94 (o_0r1[30:30], i_0r1[30:30], bna_0, reset);
  C2R I95 (o_0r1[31:31], i_0r1[31:31], bna_0, reset);
  C2R I96 (o_0r1[32:32], i_0r1[32:32], bna_0, reset);
  C2R I97 (o_0r1[33:33], i_0r1[33:33], bna_0, reset);
  C2R I98 (o_0r1[34:34], i_0r1[34:34], bna_0, reset);
  C2R I99 (o_0r1[35:35], i_0r1[35:35], bna_0, reset);
  C2R I100 (o_0r1[36:36], i_0r1[36:36], bna_0, reset);
  C2R I101 (o_0r1[37:37], i_0r1[37:37], bna_0, reset);
  C2R I102 (o_0r1[38:38], i_0r1[38:38], bna_0, reset);
  C2R I103 (o_0r1[39:39], i_0r1[39:39], bna_0, reset);
  C2R I104 (o_0r1[40:40], i_0r1[40:40], bna_0, reset);
  C2R I105 (o_0r1[41:41], i_0r1[41:41], bna_0, reset);
  C2R I106 (o_0r1[42:42], i_0r1[42:42], bna_0, reset);
  C2R I107 (o_0r1[43:43], i_0r1[43:43], bna_0, reset);
  C2R I108 (o_0r1[44:44], i_0r1[44:44], bna_0, reset);
  C2R I109 (o_0r1[45:45], i_0r1[45:45], bna_0, reset);
  C2R I110 (o_0r1[46:46], i_0r1[46:46], bna_0, reset);
  C2R I111 (o_0r1[47:47], i_0r1[47:47], bna_0, reset);
  C2R I112 (o_0r1[48:48], i_0r1[48:48], bna_0, reset);
  C2R I113 (o_0r1[49:49], i_0r1[49:49], bna_0, reset);
  C2R I114 (o_0r1[50:50], i_0r1[50:50], bna_0, reset);
  C2R I115 (o_0r1[51:51], i_0r1[51:51], bna_0, reset);
  C2R I116 (o_0r1[52:52], i_0r1[52:52], bna_0, reset);
  C2R I117 (o_0r1[53:53], i_0r1[53:53], bna_0, reset);
  C2R I118 (o_0r1[54:54], i_0r1[54:54], bna_0, reset);
  C2R I119 (o_0r1[55:55], i_0r1[55:55], bna_0, reset);
  C2R I120 (o_0r1[56:56], i_0r1[56:56], bna_0, reset);
  C2R I121 (o_0r1[57:57], i_0r1[57:57], bna_0, reset);
  C2R I122 (o_0r1[58:58], i_0r1[58:58], bna_0, reset);
  C2R I123 (o_0r1[59:59], i_0r1[59:59], bna_0, reset);
  C2R I124 (o_0r1[60:60], i_0r1[60:60], bna_0, reset);
  C2R I125 (o_0r1[61:61], i_0r1[61:61], bna_0, reset);
  C2R I126 (o_0r1[62:62], i_0r1[62:62], bna_0, reset);
  C2R I127 (o_0r1[63:63], i_0r1[63:63], bna_0, reset);
  INV I128 (bna_0, o_0a);
  OR2 I129 (bcomp_0[0:0], o_0r0[0:0], o_0r1[0:0]);
  OR2 I130 (bcomp_0[1:1], o_0r0[1:1], o_0r1[1:1]);
  OR2 I131 (bcomp_0[2:2], o_0r0[2:2], o_0r1[2:2]);
  OR2 I132 (bcomp_0[3:3], o_0r0[3:3], o_0r1[3:3]);
  OR2 I133 (bcomp_0[4:4], o_0r0[4:4], o_0r1[4:4]);
  OR2 I134 (bcomp_0[5:5], o_0r0[5:5], o_0r1[5:5]);
  OR2 I135 (bcomp_0[6:6], o_0r0[6:6], o_0r1[6:6]);
  OR2 I136 (bcomp_0[7:7], o_0r0[7:7], o_0r1[7:7]);
  OR2 I137 (bcomp_0[8:8], o_0r0[8:8], o_0r1[8:8]);
  OR2 I138 (bcomp_0[9:9], o_0r0[9:9], o_0r1[9:9]);
  OR2 I139 (bcomp_0[10:10], o_0r0[10:10], o_0r1[10:10]);
  OR2 I140 (bcomp_0[11:11], o_0r0[11:11], o_0r1[11:11]);
  OR2 I141 (bcomp_0[12:12], o_0r0[12:12], o_0r1[12:12]);
  OR2 I142 (bcomp_0[13:13], o_0r0[13:13], o_0r1[13:13]);
  OR2 I143 (bcomp_0[14:14], o_0r0[14:14], o_0r1[14:14]);
  OR2 I144 (bcomp_0[15:15], o_0r0[15:15], o_0r1[15:15]);
  OR2 I145 (bcomp_0[16:16], o_0r0[16:16], o_0r1[16:16]);
  OR2 I146 (bcomp_0[17:17], o_0r0[17:17], o_0r1[17:17]);
  OR2 I147 (bcomp_0[18:18], o_0r0[18:18], o_0r1[18:18]);
  OR2 I148 (bcomp_0[19:19], o_0r0[19:19], o_0r1[19:19]);
  OR2 I149 (bcomp_0[20:20], o_0r0[20:20], o_0r1[20:20]);
  OR2 I150 (bcomp_0[21:21], o_0r0[21:21], o_0r1[21:21]);
  OR2 I151 (bcomp_0[22:22], o_0r0[22:22], o_0r1[22:22]);
  OR2 I152 (bcomp_0[23:23], o_0r0[23:23], o_0r1[23:23]);
  OR2 I153 (bcomp_0[24:24], o_0r0[24:24], o_0r1[24:24]);
  OR2 I154 (bcomp_0[25:25], o_0r0[25:25], o_0r1[25:25]);
  OR2 I155 (bcomp_0[26:26], o_0r0[26:26], o_0r1[26:26]);
  OR2 I156 (bcomp_0[27:27], o_0r0[27:27], o_0r1[27:27]);
  OR2 I157 (bcomp_0[28:28], o_0r0[28:28], o_0r1[28:28]);
  OR2 I158 (bcomp_0[29:29], o_0r0[29:29], o_0r1[29:29]);
  OR2 I159 (bcomp_0[30:30], o_0r0[30:30], o_0r1[30:30]);
  OR2 I160 (bcomp_0[31:31], o_0r0[31:31], o_0r1[31:31]);
  OR2 I161 (bcomp_0[32:32], o_0r0[32:32], o_0r1[32:32]);
  OR2 I162 (bcomp_0[33:33], o_0r0[33:33], o_0r1[33:33]);
  OR2 I163 (bcomp_0[34:34], o_0r0[34:34], o_0r1[34:34]);
  OR2 I164 (bcomp_0[35:35], o_0r0[35:35], o_0r1[35:35]);
  OR2 I165 (bcomp_0[36:36], o_0r0[36:36], o_0r1[36:36]);
  OR2 I166 (bcomp_0[37:37], o_0r0[37:37], o_0r1[37:37]);
  OR2 I167 (bcomp_0[38:38], o_0r0[38:38], o_0r1[38:38]);
  OR2 I168 (bcomp_0[39:39], o_0r0[39:39], o_0r1[39:39]);
  OR2 I169 (bcomp_0[40:40], o_0r0[40:40], o_0r1[40:40]);
  OR2 I170 (bcomp_0[41:41], o_0r0[41:41], o_0r1[41:41]);
  OR2 I171 (bcomp_0[42:42], o_0r0[42:42], o_0r1[42:42]);
  OR2 I172 (bcomp_0[43:43], o_0r0[43:43], o_0r1[43:43]);
  OR2 I173 (bcomp_0[44:44], o_0r0[44:44], o_0r1[44:44]);
  OR2 I174 (bcomp_0[45:45], o_0r0[45:45], o_0r1[45:45]);
  OR2 I175 (bcomp_0[46:46], o_0r0[46:46], o_0r1[46:46]);
  OR2 I176 (bcomp_0[47:47], o_0r0[47:47], o_0r1[47:47]);
  OR2 I177 (bcomp_0[48:48], o_0r0[48:48], o_0r1[48:48]);
  OR2 I178 (bcomp_0[49:49], o_0r0[49:49], o_0r1[49:49]);
  OR2 I179 (bcomp_0[50:50], o_0r0[50:50], o_0r1[50:50]);
  OR2 I180 (bcomp_0[51:51], o_0r0[51:51], o_0r1[51:51]);
  OR2 I181 (bcomp_0[52:52], o_0r0[52:52], o_0r1[52:52]);
  OR2 I182 (bcomp_0[53:53], o_0r0[53:53], o_0r1[53:53]);
  OR2 I183 (bcomp_0[54:54], o_0r0[54:54], o_0r1[54:54]);
  OR2 I184 (bcomp_0[55:55], o_0r0[55:55], o_0r1[55:55]);
  OR2 I185 (bcomp_0[56:56], o_0r0[56:56], o_0r1[56:56]);
  OR2 I186 (bcomp_0[57:57], o_0r0[57:57], o_0r1[57:57]);
  OR2 I187 (bcomp_0[58:58], o_0r0[58:58], o_0r1[58:58]);
  OR2 I188 (bcomp_0[59:59], o_0r0[59:59], o_0r1[59:59]);
  OR2 I189 (bcomp_0[60:60], o_0r0[60:60], o_0r1[60:60]);
  OR2 I190 (bcomp_0[61:61], o_0r0[61:61], o_0r1[61:61]);
  OR2 I191 (bcomp_0[62:62], o_0r0[62:62], o_0r1[62:62]);
  OR2 I192 (bcomp_0[63:63], o_0r0[63:63], o_0r1[63:63]);
  C3 I193 (simp1951_0[0:0], bcomp_0[0:0], bcomp_0[1:1], bcomp_0[2:2]);
  C3 I194 (simp1951_0[1:1], bcomp_0[3:3], bcomp_0[4:4], bcomp_0[5:5]);
  C3 I195 (simp1951_0[2:2], bcomp_0[6:6], bcomp_0[7:7], bcomp_0[8:8]);
  C3 I196 (simp1951_0[3:3], bcomp_0[9:9], bcomp_0[10:10], bcomp_0[11:11]);
  C3 I197 (simp1951_0[4:4], bcomp_0[12:12], bcomp_0[13:13], bcomp_0[14:14]);
  C3 I198 (simp1951_0[5:5], bcomp_0[15:15], bcomp_0[16:16], bcomp_0[17:17]);
  C3 I199 (simp1951_0[6:6], bcomp_0[18:18], bcomp_0[19:19], bcomp_0[20:20]);
  C3 I200 (simp1951_0[7:7], bcomp_0[21:21], bcomp_0[22:22], bcomp_0[23:23]);
  C3 I201 (simp1951_0[8:8], bcomp_0[24:24], bcomp_0[25:25], bcomp_0[26:26]);
  C3 I202 (simp1951_0[9:9], bcomp_0[27:27], bcomp_0[28:28], bcomp_0[29:29]);
  C3 I203 (simp1951_0[10:10], bcomp_0[30:30], bcomp_0[31:31], bcomp_0[32:32]);
  C3 I204 (simp1951_0[11:11], bcomp_0[33:33], bcomp_0[34:34], bcomp_0[35:35]);
  C3 I205 (simp1951_0[12:12], bcomp_0[36:36], bcomp_0[37:37], bcomp_0[38:38]);
  C3 I206 (simp1951_0[13:13], bcomp_0[39:39], bcomp_0[40:40], bcomp_0[41:41]);
  C3 I207 (simp1951_0[14:14], bcomp_0[42:42], bcomp_0[43:43], bcomp_0[44:44]);
  C3 I208 (simp1951_0[15:15], bcomp_0[45:45], bcomp_0[46:46], bcomp_0[47:47]);
  C3 I209 (simp1951_0[16:16], bcomp_0[48:48], bcomp_0[49:49], bcomp_0[50:50]);
  C3 I210 (simp1951_0[17:17], bcomp_0[51:51], bcomp_0[52:52], bcomp_0[53:53]);
  C3 I211 (simp1951_0[18:18], bcomp_0[54:54], bcomp_0[55:55], bcomp_0[56:56]);
  C3 I212 (simp1951_0[19:19], bcomp_0[57:57], bcomp_0[58:58], bcomp_0[59:59]);
  C3 I213 (simp1951_0[20:20], bcomp_0[60:60], bcomp_0[61:61], bcomp_0[62:62]);
  BUFF I214 (simp1951_0[21:21], bcomp_0[63:63]);
  C3 I215 (simp1952_0[0:0], simp1951_0[0:0], simp1951_0[1:1], simp1951_0[2:2]);
  C3 I216 (simp1952_0[1:1], simp1951_0[3:3], simp1951_0[4:4], simp1951_0[5:5]);
  C3 I217 (simp1952_0[2:2], simp1951_0[6:6], simp1951_0[7:7], simp1951_0[8:8]);
  C3 I218 (simp1952_0[3:3], simp1951_0[9:9], simp1951_0[10:10], simp1951_0[11:11]);
  C3 I219 (simp1952_0[4:4], simp1951_0[12:12], simp1951_0[13:13], simp1951_0[14:14]);
  C3 I220 (simp1952_0[5:5], simp1951_0[15:15], simp1951_0[16:16], simp1951_0[17:17]);
  C3 I221 (simp1952_0[6:6], simp1951_0[18:18], simp1951_0[19:19], simp1951_0[20:20]);
  BUFF I222 (simp1952_0[7:7], simp1951_0[21:21]);
  C3 I223 (simp1953_0[0:0], simp1952_0[0:0], simp1952_0[1:1], simp1952_0[2:2]);
  C3 I224 (simp1953_0[1:1], simp1952_0[3:3], simp1952_0[4:4], simp1952_0[5:5]);
  C2 I225 (simp1953_0[2:2], simp1952_0[6:6], simp1952_0[7:7]);
  C3 I226 (i_0a, simp1953_0[0:0], simp1953_0[1:1], simp1953_0[2:2]);
endmodule

// latch tkl2x1 width = 2, depth = 1
module tkl2x1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  wire bna_0;
  wire [1:0] bcomp_0;
  C2R I0 (o_0r0[0:0], i_0r0[0:0], bna_0, reset);
  C2R I1 (o_0r0[1:1], i_0r0[1:1], bna_0, reset);
  C2R I2 (o_0r1[0:0], i_0r1[0:0], bna_0, reset);
  C2R I3 (o_0r1[1:1], i_0r1[1:1], bna_0, reset);
  INV I4 (bna_0, o_0a);
  OR2 I5 (bcomp_0[0:0], o_0r0[0:0], o_0r1[0:0]);
  OR2 I6 (bcomp_0[1:1], o_0r0[1:1], o_0r1[1:1]);
  C2 I7 (i_0a, bcomp_0[0:0], bcomp_0[1:1]);
endmodule

// latch tkl5x1 width = 5, depth = 1
module tkl5x1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [4:0] i_0r0;
  input [4:0] i_0r1;
  output i_0a;
  output [4:0] o_0r0;
  output [4:0] o_0r1;
  input o_0a;
  input reset;
  wire bna_0;
  wire [4:0] bcomp_0;
  wire [1:0] simp181_0;
  C2R I0 (o_0r0[0:0], i_0r0[0:0], bna_0, reset);
  C2R I1 (o_0r0[1:1], i_0r0[1:1], bna_0, reset);
  C2R I2 (o_0r0[2:2], i_0r0[2:2], bna_0, reset);
  C2R I3 (o_0r0[3:3], i_0r0[3:3], bna_0, reset);
  C2R I4 (o_0r0[4:4], i_0r0[4:4], bna_0, reset);
  C2R I5 (o_0r1[0:0], i_0r1[0:0], bna_0, reset);
  C2R I6 (o_0r1[1:1], i_0r1[1:1], bna_0, reset);
  C2R I7 (o_0r1[2:2], i_0r1[2:2], bna_0, reset);
  C2R I8 (o_0r1[3:3], i_0r1[3:3], bna_0, reset);
  C2R I9 (o_0r1[4:4], i_0r1[4:4], bna_0, reset);
  INV I10 (bna_0, o_0a);
  OR2 I11 (bcomp_0[0:0], o_0r0[0:0], o_0r1[0:0]);
  OR2 I12 (bcomp_0[1:1], o_0r0[1:1], o_0r1[1:1]);
  OR2 I13 (bcomp_0[2:2], o_0r0[2:2], o_0r1[2:2]);
  OR2 I14 (bcomp_0[3:3], o_0r0[3:3], o_0r1[3:3]);
  OR2 I15 (bcomp_0[4:4], o_0r0[4:4], o_0r1[4:4]);
  C3 I16 (simp181_0[0:0], bcomp_0[0:0], bcomp_0[1:1], bcomp_0[2:2]);
  C2 I17 (simp181_0[1:1], bcomp_0[3:3], bcomp_0[4:4]);
  C2 I18 (i_0a, simp181_0[0:0], simp181_0[1:1]);
endmodule

// latch tkl34x1 width = 34, depth = 1
module tkl34x1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [33:0] i_0r0;
  input [33:0] i_0r1;
  output i_0a;
  output [33:0] o_0r0;
  output [33:0] o_0r1;
  input o_0a;
  input reset;
  wire bna_0;
  wire [33:0] bcomp_0;
  wire [11:0] simp1051_0;
  wire [3:0] simp1052_0;
  wire [1:0] simp1053_0;
  C2R I0 (o_0r0[0:0], i_0r0[0:0], bna_0, reset);
  C2R I1 (o_0r0[1:1], i_0r0[1:1], bna_0, reset);
  C2R I2 (o_0r0[2:2], i_0r0[2:2], bna_0, reset);
  C2R I3 (o_0r0[3:3], i_0r0[3:3], bna_0, reset);
  C2R I4 (o_0r0[4:4], i_0r0[4:4], bna_0, reset);
  C2R I5 (o_0r0[5:5], i_0r0[5:5], bna_0, reset);
  C2R I6 (o_0r0[6:6], i_0r0[6:6], bna_0, reset);
  C2R I7 (o_0r0[7:7], i_0r0[7:7], bna_0, reset);
  C2R I8 (o_0r0[8:8], i_0r0[8:8], bna_0, reset);
  C2R I9 (o_0r0[9:9], i_0r0[9:9], bna_0, reset);
  C2R I10 (o_0r0[10:10], i_0r0[10:10], bna_0, reset);
  C2R I11 (o_0r0[11:11], i_0r0[11:11], bna_0, reset);
  C2R I12 (o_0r0[12:12], i_0r0[12:12], bna_0, reset);
  C2R I13 (o_0r0[13:13], i_0r0[13:13], bna_0, reset);
  C2R I14 (o_0r0[14:14], i_0r0[14:14], bna_0, reset);
  C2R I15 (o_0r0[15:15], i_0r0[15:15], bna_0, reset);
  C2R I16 (o_0r0[16:16], i_0r0[16:16], bna_0, reset);
  C2R I17 (o_0r0[17:17], i_0r0[17:17], bna_0, reset);
  C2R I18 (o_0r0[18:18], i_0r0[18:18], bna_0, reset);
  C2R I19 (o_0r0[19:19], i_0r0[19:19], bna_0, reset);
  C2R I20 (o_0r0[20:20], i_0r0[20:20], bna_0, reset);
  C2R I21 (o_0r0[21:21], i_0r0[21:21], bna_0, reset);
  C2R I22 (o_0r0[22:22], i_0r0[22:22], bna_0, reset);
  C2R I23 (o_0r0[23:23], i_0r0[23:23], bna_0, reset);
  C2R I24 (o_0r0[24:24], i_0r0[24:24], bna_0, reset);
  C2R I25 (o_0r0[25:25], i_0r0[25:25], bna_0, reset);
  C2R I26 (o_0r0[26:26], i_0r0[26:26], bna_0, reset);
  C2R I27 (o_0r0[27:27], i_0r0[27:27], bna_0, reset);
  C2R I28 (o_0r0[28:28], i_0r0[28:28], bna_0, reset);
  C2R I29 (o_0r0[29:29], i_0r0[29:29], bna_0, reset);
  C2R I30 (o_0r0[30:30], i_0r0[30:30], bna_0, reset);
  C2R I31 (o_0r0[31:31], i_0r0[31:31], bna_0, reset);
  C2R I32 (o_0r0[32:32], i_0r0[32:32], bna_0, reset);
  C2R I33 (o_0r0[33:33], i_0r0[33:33], bna_0, reset);
  C2R I34 (o_0r1[0:0], i_0r1[0:0], bna_0, reset);
  C2R I35 (o_0r1[1:1], i_0r1[1:1], bna_0, reset);
  C2R I36 (o_0r1[2:2], i_0r1[2:2], bna_0, reset);
  C2R I37 (o_0r1[3:3], i_0r1[3:3], bna_0, reset);
  C2R I38 (o_0r1[4:4], i_0r1[4:4], bna_0, reset);
  C2R I39 (o_0r1[5:5], i_0r1[5:5], bna_0, reset);
  C2R I40 (o_0r1[6:6], i_0r1[6:6], bna_0, reset);
  C2R I41 (o_0r1[7:7], i_0r1[7:7], bna_0, reset);
  C2R I42 (o_0r1[8:8], i_0r1[8:8], bna_0, reset);
  C2R I43 (o_0r1[9:9], i_0r1[9:9], bna_0, reset);
  C2R I44 (o_0r1[10:10], i_0r1[10:10], bna_0, reset);
  C2R I45 (o_0r1[11:11], i_0r1[11:11], bna_0, reset);
  C2R I46 (o_0r1[12:12], i_0r1[12:12], bna_0, reset);
  C2R I47 (o_0r1[13:13], i_0r1[13:13], bna_0, reset);
  C2R I48 (o_0r1[14:14], i_0r1[14:14], bna_0, reset);
  C2R I49 (o_0r1[15:15], i_0r1[15:15], bna_0, reset);
  C2R I50 (o_0r1[16:16], i_0r1[16:16], bna_0, reset);
  C2R I51 (o_0r1[17:17], i_0r1[17:17], bna_0, reset);
  C2R I52 (o_0r1[18:18], i_0r1[18:18], bna_0, reset);
  C2R I53 (o_0r1[19:19], i_0r1[19:19], bna_0, reset);
  C2R I54 (o_0r1[20:20], i_0r1[20:20], bna_0, reset);
  C2R I55 (o_0r1[21:21], i_0r1[21:21], bna_0, reset);
  C2R I56 (o_0r1[22:22], i_0r1[22:22], bna_0, reset);
  C2R I57 (o_0r1[23:23], i_0r1[23:23], bna_0, reset);
  C2R I58 (o_0r1[24:24], i_0r1[24:24], bna_0, reset);
  C2R I59 (o_0r1[25:25], i_0r1[25:25], bna_0, reset);
  C2R I60 (o_0r1[26:26], i_0r1[26:26], bna_0, reset);
  C2R I61 (o_0r1[27:27], i_0r1[27:27], bna_0, reset);
  C2R I62 (o_0r1[28:28], i_0r1[28:28], bna_0, reset);
  C2R I63 (o_0r1[29:29], i_0r1[29:29], bna_0, reset);
  C2R I64 (o_0r1[30:30], i_0r1[30:30], bna_0, reset);
  C2R I65 (o_0r1[31:31], i_0r1[31:31], bna_0, reset);
  C2R I66 (o_0r1[32:32], i_0r1[32:32], bna_0, reset);
  C2R I67 (o_0r1[33:33], i_0r1[33:33], bna_0, reset);
  INV I68 (bna_0, o_0a);
  OR2 I69 (bcomp_0[0:0], o_0r0[0:0], o_0r1[0:0]);
  OR2 I70 (bcomp_0[1:1], o_0r0[1:1], o_0r1[1:1]);
  OR2 I71 (bcomp_0[2:2], o_0r0[2:2], o_0r1[2:2]);
  OR2 I72 (bcomp_0[3:3], o_0r0[3:3], o_0r1[3:3]);
  OR2 I73 (bcomp_0[4:4], o_0r0[4:4], o_0r1[4:4]);
  OR2 I74 (bcomp_0[5:5], o_0r0[5:5], o_0r1[5:5]);
  OR2 I75 (bcomp_0[6:6], o_0r0[6:6], o_0r1[6:6]);
  OR2 I76 (bcomp_0[7:7], o_0r0[7:7], o_0r1[7:7]);
  OR2 I77 (bcomp_0[8:8], o_0r0[8:8], o_0r1[8:8]);
  OR2 I78 (bcomp_0[9:9], o_0r0[9:9], o_0r1[9:9]);
  OR2 I79 (bcomp_0[10:10], o_0r0[10:10], o_0r1[10:10]);
  OR2 I80 (bcomp_0[11:11], o_0r0[11:11], o_0r1[11:11]);
  OR2 I81 (bcomp_0[12:12], o_0r0[12:12], o_0r1[12:12]);
  OR2 I82 (bcomp_0[13:13], o_0r0[13:13], o_0r1[13:13]);
  OR2 I83 (bcomp_0[14:14], o_0r0[14:14], o_0r1[14:14]);
  OR2 I84 (bcomp_0[15:15], o_0r0[15:15], o_0r1[15:15]);
  OR2 I85 (bcomp_0[16:16], o_0r0[16:16], o_0r1[16:16]);
  OR2 I86 (bcomp_0[17:17], o_0r0[17:17], o_0r1[17:17]);
  OR2 I87 (bcomp_0[18:18], o_0r0[18:18], o_0r1[18:18]);
  OR2 I88 (bcomp_0[19:19], o_0r0[19:19], o_0r1[19:19]);
  OR2 I89 (bcomp_0[20:20], o_0r0[20:20], o_0r1[20:20]);
  OR2 I90 (bcomp_0[21:21], o_0r0[21:21], o_0r1[21:21]);
  OR2 I91 (bcomp_0[22:22], o_0r0[22:22], o_0r1[22:22]);
  OR2 I92 (bcomp_0[23:23], o_0r0[23:23], o_0r1[23:23]);
  OR2 I93 (bcomp_0[24:24], o_0r0[24:24], o_0r1[24:24]);
  OR2 I94 (bcomp_0[25:25], o_0r0[25:25], o_0r1[25:25]);
  OR2 I95 (bcomp_0[26:26], o_0r0[26:26], o_0r1[26:26]);
  OR2 I96 (bcomp_0[27:27], o_0r0[27:27], o_0r1[27:27]);
  OR2 I97 (bcomp_0[28:28], o_0r0[28:28], o_0r1[28:28]);
  OR2 I98 (bcomp_0[29:29], o_0r0[29:29], o_0r1[29:29]);
  OR2 I99 (bcomp_0[30:30], o_0r0[30:30], o_0r1[30:30]);
  OR2 I100 (bcomp_0[31:31], o_0r0[31:31], o_0r1[31:31]);
  OR2 I101 (bcomp_0[32:32], o_0r0[32:32], o_0r1[32:32]);
  OR2 I102 (bcomp_0[33:33], o_0r0[33:33], o_0r1[33:33]);
  C3 I103 (simp1051_0[0:0], bcomp_0[0:0], bcomp_0[1:1], bcomp_0[2:2]);
  C3 I104 (simp1051_0[1:1], bcomp_0[3:3], bcomp_0[4:4], bcomp_0[5:5]);
  C3 I105 (simp1051_0[2:2], bcomp_0[6:6], bcomp_0[7:7], bcomp_0[8:8]);
  C3 I106 (simp1051_0[3:3], bcomp_0[9:9], bcomp_0[10:10], bcomp_0[11:11]);
  C3 I107 (simp1051_0[4:4], bcomp_0[12:12], bcomp_0[13:13], bcomp_0[14:14]);
  C3 I108 (simp1051_0[5:5], bcomp_0[15:15], bcomp_0[16:16], bcomp_0[17:17]);
  C3 I109 (simp1051_0[6:6], bcomp_0[18:18], bcomp_0[19:19], bcomp_0[20:20]);
  C3 I110 (simp1051_0[7:7], bcomp_0[21:21], bcomp_0[22:22], bcomp_0[23:23]);
  C3 I111 (simp1051_0[8:8], bcomp_0[24:24], bcomp_0[25:25], bcomp_0[26:26]);
  C3 I112 (simp1051_0[9:9], bcomp_0[27:27], bcomp_0[28:28], bcomp_0[29:29]);
  C3 I113 (simp1051_0[10:10], bcomp_0[30:30], bcomp_0[31:31], bcomp_0[32:32]);
  BUFF I114 (simp1051_0[11:11], bcomp_0[33:33]);
  C3 I115 (simp1052_0[0:0], simp1051_0[0:0], simp1051_0[1:1], simp1051_0[2:2]);
  C3 I116 (simp1052_0[1:1], simp1051_0[3:3], simp1051_0[4:4], simp1051_0[5:5]);
  C3 I117 (simp1052_0[2:2], simp1051_0[6:6], simp1051_0[7:7], simp1051_0[8:8]);
  C3 I118 (simp1052_0[3:3], simp1051_0[9:9], simp1051_0[10:10], simp1051_0[11:11]);
  C3 I119 (simp1053_0[0:0], simp1052_0[0:0], simp1052_0[1:1], simp1052_0[2:2]);
  BUFF I120 (simp1053_0[1:1], simp1052_0[3:3]);
  C2 I121 (i_0a, simp1053_0[0:0], simp1053_0[1:1]);
endmodule

module teak_SSEM (go_0r, go_0a, done_0r, done_0a, MemA_0r0, MemA_0r1, MemA_0a, MemRNW_0r0, MemRNW_0r1, MemRNW_0a, MemR_0r0, MemR_0r1, MemR_0a, MemW_0r0, MemW_0r1, MemW_0a, halted_0r, halted_0a, reset);
  input go_0r;
  output go_0a;
  output done_0r;
  input done_0a;
  output [4:0] MemA_0r0;
  output [4:0] MemA_0r1;
  input MemA_0a;
  output MemRNW_0r0;
  output MemRNW_0r1;
  input MemRNW_0a;
  input [31:0] MemR_0r0;
  input [31:0] MemR_0r1;
  output MemR_0a;
  output [31:0] MemW_0r0;
  output [31:0] MemW_0r1;
  input MemW_0a;
  output halted_0r;
  input halted_0a;
  input reset;
  wire L3P_0r;
  wire L3P_0a;
  wire L3A_0r;
  wire L3A_0a;
  wire L5P_0r;
  wire L5P_0a;
  wire L5A_0r;
  wire L5A_0a;
  wire L9P_0r;
  wire L9P_0a;
  wire L9A_0r;
  wire L9A_0a;
  wire L10_0r;
  wire L10_0a;
  wire L12P_0r0;
  wire L12P_0r1;
  wire L12P_0a;
  wire L12A_0r0;
  wire L12A_0r1;
  wire L12A_0a;
  wire L13P_0r;
  wire L13P_0a;
  wire L13A_0r;
  wire L13A_0a;
  wire L14_0r0;
  wire L14_0r1;
  wire L14_0a;
  wire L16P_0r;
  wire L16P_0a;
  wire L16A_0r;
  wire L16A_0a;
  wire L25P_0r;
  wire L25P_0a;
  wire L25A_0r;
  wire L25A_0a;
  wire L29P_0r;
  wire L29P_0a;
  wire L29A_0r;
  wire L29A_0a;
  wire L31P_0r;
  wire L31P_0a;
  wire L31A_0r;
  wire L31A_0a;
  wire [31:0] L32P_0r0;
  wire [31:0] L32P_0r1;
  wire L32P_0a;
  wire [31:0] L32A_0r0;
  wire [31:0] L32A_0r1;
  wire L32A_0a;
  wire L34P_0r;
  wire L34P_0a;
  wire L34A_0r;
  wire L34A_0a;
  wire [2:0] L38P_0r0;
  wire [2:0] L38P_0r1;
  wire L38P_0a;
  wire [2:0] L38A_0r0;
  wire [2:0] L38A_0r1;
  wire L38A_0a;
  wire L42P_0r;
  wire L42P_0a;
  wire L42A_0r;
  wire L42A_0a;
  wire L52P_0r;
  wire L52P_0a;
  wire L52A_0r;
  wire L52A_0a;
  wire L57P_0r;
  wire L57P_0a;
  wire L57A_0r;
  wire L57A_0a;
  wire L60P_0r;
  wire L60P_0a;
  wire L60A_0r;
  wire L60A_0a;
  wire L61_0r0;
  wire L61_0r1;
  wire L61_0a;
  wire L62P_0r;
  wire L62P_0a;
  wire L62A_0r;
  wire L62A_0a;
  wire L63P_0r;
  wire L63P_0a;
  wire L63A_0r;
  wire L63A_0a;
  wire L64P_0r;
  wire L64P_0a;
  wire L64A_0r;
  wire L64A_0a;
  wire L66P_0r;
  wire L66P_0a;
  wire L66A_0r;
  wire L66A_0a;
  wire L69P_0r;
  wire L69P_0a;
  wire L69A_0r;
  wire L69A_0a;
  wire L71P_0r;
  wire L71P_0a;
  wire L71A_0r;
  wire L71A_0a;
  wire L74P_0r;
  wire L74P_0a;
  wire L74A_0r;
  wire L74A_0a;
  wire L76P_0r;
  wire L76P_0a;
  wire L76A_0r;
  wire L76A_0a;
  wire L78P_0r;
  wire L78P_0a;
  wire L78A_0r;
  wire L78A_0a;
  wire L79_0r;
  wire L79_0a;
  wire L86P_0r;
  wire L86P_0a;
  wire L86A_0r;
  wire L86A_0a;
  wire L96P_0r;
  wire L96P_0a;
  wire L96A_0r;
  wire L96A_0a;
  wire [4:0] L97_0r0;
  wire [4:0] L97_0r1;
  wire L97_0a;
  wire L98P_0r;
  wire L98P_0a;
  wire L98A_0r;
  wire L98A_0a;
  wire [4:0] L99_0r0;
  wire [4:0] L99_0r1;
  wire L99_0a;
  wire [9:0] L100P_0r0;
  wire [9:0] L100P_0r1;
  wire L100P_0a;
  wire [9:0] L100A_0r0;
  wire [9:0] L100A_0r1;
  wire L100A_0a;
  wire [5:0] L101P_0r0;
  wire [5:0] L101P_0r1;
  wire L101P_0a;
  wire [5:0] L101A_0r0;
  wire [5:0] L101A_0r1;
  wire L101A_0a;
  wire L102P_0r;
  wire L102P_0a;
  wire L102A_0r;
  wire L102A_0a;
  wire L104P_0r;
  wire L104P_0a;
  wire L104A_0r;
  wire L104A_0a;
  wire L107P_0r;
  wire L107P_0a;
  wire L107A_0r;
  wire L107A_0a;
  wire L108P_0r;
  wire L108P_0a;
  wire L108A_0r;
  wire L108A_0a;
  wire [2:0] L112P_0r0;
  wire [2:0] L112P_0r1;
  wire L112P_0a;
  wire [2:0] L112A_0r0;
  wire [2:0] L112A_0r1;
  wire L112A_0a;
  wire [2:0] L113P_0r0;
  wire [2:0] L113P_0r1;
  wire L113P_0a;
  wire [2:0] L113A_0r0;
  wire [2:0] L113A_0r1;
  wire L113A_0a;
  wire [2:0] L114P_0r0;
  wire [2:0] L114P_0r1;
  wire L114P_0a;
  wire [2:0] L114A_0r0;
  wire [2:0] L114A_0r1;
  wire L114A_0a;
  wire [2:0] L115P_0r0;
  wire [2:0] L115P_0r1;
  wire L115P_0a;
  wire [2:0] L115A_0r0;
  wire [2:0] L115A_0r1;
  wire L115A_0a;
  wire L120P_0r;
  wire L120P_0a;
  wire L120A_0r;
  wire L120A_0a;
  wire [31:0] L121_0r0;
  wire [31:0] L121_0r1;
  wire L121_0a;
  wire L122P_0r;
  wire L122P_0a;
  wire L122A_0r;
  wire L122A_0a;
  wire [31:0] L123_0r0;
  wire [31:0] L123_0r1;
  wire L123_0a;
  wire [63:0] L124P_0r0;
  wire [63:0] L124P_0r1;
  wire L124P_0a;
  wire [63:0] L124A_0r0;
  wire [63:0] L124A_0r1;
  wire L124A_0a;
  wire L126P_0r;
  wire L126P_0a;
  wire L126A_0r;
  wire L126A_0a;
  wire [31:0] L127P_0r0;
  wire [31:0] L127P_0r1;
  wire L127P_0a;
  wire [31:0] L127A_0r0;
  wire [31:0] L127A_0r1;
  wire L127A_0a;
  wire L128_0r;
  wire L128_0a;
  wire L137P_0r;
  wire L137P_0a;
  wire L137A_0r;
  wire L137A_0a;
  wire L140P_0r;
  wire L140P_0a;
  wire L140A_0r;
  wire L140A_0a;
  wire L141P_0r;
  wire L141P_0a;
  wire L141A_0r;
  wire L141A_0a;
  wire L142P_0r;
  wire L142P_0a;
  wire L142A_0r;
  wire L142A_0a;
  wire L143P_0r;
  wire L143P_0a;
  wire L143A_0r;
  wire L143A_0a;
  wire L144P_0r;
  wire L144P_0a;
  wire L144A_0r;
  wire L144A_0a;
  wire [1:0] L145P_0r0;
  wire [1:0] L145P_0r1;
  wire L145P_0a;
  wire [1:0] L145A_0r0;
  wire [1:0] L145A_0r1;
  wire L145A_0a;
  wire [1:0] L146P_0r0;
  wire [1:0] L146P_0r1;
  wire L146P_0a;
  wire [1:0] L146A_0r0;
  wire [1:0] L146A_0r1;
  wire L146A_0a;
  wire [1:0] L147P_0r0;
  wire [1:0] L147P_0r1;
  wire L147P_0a;
  wire [1:0] L147A_0r0;
  wire [1:0] L147A_0r1;
  wire L147A_0a;
  wire [1:0] L148P_0r0;
  wire [1:0] L148P_0r1;
  wire L148P_0a;
  wire [1:0] L148A_0r0;
  wire [1:0] L148A_0r1;
  wire L148A_0a;
  wire L149P_0r;
  wire L149P_0a;
  wire L149A_0r;
  wire L149A_0a;
  wire L152P_0r;
  wire L152P_0a;
  wire L152A_0r;
  wire L152A_0a;
  wire L153P_0r;
  wire L153P_0a;
  wire L153A_0r;
  wire L153A_0a;
  wire L154P_0r;
  wire L154P_0a;
  wire L154A_0r;
  wire L154A_0a;
  wire L155P_0r;
  wire L155P_0a;
  wire L155A_0r;
  wire L155A_0a;
  wire L156P_0r;
  wire L156P_0a;
  wire L156A_0r;
  wire L156A_0a;
  wire [1:0] L157P_0r0;
  wire [1:0] L157P_0r1;
  wire L157P_0a;
  wire [1:0] L157A_0r0;
  wire [1:0] L157A_0r1;
  wire L157A_0a;
  wire [1:0] L158P_0r0;
  wire [1:0] L158P_0r1;
  wire L158P_0a;
  wire [1:0] L158A_0r0;
  wire [1:0] L158A_0r1;
  wire L158A_0a;
  wire [1:0] L159P_0r0;
  wire [1:0] L159P_0r1;
  wire L159P_0a;
  wire [1:0] L159A_0r0;
  wire [1:0] L159A_0r1;
  wire L159A_0a;
  wire [1:0] L160P_0r0;
  wire [1:0] L160P_0r1;
  wire L160P_0a;
  wire [1:0] L160A_0r0;
  wire [1:0] L160A_0r1;
  wire L160A_0a;
  wire L164P_0r;
  wire L164P_0a;
  wire L164A_0r;
  wire L164A_0a;
  wire L166P_0r;
  wire L166P_0a;
  wire L166A_0r;
  wire L166A_0a;
  wire L168P_0r;
  wire L168P_0a;
  wire L168A_0r;
  wire L168A_0a;
  wire [31:0] L169P_0r0;
  wire [31:0] L169P_0r1;
  wire L169P_0a;
  wire [31:0] L169A_0r0;
  wire [31:0] L169A_0r1;
  wire L169A_0a;
  wire L170_0r;
  wire L170_0a;
  wire L171P_0r;
  wire L171P_0a;
  wire L171A_0r;
  wire L171A_0a;
  wire L177P_0r;
  wire L177P_0a;
  wire L177A_0r;
  wire L177A_0a;
  wire L178P_0r;
  wire L178P_0a;
  wire L178A_0r;
  wire L178A_0a;
  wire [2:0] L179P_0r0;
  wire [2:0] L179P_0r1;
  wire L179P_0a;
  wire [2:0] L179A_0r0;
  wire [2:0] L179A_0r1;
  wire L179A_0a;
  wire [2:0] L181P_0r0;
  wire [2:0] L181P_0r1;
  wire L181P_0a;
  wire [2:0] L181A_0r0;
  wire [2:0] L181A_0r1;
  wire L181A_0a;
  wire [2:0] L182P_0r0;
  wire [2:0] L182P_0r1;
  wire L182P_0a;
  wire [2:0] L182A_0r0;
  wire [2:0] L182A_0r1;
  wire L182A_0a;
  wire [2:0] L183P_0r0;
  wire [2:0] L183P_0r1;
  wire L183P_0a;
  wire [2:0] L183A_0r0;
  wire [2:0] L183A_0r1;
  wire L183A_0a;
  wire L187P_0r;
  wire L187P_0a;
  wire L187A_0r;
  wire L187A_0a;
  wire L189P_0r;
  wire L189P_0a;
  wire L189A_0r;
  wire L189A_0a;
  wire L193P_0r;
  wire L193P_0a;
  wire L193A_0r;
  wire L193A_0a;
  wire L194P_0r;
  wire L194P_0a;
  wire L194A_0r;
  wire L194A_0a;
  wire L196P_0r;
  wire L196P_0a;
  wire L196A_0r;
  wire L196A_0a;
  wire L199P_0r;
  wire L199P_0a;
  wire L199A_0r;
  wire L199A_0a;
  wire L200P_0r;
  wire L200P_0a;
  wire L200A_0r;
  wire L200A_0a;
  wire L201P_0r;
  wire L201P_0a;
  wire L201A_0r;
  wire L201A_0a;
  wire L202P_0r;
  wire L202P_0a;
  wire L202A_0r;
  wire L202A_0a;
  wire L203P_0r;
  wire L203P_0a;
  wire L203A_0r;
  wire L203A_0a;
  wire [1:0] L204P_0r0;
  wire [1:0] L204P_0r1;
  wire L204P_0a;
  wire [1:0] L204A_0r0;
  wire [1:0] L204A_0r1;
  wire L204A_0a;
  wire [1:0] L205P_0r0;
  wire [1:0] L205P_0r1;
  wire L205P_0a;
  wire [1:0] L205A_0r0;
  wire [1:0] L205A_0r1;
  wire L205A_0a;
  wire [1:0] L206P_0r0;
  wire [1:0] L206P_0r1;
  wire L206P_0a;
  wire [1:0] L206A_0r0;
  wire [1:0] L206A_0r1;
  wire L206A_0a;
  wire [1:0] L207P_0r0;
  wire [1:0] L207P_0r1;
  wire L207P_0a;
  wire [1:0] L207A_0r0;
  wire [1:0] L207A_0r1;
  wire L207A_0a;
  wire L208P_0r0;
  wire L208P_0r1;
  wire L208P_0a;
  wire L208A_0r0;
  wire L208A_0r1;
  wire L208A_0a;
  wire L209_0r;
  wire L209_0a;
  wire L210P_0r;
  wire L210P_0a;
  wire L210A_0r;
  wire L210A_0a;
  wire L211P_0r0;
  wire L211P_0r1;
  wire L211P_0a;
  wire L211A_0r0;
  wire L211A_0r1;
  wire L211A_0a;
  wire L212P_0r;
  wire L212P_0a;
  wire L212A_0r;
  wire L212A_0a;
  wire L213P_0r0;
  wire L213P_0r1;
  wire L213P_0a;
  wire L213A_0r0;
  wire L213A_0r1;
  wire L213A_0a;
  wire [1:0] L214P_0r0;
  wire [1:0] L214P_0r1;
  wire L214P_0a;
  wire [1:0] L214A_0r0;
  wire [1:0] L214A_0r1;
  wire L214A_0a;
  wire [1:0] L215P_0r0;
  wire [1:0] L215P_0r1;
  wire L215P_0a;
  wire [1:0] L215A_0r0;
  wire [1:0] L215A_0r1;
  wire L215A_0a;
  wire [1:0] L216P_0r0;
  wire [1:0] L216P_0r1;
  wire L216P_0a;
  wire [1:0] L216A_0r0;
  wire [1:0] L216A_0r1;
  wire L216A_0a;
  wire [1:0] L217P_0r0;
  wire [1:0] L217P_0r1;
  wire L217P_0a;
  wire [1:0] L217A_0r0;
  wire [1:0] L217A_0r1;
  wire L217A_0a;
  wire [4:0] L218P_0r0;
  wire [4:0] L218P_0r1;
  wire L218P_0a;
  wire [4:0] L218A_0r0;
  wire [4:0] L218A_0r1;
  wire L218A_0a;
  wire L219_0r;
  wire L219_0a;
  wire L220P_0r;
  wire L220P_0a;
  wire L220A_0r;
  wire L220A_0a;
  wire [4:0] L221_0r0;
  wire [4:0] L221_0r1;
  wire L221_0a;
  wire L222P_0r;
  wire L222P_0a;
  wire L222A_0r;
  wire L222A_0a;
  wire [4:0] L223P_0r0;
  wire [4:0] L223P_0r1;
  wire L223P_0a;
  wire [4:0] L223A_0r0;
  wire [4:0] L223A_0r1;
  wire L223A_0a;
  wire [1:0] L224P_0r0;
  wire [1:0] L224P_0r1;
  wire L224P_0a;
  wire [1:0] L224A_0r0;
  wire [1:0] L224A_0r1;
  wire L224A_0a;
  wire [1:0] L225P_0r0;
  wire [1:0] L225P_0r1;
  wire L225P_0a;
  wire [1:0] L225A_0r0;
  wire [1:0] L225A_0r1;
  wire L225A_0a;
  wire [1:0] L226P_0r0;
  wire [1:0] L226P_0r1;
  wire L226P_0a;
  wire [1:0] L226A_0r0;
  wire [1:0] L226A_0r1;
  wire L226A_0a;
  wire [4:0] L228P_0r0;
  wire [4:0] L228P_0r1;
  wire L228P_0a;
  wire [4:0] L228A_0r0;
  wire [4:0] L228A_0r1;
  wire L228A_0a;
  wire L229_0r;
  wire L229_0a;
  wire L230P_0r;
  wire L230P_0a;
  wire L230A_0r;
  wire L230A_0a;
  wire [4:0] L231P_0r0;
  wire [4:0] L231P_0r1;
  wire L231P_0a;
  wire [4:0] L231A_0r0;
  wire [4:0] L231A_0r1;
  wire L231A_0a;
  wire L232P_0r;
  wire L232P_0a;
  wire L232A_0r;
  wire L232A_0a;
  wire [4:0] L233P_0r0;
  wire [4:0] L233P_0r1;
  wire L233P_0a;
  wire [4:0] L233A_0r0;
  wire [4:0] L233A_0r1;
  wire L233A_0a;
  wire [1:0] L234P_0r0;
  wire [1:0] L234P_0r1;
  wire L234P_0a;
  wire [1:0] L234A_0r0;
  wire [1:0] L234A_0r1;
  wire L234A_0a;
  wire [1:0] L235P_0r0;
  wire [1:0] L235P_0r1;
  wire L235P_0a;
  wire [1:0] L235A_0r0;
  wire [1:0] L235A_0r1;
  wire L235A_0a;
  wire [1:0] L236P_0r0;
  wire [1:0] L236P_0r1;
  wire L236P_0a;
  wire [1:0] L236A_0r0;
  wire [1:0] L236A_0r1;
  wire L236A_0a;
  wire [1:0] L237P_0r0;
  wire [1:0] L237P_0r1;
  wire L237P_0a;
  wire [1:0] L237A_0r0;
  wire [1:0] L237A_0r1;
  wire L237A_0a;
  wire [31:0] L238P_0r0;
  wire [31:0] L238P_0r1;
  wire L238P_0a;
  wire [31:0] L238A_0r0;
  wire [31:0] L238A_0r1;
  wire L238A_0a;
  wire L239_0r;
  wire L239_0a;
  wire L240P_0r;
  wire L240P_0a;
  wire L240A_0r;
  wire L240A_0a;
  wire [31:0] L241P_0r0;
  wire [31:0] L241P_0r1;
  wire L241P_0a;
  wire [31:0] L241A_0r0;
  wire [31:0] L241A_0r1;
  wire L241A_0a;
  wire L242P_0r;
  wire L242P_0a;
  wire L242A_0r;
  wire L242A_0a;
  wire [31:0] L243_0r0;
  wire [31:0] L243_0r1;
  wire L243_0a;
  wire [1:0] L244P_0r0;
  wire [1:0] L244P_0r1;
  wire L244P_0a;
  wire [1:0] L244A_0r0;
  wire [1:0] L244A_0r1;
  wire L244A_0a;
  wire [1:0] L245P_0r0;
  wire [1:0] L245P_0r1;
  wire L245P_0a;
  wire [1:0] L245A_0r0;
  wire [1:0] L245A_0r1;
  wire L245A_0a;
  wire [1:0] L246P_0r0;
  wire [1:0] L246P_0r1;
  wire L246P_0a;
  wire [1:0] L246A_0r0;
  wire [1:0] L246A_0r1;
  wire L246A_0a;
  wire [1:0] L247P_0r0;
  wire [1:0] L247P_0r1;
  wire L247P_0a;
  wire [1:0] L247A_0r0;
  wire [1:0] L247A_0r1;
  wire L247A_0a;
  wire L248P_0r;
  wire L248P_0a;
  wire L248A_0r;
  wire L248A_0a;
  wire [4:0] L249_0r0;
  wire [4:0] L249_0r1;
  wire L249_0a;
  wire L250P_0r;
  wire L250P_0a;
  wire L250A_0r;
  wire L250A_0a;
  wire [4:0] L251_0r0;
  wire [4:0] L251_0r1;
  wire L251_0a;
  wire [4:0] L252P_0r0;
  wire [4:0] L252P_0r1;
  wire L252P_0a;
  wire [4:0] L252A_0r0;
  wire [4:0] L252A_0r1;
  wire L252A_0a;
  wire L253P_0r;
  wire L253P_0a;
  wire L253A_0r;
  wire L253A_0a;
  wire [4:0] L254_0r0;
  wire [4:0] L254_0r1;
  wire L254_0a;
  wire [1:0] L255P_0r0;
  wire [1:0] L255P_0r1;
  wire L255P_0a;
  wire [1:0] L255A_0r0;
  wire [1:0] L255A_0r1;
  wire L255A_0a;
  wire [1:0] L256P_0r0;
  wire [1:0] L256P_0r1;
  wire L256P_0a;
  wire [1:0] L256A_0r0;
  wire [1:0] L256A_0r1;
  wire L256A_0a;
  wire [1:0] L257P_0r0;
  wire [1:0] L257P_0r1;
  wire L257P_0a;
  wire [1:0] L257A_0r0;
  wire [1:0] L257A_0r1;
  wire L257A_0a;
  wire [1:0] L258P_0r0;
  wire [1:0] L258P_0r1;
  wire L258P_0a;
  wire [1:0] L258A_0r0;
  wire [1:0] L258A_0r1;
  wire L258A_0a;
  wire L259P_0r;
  wire L259P_0a;
  wire L259A_0r;
  wire L259A_0a;
  wire L260P_0r0;
  wire L260P_0r1;
  wire L260P_0a;
  wire L260A_0r0;
  wire L260A_0r1;
  wire L260A_0a;
  wire L261P_0r;
  wire L261P_0a;
  wire L261A_0r;
  wire L261A_0a;
  wire L262P_0r0;
  wire L262P_0r1;
  wire L262P_0a;
  wire L262A_0r0;
  wire L262A_0r1;
  wire L262A_0a;
  wire L263P_0r;
  wire L263P_0a;
  wire L263A_0r;
  wire L263A_0a;
  wire L264P_0r0;
  wire L264P_0r1;
  wire L264P_0a;
  wire L264A_0r0;
  wire L264A_0r1;
  wire L264A_0a;
  wire L265P_0r0;
  wire L265P_0r1;
  wire L265P_0a;
  wire L265A_0r0;
  wire L265A_0r1;
  wire L265A_0a;
  wire L266P_0r;
  wire L266P_0a;
  wire L266A_0r;
  wire L266A_0a;
  wire L267_0r0;
  wire L267_0r1;
  wire L267_0a;
  wire [2:0] L268P_0r0;
  wire [2:0] L268P_0r1;
  wire L268P_0a;
  wire [2:0] L268A_0r0;
  wire [2:0] L268A_0r1;
  wire L268A_0a;
  wire [2:0] L269P_0r0;
  wire [2:0] L269P_0r1;
  wire L269P_0a;
  wire [2:0] L269A_0r0;
  wire [2:0] L269A_0r1;
  wire L269A_0a;
  wire [2:0] L270P_0r0;
  wire [2:0] L270P_0r1;
  wire L270P_0a;
  wire [2:0] L270A_0r0;
  wire [2:0] L270A_0r1;
  wire L270A_0a;
  wire [2:0] L271P_0r0;
  wire [2:0] L271P_0r1;
  wire L271P_0a;
  wire [2:0] L271A_0r0;
  wire [2:0] L271A_0r1;
  wire L271A_0a;
  wire [2:0] L272P_0r0;
  wire [2:0] L272P_0r1;
  wire L272P_0a;
  wire [2:0] L272A_0r0;
  wire [2:0] L272A_0r1;
  wire L272A_0a;
  wire [31:0] L273_0r0;
  wire [31:0] L273_0r1;
  wire L273_0a;
  wire [1:0] L274P_0r0;
  wire [1:0] L274P_0r1;
  wire L274P_0a;
  wire [1:0] L274A_0r0;
  wire [1:0] L274A_0r1;
  wire L274A_0a;
  wire [1:0] L275P_0r0;
  wire [1:0] L275P_0r1;
  wire L275P_0a;
  wire [1:0] L275A_0r0;
  wire [1:0] L275A_0r1;
  wire L275A_0a;
  wire [1:0] L276P_0r0;
  wire [1:0] L276P_0r1;
  wire L276P_0a;
  wire [1:0] L276A_0r0;
  wire [1:0] L276A_0r1;
  wire L276A_0a;
  wire [33:0] L277P_0r0;
  wire [33:0] L277P_0r1;
  wire L277P_0a;
  wire [33:0] L277A_0r0;
  wire [33:0] L277A_0r1;
  wire L277A_0a;
  wire L279_0r;
  wire L279_0a;
  wire L280P_0r;
  wire L280P_0a;
  wire L280A_0r;
  wire L280A_0a;
  wire L281P_0r;
  wire L281P_0a;
  wire L281A_0r;
  wire L281A_0a;
  wire L283_0r;
  wire L283_0a;
  wire [31:0] L284P_0r0;
  wire [31:0] L284P_0r1;
  wire L284P_0a;
  wire [31:0] L284A_0r0;
  wire [31:0] L284A_0r1;
  wire L284A_0a;
  wire [2:0] L285P_0r0;
  wire [2:0] L285P_0r1;
  wire L285P_0a;
  wire [2:0] L285A_0r0;
  wire [2:0] L285A_0r1;
  wire L285A_0a;
  wire L286P_0r;
  wire L286P_0a;
  wire L286A_0r;
  wire L286A_0a;
  wire L287P_0r;
  wire L287P_0a;
  wire L287A_0r;
  wire L287A_0a;
  wire L288P_0r;
  wire L288P_0a;
  wire L288A_0r;
  wire L288A_0a;
  wire L289P_0r;
  wire L289P_0a;
  wire L289A_0r;
  wire L289A_0a;
  wire L290P_0r;
  wire L290P_0a;
  wire L290A_0r;
  wire L290A_0a;
  wire L291P_0r;
  wire L291P_0a;
  wire L291A_0r;
  wire L291A_0a;
  wire L292P_0r;
  wire L292P_0a;
  wire L292A_0r;
  wire L292A_0a;
  wire L293P_0r;
  wire L293P_0a;
  wire L293A_0r;
  wire L293A_0a;
  wire L294P_0r;
  wire L294P_0a;
  wire L294A_0r;
  wire L294A_0a;
  wire L295P_0r;
  wire L295P_0a;
  wire L295A_0r;
  wire L295A_0a;
  wire L296P_0r;
  wire L296P_0a;
  wire L296A_0r;
  wire L296A_0a;
  wire L297P_0r;
  wire L297P_0a;
  wire L297A_0r;
  wire L297A_0a;
  wire L298P_0r;
  wire L298P_0a;
  wire L298A_0r;
  wire L298A_0a;
  wire [2:0] L299P_0r0;
  wire [2:0] L299P_0r1;
  wire L299P_0a;
  wire [2:0] L299A_0r0;
  wire [2:0] L299A_0r1;
  wire L299A_0a;
  wire L301P_0r;
  wire L301P_0a;
  wire L301A_0r;
  wire L301A_0a;
  wire [1:0] L302P_0r0;
  wire [1:0] L302P_0r1;
  wire L302P_0a;
  wire [1:0] L302A_0r0;
  wire [1:0] L302A_0r1;
  wire L302A_0a;
  wire L304P_0r;
  wire L304P_0a;
  wire L304A_0r;
  wire L304A_0a;
  wire L306P_0r;
  wire L306P_0a;
  wire L306A_0r;
  wire L306A_0a;
  wire L308P_0r;
  wire L308P_0a;
  wire L308A_0r;
  wire L308A_0a;
  wire [2:0] L309P_0r0;
  wire [2:0] L309P_0r1;
  wire L309P_0a;
  wire [2:0] L309A_0r0;
  wire [2:0] L309A_0r1;
  wire L309A_0a;
  wire [1:0] L310P_0r0;
  wire [1:0] L310P_0r1;
  wire L310P_0a;
  wire [1:0] L310A_0r0;
  wire [1:0] L310A_0r1;
  wire L310A_0a;
  wire L311P_0r;
  wire L311P_0a;
  wire L311A_0r;
  wire L311A_0a;
  wire L312P_0r;
  wire L312P_0a;
  wire L312A_0r;
  wire L312A_0a;
  wire L313P_0r;
  wire L313P_0a;
  wire L313A_0r;
  wire L313A_0a;
  wire L314P_0r;
  wire L314P_0a;
  wire L314A_0r;
  wire L314A_0a;
  wire L315P_0r;
  wire L315P_0a;
  wire L315A_0r;
  wire L315A_0a;
  wire L318P_0r;
  wire L318P_0a;
  wire L318A_0r;
  wire L318A_0a;
  tko0m1_1nm1b0 I0 (L286P_0r, L286P_0a, L213A_0r0, L213A_0r1, L213A_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0 I1 (L10_0r, L10_0a, L153A_0r, L153A_0a, L154A_0r, L154A_0a, L141A_0r, L141A_0a, L142A_0r, L142A_0a, L212A_0r, L212A_0a, L286A_0r, L286A_0a, reset);
  tkj0m0_0_0 I2 (L3P_0r, L3P_0a, L5P_0r, L5P_0a, L9P_0r, L9P_0a, L76A_0r, L76A_0a, reset);
  tko1m1_1noti0w1b I3 (L14_0r0, L14_0r1, L14_0a, L12A_0r0, L12A_0r1, L12A_0a, reset);
  tko0m5_1nm5b1 I4 (L287P_0r, L287P_0a, L223A_0r0[4:0], L223A_0r1[4:0], L223A_0a, reset);
  tko0m1_1nm1b1 I5 (L288P_0r, L288P_0a, L260A_0r0, L260A_0r1, L260A_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0_o0w0 I6 (L34P_0r, L34P_0a, L259A_0r, L259A_0a, L288A_0r, L288A_0a, L296A_0r, L296A_0a, L248A_0r, L248A_0a, L31A_0r, L31A_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I7 (L61_0r0, L61_0r1, L61_0a, L62A_0r, L62A_0a, L63A_0r, L63A_0a, reset);
  tko0m1_1nm1b1 I8 (L289P_0r, L289P_0a, L211A_0r0, L211A_0r1, L211A_0a, reset);
  tks3_o0w3_2o0w0_3o0w0_4c1o0w0_6o0w0_7o0w0_0m1o0w3 I9 (L38P_0r0[2:0], L38P_0r1[2:0], L38P_0a, L52A_0r, L52A_0a, L194A_0r, L194A_0a, L314A_0r, L314A_0a, L60A_0r, L60A_0a, L66A_0r, L66A_0a, L299A_0r0[2:0], L299A_0r1[2:0], L299A_0a, reset);
  tkm6x0b I10 (L281P_0r, L281P_0a, L280P_0r, L280P_0a, L57P_0r, L57P_0a, L62P_0r, L62P_0a, L64P_0r, L64P_0a, L69P_0r, L69P_0a, L71A_0r, L71A_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I11 (L12P_0r0, L12P_0r1, L12P_0a, L78A_0r, L78A_0a, L16A_0r, L16A_0a, reset);
  tkm2x0b I12 (L76P_0r, L76P_0a, L74P_0r, L74P_0a, L13A_0r, L13A_0a, reset);
  tkj0m0_0 I13 (L86P_0r, L86P_0a, L306P_0r, L306P_0a, L280A_0r, L280A_0a, reset);
  tkj10m5_5 I14 (L97_0r0[4:0], L97_0r1[4:0], L97_0a, L99_0r0[4:0], L99_0r1[4:0], L99_0a, L100A_0r0[9:0], L100A_0r1[9:0], L100A_0a, reset);
  tko10m6_1nm1b0_2api0w5bt1o0w1b_3nm1b0_4api5w5bt3o0w1b_5addt2o0w6bt4o0w6b I15 (L100P_0r0[9:0], L100P_0r1[9:0], L100P_0a, L101A_0r0[5:0], L101A_0r1[5:0], L101A_0a, reset);
  tkf6mo0w0_o0w5 I16 (L101P_0r0[5:0], L101P_0r1[5:0], L101P_0a, L232A_0r, L232A_0a, L233A_0r0[4:0], L233A_0r1[4:0], L233A_0a, reset);
  tkf0mo0w0_o0w0 I17 (L102P_0r, L102P_0a, L96A_0r, L96A_0a, L98A_0r, L98A_0a, reset);
  tkf0mo0w0_o0w0 I18 (L63P_0r, L63P_0a, L107A_0r, L107A_0a, L108A_0r, L108A_0a, reset);
  tkm2x0b I19 (L107P_0r, L107P_0a, L304P_0r, L304P_0a, L102A_0r, L102A_0a, reset);
  tko0m3_1nm3b2 I20 (L108P_0r, L108P_0a, L112A_0r0[2:0], L112A_0r1[2:0], L112A_0a, reset);
  tkm2x3b I21 (L113P_0r0[2:0], L113P_0r1[2:0], L113P_0a, L112P_0r0[2:0], L112P_0r1[2:0], L112P_0a, L114A_0r0[2:0], L114A_0r1[2:0], L114A_0a, reset);
  tkj3m0_3 I22 (L104P_0r, L104P_0a, L114P_0r0[2:0], L114P_0r1[2:0], L114P_0a, L115A_0r0[2:0], L115A_0r1[2:0], L115A_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_4o0w0 I23 (L115P_0r0[2:0], L115P_0r1[2:0], L115P_0a, L34A_0r, L34A_0a, L64A_0r, L64A_0a, L86A_0r, L86A_0a, reset);
  tkj64m32_32 I24 (L121_0r0[31:0], L121_0r1[31:0], L121_0a, L123_0r0[31:0], L123_0r1[31:0], L123_0a, L124A_0r0[63:0], L124A_0r1[63:0], L124A_0a, reset);
  tkf0mo0w0_o0w0 I25 (L126P_0r, L126P_0a, L120A_0r, L120A_0a, L122A_0r, L122A_0a, reset);
  tkj0m0_0 I26 (L128_0r, L128_0a, L308P_0r, L308P_0a, L281A_0r, L281A_0a, reset);
  tko0m5_1nm5b0 I27 (L290P_0r, L290P_0a, L231A_0r0[4:0], L231A_0r1[4:0], L231A_0a, reset);
  tkf0mo0w0_o0w0 I28 (L42P_0r, L42P_0a, L143A_0r, L143A_0a, L144A_0r, L144A_0a, reset);
  tkm2x0b I29 (L141P_0r, L141P_0a, L143P_0r, L143P_0a, L137A_0r, L137A_0a, reset);
  tko0m2_1nm2b1 I30 (L142P_0r, L142P_0a, L145A_0r0[1:0], L145A_0r1[1:0], L145A_0a, reset);
  tko0m2_1nm2b2 I31 (L144P_0r, L144P_0a, L146A_0r0[1:0], L146A_0r1[1:0], L146A_0a, reset);
  tkm2x2b I32 (L145P_0r0[1:0], L145P_0r1[1:0], L145P_0a, L146P_0r0[1:0], L146P_0r1[1:0], L146P_0a, L147A_0r0[1:0], L147A_0r1[1:0], L147A_0a, reset);
  tkj2m0_2 I33 (L140P_0r, L140P_0a, L147P_0r0[1:0], L147P_0r1[1:0], L147P_0a, L148A_0r0[1:0], L148A_0r1[1:0], L148A_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I34 (L148P_0r0[1:0], L148P_0r1[1:0], L148P_0a, L5A_0r, L5A_0a, L311A_0r, L311A_0a, reset);
  tko0m32_1nm32b0 I35 (L291P_0r, L291P_0a, L241A_0r0[31:0], L241A_0r1[31:0], L241A_0a, reset);
  tkf0mo0w0_o0w0 I36 (L52P_0r, L52P_0a, L155A_0r, L155A_0a, L156A_0r, L156A_0a, reset);
  tkm2x0b I37 (L153P_0r, L153P_0a, L155P_0r, L155P_0a, L149A_0r, L149A_0a, reset);
  tko0m2_1nm2b1 I38 (L154P_0r, L154P_0a, L157A_0r0[1:0], L157A_0r1[1:0], L157A_0a, reset);
  tko0m2_1nm2b2 I39 (L156P_0r, L156P_0a, L158A_0r0[1:0], L158A_0r1[1:0], L158A_0a, reset);
  tkm2x2b I40 (L157P_0r0[1:0], L157P_0r1[1:0], L157P_0a, L158P_0r0[1:0], L158P_0r1[1:0], L158P_0a, L159A_0r0[1:0], L159A_0r1[1:0], L159A_0a, reset);
  tkj2m0_2 I41 (L152P_0r, L152P_0a, L159P_0r0[1:0], L159P_0r1[1:0], L159P_0a, L160A_0r0[1:0], L160A_0r1[1:0], L160A_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I42 (L160P_0r0[1:0], L160P_0r1[1:0], L160P_0a, L3A_0r, L3A_0a, L313A_0r, L313A_0a, reset);
  tko0m1_1nm1b1 I43 (L292P_0r, L292P_0a, L262A_0r0, L262A_0r1, L262A_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0_o0w0 I44 (L171P_0r, L171P_0a, L261A_0r, L261A_0a, L292A_0r, L292A_0a, L200A_0r, L200A_0a, L201A_0r, L201A_0a, L168A_0r, L168A_0a, reset);
  tkm2x0b I45 (L177P_0r, L177P_0a, L301P_0r, L301P_0a, L171A_0r, L171A_0a, reset);
  tko0m3_1nm3b4 I46 (L178P_0r, L178P_0a, L181A_0r0[2:0], L181A_0r1[2:0], L181A_0a, reset);
  tkm2x3b I47 (L179P_0r0[2:0], L179P_0r1[2:0], L179P_0a, L181P_0r0[2:0], L181P_0r1[2:0], L181P_0a, L182A_0r0[2:0], L182A_0r1[2:0], L182A_0a, reset);
  tkj3m0_0_0_3 I48 (L164P_0r, L164P_0a, L166P_0r, L166P_0a, L170_0r, L170_0a, L182P_0r0[2:0], L182P_0r1[2:0], L182P_0a, L183A_0r0[2:0], L183A_0r1[2:0], L183A_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_4o0w0 I49 (L183P_0r0[2:0], L183P_0r1[2:0], L183P_0a, L42A_0r, L42A_0a, L312A_0r, L312A_0a, L126A_0r, L126A_0a, reset);
  tko0m1_1nm1b0 I50 (L293P_0r, L293P_0a, L264A_0r0, L264A_0r1, L264A_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0 I51 (L194P_0r, L194P_0a, L263A_0r, L263A_0a, L293A_0r, L293A_0a, L202A_0r, L202A_0a, L203A_0r, L203A_0a, L298A_0r, L298A_0a, L193A_0r, L193A_0a, reset);
  tkj0m0_0_0 I52 (L187P_0r, L187P_0a, L189P_0r, L189P_0a, L193P_0r, L193P_0a, L57A_0r, L57A_0a, reset);
  tkm2x0b I53 (L200P_0r, L200P_0a, L202P_0r, L202P_0a, L196A_0r, L196A_0a, reset);
  tko0m2_1nm2b1 I54 (L201P_0r, L201P_0a, L204A_0r0[1:0], L204A_0r1[1:0], L204A_0a, reset);
  tko0m2_1nm2b2 I55 (L203P_0r, L203P_0a, L205A_0r0[1:0], L205A_0r1[1:0], L205A_0a, reset);
  tkm2x2b I56 (L204P_0r0[1:0], L204P_0r1[1:0], L204P_0a, L205P_0r0[1:0], L205P_0r1[1:0], L205P_0a, L206A_0r0[1:0], L206A_0r1[1:0], L206A_0a, reset);
  tkj2m0_2 I57 (L199P_0r, L199P_0a, L206P_0r0[1:0], L206P_0r1[1:0], L206P_0a, L207A_0r0[1:0], L207A_0r1[1:0], L207A_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I58 (L207P_0r0[1:0], L207P_0r1[1:0], L207P_0a, L166A_0r, L166A_0a, L189A_0r, L189A_0a, reset);
  tkf0mo0w0_o0w0 I59 (L66P_0r, L66P_0a, L210A_0r, L210A_0a, L289A_0r, L289A_0a, reset);
  tkm2x1b I60 (L211P_0r0, L211P_0r1, L211P_0a, L213P_0r0, L213P_0r1, L213P_0a, L208A_0r0, L208A_0r1, L208A_0a, reset);
  tko0m2_1nm2b1 I61 (L210P_0r, L210P_0a, L214A_0r0[1:0], L214A_0r1[1:0], L214A_0a, reset);
  tko0m2_1nm2b2 I62 (L212P_0r, L212P_0a, L215A_0r0[1:0], L215A_0r1[1:0], L215A_0a, reset);
  tkm2x2b I63 (L214P_0r0[1:0], L214P_0r1[1:0], L214P_0a, L215P_0r0[1:0], L215P_0r1[1:0], L215P_0a, L216A_0r0[1:0], L216A_0r1[1:0], L216A_0a, reset);
  tkj2m0_2 I64 (L209_0r, L209_0a, L216P_0r0[1:0], L216P_0r1[1:0], L216P_0a, L217A_0r0[1:0], L217A_0r1[1:0], L217A_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I65 (L217P_0r0[1:0], L217P_0r1[1:0], L217P_0a, L69A_0r, L69A_0a, L9A_0r, L9A_0a, reset);
  tkvStopped1_wo0w1_ro0w1 I66 (L208P_0r0, L208P_0r1, L208P_0a, L209_0r, L209_0a, L13P_0r, L13P_0a, L14_0r0, L14_0r1, L14_0a, reset);
  tkvMDR32_wo0w32_ro0w32o0w5 I67 (L169P_0r0[31:0], L169P_0r1[31:0], L169P_0a, L170_0r, L170_0a, L122P_0r, L122P_0a, L294P_0r, L294P_0a, L123_0r0[31:0], L123_0r1[31:0], L123_0a, L221_0r0[4:0], L221_0r1[4:0], L221_0a, reset);
  tkf0mo0w0_o0w0 I68 (L16P_0r, L16P_0a, L222A_0r, L222A_0a, L287A_0r, L287A_0a, reset);
  tkm2x5b I69 (L221_0r0[4:0], L221_0r1[4:0], L221_0a, L223P_0r0[4:0], L223P_0r1[4:0], L223P_0a, L218A_0r0[4:0], L218A_0r1[4:0], L218A_0a, reset);
  tko0m2_1nm2b1 I70 (L220P_0r, L220P_0a, L224A_0r0[1:0], L224A_0r1[1:0], L224A_0a, reset);
  tko0m2_1nm2b2 I71 (L222P_0r, L222P_0a, L225A_0r0[1:0], L225A_0r1[1:0], L225A_0a, reset);
  tkm2x2b I72 (L224P_0r0[1:0], L224P_0r1[1:0], L224P_0a, L225P_0r0[1:0], L225P_0r1[1:0], L225P_0a, L226A_0r0[1:0], L226A_0r1[1:0], L226A_0a, reset);
  tkj2m0_2 I73 (L219_0r, L219_0a, L226P_0r0[1:0], L226P_0r1[1:0], L226P_0a, L302A_0r0[1:0], L302A_0r1[1:0], L302A_0a, reset);
  tkvPCstep5_wo0w5_ro0w5 I74 (L218P_0r0[4:0], L218P_0r1[4:0], L218P_0a, L219_0r, L219_0a, L98P_0r, L98P_0a, L99_0r0[4:0], L99_0r1[4:0], L99_0a, reset);
  tkf0mo0w0_o0w0 I75 (L137P_0r, L137P_0a, L230A_0r, L230A_0a, L290A_0r, L290A_0a, reset);
  tkm2x5b I76 (L231P_0r0[4:0], L231P_0r1[4:0], L231P_0a, L233P_0r0[4:0], L233P_0r1[4:0], L233P_0a, L228A_0r0[4:0], L228A_0r1[4:0], L228A_0a, reset);
  tko0m2_1nm2b1 I77 (L230P_0r, L230P_0a, L234A_0r0[1:0], L234A_0r1[1:0], L234A_0a, reset);
  tko0m2_1nm2b2 I78 (L232P_0r, L232P_0a, L235A_0r0[1:0], L235A_0r1[1:0], L235A_0a, reset);
  tkm2x2b I79 (L234P_0r0[1:0], L234P_0r1[1:0], L234P_0a, L235P_0r0[1:0], L235P_0r1[1:0], L235P_0a, L236A_0r0[1:0], L236A_0r1[1:0], L236A_0a, reset);
  tkj2m0_2 I80 (L229_0r, L229_0a, L236P_0r0[1:0], L236P_0r1[1:0], L236P_0a, L237A_0r0[1:0], L237A_0r1[1:0], L237A_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I81 (L237P_0r0[1:0], L237P_0r1[1:0], L237P_0a, L140A_0r, L140A_0a, L104A_0r, L104A_0a, reset);
  tkvPC5_wo0w5_ro0w5o0w5 I82 (L228P_0r0[4:0], L228P_0r1[4:0], L228P_0a, L229_0r, L229_0a, L96P_0r, L96P_0a, L296P_0r, L296P_0a, L97_0r0[4:0], L97_0r1[4:0], L97_0a, L249_0r0[4:0], L249_0r1[4:0], L249_0a, reset);
  tkvIR32_wo0w32_ro0w5 I83 (L284P_0r0[31:0], L284P_0r1[31:0], L284P_0a, L283_0r, L283_0a, L297P_0r, L297P_0a, L251_0r0[4:0], L251_0r1[4:0], L251_0a, reset);
  tkvACCslave32_wo0w32_ro0w32o0w32 I84 (L127P_0r0[31:0], L127P_0r1[31:0], L127P_0a, L128_0r, L128_0a, L298P_0r, L298P_0a, L295P_0r, L295P_0a, MemW_0r0[31:0], MemW_0r1[31:0], MemW_0a, L243_0r0[31:0], L243_0r1[31:0], L243_0a, reset);
  tkf0mo0w0_o0w0 I85 (L149P_0r, L149P_0a, L240A_0r, L240A_0a, L291A_0r, L291A_0a, reset);
  tkm2x32b I86 (L241P_0r0[31:0], L241P_0r1[31:0], L241P_0a, L243_0r0[31:0], L243_0r1[31:0], L243_0a, L238A_0r0[31:0], L238A_0r1[31:0], L238A_0a, reset);
  tko0m2_1nm2b1 I87 (L240P_0r, L240P_0a, L244A_0r0[1:0], L244A_0r1[1:0], L244A_0a, reset);
  tko0m2_1nm2b2 I88 (L242P_0r, L242P_0a, L245A_0r0[1:0], L245A_0r1[1:0], L245A_0a, reset);
  tkm2x2b I89 (L244P_0r0[1:0], L244P_0r1[1:0], L244P_0a, L245P_0r0[1:0], L245P_0r1[1:0], L245P_0a, L246A_0r0[1:0], L246A_0r1[1:0], L246A_0a, reset);
  tkj2m0_2 I90 (L239_0r, L239_0a, L246P_0r0[1:0], L246P_0r1[1:0], L246P_0a, L247A_0r0[1:0], L247A_0r1[1:0], L247A_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I91 (L247P_0r0[1:0], L247P_0r1[1:0], L247P_0a, L152A_0r, L152A_0a, L74A_0r, L74A_0a, reset);
  tkvACC32_wo0w32_ro0w32o31w1 I92 (L238P_0r0[31:0], L238P_0r1[31:0], L238P_0a, L239_0r, L239_0a, L120P_0r, L120P_0a, L60P_0r, L60P_0a, L121_0r0[31:0], L121_0r1[31:0], L121_0a, L61_0r0, L61_0r1, L61_0a, reset);
  tkm2x5b I93 (L249_0r0[4:0], L249_0r1[4:0], L249_0a, L251_0r0[4:0], L251_0r1[4:0], L251_0a, L252A_0r0[4:0], L252A_0r1[4:0], L252A_0a, reset);
  tkf5mo0w0_o0w5 I94 (L252P_0r0[4:0], L252P_0r1[4:0], L252P_0a, L253A_0r, L253A_0a, L254_0r0[4:0], L254_0r1[4:0], L254_0a, reset);
  tko0m2_1nm2b1 I95 (L248P_0r, L248P_0a, L255A_0r0[1:0], L255A_0r1[1:0], L255A_0a, reset);
  tko0m2_1nm2b2 I96 (L250P_0r, L250P_0a, L256A_0r0[1:0], L256A_0r1[1:0], L256A_0a, reset);
  tkm2x2b I97 (L255P_0r0[1:0], L255P_0r1[1:0], L255P_0a, L256P_0r0[1:0], L256P_0r1[1:0], L256P_0a, L257A_0r0[1:0], L257A_0r1[1:0], L257A_0a, reset);
  tkj2m0_2 I98 (L253P_0r, L253P_0a, L257P_0r0[1:0], L257P_0r1[1:0], L257P_0a, L258A_0r0[1:0], L258A_0r1[1:0], L258A_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I99 (L258P_0r0[1:0], L258P_0r1[1:0], L258P_0a, L29A_0r, L29A_0a, L199A_0r, L199A_0a, reset);
  tkm3x1b I100 (L260P_0r0, L260P_0r1, L260P_0a, L262P_0r0, L262P_0r1, L262P_0a, L264P_0r0, L264P_0r1, L264P_0a, L265A_0r0, L265A_0r1, L265A_0a, reset);
  tkf1mo0w0_o0w1 I101 (L265P_0r0, L265P_0r1, L265P_0a, L266A_0r, L266A_0a, L267_0r0, L267_0r1, L267_0a, reset);
  tko0m3_1nm3b1 I102 (L259P_0r, L259P_0a, L268A_0r0[2:0], L268A_0r1[2:0], L268A_0a, reset);
  tko0m3_1nm3b2 I103 (L261P_0r, L261P_0a, L269A_0r0[2:0], L269A_0r1[2:0], L269A_0a, reset);
  tko0m3_1nm3b4 I104 (L263P_0r, L263P_0a, L270A_0r0[2:0], L270A_0r1[2:0], L270A_0a, reset);
  tkm3x3b I105 (L268P_0r0[2:0], L268P_0r1[2:0], L268P_0a, L269P_0r0[2:0], L269P_0r1[2:0], L269P_0a, L270P_0r0[2:0], L270P_0r1[2:0], L270P_0a, L271A_0r0[2:0], L271A_0r1[2:0], L271A_0a, reset);
  tkj3m0_3 I106 (L266P_0r, L266P_0a, L271P_0r0[2:0], L271P_0r1[2:0], L271P_0a, L272A_0r0[2:0], L272A_0r1[2:0], L272A_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_4o0w0 I107 (L272P_0r0[2:0], L272P_0r1[2:0], L272P_0a, L25A_0r, L25A_0a, L164A_0r, L164A_0a, L187A_0r, L187A_0a, reset);
  tko0m2_1nm2b1 I108 (L31P_0r, L31P_0a, L274A_0r0[1:0], L274A_0r1[1:0], L274A_0a, reset);
  tko0m2_1nm2b2 I109 (L168P_0r, L168P_0a, L275A_0r0[1:0], L275A_0r1[1:0], L275A_0a, reset);
  tkm2x2b I110 (L274P_0r0[1:0], L274P_0r1[1:0], L274P_0a, L275P_0r0[1:0], L275P_0r1[1:0], L275P_0a, L276A_0r0[1:0], L276A_0r1[1:0], L276A_0a, reset);
  tkj34m32_2 I111 (L273_0r0[31:0], L273_0r1[31:0], L273_0a, L276P_0r0[1:0], L276P_0r1[1:0], L276P_0a, L277A_0r0[33:0], L277A_0r1[33:0], L277A_0a, reset);
  tks34_o32w2_1o0w32_2o0w32 I112 (L277P_0r0[33:0], L277P_0r1[33:0], L277P_0a, L32A_0r0[31:0], L32A_0r1[31:0], L32A_0a, L169A_0r0[31:0], L169A_0r1[31:0], L169A_0a, reset);
  tkf0mo0w0_o0w0 I113 (L78P_0r, L78P_0a, L79_0r, L79_0a, L279_0r, L279_0a, reset);
  tkf32mo0w32_o13w3 I114 (L32P_0r0[31:0], L32P_0r1[31:0], L32P_0a, L284A_0r0[31:0], L284A_0r1[31:0], L284A_0a, L285A_0r0[2:0], L285A_0r1[2:0], L285A_0a, reset);
  tkj3m3_0_0_0 I115 (L285P_0r0[2:0], L285P_0r1[2:0], L285P_0a, L25P_0r, L25P_0a, L29P_0r, L29P_0a, L283_0r, L283_0a, L38A_0r0[2:0], L38A_0r1[2:0], L38A_0a, reset);
  tkf0mo0w0_o0w0 I116 (L71P_0r, L71P_0a, L295A_0r, L295A_0a, L242A_0r, L242A_0a, reset);
  tkf0mo0w0_o0w0 I117 (L196P_0r, L196P_0a, L297A_0r, L297A_0a, L250A_0r, L250A_0a, reset);
  tkf3mo0w3_o0w0 I118 (L299P_0r0[2:0], L299P_0r1[2:0], L299P_0a, L309A_0r0[2:0], L309A_0r1[2:0], L309A_0a, L301A_0r, L301A_0a, reset);
  tkf2mo0w2_o0w0 I119 (L302P_0r0[1:0], L302P_0r1[1:0], L302P_0a, L310A_0r0[1:0], L310A_0r1[1:0], L310A_0a, L304A_0r, L304A_0a, reset);
  tko64m32_1nm2b0_2api0w32bt1o0w2b_3nm2b0_4api32w32bt3o0w2b_5subt2o0w34bt4o0w34b_6apt5o0w32b I120 (L124P_0r0[63:0], L124P_0r1[63:0], L124P_0a, L127A_0r0[31:0], L127A_0r1[31:0], L127A_0a, reset);
  tko3m3_1nm3b1_2nm3b2_3mx0_1_i0w3bt1o0w3bt2o0w3b I121 (L309P_0r0[2:0], L309P_0r1[2:0], L309P_0a, L179A_0r0[2:0], L179A_0r1[2:0], L179A_0a, reset);
  tko2m3_1nm3b4_2nm3b1_3mx1_2_i0w2bt1o0w3bt2o0w3b I122 (L310P_0r0[1:0], L310P_0r1[1:0], L310P_0a, L113A_0r0[2:0], L113A_0r1[2:0], L113A_0a, reset);
  tkm2x0b I123 (L311P_0r, L311P_0a, L312P_0r, L312P_0a, L315A_0r, L315A_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I124 (L315P_0r, L315P_0a, L294A_0r, L294A_0a, L220A_0r, L220A_0a, L306A_0r, L306A_0a, reset);
  tkm2x0b I125 (L313P_0r, L313P_0a, L314P_0r, L314P_0a, L318A_0r, L318A_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I126 (L318P_0r, L318P_0a, L177A_0r, L177A_0a, L178A_0r, L178A_0a, L308A_0r, L308A_0a, reset);
  tkl0x1 I127 (L3A_0r, L3A_0a, L3P_0r, L3P_0a, reset);
  tkl0x1 I128 (L5A_0r, L5A_0a, L5P_0r, L5P_0a, reset);
  tkl0x1 I129 (L9A_0r, L9A_0a, L9P_0r, L9P_0a, reset);
  tkl0x1 I130 (go_0r, go_0a, L10_0r, L10_0a, reset);
  tkl1x1 I131 (L12A_0r0, L12A_0r1, L12A_0a, L12P_0r0, L12P_0r1, L12P_0a, reset);
  tkl0x1 I132 (L13A_0r, L13A_0a, L13P_0r, L13P_0a, reset);
  tkl0x1 I133 (L16A_0r, L16A_0a, L16P_0r, L16P_0a, reset);
  tkl0x1 I134 (L25A_0r, L25A_0a, L25P_0r, L25P_0a, reset);
  tkl0x1 I135 (L29A_0r, L29A_0a, L29P_0r, L29P_0a, reset);
  tkl0x1 I136 (L31A_0r, L31A_0a, L31P_0r, L31P_0a, reset);
  tkl32x1 I137 (L32A_0r0[31:0], L32A_0r1[31:0], L32A_0a, L32P_0r0[31:0], L32P_0r1[31:0], L32P_0a, reset);
  tkl0x1 I138 (L34A_0r, L34A_0a, L34P_0r, L34P_0a, reset);
  tkl3x1 I139 (L38A_0r0[2:0], L38A_0r1[2:0], L38A_0a, L38P_0r0[2:0], L38P_0r1[2:0], L38P_0a, reset);
  tkl0x1 I140 (L42A_0r, L42A_0a, L42P_0r, L42P_0a, reset);
  tkl0x1 I141 (L52A_0r, L52A_0a, L52P_0r, L52P_0a, reset);
  tkl0x1 I142 (L57A_0r, L57A_0a, L57P_0r, L57P_0a, reset);
  tkl0x1 I143 (L60A_0r, L60A_0a, L60P_0r, L60P_0a, reset);
  tkl0x1 I144 (L62A_0r, L62A_0a, L62P_0r, L62P_0a, reset);
  tkl0x1 I145 (L63A_0r, L63A_0a, L63P_0r, L63P_0a, reset);
  tkl0x1 I146 (L64A_0r, L64A_0a, L64P_0r, L64P_0a, reset);
  tkl0x1 I147 (L66A_0r, L66A_0a, L66P_0r, L66P_0a, reset);
  tkl0x1 I148 (L69A_0r, L69A_0a, L69P_0r, L69P_0a, reset);
  tkl0x1 I149 (L71A_0r, L71A_0a, L71P_0r, L71P_0a, reset);
  tkl0x1 I150 (L74A_0r, L74A_0a, L74P_0r, L74P_0a, reset);
  tkl0x1 I151 (L76A_0r, L76A_0a, L76P_0r, L76P_0a, reset);
  tkl0x1 I152 (L78A_0r, L78A_0a, L78P_0r, L78P_0a, reset);
  tkl0x1 I153 (L79_0r, L79_0a, done_0r, done_0a, reset);
  tkl0x1 I154 (L86A_0r, L86A_0a, L86P_0r, L86P_0a, reset);
  tkl0x1 I155 (L96A_0r, L96A_0a, L96P_0r, L96P_0a, reset);
  tkl0x1 I156 (L98A_0r, L98A_0a, L98P_0r, L98P_0a, reset);
  tkl10x1 I157 (L100A_0r0[9:0], L100A_0r1[9:0], L100A_0a, L100P_0r0[9:0], L100P_0r1[9:0], L100P_0a, reset);
  tkl6x1 I158 (L101A_0r0[5:0], L101A_0r1[5:0], L101A_0a, L101P_0r0[5:0], L101P_0r1[5:0], L101P_0a, reset);
  tkl0x1 I159 (L102A_0r, L102A_0a, L102P_0r, L102P_0a, reset);
  tkl0x1 I160 (L104A_0r, L104A_0a, L104P_0r, L104P_0a, reset);
  tkl0x1 I161 (L107A_0r, L107A_0a, L107P_0r, L107P_0a, reset);
  tkl0x1 I162 (L108A_0r, L108A_0a, L108P_0r, L108P_0a, reset);
  tkl3x1 I163 (L112A_0r0[2:0], L112A_0r1[2:0], L112A_0a, L112P_0r0[2:0], L112P_0r1[2:0], L112P_0a, reset);
  tkl3x1 I164 (L113A_0r0[2:0], L113A_0r1[2:0], L113A_0a, L113P_0r0[2:0], L113P_0r1[2:0], L113P_0a, reset);
  tkl3x1 I165 (L114A_0r0[2:0], L114A_0r1[2:0], L114A_0a, L114P_0r0[2:0], L114P_0r1[2:0], L114P_0a, reset);
  tkl3x1 I166 (L115A_0r0[2:0], L115A_0r1[2:0], L115A_0a, L115P_0r0[2:0], L115P_0r1[2:0], L115P_0a, reset);
  tkl0x1 I167 (L120A_0r, L120A_0a, L120P_0r, L120P_0a, reset);
  tkl0x1 I168 (L122A_0r, L122A_0a, L122P_0r, L122P_0a, reset);
  tkl64x1 I169 (L124A_0r0[63:0], L124A_0r1[63:0], L124A_0a, L124P_0r0[63:0], L124P_0r1[63:0], L124P_0a, reset);
  tkl0x1 I170 (L126A_0r, L126A_0a, L126P_0r, L126P_0a, reset);
  tkl32x1 I171 (L127A_0r0[31:0], L127A_0r1[31:0], L127A_0a, L127P_0r0[31:0], L127P_0r1[31:0], L127P_0a, reset);
  tkl0x1 I172 (L137A_0r, L137A_0a, L137P_0r, L137P_0a, reset);
  tkl0x1 I173 (L140A_0r, L140A_0a, L140P_0r, L140P_0a, reset);
  tkl0x1 I174 (L141A_0r, L141A_0a, L141P_0r, L141P_0a, reset);
  tkl0x1 I175 (L142A_0r, L142A_0a, L142P_0r, L142P_0a, reset);
  tkl0x1 I176 (L143A_0r, L143A_0a, L143P_0r, L143P_0a, reset);
  tkl0x1 I177 (L144A_0r, L144A_0a, L144P_0r, L144P_0a, reset);
  tkl2x1 I178 (L145A_0r0[1:0], L145A_0r1[1:0], L145A_0a, L145P_0r0[1:0], L145P_0r1[1:0], L145P_0a, reset);
  tkl2x1 I179 (L146A_0r0[1:0], L146A_0r1[1:0], L146A_0a, L146P_0r0[1:0], L146P_0r1[1:0], L146P_0a, reset);
  tkl2x1 I180 (L147A_0r0[1:0], L147A_0r1[1:0], L147A_0a, L147P_0r0[1:0], L147P_0r1[1:0], L147P_0a, reset);
  tkl2x1 I181 (L148A_0r0[1:0], L148A_0r1[1:0], L148A_0a, L148P_0r0[1:0], L148P_0r1[1:0], L148P_0a, reset);
  tkl0x1 I182 (L149A_0r, L149A_0a, L149P_0r, L149P_0a, reset);
  tkl0x1 I183 (L152A_0r, L152A_0a, L152P_0r, L152P_0a, reset);
  tkl0x1 I184 (L153A_0r, L153A_0a, L153P_0r, L153P_0a, reset);
  tkl0x1 I185 (L154A_0r, L154A_0a, L154P_0r, L154P_0a, reset);
  tkl0x1 I186 (L155A_0r, L155A_0a, L155P_0r, L155P_0a, reset);
  tkl0x1 I187 (L156A_0r, L156A_0a, L156P_0r, L156P_0a, reset);
  tkl2x1 I188 (L157A_0r0[1:0], L157A_0r1[1:0], L157A_0a, L157P_0r0[1:0], L157P_0r1[1:0], L157P_0a, reset);
  tkl2x1 I189 (L158A_0r0[1:0], L158A_0r1[1:0], L158A_0a, L158P_0r0[1:0], L158P_0r1[1:0], L158P_0a, reset);
  tkl2x1 I190 (L159A_0r0[1:0], L159A_0r1[1:0], L159A_0a, L159P_0r0[1:0], L159P_0r1[1:0], L159P_0a, reset);
  tkl2x1 I191 (L160A_0r0[1:0], L160A_0r1[1:0], L160A_0a, L160P_0r0[1:0], L160P_0r1[1:0], L160P_0a, reset);
  tkl0x1 I192 (L164A_0r, L164A_0a, L164P_0r, L164P_0a, reset);
  tkl0x1 I193 (L166A_0r, L166A_0a, L166P_0r, L166P_0a, reset);
  tkl0x1 I194 (L168A_0r, L168A_0a, L168P_0r, L168P_0a, reset);
  tkl32x1 I195 (L169A_0r0[31:0], L169A_0r1[31:0], L169A_0a, L169P_0r0[31:0], L169P_0r1[31:0], L169P_0a, reset);
  tkl0x1 I196 (L171A_0r, L171A_0a, L171P_0r, L171P_0a, reset);
  tkl0x1 I197 (L177A_0r, L177A_0a, L177P_0r, L177P_0a, reset);
  tkl0x1 I198 (L178A_0r, L178A_0a, L178P_0r, L178P_0a, reset);
  tkl3x1 I199 (L179A_0r0[2:0], L179A_0r1[2:0], L179A_0a, L179P_0r0[2:0], L179P_0r1[2:0], L179P_0a, reset);
  tkl3x1 I200 (L181A_0r0[2:0], L181A_0r1[2:0], L181A_0a, L181P_0r0[2:0], L181P_0r1[2:0], L181P_0a, reset);
  tkl3x1 I201 (L182A_0r0[2:0], L182A_0r1[2:0], L182A_0a, L182P_0r0[2:0], L182P_0r1[2:0], L182P_0a, reset);
  tkl3x1 I202 (L183A_0r0[2:0], L183A_0r1[2:0], L183A_0a, L183P_0r0[2:0], L183P_0r1[2:0], L183P_0a, reset);
  tkl0x1 I203 (L187A_0r, L187A_0a, L187P_0r, L187P_0a, reset);
  tkl0x1 I204 (L189A_0r, L189A_0a, L189P_0r, L189P_0a, reset);
  tkl0x1 I205 (L193A_0r, L193A_0a, L193P_0r, L193P_0a, reset);
  tkl0x1 I206 (L194A_0r, L194A_0a, L194P_0r, L194P_0a, reset);
  tkl0x1 I207 (L196A_0r, L196A_0a, L196P_0r, L196P_0a, reset);
  tkl0x1 I208 (L199A_0r, L199A_0a, L199P_0r, L199P_0a, reset);
  tkl0x1 I209 (L200A_0r, L200A_0a, L200P_0r, L200P_0a, reset);
  tkl0x1 I210 (L201A_0r, L201A_0a, L201P_0r, L201P_0a, reset);
  tkl0x1 I211 (L202A_0r, L202A_0a, L202P_0r, L202P_0a, reset);
  tkl0x1 I212 (L203A_0r, L203A_0a, L203P_0r, L203P_0a, reset);
  tkl2x1 I213 (L204A_0r0[1:0], L204A_0r1[1:0], L204A_0a, L204P_0r0[1:0], L204P_0r1[1:0], L204P_0a, reset);
  tkl2x1 I214 (L205A_0r0[1:0], L205A_0r1[1:0], L205A_0a, L205P_0r0[1:0], L205P_0r1[1:0], L205P_0a, reset);
  tkl2x1 I215 (L206A_0r0[1:0], L206A_0r1[1:0], L206A_0a, L206P_0r0[1:0], L206P_0r1[1:0], L206P_0a, reset);
  tkl2x1 I216 (L207A_0r0[1:0], L207A_0r1[1:0], L207A_0a, L207P_0r0[1:0], L207P_0r1[1:0], L207P_0a, reset);
  tkl1x1 I217 (L208A_0r0, L208A_0r1, L208A_0a, L208P_0r0, L208P_0r1, L208P_0a, reset);
  tkl0x1 I218 (L210A_0r, L210A_0a, L210P_0r, L210P_0a, reset);
  tkl1x1 I219 (L211A_0r0, L211A_0r1, L211A_0a, L211P_0r0, L211P_0r1, L211P_0a, reset);
  tkl0x1 I220 (L212A_0r, L212A_0a, L212P_0r, L212P_0a, reset);
  tkl1x1 I221 (L213A_0r0, L213A_0r1, L213A_0a, L213P_0r0, L213P_0r1, L213P_0a, reset);
  tkl2x1 I222 (L214A_0r0[1:0], L214A_0r1[1:0], L214A_0a, L214P_0r0[1:0], L214P_0r1[1:0], L214P_0a, reset);
  tkl2x1 I223 (L215A_0r0[1:0], L215A_0r1[1:0], L215A_0a, L215P_0r0[1:0], L215P_0r1[1:0], L215P_0a, reset);
  tkl2x1 I224 (L216A_0r0[1:0], L216A_0r1[1:0], L216A_0a, L216P_0r0[1:0], L216P_0r1[1:0], L216P_0a, reset);
  tkl2x1 I225 (L217A_0r0[1:0], L217A_0r1[1:0], L217A_0a, L217P_0r0[1:0], L217P_0r1[1:0], L217P_0a, reset);
  tkl5x1 I226 (L218A_0r0[4:0], L218A_0r1[4:0], L218A_0a, L218P_0r0[4:0], L218P_0r1[4:0], L218P_0a, reset);
  tkl0x1 I227 (L220A_0r, L220A_0a, L220P_0r, L220P_0a, reset);
  tkl0x1 I228 (L222A_0r, L222A_0a, L222P_0r, L222P_0a, reset);
  tkl5x1 I229 (L223A_0r0[4:0], L223A_0r1[4:0], L223A_0a, L223P_0r0[4:0], L223P_0r1[4:0], L223P_0a, reset);
  tkl2x1 I230 (L224A_0r0[1:0], L224A_0r1[1:0], L224A_0a, L224P_0r0[1:0], L224P_0r1[1:0], L224P_0a, reset);
  tkl2x1 I231 (L225A_0r0[1:0], L225A_0r1[1:0], L225A_0a, L225P_0r0[1:0], L225P_0r1[1:0], L225P_0a, reset);
  tkl2x1 I232 (L226A_0r0[1:0], L226A_0r1[1:0], L226A_0a, L226P_0r0[1:0], L226P_0r1[1:0], L226P_0a, reset);
  tkl5x1 I233 (L228A_0r0[4:0], L228A_0r1[4:0], L228A_0a, L228P_0r0[4:0], L228P_0r1[4:0], L228P_0a, reset);
  tkl0x1 I234 (L230A_0r, L230A_0a, L230P_0r, L230P_0a, reset);
  tkl5x1 I235 (L231A_0r0[4:0], L231A_0r1[4:0], L231A_0a, L231P_0r0[4:0], L231P_0r1[4:0], L231P_0a, reset);
  tkl0x1 I236 (L232A_0r, L232A_0a, L232P_0r, L232P_0a, reset);
  tkl5x1 I237 (L233A_0r0[4:0], L233A_0r1[4:0], L233A_0a, L233P_0r0[4:0], L233P_0r1[4:0], L233P_0a, reset);
  tkl2x1 I238 (L234A_0r0[1:0], L234A_0r1[1:0], L234A_0a, L234P_0r0[1:0], L234P_0r1[1:0], L234P_0a, reset);
  tkl2x1 I239 (L235A_0r0[1:0], L235A_0r1[1:0], L235A_0a, L235P_0r0[1:0], L235P_0r1[1:0], L235P_0a, reset);
  tkl2x1 I240 (L236A_0r0[1:0], L236A_0r1[1:0], L236A_0a, L236P_0r0[1:0], L236P_0r1[1:0], L236P_0a, reset);
  tkl2x1 I241 (L237A_0r0[1:0], L237A_0r1[1:0], L237A_0a, L237P_0r0[1:0], L237P_0r1[1:0], L237P_0a, reset);
  tkl32x1 I242 (L238A_0r0[31:0], L238A_0r1[31:0], L238A_0a, L238P_0r0[31:0], L238P_0r1[31:0], L238P_0a, reset);
  tkl0x1 I243 (L240A_0r, L240A_0a, L240P_0r, L240P_0a, reset);
  tkl32x1 I244 (L241A_0r0[31:0], L241A_0r1[31:0], L241A_0a, L241P_0r0[31:0], L241P_0r1[31:0], L241P_0a, reset);
  tkl0x1 I245 (L242A_0r, L242A_0a, L242P_0r, L242P_0a, reset);
  tkl2x1 I246 (L244A_0r0[1:0], L244A_0r1[1:0], L244A_0a, L244P_0r0[1:0], L244P_0r1[1:0], L244P_0a, reset);
  tkl2x1 I247 (L245A_0r0[1:0], L245A_0r1[1:0], L245A_0a, L245P_0r0[1:0], L245P_0r1[1:0], L245P_0a, reset);
  tkl2x1 I248 (L246A_0r0[1:0], L246A_0r1[1:0], L246A_0a, L246P_0r0[1:0], L246P_0r1[1:0], L246P_0a, reset);
  tkl2x1 I249 (L247A_0r0[1:0], L247A_0r1[1:0], L247A_0a, L247P_0r0[1:0], L247P_0r1[1:0], L247P_0a, reset);
  tkl0x1 I250 (L248A_0r, L248A_0a, L248P_0r, L248P_0a, reset);
  tkl0x1 I251 (L250A_0r, L250A_0a, L250P_0r, L250P_0a, reset);
  tkl5x1 I252 (L252A_0r0[4:0], L252A_0r1[4:0], L252A_0a, L252P_0r0[4:0], L252P_0r1[4:0], L252P_0a, reset);
  tkl0x1 I253 (L253A_0r, L253A_0a, L253P_0r, L253P_0a, reset);
  tkl5x1 I254 (L254_0r0[4:0], L254_0r1[4:0], L254_0a, MemA_0r0[4:0], MemA_0r1[4:0], MemA_0a, reset);
  tkl2x1 I255 (L255A_0r0[1:0], L255A_0r1[1:0], L255A_0a, L255P_0r0[1:0], L255P_0r1[1:0], L255P_0a, reset);
  tkl2x1 I256 (L256A_0r0[1:0], L256A_0r1[1:0], L256A_0a, L256P_0r0[1:0], L256P_0r1[1:0], L256P_0a, reset);
  tkl2x1 I257 (L257A_0r0[1:0], L257A_0r1[1:0], L257A_0a, L257P_0r0[1:0], L257P_0r1[1:0], L257P_0a, reset);
  tkl2x1 I258 (L258A_0r0[1:0], L258A_0r1[1:0], L258A_0a, L258P_0r0[1:0], L258P_0r1[1:0], L258P_0a, reset);
  tkl0x1 I259 (L259A_0r, L259A_0a, L259P_0r, L259P_0a, reset);
  tkl1x1 I260 (L260A_0r0, L260A_0r1, L260A_0a, L260P_0r0, L260P_0r1, L260P_0a, reset);
  tkl0x1 I261 (L261A_0r, L261A_0a, L261P_0r, L261P_0a, reset);
  tkl1x1 I262 (L262A_0r0, L262A_0r1, L262A_0a, L262P_0r0, L262P_0r1, L262P_0a, reset);
  tkl0x1 I263 (L263A_0r, L263A_0a, L263P_0r, L263P_0a, reset);
  tkl1x1 I264 (L264A_0r0, L264A_0r1, L264A_0a, L264P_0r0, L264P_0r1, L264P_0a, reset);
  tkl1x1 I265 (L265A_0r0, L265A_0r1, L265A_0a, L265P_0r0, L265P_0r1, L265P_0a, reset);
  tkl0x1 I266 (L266A_0r, L266A_0a, L266P_0r, L266P_0a, reset);
  tkl1x1 I267 (L267_0r0, L267_0r1, L267_0a, MemRNW_0r0, MemRNW_0r1, MemRNW_0a, reset);
  tkl3x1 I268 (L268A_0r0[2:0], L268A_0r1[2:0], L268A_0a, L268P_0r0[2:0], L268P_0r1[2:0], L268P_0a, reset);
  tkl3x1 I269 (L269A_0r0[2:0], L269A_0r1[2:0], L269A_0a, L269P_0r0[2:0], L269P_0r1[2:0], L269P_0a, reset);
  tkl3x1 I270 (L270A_0r0[2:0], L270A_0r1[2:0], L270A_0a, L270P_0r0[2:0], L270P_0r1[2:0], L270P_0a, reset);
  tkl3x1 I271 (L271A_0r0[2:0], L271A_0r1[2:0], L271A_0a, L271P_0r0[2:0], L271P_0r1[2:0], L271P_0a, reset);
  tkl3x1 I272 (L272A_0r0[2:0], L272A_0r1[2:0], L272A_0a, L272P_0r0[2:0], L272P_0r1[2:0], L272P_0a, reset);
  tkl32x1 I273 (MemR_0r0[31:0], MemR_0r1[31:0], MemR_0a, L273_0r0[31:0], L273_0r1[31:0], L273_0a, reset);
  tkl2x1 I274 (L274A_0r0[1:0], L274A_0r1[1:0], L274A_0a, L274P_0r0[1:0], L274P_0r1[1:0], L274P_0a, reset);
  tkl2x1 I275 (L275A_0r0[1:0], L275A_0r1[1:0], L275A_0a, L275P_0r0[1:0], L275P_0r1[1:0], L275P_0a, reset);
  tkl2x1 I276 (L276A_0r0[1:0], L276A_0r1[1:0], L276A_0a, L276P_0r0[1:0], L276P_0r1[1:0], L276P_0a, reset);
  tkl34x1 I277 (L277A_0r0[33:0], L277A_0r1[33:0], L277A_0a, L277P_0r0[33:0], L277P_0r1[33:0], L277P_0a, reset);
  tkl0x1 I278 (L279_0r, L279_0a, halted_0r, halted_0a, reset);
  tkl0x1 I279 (L280A_0r, L280A_0a, L280P_0r, L280P_0a, reset);
  tkl0x1 I280 (L281A_0r, L281A_0a, L281P_0r, L281P_0a, reset);
  tkl32x1 I281 (L284A_0r0[31:0], L284A_0r1[31:0], L284A_0a, L284P_0r0[31:0], L284P_0r1[31:0], L284P_0a, reset);
  tkl3x1 I282 (L285A_0r0[2:0], L285A_0r1[2:0], L285A_0a, L285P_0r0[2:0], L285P_0r1[2:0], L285P_0a, reset);
  tkl0x1 I283 (L286A_0r, L286A_0a, L286P_0r, L286P_0a, reset);
  tkl0x1 I284 (L287A_0r, L287A_0a, L287P_0r, L287P_0a, reset);
  tkl0x1 I285 (L288A_0r, L288A_0a, L288P_0r, L288P_0a, reset);
  tkl0x1 I286 (L289A_0r, L289A_0a, L289P_0r, L289P_0a, reset);
  tkl0x1 I287 (L290A_0r, L290A_0a, L290P_0r, L290P_0a, reset);
  tkl0x1 I288 (L291A_0r, L291A_0a, L291P_0r, L291P_0a, reset);
  tkl0x1 I289 (L292A_0r, L292A_0a, L292P_0r, L292P_0a, reset);
  tkl0x1 I290 (L293A_0r, L293A_0a, L293P_0r, L293P_0a, reset);
  tkl0x1 I291 (L294A_0r, L294A_0a, L294P_0r, L294P_0a, reset);
  tkl0x1 I292 (L295A_0r, L295A_0a, L295P_0r, L295P_0a, reset);
  tkl0x1 I293 (L296A_0r, L296A_0a, L296P_0r, L296P_0a, reset);
  tkl0x1 I294 (L297A_0r, L297A_0a, L297P_0r, L297P_0a, reset);
  tkl0x1 I295 (L298A_0r, L298A_0a, L298P_0r, L298P_0a, reset);
  tkl3x1 I296 (L299A_0r0[2:0], L299A_0r1[2:0], L299A_0a, L299P_0r0[2:0], L299P_0r1[2:0], L299P_0a, reset);
  tkl0x1 I297 (L301A_0r, L301A_0a, L301P_0r, L301P_0a, reset);
  tkl2x1 I298 (L302A_0r0[1:0], L302A_0r1[1:0], L302A_0a, L302P_0r0[1:0], L302P_0r1[1:0], L302P_0a, reset);
  tkl0x1 I299 (L304A_0r, L304A_0a, L304P_0r, L304P_0a, reset);
  tkl0x1 I300 (L306A_0r, L306A_0a, L306P_0r, L306P_0a, reset);
  tkl0x1 I301 (L308A_0r, L308A_0a, L308P_0r, L308P_0a, reset);
  tkl3x1 I302 (L309A_0r0[2:0], L309A_0r1[2:0], L309A_0a, L309P_0r0[2:0], L309P_0r1[2:0], L309P_0a, reset);
  tkl2x1 I303 (L310A_0r0[1:0], L310A_0r1[1:0], L310A_0a, L310P_0r0[1:0], L310P_0r1[1:0], L310P_0a, reset);
  tkl0x1 I304 (L311A_0r, L311A_0a, L311P_0r, L311P_0a, reset);
  tkl0x1 I305 (L312A_0r, L312A_0a, L312P_0r, L312P_0a, reset);
  tkl0x1 I306 (L313A_0r, L313A_0a, L313P_0r, L313P_0a, reset);
  tkl0x1 I307 (L314A_0r, L314A_0a, L314P_0r, L314P_0a, reset);
  tkl0x1 I308 (L315A_0r, L315A_0a, L315P_0r, L315P_0a, reset);
  tkl0x1 I309 (L318A_0r, L318A_0a, L318P_0r, L318P_0a, reset);
endmodule

// Netlist costs:
// teak_SSEM: AND2*1317 AO22*146 AO222*76 BUFF*1777 C2*415 C2R*1261 C3*740 GND*116 INV*270 NAND2*82 NOR2*173 NOR3*223 OR2*1166 OR3*15
// tkf0mo0w0_o0w0: BUFF*2 C2*1
// tkf0mo0w0_o0w0_o0w0: BUFF*3 C3*1
// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0: BUFF*5 C2*2 C3*1
// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0: BUFF*6 C2*1 C3*2
// tkf1mo0w0_o0w1: BUFF*4 C3*1 OR2*1
// tkf2mo0w2_o0w0: BUFF*6 C3*1 OR2*1
// tkf32mo0w32_o13w3: BUFF*69 C2*2 C3*1 OR2*1
// tkf3mo0w3_o0w0: BUFF*8 C3*1 OR2*1
// tkf5mo0w0_o0w5: BUFF*12 C3*1 OR2*1
// tkf6mo0w0_o0w5: BUFF*10 C2*3 C3*1 OR2*2
// tkj0m0_0: BUFF*2 C2*1
// tkj0m0_0_0: BUFF*3 C3*1
// tkj10m5_5: BUFF*41 C2*2 OR2*1
// tkj2m0_2: BUFF*9 C2*2
// tkj34m32_2: BUFF*137 C2*2 OR2*1
// tkj3m0_0_0_3: BUFF*14 C2*2 C3*1
// tkj3m0_3: BUFF*13 C2*2
// tkj3m3_0_0_0: BUFF*14 C2*2 C3*1
// tkj64m32_32: BUFF*257 C2*2 OR2*1
// tkl0x1: BUFF*1 C2R*1 INV*1
// tkl10x1: BUFF*2 C2*1 C2R*20 C3*4 INV*1 OR2*10
// tkl1x1: BUFF*1 C2R*2 INV*1 OR2*1
// tkl2x1: C2*1 C2R*4 INV*1 OR2*2
// tkl32x1: BUFF*1 C2*3 C2R*64 C3*14 INV*1 OR2*32
// tkl34x1: BUFF*2 C2*1 C2R*68 C3*16 INV*1 OR2*34
// tkl3x1: C2R*6 C3*1 INV*1 OR2*3
// tkl5x1: C2*2 C2R*10 C3*1 INV*1 OR2*5
// tkl64x1: BUFF*2 C2*1 C2R*128 C3*31 INV*1 OR2*64
// tkl6x1: C2*1 C2R*12 C3*2 INV*1 OR2*6
// tkm2x0b: C2R*4 NOR2*1 OR2*1
// tkm2x1b: AND2*4 BUFF*2 C2R*4 NOR2*1 OR2*5
// tkm2x2b: AND2*8 C2*2 C2R*4 NOR2*1 OR2*9
// tkm2x32b: AND2*128 BUFF*2 C2*6 C2R*4 C3*28 NOR2*1 OR2*129
// tkm2x3b: AND2*12 C2R*4 C3*2 NOR2*1 OR2*13
// tkm2x5b: AND2*20 C2*4 C2R*4 C3*2 NOR2*1 OR2*21
// tkm3x1b: AND2*6 BUFF*3 C2R*6 NOR2*1 OR2*3 OR3*3
// tkm3x3b: AND2*18 C2R*6 C3*3 NOR2*1 OR2*9 OR3*7
// tkm6x0b: C2R*12 NAND2*1 NOR2*1 NOR3*2
// tko0m1_1nm1b0: BUFF*2 GND*1
// tko0m1_1nm1b1: BUFF*2 GND*1
// tko0m2_1nm2b1: BUFF*3 GND*2
// tko0m2_1nm2b2: BUFF*3 GND*2
// tko0m32_1nm32b0: BUFF*33 GND*32
// tko0m3_1nm3b1: BUFF*4 GND*3
// tko0m3_1nm3b2: BUFF*4 GND*3
// tko0m3_1nm3b4: BUFF*4 GND*3
// tko0m5_1nm5b0: BUFF*6 GND*5
// tko0m5_1nm5b1: BUFF*6 GND*5
// tko10m6_1nm1b0_2api0w5bt1o0w1b_3nm1b0_4api5w5bt3o0w1b_5addt2o0w6bt4o0w6b: AO222*10 BUFF*30 C2*5 C3*44 GND*2 INV*10 NAND2*10 NOR3*10 OR2*12 OR3*1
// tko1m1_1noti0w1b: BUFF*3
// tko2m3_1nm3b4_2nm3b1_3mx1_2_i0w2bt1o0w3bt2o0w3b: BUFF*9 C2*4 C2R*14 C3*3 GND*6 OR2*16
// tko3m3_1nm3b1_2nm3b2_3mx0_1_i0w3bt1o0w3bt2o0w3b: BUFF*9 C2R*14 C3*7 GND*6 OR2*18
// tko64m32_1nm2b0_2api0w32bt1o0w2b_3nm2b0_4api32w32bt3o0w2b_5subt2o0w34bt4o0w34b_6apt5o0w32b: AO222*66 BUFF*208 C2*5 C3*295 GND*4 INV*66 NAND2*66 NOR3*66 OR2*66 OR3*1
// tks1_o0w1_0o0w0_1o0w0: BUFF*7 C2*3 OR2*2
// tks2_o0w2_1o0w0_2o0w0: BUFF*4 C2*6 OR2*3
// tks34_o32w2_1o0w32_2o0w32: BUFF*4 C2*134 C3*16 OR2*35
// tks3_o0w3_1o0w0_2o0w0_4o0w0: BUFF*6 C2*4 C3*4 OR2*3 OR3*1
// tks3_o0w3_2o0w0_3o0w0_4c1o0w0_6o0w0_7o0w0_0m1o0w3: BUFF*10 C2*14 C3*7 NAND2*1 NOR3*2 OR2*4
// tkvACC32_wo0w32_ro0w32o31w1: AND2*226 AO22*33 BUFF*102 C2*5 C3*29 INV*2 NAND2*1 NOR2*33 NOR3*33 OR2*32
// tkvACCslave32_wo0w32_ro0w32o0w32: AND2*288 AO22*33 BUFF*102 C2*5 C3*29 INV*2 NAND2*1 NOR2*33 NOR3*33 OR2*32
// tkvIR32_wo0w32_ro0w5: AND2*170 AO22*33 BUFF*101 C2*5 C3*29 INV*1 NOR2*33 NOR3*32 OR2*33
// tkvMDR32_wo0w32_ro0w32o0w5: AND2*234 AO22*33 BUFF*102 C2*5 C3*29 INV*2 NAND2*1 NOR2*33 NOR3*33 OR2*32
// tkvPC5_wo0w5_ro0w5o0w5: AND2*45 AO22*6 BUFF*19 C2*3 C3*3 INV*2 NAND2*1 NOR2*6 NOR3*6 OR2*5
// tkvPCstep5_wo0w5_ro0w5: AND2*35 AO22*6 BUFF*18 C2*3 C3*3 INV*1 NOR2*6 NOR3*5 OR2*6
// tkvStopped1_wo0w1_ro0w1: AND2*7 AO22*2 BUFF*7 C2*1 INV*1 NOR2*2 NOR3*1 OR2*2
