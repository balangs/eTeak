/*
    `nanoMultiplierPush.v'
    Balsa Verilog netlist file
    Created: Mon Nov  3 15:02:23 GMT 2008
    By: tarazonl@royaloak.cs.man.ac.uk (Linux)
    With net-verilog (balsa-netlist) version: 3.5.1
    Using technology: example/dual_b
    Command line : (balsa-netlist -bsdi helper nanoMultiplierPush)

    Using `simulation-initialise'
    You must set the following preprocessor directives to use this file:
        balsa_simulate: set if you wish to initialise signal values during sim.
        balsa_init_time: duration of forced initialisation
*/

module BALSA_TELEM (
  Ar,
  Aa,
  Br,
  Ba
);
  input Ar;
  output Aa;
  output Br;
  input Ba;
  wire s;
  AND2 I0 (Br, Ar, s);
  INV I1 (s, Aa);
  C2N I2 (Aa, Ba, Ar);
endmodule

module BrzActiveEagerFalseVariable_1_1_s0_ (
  trigger_0r, trigger_0a,
  write_0r, write_0a0d, write_0a1d,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d
);
  input trigger_0r;
  output trigger_0a;
  output write_0r;
  input write_0a0d;
  input write_0a1d;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output read_0a0d;
  output read_0a1d;
  wire cd_0n;
  wire partCD_0n;
  wire store_0n;
  wire store_1n;
  wire readReq_0n;
  wire writeAck_0n;
  wire sigAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_0a1d, store_1n, readReq_0n);
  AND2 I1 (read_0a0d, store_0n, readReq_0n);
  BUFF I2 (readReq_0n, read_0r);
  BUFF I3 (store_1n, write_0a1d);
  BUFF I4 (store_0n, write_0a0d);
  C2 I5 (trigger_0a, writeAck_0n, cd_0n);
  AND2 I6 (writeAck_0n, sigAck_0n, rReqOr_0n);
  INV I7 (rReqOr_0n, readReq_0n);
  BALSA_TELEM I8 (trigger_0r, sigAck_0n, signal_0r, signal_0a);
  BUFF I9 (cd_0n, partCD_0n);
  OR2 I10 (partCD_0n, store_0n, store_1n);
  BUFF I11 (write_0r, trigger_0r);
endmodule

module BrzActiveEagerFalseVariable_1_2_s0_ (
  trigger_0r, trigger_0a,
  write_0r, write_0a0d, write_0a1d,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d
);
  input trigger_0r;
  output trigger_0a;
  output write_0r;
  input write_0a0d;
  input write_0a1d;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output read_0a0d;
  output read_0a1d;
  input read_1r;
  output read_1a0d;
  output read_1a1d;
  wire cd_0n;
  wire partCD_0n;
  wire store_0n;
  wire store_1n;
  wire readReq_0n;
  wire readReq_1n;
  wire writeAck_0n;
  wire sigAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_1a1d, store_1n, readReq_1n);
  AND2 I1 (read_1a0d, store_0n, readReq_1n);
  AND2 I2 (read_0a1d, store_1n, readReq_0n);
  AND2 I3 (read_0a0d, store_0n, readReq_0n);
  BUFF I4 (readReq_0n, read_0r);
  BUFF I5 (readReq_1n, read_1r);
  BUFF I6 (store_1n, write_0a1d);
  BUFF I7 (store_0n, write_0a0d);
  C2 I8 (trigger_0a, writeAck_0n, cd_0n);
  AND2 I9 (writeAck_0n, sigAck_0n, rReqOr_0n);
  NOR2 I10 (rReqOr_0n, readReq_0n, readReq_1n);
  BALSA_TELEM I11 (trigger_0r, sigAck_0n, signal_0r, signal_0a);
  BUFF I12 (cd_0n, partCD_0n);
  OR2 I13 (partCD_0n, store_0n, store_1n);
  BUFF I14 (write_0r, trigger_0r);
endmodule

module BrzActiveEagerFalseVariable_3_3_s0_ (
  trigger_0r, trigger_0a,
  write_0r, write_0a0d, write_0a1d,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d,
  read_2r, read_2a0d, read_2a1d
);
  input trigger_0r;
  output trigger_0a;
  output write_0r;
  input [2:0] write_0a0d;
  input [2:0] write_0a1d;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output [2:0] read_0a0d;
  output [2:0] read_0a1d;
  input read_1r;
  output [2:0] read_1a0d;
  output [2:0] read_1a1d;
  input read_2r;
  output [2:0] read_2a0d;
  output [2:0] read_2a1d;
  wire cd_0n;
  wire [2:0] partCD_0n;
  wire [2:0] store_0n;
  wire [2:0] store_1n;
  wire readReq_0n;
  wire readReq_1n;
  wire readReq_2n;
  wire writeAck_0n;
  wire sigAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_2a1d[0], store_1n[0], readReq_2n);
  AND2 I1 (read_2a1d[1], store_1n[1], readReq_2n);
  AND2 I2 (read_2a1d[2], store_1n[2], readReq_2n);
  AND2 I3 (read_2a0d[0], store_0n[0], readReq_2n);
  AND2 I4 (read_2a0d[1], store_0n[1], readReq_2n);
  AND2 I5 (read_2a0d[2], store_0n[2], readReq_2n);
  AND2 I6 (read_1a1d[0], store_1n[0], readReq_1n);
  AND2 I7 (read_1a1d[1], store_1n[1], readReq_1n);
  AND2 I8 (read_1a1d[2], store_1n[2], readReq_1n);
  AND2 I9 (read_1a0d[0], store_0n[0], readReq_1n);
  AND2 I10 (read_1a0d[1], store_0n[1], readReq_1n);
  AND2 I11 (read_1a0d[2], store_0n[2], readReq_1n);
  AND2 I12 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I13 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I14 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I15 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I16 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I17 (read_0a0d[2], store_0n[2], readReq_0n);
  BUFF I18 (readReq_0n, read_0r);
  BUFF I19 (readReq_1n, read_1r);
  BUFF I20 (readReq_2n, read_2r);
  BUFF I21 (store_1n[0], write_0a1d[0]);
  BUFF I22 (store_1n[1], write_0a1d[1]);
  BUFF I23 (store_1n[2], write_0a1d[2]);
  BUFF I24 (store_0n[0], write_0a0d[0]);
  BUFF I25 (store_0n[1], write_0a0d[1]);
  BUFF I26 (store_0n[2], write_0a0d[2]);
  C2 I27 (trigger_0a, writeAck_0n, cd_0n);
  AND2 I28 (writeAck_0n, sigAck_0n, rReqOr_0n);
  NOR3 I29 (rReqOr_0n, readReq_0n, readReq_1n, readReq_2n);
  BALSA_TELEM I30 (trigger_0r, sigAck_0n, signal_0r, signal_0a);
  C3 I31 (cd_0n, partCD_0n[0], partCD_0n[1], partCD_0n[2]);
  OR2 I32 (partCD_0n[0], store_0n[0], store_1n[0]);
  OR2 I33 (partCD_0n[1], store_0n[1], store_1n[1]);
  OR2 I34 (partCD_0n[2], store_0n[2], store_1n[2]);
  BUFF I35 (write_0r, trigger_0r);
endmodule

module BrzActiveEagerFalseVariable_3_3_s22__3b2_2_m1m (
  trigger_0r, trigger_0a,
  write_0r, write_0a0d, write_0a1d,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d,
  read_2r, read_2a0d, read_2a1d
);
  input trigger_0r;
  output trigger_0a;
  output write_0r;
  input [2:0] write_0a0d;
  input [2:0] write_0a1d;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output [2:0] read_0a0d;
  output [2:0] read_0a1d;
  input read_1r;
  output read_1a0d;
  output read_1a1d;
  input read_2r;
  output read_2a0d;
  output read_2a1d;
  wire cd_0n;
  wire [2:0] partCD_0n;
  wire [2:0] store_0n;
  wire [2:0] store_1n;
  wire readReq_0n;
  wire readReq_1n;
  wire readReq_2n;
  wire writeAck_0n;
  wire sigAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_2a1d, store_1n[0], readReq_2n);
  AND2 I1 (read_2a0d, store_0n[0], readReq_2n);
  AND2 I2 (read_1a1d, store_1n[2], readReq_1n);
  AND2 I3 (read_1a0d, store_0n[2], readReq_1n);
  AND2 I4 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I5 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I6 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I7 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I8 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I9 (read_0a0d[2], store_0n[2], readReq_0n);
  BUFF I10 (readReq_0n, read_0r);
  BUFF I11 (readReq_1n, read_1r);
  BUFF I12 (readReq_2n, read_2r);
  BUFF I13 (store_1n[0], write_0a1d[0]);
  BUFF I14 (store_1n[1], write_0a1d[1]);
  BUFF I15 (store_1n[2], write_0a1d[2]);
  BUFF I16 (store_0n[0], write_0a0d[0]);
  BUFF I17 (store_0n[1], write_0a0d[1]);
  BUFF I18 (store_0n[2], write_0a0d[2]);
  C2 I19 (trigger_0a, writeAck_0n, cd_0n);
  AND2 I20 (writeAck_0n, sigAck_0n, rReqOr_0n);
  NOR3 I21 (rReqOr_0n, readReq_0n, readReq_1n, readReq_2n);
  BALSA_TELEM I22 (trigger_0r, sigAck_0n, signal_0r, signal_0a);
  C3 I23 (cd_0n, partCD_0n[0], partCD_0n[1], partCD_0n[2]);
  OR2 I24 (partCD_0n[0], store_0n[0], store_1n[0]);
  OR2 I25 (partCD_0n[1], store_0n[1], store_1n[1]);
  OR2 I26 (partCD_0n[2], store_0n[2], store_1n[2]);
  BUFF I27 (write_0r, trigger_0r);
endmodule

module BrzActiveEagerFalseVariable_32_1_s0_ (
  trigger_0r, trigger_0a,
  write_0r, write_0a0d, write_0a1d,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d
);
  input trigger_0r;
  output trigger_0a;
  output write_0r;
  input [31:0] write_0a0d;
  input [31:0] write_0a1d;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output [31:0] read_0a0d;
  output [31:0] read_0a1d;
  wire [16:0] internal_0n;
  wire cd_0n;
  wire [31:0] partCD_0n;
  wire [31:0] store_0n;
  wire [31:0] store_1n;
  wire readReq_0n;
  wire writeAck_0n;
  wire sigAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I1 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I2 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I3 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I4 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I5 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I6 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I7 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I8 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I9 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I10 (read_0a1d[10], store_1n[10], readReq_0n);
  AND2 I11 (read_0a1d[11], store_1n[11], readReq_0n);
  AND2 I12 (read_0a1d[12], store_1n[12], readReq_0n);
  AND2 I13 (read_0a1d[13], store_1n[13], readReq_0n);
  AND2 I14 (read_0a1d[14], store_1n[14], readReq_0n);
  AND2 I15 (read_0a1d[15], store_1n[15], readReq_0n);
  AND2 I16 (read_0a1d[16], store_1n[16], readReq_0n);
  AND2 I17 (read_0a1d[17], store_1n[17], readReq_0n);
  AND2 I18 (read_0a1d[18], store_1n[18], readReq_0n);
  AND2 I19 (read_0a1d[19], store_1n[19], readReq_0n);
  AND2 I20 (read_0a1d[20], store_1n[20], readReq_0n);
  AND2 I21 (read_0a1d[21], store_1n[21], readReq_0n);
  AND2 I22 (read_0a1d[22], store_1n[22], readReq_0n);
  AND2 I23 (read_0a1d[23], store_1n[23], readReq_0n);
  AND2 I24 (read_0a1d[24], store_1n[24], readReq_0n);
  AND2 I25 (read_0a1d[25], store_1n[25], readReq_0n);
  AND2 I26 (read_0a1d[26], store_1n[26], readReq_0n);
  AND2 I27 (read_0a1d[27], store_1n[27], readReq_0n);
  AND2 I28 (read_0a1d[28], store_1n[28], readReq_0n);
  AND2 I29 (read_0a1d[29], store_1n[29], readReq_0n);
  AND2 I30 (read_0a1d[30], store_1n[30], readReq_0n);
  AND2 I31 (read_0a1d[31], store_1n[31], readReq_0n);
  AND2 I32 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I33 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I34 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I35 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I36 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I37 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I38 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I39 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I40 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I41 (read_0a0d[9], store_0n[9], readReq_0n);
  AND2 I42 (read_0a0d[10], store_0n[10], readReq_0n);
  AND2 I43 (read_0a0d[11], store_0n[11], readReq_0n);
  AND2 I44 (read_0a0d[12], store_0n[12], readReq_0n);
  AND2 I45 (read_0a0d[13], store_0n[13], readReq_0n);
  AND2 I46 (read_0a0d[14], store_0n[14], readReq_0n);
  AND2 I47 (read_0a0d[15], store_0n[15], readReq_0n);
  AND2 I48 (read_0a0d[16], store_0n[16], readReq_0n);
  AND2 I49 (read_0a0d[17], store_0n[17], readReq_0n);
  AND2 I50 (read_0a0d[18], store_0n[18], readReq_0n);
  AND2 I51 (read_0a0d[19], store_0n[19], readReq_0n);
  AND2 I52 (read_0a0d[20], store_0n[20], readReq_0n);
  AND2 I53 (read_0a0d[21], store_0n[21], readReq_0n);
  AND2 I54 (read_0a0d[22], store_0n[22], readReq_0n);
  AND2 I55 (read_0a0d[23], store_0n[23], readReq_0n);
  AND2 I56 (read_0a0d[24], store_0n[24], readReq_0n);
  AND2 I57 (read_0a0d[25], store_0n[25], readReq_0n);
  AND2 I58 (read_0a0d[26], store_0n[26], readReq_0n);
  AND2 I59 (read_0a0d[27], store_0n[27], readReq_0n);
  AND2 I60 (read_0a0d[28], store_0n[28], readReq_0n);
  AND2 I61 (read_0a0d[29], store_0n[29], readReq_0n);
  AND2 I62 (read_0a0d[30], store_0n[30], readReq_0n);
  AND2 I63 (read_0a0d[31], store_0n[31], readReq_0n);
  BUFF I64 (readReq_0n, read_0r);
  BUFF I65 (store_1n[0], write_0a1d[0]);
  BUFF I66 (store_1n[1], write_0a1d[1]);
  BUFF I67 (store_1n[2], write_0a1d[2]);
  BUFF I68 (store_1n[3], write_0a1d[3]);
  BUFF I69 (store_1n[4], write_0a1d[4]);
  BUFF I70 (store_1n[5], write_0a1d[5]);
  BUFF I71 (store_1n[6], write_0a1d[6]);
  BUFF I72 (store_1n[7], write_0a1d[7]);
  BUFF I73 (store_1n[8], write_0a1d[8]);
  BUFF I74 (store_1n[9], write_0a1d[9]);
  BUFF I75 (store_1n[10], write_0a1d[10]);
  BUFF I76 (store_1n[11], write_0a1d[11]);
  BUFF I77 (store_1n[12], write_0a1d[12]);
  BUFF I78 (store_1n[13], write_0a1d[13]);
  BUFF I79 (store_1n[14], write_0a1d[14]);
  BUFF I80 (store_1n[15], write_0a1d[15]);
  BUFF I81 (store_1n[16], write_0a1d[16]);
  BUFF I82 (store_1n[17], write_0a1d[17]);
  BUFF I83 (store_1n[18], write_0a1d[18]);
  BUFF I84 (store_1n[19], write_0a1d[19]);
  BUFF I85 (store_1n[20], write_0a1d[20]);
  BUFF I86 (store_1n[21], write_0a1d[21]);
  BUFF I87 (store_1n[22], write_0a1d[22]);
  BUFF I88 (store_1n[23], write_0a1d[23]);
  BUFF I89 (store_1n[24], write_0a1d[24]);
  BUFF I90 (store_1n[25], write_0a1d[25]);
  BUFF I91 (store_1n[26], write_0a1d[26]);
  BUFF I92 (store_1n[27], write_0a1d[27]);
  BUFF I93 (store_1n[28], write_0a1d[28]);
  BUFF I94 (store_1n[29], write_0a1d[29]);
  BUFF I95 (store_1n[30], write_0a1d[30]);
  BUFF I96 (store_1n[31], write_0a1d[31]);
  BUFF I97 (store_0n[0], write_0a0d[0]);
  BUFF I98 (store_0n[1], write_0a0d[1]);
  BUFF I99 (store_0n[2], write_0a0d[2]);
  BUFF I100 (store_0n[3], write_0a0d[3]);
  BUFF I101 (store_0n[4], write_0a0d[4]);
  BUFF I102 (store_0n[5], write_0a0d[5]);
  BUFF I103 (store_0n[6], write_0a0d[6]);
  BUFF I104 (store_0n[7], write_0a0d[7]);
  BUFF I105 (store_0n[8], write_0a0d[8]);
  BUFF I106 (store_0n[9], write_0a0d[9]);
  BUFF I107 (store_0n[10], write_0a0d[10]);
  BUFF I108 (store_0n[11], write_0a0d[11]);
  BUFF I109 (store_0n[12], write_0a0d[12]);
  BUFF I110 (store_0n[13], write_0a0d[13]);
  BUFF I111 (store_0n[14], write_0a0d[14]);
  BUFF I112 (store_0n[15], write_0a0d[15]);
  BUFF I113 (store_0n[16], write_0a0d[16]);
  BUFF I114 (store_0n[17], write_0a0d[17]);
  BUFF I115 (store_0n[18], write_0a0d[18]);
  BUFF I116 (store_0n[19], write_0a0d[19]);
  BUFF I117 (store_0n[20], write_0a0d[20]);
  BUFF I118 (store_0n[21], write_0a0d[21]);
  BUFF I119 (store_0n[22], write_0a0d[22]);
  BUFF I120 (store_0n[23], write_0a0d[23]);
  BUFF I121 (store_0n[24], write_0a0d[24]);
  BUFF I122 (store_0n[25], write_0a0d[25]);
  BUFF I123 (store_0n[26], write_0a0d[26]);
  BUFF I124 (store_0n[27], write_0a0d[27]);
  BUFF I125 (store_0n[28], write_0a0d[28]);
  BUFF I126 (store_0n[29], write_0a0d[29]);
  BUFF I127 (store_0n[30], write_0a0d[30]);
  BUFF I128 (store_0n[31], write_0a0d[31]);
  C2 I129 (trigger_0a, writeAck_0n, cd_0n);
  AND2 I130 (writeAck_0n, sigAck_0n, rReqOr_0n);
  INV I131 (rReqOr_0n, readReq_0n);
  BALSA_TELEM I132 (trigger_0r, sigAck_0n, signal_0r, signal_0a);
  C3 I133 (internal_0n[0], partCD_0n[0], partCD_0n[1], partCD_0n[2]);
  C3 I134 (internal_0n[1], partCD_0n[3], partCD_0n[4], partCD_0n[5]);
  C3 I135 (internal_0n[2], partCD_0n[6], partCD_0n[7], partCD_0n[8]);
  C3 I136 (internal_0n[3], partCD_0n[9], partCD_0n[10], partCD_0n[11]);
  C3 I137 (internal_0n[4], partCD_0n[12], partCD_0n[13], partCD_0n[14]);
  C3 I138 (internal_0n[5], partCD_0n[15], partCD_0n[16], partCD_0n[17]);
  C3 I139 (internal_0n[6], partCD_0n[18], partCD_0n[19], partCD_0n[20]);
  C3 I140 (internal_0n[7], partCD_0n[21], partCD_0n[22], partCD_0n[23]);
  C3 I141 (internal_0n[8], partCD_0n[24], partCD_0n[25], partCD_0n[26]);
  C3 I142 (internal_0n[9], partCD_0n[27], partCD_0n[28], partCD_0n[29]);
  C2 I143 (internal_0n[10], partCD_0n[30], partCD_0n[31]);
  C3 I144 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I145 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I146 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I147 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I148 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I149 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I150 (cd_0n, internal_0n[15], internal_0n[16]);
  OR2 I151 (partCD_0n[0], store_0n[0], store_1n[0]);
  OR2 I152 (partCD_0n[1], store_0n[1], store_1n[1]);
  OR2 I153 (partCD_0n[2], store_0n[2], store_1n[2]);
  OR2 I154 (partCD_0n[3], store_0n[3], store_1n[3]);
  OR2 I155 (partCD_0n[4], store_0n[4], store_1n[4]);
  OR2 I156 (partCD_0n[5], store_0n[5], store_1n[5]);
  OR2 I157 (partCD_0n[6], store_0n[6], store_1n[6]);
  OR2 I158 (partCD_0n[7], store_0n[7], store_1n[7]);
  OR2 I159 (partCD_0n[8], store_0n[8], store_1n[8]);
  OR2 I160 (partCD_0n[9], store_0n[9], store_1n[9]);
  OR2 I161 (partCD_0n[10], store_0n[10], store_1n[10]);
  OR2 I162 (partCD_0n[11], store_0n[11], store_1n[11]);
  OR2 I163 (partCD_0n[12], store_0n[12], store_1n[12]);
  OR2 I164 (partCD_0n[13], store_0n[13], store_1n[13]);
  OR2 I165 (partCD_0n[14], store_0n[14], store_1n[14]);
  OR2 I166 (partCD_0n[15], store_0n[15], store_1n[15]);
  OR2 I167 (partCD_0n[16], store_0n[16], store_1n[16]);
  OR2 I168 (partCD_0n[17], store_0n[17], store_1n[17]);
  OR2 I169 (partCD_0n[18], store_0n[18], store_1n[18]);
  OR2 I170 (partCD_0n[19], store_0n[19], store_1n[19]);
  OR2 I171 (partCD_0n[20], store_0n[20], store_1n[20]);
  OR2 I172 (partCD_0n[21], store_0n[21], store_1n[21]);
  OR2 I173 (partCD_0n[22], store_0n[22], store_1n[22]);
  OR2 I174 (partCD_0n[23], store_0n[23], store_1n[23]);
  OR2 I175 (partCD_0n[24], store_0n[24], store_1n[24]);
  OR2 I176 (partCD_0n[25], store_0n[25], store_1n[25]);
  OR2 I177 (partCD_0n[26], store_0n[26], store_1n[26]);
  OR2 I178 (partCD_0n[27], store_0n[27], store_1n[27]);
  OR2 I179 (partCD_0n[28], store_0n[28], store_1n[28]);
  OR2 I180 (partCD_0n[29], store_0n[29], store_1n[29]);
  OR2 I181 (partCD_0n[30], store_0n[30], store_1n[30]);
  OR2 I182 (partCD_0n[31], store_0n[31], store_1n[31]);
  BUFF I183 (write_0r, trigger_0r);
endmodule

module BrzActiveEagerFalseVariable_32_2_s0_ (
  trigger_0r, trigger_0a,
  write_0r, write_0a0d, write_0a1d,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d
);
  input trigger_0r;
  output trigger_0a;
  output write_0r;
  input [31:0] write_0a0d;
  input [31:0] write_0a1d;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output [31:0] read_0a0d;
  output [31:0] read_0a1d;
  input read_1r;
  output [31:0] read_1a0d;
  output [31:0] read_1a1d;
  wire [16:0] internal_0n;
  wire cd_0n;
  wire [31:0] partCD_0n;
  wire [31:0] store_0n;
  wire [31:0] store_1n;
  wire readReq_0n;
  wire readReq_1n;
  wire writeAck_0n;
  wire sigAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_1a1d[0], store_1n[0], readReq_1n);
  AND2 I1 (read_1a1d[1], store_1n[1], readReq_1n);
  AND2 I2 (read_1a1d[2], store_1n[2], readReq_1n);
  AND2 I3 (read_1a1d[3], store_1n[3], readReq_1n);
  AND2 I4 (read_1a1d[4], store_1n[4], readReq_1n);
  AND2 I5 (read_1a1d[5], store_1n[5], readReq_1n);
  AND2 I6 (read_1a1d[6], store_1n[6], readReq_1n);
  AND2 I7 (read_1a1d[7], store_1n[7], readReq_1n);
  AND2 I8 (read_1a1d[8], store_1n[8], readReq_1n);
  AND2 I9 (read_1a1d[9], store_1n[9], readReq_1n);
  AND2 I10 (read_1a1d[10], store_1n[10], readReq_1n);
  AND2 I11 (read_1a1d[11], store_1n[11], readReq_1n);
  AND2 I12 (read_1a1d[12], store_1n[12], readReq_1n);
  AND2 I13 (read_1a1d[13], store_1n[13], readReq_1n);
  AND2 I14 (read_1a1d[14], store_1n[14], readReq_1n);
  AND2 I15 (read_1a1d[15], store_1n[15], readReq_1n);
  AND2 I16 (read_1a1d[16], store_1n[16], readReq_1n);
  AND2 I17 (read_1a1d[17], store_1n[17], readReq_1n);
  AND2 I18 (read_1a1d[18], store_1n[18], readReq_1n);
  AND2 I19 (read_1a1d[19], store_1n[19], readReq_1n);
  AND2 I20 (read_1a1d[20], store_1n[20], readReq_1n);
  AND2 I21 (read_1a1d[21], store_1n[21], readReq_1n);
  AND2 I22 (read_1a1d[22], store_1n[22], readReq_1n);
  AND2 I23 (read_1a1d[23], store_1n[23], readReq_1n);
  AND2 I24 (read_1a1d[24], store_1n[24], readReq_1n);
  AND2 I25 (read_1a1d[25], store_1n[25], readReq_1n);
  AND2 I26 (read_1a1d[26], store_1n[26], readReq_1n);
  AND2 I27 (read_1a1d[27], store_1n[27], readReq_1n);
  AND2 I28 (read_1a1d[28], store_1n[28], readReq_1n);
  AND2 I29 (read_1a1d[29], store_1n[29], readReq_1n);
  AND2 I30 (read_1a1d[30], store_1n[30], readReq_1n);
  AND2 I31 (read_1a1d[31], store_1n[31], readReq_1n);
  AND2 I32 (read_1a0d[0], store_0n[0], readReq_1n);
  AND2 I33 (read_1a0d[1], store_0n[1], readReq_1n);
  AND2 I34 (read_1a0d[2], store_0n[2], readReq_1n);
  AND2 I35 (read_1a0d[3], store_0n[3], readReq_1n);
  AND2 I36 (read_1a0d[4], store_0n[4], readReq_1n);
  AND2 I37 (read_1a0d[5], store_0n[5], readReq_1n);
  AND2 I38 (read_1a0d[6], store_0n[6], readReq_1n);
  AND2 I39 (read_1a0d[7], store_0n[7], readReq_1n);
  AND2 I40 (read_1a0d[8], store_0n[8], readReq_1n);
  AND2 I41 (read_1a0d[9], store_0n[9], readReq_1n);
  AND2 I42 (read_1a0d[10], store_0n[10], readReq_1n);
  AND2 I43 (read_1a0d[11], store_0n[11], readReq_1n);
  AND2 I44 (read_1a0d[12], store_0n[12], readReq_1n);
  AND2 I45 (read_1a0d[13], store_0n[13], readReq_1n);
  AND2 I46 (read_1a0d[14], store_0n[14], readReq_1n);
  AND2 I47 (read_1a0d[15], store_0n[15], readReq_1n);
  AND2 I48 (read_1a0d[16], store_0n[16], readReq_1n);
  AND2 I49 (read_1a0d[17], store_0n[17], readReq_1n);
  AND2 I50 (read_1a0d[18], store_0n[18], readReq_1n);
  AND2 I51 (read_1a0d[19], store_0n[19], readReq_1n);
  AND2 I52 (read_1a0d[20], store_0n[20], readReq_1n);
  AND2 I53 (read_1a0d[21], store_0n[21], readReq_1n);
  AND2 I54 (read_1a0d[22], store_0n[22], readReq_1n);
  AND2 I55 (read_1a0d[23], store_0n[23], readReq_1n);
  AND2 I56 (read_1a0d[24], store_0n[24], readReq_1n);
  AND2 I57 (read_1a0d[25], store_0n[25], readReq_1n);
  AND2 I58 (read_1a0d[26], store_0n[26], readReq_1n);
  AND2 I59 (read_1a0d[27], store_0n[27], readReq_1n);
  AND2 I60 (read_1a0d[28], store_0n[28], readReq_1n);
  AND2 I61 (read_1a0d[29], store_0n[29], readReq_1n);
  AND2 I62 (read_1a0d[30], store_0n[30], readReq_1n);
  AND2 I63 (read_1a0d[31], store_0n[31], readReq_1n);
  AND2 I64 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I65 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I66 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I67 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I68 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I69 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I70 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I71 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I72 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I73 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I74 (read_0a1d[10], store_1n[10], readReq_0n);
  AND2 I75 (read_0a1d[11], store_1n[11], readReq_0n);
  AND2 I76 (read_0a1d[12], store_1n[12], readReq_0n);
  AND2 I77 (read_0a1d[13], store_1n[13], readReq_0n);
  AND2 I78 (read_0a1d[14], store_1n[14], readReq_0n);
  AND2 I79 (read_0a1d[15], store_1n[15], readReq_0n);
  AND2 I80 (read_0a1d[16], store_1n[16], readReq_0n);
  AND2 I81 (read_0a1d[17], store_1n[17], readReq_0n);
  AND2 I82 (read_0a1d[18], store_1n[18], readReq_0n);
  AND2 I83 (read_0a1d[19], store_1n[19], readReq_0n);
  AND2 I84 (read_0a1d[20], store_1n[20], readReq_0n);
  AND2 I85 (read_0a1d[21], store_1n[21], readReq_0n);
  AND2 I86 (read_0a1d[22], store_1n[22], readReq_0n);
  AND2 I87 (read_0a1d[23], store_1n[23], readReq_0n);
  AND2 I88 (read_0a1d[24], store_1n[24], readReq_0n);
  AND2 I89 (read_0a1d[25], store_1n[25], readReq_0n);
  AND2 I90 (read_0a1d[26], store_1n[26], readReq_0n);
  AND2 I91 (read_0a1d[27], store_1n[27], readReq_0n);
  AND2 I92 (read_0a1d[28], store_1n[28], readReq_0n);
  AND2 I93 (read_0a1d[29], store_1n[29], readReq_0n);
  AND2 I94 (read_0a1d[30], store_1n[30], readReq_0n);
  AND2 I95 (read_0a1d[31], store_1n[31], readReq_0n);
  AND2 I96 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I97 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I98 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I99 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I100 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I101 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I102 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I103 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I104 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I105 (read_0a0d[9], store_0n[9], readReq_0n);
  AND2 I106 (read_0a0d[10], store_0n[10], readReq_0n);
  AND2 I107 (read_0a0d[11], store_0n[11], readReq_0n);
  AND2 I108 (read_0a0d[12], store_0n[12], readReq_0n);
  AND2 I109 (read_0a0d[13], store_0n[13], readReq_0n);
  AND2 I110 (read_0a0d[14], store_0n[14], readReq_0n);
  AND2 I111 (read_0a0d[15], store_0n[15], readReq_0n);
  AND2 I112 (read_0a0d[16], store_0n[16], readReq_0n);
  AND2 I113 (read_0a0d[17], store_0n[17], readReq_0n);
  AND2 I114 (read_0a0d[18], store_0n[18], readReq_0n);
  AND2 I115 (read_0a0d[19], store_0n[19], readReq_0n);
  AND2 I116 (read_0a0d[20], store_0n[20], readReq_0n);
  AND2 I117 (read_0a0d[21], store_0n[21], readReq_0n);
  AND2 I118 (read_0a0d[22], store_0n[22], readReq_0n);
  AND2 I119 (read_0a0d[23], store_0n[23], readReq_0n);
  AND2 I120 (read_0a0d[24], store_0n[24], readReq_0n);
  AND2 I121 (read_0a0d[25], store_0n[25], readReq_0n);
  AND2 I122 (read_0a0d[26], store_0n[26], readReq_0n);
  AND2 I123 (read_0a0d[27], store_0n[27], readReq_0n);
  AND2 I124 (read_0a0d[28], store_0n[28], readReq_0n);
  AND2 I125 (read_0a0d[29], store_0n[29], readReq_0n);
  AND2 I126 (read_0a0d[30], store_0n[30], readReq_0n);
  AND2 I127 (read_0a0d[31], store_0n[31], readReq_0n);
  BUFF I128 (readReq_0n, read_0r);
  BUFF I129 (readReq_1n, read_1r);
  BUFF I130 (store_1n[0], write_0a1d[0]);
  BUFF I131 (store_1n[1], write_0a1d[1]);
  BUFF I132 (store_1n[2], write_0a1d[2]);
  BUFF I133 (store_1n[3], write_0a1d[3]);
  BUFF I134 (store_1n[4], write_0a1d[4]);
  BUFF I135 (store_1n[5], write_0a1d[5]);
  BUFF I136 (store_1n[6], write_0a1d[6]);
  BUFF I137 (store_1n[7], write_0a1d[7]);
  BUFF I138 (store_1n[8], write_0a1d[8]);
  BUFF I139 (store_1n[9], write_0a1d[9]);
  BUFF I140 (store_1n[10], write_0a1d[10]);
  BUFF I141 (store_1n[11], write_0a1d[11]);
  BUFF I142 (store_1n[12], write_0a1d[12]);
  BUFF I143 (store_1n[13], write_0a1d[13]);
  BUFF I144 (store_1n[14], write_0a1d[14]);
  BUFF I145 (store_1n[15], write_0a1d[15]);
  BUFF I146 (store_1n[16], write_0a1d[16]);
  BUFF I147 (store_1n[17], write_0a1d[17]);
  BUFF I148 (store_1n[18], write_0a1d[18]);
  BUFF I149 (store_1n[19], write_0a1d[19]);
  BUFF I150 (store_1n[20], write_0a1d[20]);
  BUFF I151 (store_1n[21], write_0a1d[21]);
  BUFF I152 (store_1n[22], write_0a1d[22]);
  BUFF I153 (store_1n[23], write_0a1d[23]);
  BUFF I154 (store_1n[24], write_0a1d[24]);
  BUFF I155 (store_1n[25], write_0a1d[25]);
  BUFF I156 (store_1n[26], write_0a1d[26]);
  BUFF I157 (store_1n[27], write_0a1d[27]);
  BUFF I158 (store_1n[28], write_0a1d[28]);
  BUFF I159 (store_1n[29], write_0a1d[29]);
  BUFF I160 (store_1n[30], write_0a1d[30]);
  BUFF I161 (store_1n[31], write_0a1d[31]);
  BUFF I162 (store_0n[0], write_0a0d[0]);
  BUFF I163 (store_0n[1], write_0a0d[1]);
  BUFF I164 (store_0n[2], write_0a0d[2]);
  BUFF I165 (store_0n[3], write_0a0d[3]);
  BUFF I166 (store_0n[4], write_0a0d[4]);
  BUFF I167 (store_0n[5], write_0a0d[5]);
  BUFF I168 (store_0n[6], write_0a0d[6]);
  BUFF I169 (store_0n[7], write_0a0d[7]);
  BUFF I170 (store_0n[8], write_0a0d[8]);
  BUFF I171 (store_0n[9], write_0a0d[9]);
  BUFF I172 (store_0n[10], write_0a0d[10]);
  BUFF I173 (store_0n[11], write_0a0d[11]);
  BUFF I174 (store_0n[12], write_0a0d[12]);
  BUFF I175 (store_0n[13], write_0a0d[13]);
  BUFF I176 (store_0n[14], write_0a0d[14]);
  BUFF I177 (store_0n[15], write_0a0d[15]);
  BUFF I178 (store_0n[16], write_0a0d[16]);
  BUFF I179 (store_0n[17], write_0a0d[17]);
  BUFF I180 (store_0n[18], write_0a0d[18]);
  BUFF I181 (store_0n[19], write_0a0d[19]);
  BUFF I182 (store_0n[20], write_0a0d[20]);
  BUFF I183 (store_0n[21], write_0a0d[21]);
  BUFF I184 (store_0n[22], write_0a0d[22]);
  BUFF I185 (store_0n[23], write_0a0d[23]);
  BUFF I186 (store_0n[24], write_0a0d[24]);
  BUFF I187 (store_0n[25], write_0a0d[25]);
  BUFF I188 (store_0n[26], write_0a0d[26]);
  BUFF I189 (store_0n[27], write_0a0d[27]);
  BUFF I190 (store_0n[28], write_0a0d[28]);
  BUFF I191 (store_0n[29], write_0a0d[29]);
  BUFF I192 (store_0n[30], write_0a0d[30]);
  BUFF I193 (store_0n[31], write_0a0d[31]);
  C2 I194 (trigger_0a, writeAck_0n, cd_0n);
  AND2 I195 (writeAck_0n, sigAck_0n, rReqOr_0n);
  NOR2 I196 (rReqOr_0n, readReq_0n, readReq_1n);
  BALSA_TELEM I197 (trigger_0r, sigAck_0n, signal_0r, signal_0a);
  C3 I198 (internal_0n[0], partCD_0n[0], partCD_0n[1], partCD_0n[2]);
  C3 I199 (internal_0n[1], partCD_0n[3], partCD_0n[4], partCD_0n[5]);
  C3 I200 (internal_0n[2], partCD_0n[6], partCD_0n[7], partCD_0n[8]);
  C3 I201 (internal_0n[3], partCD_0n[9], partCD_0n[10], partCD_0n[11]);
  C3 I202 (internal_0n[4], partCD_0n[12], partCD_0n[13], partCD_0n[14]);
  C3 I203 (internal_0n[5], partCD_0n[15], partCD_0n[16], partCD_0n[17]);
  C3 I204 (internal_0n[6], partCD_0n[18], partCD_0n[19], partCD_0n[20]);
  C3 I205 (internal_0n[7], partCD_0n[21], partCD_0n[22], partCD_0n[23]);
  C3 I206 (internal_0n[8], partCD_0n[24], partCD_0n[25], partCD_0n[26]);
  C3 I207 (internal_0n[9], partCD_0n[27], partCD_0n[28], partCD_0n[29]);
  C2 I208 (internal_0n[10], partCD_0n[30], partCD_0n[31]);
  C3 I209 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I210 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I211 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I212 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I213 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I214 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I215 (cd_0n, internal_0n[15], internal_0n[16]);
  OR2 I216 (partCD_0n[0], store_0n[0], store_1n[0]);
  OR2 I217 (partCD_0n[1], store_0n[1], store_1n[1]);
  OR2 I218 (partCD_0n[2], store_0n[2], store_1n[2]);
  OR2 I219 (partCD_0n[3], store_0n[3], store_1n[3]);
  OR2 I220 (partCD_0n[4], store_0n[4], store_1n[4]);
  OR2 I221 (partCD_0n[5], store_0n[5], store_1n[5]);
  OR2 I222 (partCD_0n[6], store_0n[6], store_1n[6]);
  OR2 I223 (partCD_0n[7], store_0n[7], store_1n[7]);
  OR2 I224 (partCD_0n[8], store_0n[8], store_1n[8]);
  OR2 I225 (partCD_0n[9], store_0n[9], store_1n[9]);
  OR2 I226 (partCD_0n[10], store_0n[10], store_1n[10]);
  OR2 I227 (partCD_0n[11], store_0n[11], store_1n[11]);
  OR2 I228 (partCD_0n[12], store_0n[12], store_1n[12]);
  OR2 I229 (partCD_0n[13], store_0n[13], store_1n[13]);
  OR2 I230 (partCD_0n[14], store_0n[14], store_1n[14]);
  OR2 I231 (partCD_0n[15], store_0n[15], store_1n[15]);
  OR2 I232 (partCD_0n[16], store_0n[16], store_1n[16]);
  OR2 I233 (partCD_0n[17], store_0n[17], store_1n[17]);
  OR2 I234 (partCD_0n[18], store_0n[18], store_1n[18]);
  OR2 I235 (partCD_0n[19], store_0n[19], store_1n[19]);
  OR2 I236 (partCD_0n[20], store_0n[20], store_1n[20]);
  OR2 I237 (partCD_0n[21], store_0n[21], store_1n[21]);
  OR2 I238 (partCD_0n[22], store_0n[22], store_1n[22]);
  OR2 I239 (partCD_0n[23], store_0n[23], store_1n[23]);
  OR2 I240 (partCD_0n[24], store_0n[24], store_1n[24]);
  OR2 I241 (partCD_0n[25], store_0n[25], store_1n[25]);
  OR2 I242 (partCD_0n[26], store_0n[26], store_1n[26]);
  OR2 I243 (partCD_0n[27], store_0n[27], store_1n[27]);
  OR2 I244 (partCD_0n[28], store_0n[28], store_1n[28]);
  OR2 I245 (partCD_0n[29], store_0n[29], store_1n[29]);
  OR2 I246 (partCD_0n[30], store_0n[30], store_1n[30]);
  OR2 I247 (partCD_0n[31], store_0n[31], store_1n[31]);
  BUFF I248 (write_0r, trigger_0r);
endmodule

module BrzActiveEagerFalseVariable_32_3_s13__3b31_m3m (
  trigger_0r, trigger_0a,
  write_0r, write_0a0d, write_0a1d,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d,
  read_2r, read_2a0d, read_2a1d
);
  input trigger_0r;
  output trigger_0a;
  output write_0r;
  input [31:0] write_0a0d;
  input [31:0] write_0a1d;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output [31:0] read_0a0d;
  output [31:0] read_0a1d;
  input read_1r;
  output read_1a0d;
  output read_1a1d;
  input read_2r;
  output [31:0] read_2a0d;
  output [31:0] read_2a1d;
  wire [16:0] internal_0n;
  wire cd_0n;
  wire [31:0] partCD_0n;
  wire [31:0] store_0n;
  wire [31:0] store_1n;
  wire readReq_0n;
  wire readReq_1n;
  wire readReq_2n;
  wire writeAck_0n;
  wire sigAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_2a1d[0], store_1n[0], readReq_2n);
  AND2 I1 (read_2a1d[1], store_1n[1], readReq_2n);
  AND2 I2 (read_2a1d[2], store_1n[2], readReq_2n);
  AND2 I3 (read_2a1d[3], store_1n[3], readReq_2n);
  AND2 I4 (read_2a1d[4], store_1n[4], readReq_2n);
  AND2 I5 (read_2a1d[5], store_1n[5], readReq_2n);
  AND2 I6 (read_2a1d[6], store_1n[6], readReq_2n);
  AND2 I7 (read_2a1d[7], store_1n[7], readReq_2n);
  AND2 I8 (read_2a1d[8], store_1n[8], readReq_2n);
  AND2 I9 (read_2a1d[9], store_1n[9], readReq_2n);
  AND2 I10 (read_2a1d[10], store_1n[10], readReq_2n);
  AND2 I11 (read_2a1d[11], store_1n[11], readReq_2n);
  AND2 I12 (read_2a1d[12], store_1n[12], readReq_2n);
  AND2 I13 (read_2a1d[13], store_1n[13], readReq_2n);
  AND2 I14 (read_2a1d[14], store_1n[14], readReq_2n);
  AND2 I15 (read_2a1d[15], store_1n[15], readReq_2n);
  AND2 I16 (read_2a1d[16], store_1n[16], readReq_2n);
  AND2 I17 (read_2a1d[17], store_1n[17], readReq_2n);
  AND2 I18 (read_2a1d[18], store_1n[18], readReq_2n);
  AND2 I19 (read_2a1d[19], store_1n[19], readReq_2n);
  AND2 I20 (read_2a1d[20], store_1n[20], readReq_2n);
  AND2 I21 (read_2a1d[21], store_1n[21], readReq_2n);
  AND2 I22 (read_2a1d[22], store_1n[22], readReq_2n);
  AND2 I23 (read_2a1d[23], store_1n[23], readReq_2n);
  AND2 I24 (read_2a1d[24], store_1n[24], readReq_2n);
  AND2 I25 (read_2a1d[25], store_1n[25], readReq_2n);
  AND2 I26 (read_2a1d[26], store_1n[26], readReq_2n);
  AND2 I27 (read_2a1d[27], store_1n[27], readReq_2n);
  AND2 I28 (read_2a1d[28], store_1n[28], readReq_2n);
  AND2 I29 (read_2a1d[29], store_1n[29], readReq_2n);
  AND2 I30 (read_2a1d[30], store_1n[30], readReq_2n);
  AND2 I31 (read_2a1d[31], store_1n[31], readReq_2n);
  AND2 I32 (read_2a0d[0], store_0n[0], readReq_2n);
  AND2 I33 (read_2a0d[1], store_0n[1], readReq_2n);
  AND2 I34 (read_2a0d[2], store_0n[2], readReq_2n);
  AND2 I35 (read_2a0d[3], store_0n[3], readReq_2n);
  AND2 I36 (read_2a0d[4], store_0n[4], readReq_2n);
  AND2 I37 (read_2a0d[5], store_0n[5], readReq_2n);
  AND2 I38 (read_2a0d[6], store_0n[6], readReq_2n);
  AND2 I39 (read_2a0d[7], store_0n[7], readReq_2n);
  AND2 I40 (read_2a0d[8], store_0n[8], readReq_2n);
  AND2 I41 (read_2a0d[9], store_0n[9], readReq_2n);
  AND2 I42 (read_2a0d[10], store_0n[10], readReq_2n);
  AND2 I43 (read_2a0d[11], store_0n[11], readReq_2n);
  AND2 I44 (read_2a0d[12], store_0n[12], readReq_2n);
  AND2 I45 (read_2a0d[13], store_0n[13], readReq_2n);
  AND2 I46 (read_2a0d[14], store_0n[14], readReq_2n);
  AND2 I47 (read_2a0d[15], store_0n[15], readReq_2n);
  AND2 I48 (read_2a0d[16], store_0n[16], readReq_2n);
  AND2 I49 (read_2a0d[17], store_0n[17], readReq_2n);
  AND2 I50 (read_2a0d[18], store_0n[18], readReq_2n);
  AND2 I51 (read_2a0d[19], store_0n[19], readReq_2n);
  AND2 I52 (read_2a0d[20], store_0n[20], readReq_2n);
  AND2 I53 (read_2a0d[21], store_0n[21], readReq_2n);
  AND2 I54 (read_2a0d[22], store_0n[22], readReq_2n);
  AND2 I55 (read_2a0d[23], store_0n[23], readReq_2n);
  AND2 I56 (read_2a0d[24], store_0n[24], readReq_2n);
  AND2 I57 (read_2a0d[25], store_0n[25], readReq_2n);
  AND2 I58 (read_2a0d[26], store_0n[26], readReq_2n);
  AND2 I59 (read_2a0d[27], store_0n[27], readReq_2n);
  AND2 I60 (read_2a0d[28], store_0n[28], readReq_2n);
  AND2 I61 (read_2a0d[29], store_0n[29], readReq_2n);
  AND2 I62 (read_2a0d[30], store_0n[30], readReq_2n);
  AND2 I63 (read_2a0d[31], store_0n[31], readReq_2n);
  AND2 I64 (read_1a1d, store_1n[31], readReq_1n);
  AND2 I65 (read_1a0d, store_0n[31], readReq_1n);
  AND2 I66 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I67 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I68 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I69 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I70 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I71 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I72 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I73 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I74 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I75 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I76 (read_0a1d[10], store_1n[10], readReq_0n);
  AND2 I77 (read_0a1d[11], store_1n[11], readReq_0n);
  AND2 I78 (read_0a1d[12], store_1n[12], readReq_0n);
  AND2 I79 (read_0a1d[13], store_1n[13], readReq_0n);
  AND2 I80 (read_0a1d[14], store_1n[14], readReq_0n);
  AND2 I81 (read_0a1d[15], store_1n[15], readReq_0n);
  AND2 I82 (read_0a1d[16], store_1n[16], readReq_0n);
  AND2 I83 (read_0a1d[17], store_1n[17], readReq_0n);
  AND2 I84 (read_0a1d[18], store_1n[18], readReq_0n);
  AND2 I85 (read_0a1d[19], store_1n[19], readReq_0n);
  AND2 I86 (read_0a1d[20], store_1n[20], readReq_0n);
  AND2 I87 (read_0a1d[21], store_1n[21], readReq_0n);
  AND2 I88 (read_0a1d[22], store_1n[22], readReq_0n);
  AND2 I89 (read_0a1d[23], store_1n[23], readReq_0n);
  AND2 I90 (read_0a1d[24], store_1n[24], readReq_0n);
  AND2 I91 (read_0a1d[25], store_1n[25], readReq_0n);
  AND2 I92 (read_0a1d[26], store_1n[26], readReq_0n);
  AND2 I93 (read_0a1d[27], store_1n[27], readReq_0n);
  AND2 I94 (read_0a1d[28], store_1n[28], readReq_0n);
  AND2 I95 (read_0a1d[29], store_1n[29], readReq_0n);
  AND2 I96 (read_0a1d[30], store_1n[30], readReq_0n);
  AND2 I97 (read_0a1d[31], store_1n[31], readReq_0n);
  AND2 I98 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I99 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I100 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I101 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I102 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I103 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I104 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I105 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I106 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I107 (read_0a0d[9], store_0n[9], readReq_0n);
  AND2 I108 (read_0a0d[10], store_0n[10], readReq_0n);
  AND2 I109 (read_0a0d[11], store_0n[11], readReq_0n);
  AND2 I110 (read_0a0d[12], store_0n[12], readReq_0n);
  AND2 I111 (read_0a0d[13], store_0n[13], readReq_0n);
  AND2 I112 (read_0a0d[14], store_0n[14], readReq_0n);
  AND2 I113 (read_0a0d[15], store_0n[15], readReq_0n);
  AND2 I114 (read_0a0d[16], store_0n[16], readReq_0n);
  AND2 I115 (read_0a0d[17], store_0n[17], readReq_0n);
  AND2 I116 (read_0a0d[18], store_0n[18], readReq_0n);
  AND2 I117 (read_0a0d[19], store_0n[19], readReq_0n);
  AND2 I118 (read_0a0d[20], store_0n[20], readReq_0n);
  AND2 I119 (read_0a0d[21], store_0n[21], readReq_0n);
  AND2 I120 (read_0a0d[22], store_0n[22], readReq_0n);
  AND2 I121 (read_0a0d[23], store_0n[23], readReq_0n);
  AND2 I122 (read_0a0d[24], store_0n[24], readReq_0n);
  AND2 I123 (read_0a0d[25], store_0n[25], readReq_0n);
  AND2 I124 (read_0a0d[26], store_0n[26], readReq_0n);
  AND2 I125 (read_0a0d[27], store_0n[27], readReq_0n);
  AND2 I126 (read_0a0d[28], store_0n[28], readReq_0n);
  AND2 I127 (read_0a0d[29], store_0n[29], readReq_0n);
  AND2 I128 (read_0a0d[30], store_0n[30], readReq_0n);
  AND2 I129 (read_0a0d[31], store_0n[31], readReq_0n);
  BUFF I130 (readReq_0n, read_0r);
  BUFF I131 (readReq_1n, read_1r);
  BUFF I132 (readReq_2n, read_2r);
  BUFF I133 (store_1n[0], write_0a1d[0]);
  BUFF I134 (store_1n[1], write_0a1d[1]);
  BUFF I135 (store_1n[2], write_0a1d[2]);
  BUFF I136 (store_1n[3], write_0a1d[3]);
  BUFF I137 (store_1n[4], write_0a1d[4]);
  BUFF I138 (store_1n[5], write_0a1d[5]);
  BUFF I139 (store_1n[6], write_0a1d[6]);
  BUFF I140 (store_1n[7], write_0a1d[7]);
  BUFF I141 (store_1n[8], write_0a1d[8]);
  BUFF I142 (store_1n[9], write_0a1d[9]);
  BUFF I143 (store_1n[10], write_0a1d[10]);
  BUFF I144 (store_1n[11], write_0a1d[11]);
  BUFF I145 (store_1n[12], write_0a1d[12]);
  BUFF I146 (store_1n[13], write_0a1d[13]);
  BUFF I147 (store_1n[14], write_0a1d[14]);
  BUFF I148 (store_1n[15], write_0a1d[15]);
  BUFF I149 (store_1n[16], write_0a1d[16]);
  BUFF I150 (store_1n[17], write_0a1d[17]);
  BUFF I151 (store_1n[18], write_0a1d[18]);
  BUFF I152 (store_1n[19], write_0a1d[19]);
  BUFF I153 (store_1n[20], write_0a1d[20]);
  BUFF I154 (store_1n[21], write_0a1d[21]);
  BUFF I155 (store_1n[22], write_0a1d[22]);
  BUFF I156 (store_1n[23], write_0a1d[23]);
  BUFF I157 (store_1n[24], write_0a1d[24]);
  BUFF I158 (store_1n[25], write_0a1d[25]);
  BUFF I159 (store_1n[26], write_0a1d[26]);
  BUFF I160 (store_1n[27], write_0a1d[27]);
  BUFF I161 (store_1n[28], write_0a1d[28]);
  BUFF I162 (store_1n[29], write_0a1d[29]);
  BUFF I163 (store_1n[30], write_0a1d[30]);
  BUFF I164 (store_1n[31], write_0a1d[31]);
  BUFF I165 (store_0n[0], write_0a0d[0]);
  BUFF I166 (store_0n[1], write_0a0d[1]);
  BUFF I167 (store_0n[2], write_0a0d[2]);
  BUFF I168 (store_0n[3], write_0a0d[3]);
  BUFF I169 (store_0n[4], write_0a0d[4]);
  BUFF I170 (store_0n[5], write_0a0d[5]);
  BUFF I171 (store_0n[6], write_0a0d[6]);
  BUFF I172 (store_0n[7], write_0a0d[7]);
  BUFF I173 (store_0n[8], write_0a0d[8]);
  BUFF I174 (store_0n[9], write_0a0d[9]);
  BUFF I175 (store_0n[10], write_0a0d[10]);
  BUFF I176 (store_0n[11], write_0a0d[11]);
  BUFF I177 (store_0n[12], write_0a0d[12]);
  BUFF I178 (store_0n[13], write_0a0d[13]);
  BUFF I179 (store_0n[14], write_0a0d[14]);
  BUFF I180 (store_0n[15], write_0a0d[15]);
  BUFF I181 (store_0n[16], write_0a0d[16]);
  BUFF I182 (store_0n[17], write_0a0d[17]);
  BUFF I183 (store_0n[18], write_0a0d[18]);
  BUFF I184 (store_0n[19], write_0a0d[19]);
  BUFF I185 (store_0n[20], write_0a0d[20]);
  BUFF I186 (store_0n[21], write_0a0d[21]);
  BUFF I187 (store_0n[22], write_0a0d[22]);
  BUFF I188 (store_0n[23], write_0a0d[23]);
  BUFF I189 (store_0n[24], write_0a0d[24]);
  BUFF I190 (store_0n[25], write_0a0d[25]);
  BUFF I191 (store_0n[26], write_0a0d[26]);
  BUFF I192 (store_0n[27], write_0a0d[27]);
  BUFF I193 (store_0n[28], write_0a0d[28]);
  BUFF I194 (store_0n[29], write_0a0d[29]);
  BUFF I195 (store_0n[30], write_0a0d[30]);
  BUFF I196 (store_0n[31], write_0a0d[31]);
  C2 I197 (trigger_0a, writeAck_0n, cd_0n);
  AND2 I198 (writeAck_0n, sigAck_0n, rReqOr_0n);
  NOR3 I199 (rReqOr_0n, readReq_0n, readReq_1n, readReq_2n);
  BALSA_TELEM I200 (trigger_0r, sigAck_0n, signal_0r, signal_0a);
  C3 I201 (internal_0n[0], partCD_0n[0], partCD_0n[1], partCD_0n[2]);
  C3 I202 (internal_0n[1], partCD_0n[3], partCD_0n[4], partCD_0n[5]);
  C3 I203 (internal_0n[2], partCD_0n[6], partCD_0n[7], partCD_0n[8]);
  C3 I204 (internal_0n[3], partCD_0n[9], partCD_0n[10], partCD_0n[11]);
  C3 I205 (internal_0n[4], partCD_0n[12], partCD_0n[13], partCD_0n[14]);
  C3 I206 (internal_0n[5], partCD_0n[15], partCD_0n[16], partCD_0n[17]);
  C3 I207 (internal_0n[6], partCD_0n[18], partCD_0n[19], partCD_0n[20]);
  C3 I208 (internal_0n[7], partCD_0n[21], partCD_0n[22], partCD_0n[23]);
  C3 I209 (internal_0n[8], partCD_0n[24], partCD_0n[25], partCD_0n[26]);
  C3 I210 (internal_0n[9], partCD_0n[27], partCD_0n[28], partCD_0n[29]);
  C2 I211 (internal_0n[10], partCD_0n[30], partCD_0n[31]);
  C3 I212 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I213 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I214 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I215 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I216 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I217 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I218 (cd_0n, internal_0n[15], internal_0n[16]);
  OR2 I219 (partCD_0n[0], store_0n[0], store_1n[0]);
  OR2 I220 (partCD_0n[1], store_0n[1], store_1n[1]);
  OR2 I221 (partCD_0n[2], store_0n[2], store_1n[2]);
  OR2 I222 (partCD_0n[3], store_0n[3], store_1n[3]);
  OR2 I223 (partCD_0n[4], store_0n[4], store_1n[4]);
  OR2 I224 (partCD_0n[5], store_0n[5], store_1n[5]);
  OR2 I225 (partCD_0n[6], store_0n[6], store_1n[6]);
  OR2 I226 (partCD_0n[7], store_0n[7], store_1n[7]);
  OR2 I227 (partCD_0n[8], store_0n[8], store_1n[8]);
  OR2 I228 (partCD_0n[9], store_0n[9], store_1n[9]);
  OR2 I229 (partCD_0n[10], store_0n[10], store_1n[10]);
  OR2 I230 (partCD_0n[11], store_0n[11], store_1n[11]);
  OR2 I231 (partCD_0n[12], store_0n[12], store_1n[12]);
  OR2 I232 (partCD_0n[13], store_0n[13], store_1n[13]);
  OR2 I233 (partCD_0n[14], store_0n[14], store_1n[14]);
  OR2 I234 (partCD_0n[15], store_0n[15], store_1n[15]);
  OR2 I235 (partCD_0n[16], store_0n[16], store_1n[16]);
  OR2 I236 (partCD_0n[17], store_0n[17], store_1n[17]);
  OR2 I237 (partCD_0n[18], store_0n[18], store_1n[18]);
  OR2 I238 (partCD_0n[19], store_0n[19], store_1n[19]);
  OR2 I239 (partCD_0n[20], store_0n[20], store_1n[20]);
  OR2 I240 (partCD_0n[21], store_0n[21], store_1n[21]);
  OR2 I241 (partCD_0n[22], store_0n[22], store_1n[22]);
  OR2 I242 (partCD_0n[23], store_0n[23], store_1n[23]);
  OR2 I243 (partCD_0n[24], store_0n[24], store_1n[24]);
  OR2 I244 (partCD_0n[25], store_0n[25], store_1n[25]);
  OR2 I245 (partCD_0n[26], store_0n[26], store_1n[26]);
  OR2 I246 (partCD_0n[27], store_0n[27], store_1n[27]);
  OR2 I247 (partCD_0n[28], store_0n[28], store_1n[28]);
  OR2 I248 (partCD_0n[29], store_0n[29], store_1n[29]);
  OR2 I249 (partCD_0n[30], store_0n[30], store_1n[30]);
  OR2 I250 (partCD_0n[31], store_0n[31], store_1n[31]);
  BUFF I251 (write_0r, trigger_0r);
endmodule

module BrzActiveEagerFalseVariable_33_1_s0_ (
  trigger_0r, trigger_0a,
  write_0r, write_0a0d, write_0a1d,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d
);
  input trigger_0r;
  output trigger_0a;
  output write_0r;
  input [32:0] write_0a0d;
  input [32:0] write_0a1d;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output [32:0] read_0a0d;
  output [32:0] read_0a1d;
  wire [16:0] internal_0n;
  wire cd_0n;
  wire [32:0] partCD_0n;
  wire [32:0] store_0n;
  wire [32:0] store_1n;
  wire readReq_0n;
  wire writeAck_0n;
  wire sigAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I1 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I2 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I3 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I4 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I5 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I6 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I7 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I8 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I9 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I10 (read_0a1d[10], store_1n[10], readReq_0n);
  AND2 I11 (read_0a1d[11], store_1n[11], readReq_0n);
  AND2 I12 (read_0a1d[12], store_1n[12], readReq_0n);
  AND2 I13 (read_0a1d[13], store_1n[13], readReq_0n);
  AND2 I14 (read_0a1d[14], store_1n[14], readReq_0n);
  AND2 I15 (read_0a1d[15], store_1n[15], readReq_0n);
  AND2 I16 (read_0a1d[16], store_1n[16], readReq_0n);
  AND2 I17 (read_0a1d[17], store_1n[17], readReq_0n);
  AND2 I18 (read_0a1d[18], store_1n[18], readReq_0n);
  AND2 I19 (read_0a1d[19], store_1n[19], readReq_0n);
  AND2 I20 (read_0a1d[20], store_1n[20], readReq_0n);
  AND2 I21 (read_0a1d[21], store_1n[21], readReq_0n);
  AND2 I22 (read_0a1d[22], store_1n[22], readReq_0n);
  AND2 I23 (read_0a1d[23], store_1n[23], readReq_0n);
  AND2 I24 (read_0a1d[24], store_1n[24], readReq_0n);
  AND2 I25 (read_0a1d[25], store_1n[25], readReq_0n);
  AND2 I26 (read_0a1d[26], store_1n[26], readReq_0n);
  AND2 I27 (read_0a1d[27], store_1n[27], readReq_0n);
  AND2 I28 (read_0a1d[28], store_1n[28], readReq_0n);
  AND2 I29 (read_0a1d[29], store_1n[29], readReq_0n);
  AND2 I30 (read_0a1d[30], store_1n[30], readReq_0n);
  AND2 I31 (read_0a1d[31], store_1n[31], readReq_0n);
  AND2 I32 (read_0a1d[32], store_1n[32], readReq_0n);
  AND2 I33 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I34 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I35 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I36 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I37 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I38 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I39 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I40 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I41 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I42 (read_0a0d[9], store_0n[9], readReq_0n);
  AND2 I43 (read_0a0d[10], store_0n[10], readReq_0n);
  AND2 I44 (read_0a0d[11], store_0n[11], readReq_0n);
  AND2 I45 (read_0a0d[12], store_0n[12], readReq_0n);
  AND2 I46 (read_0a0d[13], store_0n[13], readReq_0n);
  AND2 I47 (read_0a0d[14], store_0n[14], readReq_0n);
  AND2 I48 (read_0a0d[15], store_0n[15], readReq_0n);
  AND2 I49 (read_0a0d[16], store_0n[16], readReq_0n);
  AND2 I50 (read_0a0d[17], store_0n[17], readReq_0n);
  AND2 I51 (read_0a0d[18], store_0n[18], readReq_0n);
  AND2 I52 (read_0a0d[19], store_0n[19], readReq_0n);
  AND2 I53 (read_0a0d[20], store_0n[20], readReq_0n);
  AND2 I54 (read_0a0d[21], store_0n[21], readReq_0n);
  AND2 I55 (read_0a0d[22], store_0n[22], readReq_0n);
  AND2 I56 (read_0a0d[23], store_0n[23], readReq_0n);
  AND2 I57 (read_0a0d[24], store_0n[24], readReq_0n);
  AND2 I58 (read_0a0d[25], store_0n[25], readReq_0n);
  AND2 I59 (read_0a0d[26], store_0n[26], readReq_0n);
  AND2 I60 (read_0a0d[27], store_0n[27], readReq_0n);
  AND2 I61 (read_0a0d[28], store_0n[28], readReq_0n);
  AND2 I62 (read_0a0d[29], store_0n[29], readReq_0n);
  AND2 I63 (read_0a0d[30], store_0n[30], readReq_0n);
  AND2 I64 (read_0a0d[31], store_0n[31], readReq_0n);
  AND2 I65 (read_0a0d[32], store_0n[32], readReq_0n);
  BUFF I66 (readReq_0n, read_0r);
  BUFF I67 (store_1n[0], write_0a1d[0]);
  BUFF I68 (store_1n[1], write_0a1d[1]);
  BUFF I69 (store_1n[2], write_0a1d[2]);
  BUFF I70 (store_1n[3], write_0a1d[3]);
  BUFF I71 (store_1n[4], write_0a1d[4]);
  BUFF I72 (store_1n[5], write_0a1d[5]);
  BUFF I73 (store_1n[6], write_0a1d[6]);
  BUFF I74 (store_1n[7], write_0a1d[7]);
  BUFF I75 (store_1n[8], write_0a1d[8]);
  BUFF I76 (store_1n[9], write_0a1d[9]);
  BUFF I77 (store_1n[10], write_0a1d[10]);
  BUFF I78 (store_1n[11], write_0a1d[11]);
  BUFF I79 (store_1n[12], write_0a1d[12]);
  BUFF I80 (store_1n[13], write_0a1d[13]);
  BUFF I81 (store_1n[14], write_0a1d[14]);
  BUFF I82 (store_1n[15], write_0a1d[15]);
  BUFF I83 (store_1n[16], write_0a1d[16]);
  BUFF I84 (store_1n[17], write_0a1d[17]);
  BUFF I85 (store_1n[18], write_0a1d[18]);
  BUFF I86 (store_1n[19], write_0a1d[19]);
  BUFF I87 (store_1n[20], write_0a1d[20]);
  BUFF I88 (store_1n[21], write_0a1d[21]);
  BUFF I89 (store_1n[22], write_0a1d[22]);
  BUFF I90 (store_1n[23], write_0a1d[23]);
  BUFF I91 (store_1n[24], write_0a1d[24]);
  BUFF I92 (store_1n[25], write_0a1d[25]);
  BUFF I93 (store_1n[26], write_0a1d[26]);
  BUFF I94 (store_1n[27], write_0a1d[27]);
  BUFF I95 (store_1n[28], write_0a1d[28]);
  BUFF I96 (store_1n[29], write_0a1d[29]);
  BUFF I97 (store_1n[30], write_0a1d[30]);
  BUFF I98 (store_1n[31], write_0a1d[31]);
  BUFF I99 (store_1n[32], write_0a1d[32]);
  BUFF I100 (store_0n[0], write_0a0d[0]);
  BUFF I101 (store_0n[1], write_0a0d[1]);
  BUFF I102 (store_0n[2], write_0a0d[2]);
  BUFF I103 (store_0n[3], write_0a0d[3]);
  BUFF I104 (store_0n[4], write_0a0d[4]);
  BUFF I105 (store_0n[5], write_0a0d[5]);
  BUFF I106 (store_0n[6], write_0a0d[6]);
  BUFF I107 (store_0n[7], write_0a0d[7]);
  BUFF I108 (store_0n[8], write_0a0d[8]);
  BUFF I109 (store_0n[9], write_0a0d[9]);
  BUFF I110 (store_0n[10], write_0a0d[10]);
  BUFF I111 (store_0n[11], write_0a0d[11]);
  BUFF I112 (store_0n[12], write_0a0d[12]);
  BUFF I113 (store_0n[13], write_0a0d[13]);
  BUFF I114 (store_0n[14], write_0a0d[14]);
  BUFF I115 (store_0n[15], write_0a0d[15]);
  BUFF I116 (store_0n[16], write_0a0d[16]);
  BUFF I117 (store_0n[17], write_0a0d[17]);
  BUFF I118 (store_0n[18], write_0a0d[18]);
  BUFF I119 (store_0n[19], write_0a0d[19]);
  BUFF I120 (store_0n[20], write_0a0d[20]);
  BUFF I121 (store_0n[21], write_0a0d[21]);
  BUFF I122 (store_0n[22], write_0a0d[22]);
  BUFF I123 (store_0n[23], write_0a0d[23]);
  BUFF I124 (store_0n[24], write_0a0d[24]);
  BUFF I125 (store_0n[25], write_0a0d[25]);
  BUFF I126 (store_0n[26], write_0a0d[26]);
  BUFF I127 (store_0n[27], write_0a0d[27]);
  BUFF I128 (store_0n[28], write_0a0d[28]);
  BUFF I129 (store_0n[29], write_0a0d[29]);
  BUFF I130 (store_0n[30], write_0a0d[30]);
  BUFF I131 (store_0n[31], write_0a0d[31]);
  BUFF I132 (store_0n[32], write_0a0d[32]);
  C2 I133 (trigger_0a, writeAck_0n, cd_0n);
  AND2 I134 (writeAck_0n, sigAck_0n, rReqOr_0n);
  INV I135 (rReqOr_0n, readReq_0n);
  BALSA_TELEM I136 (trigger_0r, sigAck_0n, signal_0r, signal_0a);
  C3 I137 (internal_0n[0], partCD_0n[0], partCD_0n[1], partCD_0n[2]);
  C3 I138 (internal_0n[1], partCD_0n[3], partCD_0n[4], partCD_0n[5]);
  C3 I139 (internal_0n[2], partCD_0n[6], partCD_0n[7], partCD_0n[8]);
  C3 I140 (internal_0n[3], partCD_0n[9], partCD_0n[10], partCD_0n[11]);
  C3 I141 (internal_0n[4], partCD_0n[12], partCD_0n[13], partCD_0n[14]);
  C3 I142 (internal_0n[5], partCD_0n[15], partCD_0n[16], partCD_0n[17]);
  C3 I143 (internal_0n[6], partCD_0n[18], partCD_0n[19], partCD_0n[20]);
  C3 I144 (internal_0n[7], partCD_0n[21], partCD_0n[22], partCD_0n[23]);
  C3 I145 (internal_0n[8], partCD_0n[24], partCD_0n[25], partCD_0n[26]);
  C3 I146 (internal_0n[9], partCD_0n[27], partCD_0n[28], partCD_0n[29]);
  C3 I147 (internal_0n[10], partCD_0n[30], partCD_0n[31], partCD_0n[32]);
  C3 I148 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I149 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I150 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I151 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I152 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I153 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I154 (cd_0n, internal_0n[15], internal_0n[16]);
  OR2 I155 (partCD_0n[0], store_0n[0], store_1n[0]);
  OR2 I156 (partCD_0n[1], store_0n[1], store_1n[1]);
  OR2 I157 (partCD_0n[2], store_0n[2], store_1n[2]);
  OR2 I158 (partCD_0n[3], store_0n[3], store_1n[3]);
  OR2 I159 (partCD_0n[4], store_0n[4], store_1n[4]);
  OR2 I160 (partCD_0n[5], store_0n[5], store_1n[5]);
  OR2 I161 (partCD_0n[6], store_0n[6], store_1n[6]);
  OR2 I162 (partCD_0n[7], store_0n[7], store_1n[7]);
  OR2 I163 (partCD_0n[8], store_0n[8], store_1n[8]);
  OR2 I164 (partCD_0n[9], store_0n[9], store_1n[9]);
  OR2 I165 (partCD_0n[10], store_0n[10], store_1n[10]);
  OR2 I166 (partCD_0n[11], store_0n[11], store_1n[11]);
  OR2 I167 (partCD_0n[12], store_0n[12], store_1n[12]);
  OR2 I168 (partCD_0n[13], store_0n[13], store_1n[13]);
  OR2 I169 (partCD_0n[14], store_0n[14], store_1n[14]);
  OR2 I170 (partCD_0n[15], store_0n[15], store_1n[15]);
  OR2 I171 (partCD_0n[16], store_0n[16], store_1n[16]);
  OR2 I172 (partCD_0n[17], store_0n[17], store_1n[17]);
  OR2 I173 (partCD_0n[18], store_0n[18], store_1n[18]);
  OR2 I174 (partCD_0n[19], store_0n[19], store_1n[19]);
  OR2 I175 (partCD_0n[20], store_0n[20], store_1n[20]);
  OR2 I176 (partCD_0n[21], store_0n[21], store_1n[21]);
  OR2 I177 (partCD_0n[22], store_0n[22], store_1n[22]);
  OR2 I178 (partCD_0n[23], store_0n[23], store_1n[23]);
  OR2 I179 (partCD_0n[24], store_0n[24], store_1n[24]);
  OR2 I180 (partCD_0n[25], store_0n[25], store_1n[25]);
  OR2 I181 (partCD_0n[26], store_0n[26], store_1n[26]);
  OR2 I182 (partCD_0n[27], store_0n[27], store_1n[27]);
  OR2 I183 (partCD_0n[28], store_0n[28], store_1n[28]);
  OR2 I184 (partCD_0n[29], store_0n[29], store_1n[29]);
  OR2 I185 (partCD_0n[30], store_0n[30], store_1n[30]);
  OR2 I186 (partCD_0n[31], store_0n[31], store_1n[31]);
  OR2 I187 (partCD_0n[32], store_0n[32], store_1n[32]);
  BUFF I188 (write_0r, trigger_0r);
endmodule

module BrzActiveEagerFalseVariable_34_2_s22_1_2e__m5m (
  trigger_0r, trigger_0a,
  write_0r, write_0a0d, write_0a1d,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d
);
  input trigger_0r;
  output trigger_0a;
  output write_0r;
  input [33:0] write_0a0d;
  input [33:0] write_0a1d;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output [31:0] read_0a0d;
  output [31:0] read_0a1d;
  input read_1r;
  output read_1a0d;
  output read_1a1d;
  wire [17:0] internal_0n;
  wire cd_0n;
  wire [33:0] partCD_0n;
  wire [33:0] store_0n;
  wire [33:0] store_1n;
  wire readReq_0n;
  wire readReq_1n;
  wire writeAck_0n;
  wire sigAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_1a1d, store_1n[33], readReq_1n);
  AND2 I1 (read_1a0d, store_0n[33], readReq_1n);
  AND2 I2 (read_0a1d[0], store_1n[1], readReq_0n);
  AND2 I3 (read_0a1d[1], store_1n[2], readReq_0n);
  AND2 I4 (read_0a1d[2], store_1n[3], readReq_0n);
  AND2 I5 (read_0a1d[3], store_1n[4], readReq_0n);
  AND2 I6 (read_0a1d[4], store_1n[5], readReq_0n);
  AND2 I7 (read_0a1d[5], store_1n[6], readReq_0n);
  AND2 I8 (read_0a1d[6], store_1n[7], readReq_0n);
  AND2 I9 (read_0a1d[7], store_1n[8], readReq_0n);
  AND2 I10 (read_0a1d[8], store_1n[9], readReq_0n);
  AND2 I11 (read_0a1d[9], store_1n[10], readReq_0n);
  AND2 I12 (read_0a1d[10], store_1n[11], readReq_0n);
  AND2 I13 (read_0a1d[11], store_1n[12], readReq_0n);
  AND2 I14 (read_0a1d[12], store_1n[13], readReq_0n);
  AND2 I15 (read_0a1d[13], store_1n[14], readReq_0n);
  AND2 I16 (read_0a1d[14], store_1n[15], readReq_0n);
  AND2 I17 (read_0a1d[15], store_1n[16], readReq_0n);
  AND2 I18 (read_0a1d[16], store_1n[17], readReq_0n);
  AND2 I19 (read_0a1d[17], store_1n[18], readReq_0n);
  AND2 I20 (read_0a1d[18], store_1n[19], readReq_0n);
  AND2 I21 (read_0a1d[19], store_1n[20], readReq_0n);
  AND2 I22 (read_0a1d[20], store_1n[21], readReq_0n);
  AND2 I23 (read_0a1d[21], store_1n[22], readReq_0n);
  AND2 I24 (read_0a1d[22], store_1n[23], readReq_0n);
  AND2 I25 (read_0a1d[23], store_1n[24], readReq_0n);
  AND2 I26 (read_0a1d[24], store_1n[25], readReq_0n);
  AND2 I27 (read_0a1d[25], store_1n[26], readReq_0n);
  AND2 I28 (read_0a1d[26], store_1n[27], readReq_0n);
  AND2 I29 (read_0a1d[27], store_1n[28], readReq_0n);
  AND2 I30 (read_0a1d[28], store_1n[29], readReq_0n);
  AND2 I31 (read_0a1d[29], store_1n[30], readReq_0n);
  AND2 I32 (read_0a1d[30], store_1n[31], readReq_0n);
  AND2 I33 (read_0a1d[31], store_1n[32], readReq_0n);
  AND2 I34 (read_0a0d[0], store_0n[1], readReq_0n);
  AND2 I35 (read_0a0d[1], store_0n[2], readReq_0n);
  AND2 I36 (read_0a0d[2], store_0n[3], readReq_0n);
  AND2 I37 (read_0a0d[3], store_0n[4], readReq_0n);
  AND2 I38 (read_0a0d[4], store_0n[5], readReq_0n);
  AND2 I39 (read_0a0d[5], store_0n[6], readReq_0n);
  AND2 I40 (read_0a0d[6], store_0n[7], readReq_0n);
  AND2 I41 (read_0a0d[7], store_0n[8], readReq_0n);
  AND2 I42 (read_0a0d[8], store_0n[9], readReq_0n);
  AND2 I43 (read_0a0d[9], store_0n[10], readReq_0n);
  AND2 I44 (read_0a0d[10], store_0n[11], readReq_0n);
  AND2 I45 (read_0a0d[11], store_0n[12], readReq_0n);
  AND2 I46 (read_0a0d[12], store_0n[13], readReq_0n);
  AND2 I47 (read_0a0d[13], store_0n[14], readReq_0n);
  AND2 I48 (read_0a0d[14], store_0n[15], readReq_0n);
  AND2 I49 (read_0a0d[15], store_0n[16], readReq_0n);
  AND2 I50 (read_0a0d[16], store_0n[17], readReq_0n);
  AND2 I51 (read_0a0d[17], store_0n[18], readReq_0n);
  AND2 I52 (read_0a0d[18], store_0n[19], readReq_0n);
  AND2 I53 (read_0a0d[19], store_0n[20], readReq_0n);
  AND2 I54 (read_0a0d[20], store_0n[21], readReq_0n);
  AND2 I55 (read_0a0d[21], store_0n[22], readReq_0n);
  AND2 I56 (read_0a0d[22], store_0n[23], readReq_0n);
  AND2 I57 (read_0a0d[23], store_0n[24], readReq_0n);
  AND2 I58 (read_0a0d[24], store_0n[25], readReq_0n);
  AND2 I59 (read_0a0d[25], store_0n[26], readReq_0n);
  AND2 I60 (read_0a0d[26], store_0n[27], readReq_0n);
  AND2 I61 (read_0a0d[27], store_0n[28], readReq_0n);
  AND2 I62 (read_0a0d[28], store_0n[29], readReq_0n);
  AND2 I63 (read_0a0d[29], store_0n[30], readReq_0n);
  AND2 I64 (read_0a0d[30], store_0n[31], readReq_0n);
  AND2 I65 (read_0a0d[31], store_0n[32], readReq_0n);
  BUFF I66 (readReq_0n, read_0r);
  BUFF I67 (readReq_1n, read_1r);
  BUFF I68 (store_1n[0], write_0a1d[0]);
  BUFF I69 (store_1n[1], write_0a1d[1]);
  BUFF I70 (store_1n[2], write_0a1d[2]);
  BUFF I71 (store_1n[3], write_0a1d[3]);
  BUFF I72 (store_1n[4], write_0a1d[4]);
  BUFF I73 (store_1n[5], write_0a1d[5]);
  BUFF I74 (store_1n[6], write_0a1d[6]);
  BUFF I75 (store_1n[7], write_0a1d[7]);
  BUFF I76 (store_1n[8], write_0a1d[8]);
  BUFF I77 (store_1n[9], write_0a1d[9]);
  BUFF I78 (store_1n[10], write_0a1d[10]);
  BUFF I79 (store_1n[11], write_0a1d[11]);
  BUFF I80 (store_1n[12], write_0a1d[12]);
  BUFF I81 (store_1n[13], write_0a1d[13]);
  BUFF I82 (store_1n[14], write_0a1d[14]);
  BUFF I83 (store_1n[15], write_0a1d[15]);
  BUFF I84 (store_1n[16], write_0a1d[16]);
  BUFF I85 (store_1n[17], write_0a1d[17]);
  BUFF I86 (store_1n[18], write_0a1d[18]);
  BUFF I87 (store_1n[19], write_0a1d[19]);
  BUFF I88 (store_1n[20], write_0a1d[20]);
  BUFF I89 (store_1n[21], write_0a1d[21]);
  BUFF I90 (store_1n[22], write_0a1d[22]);
  BUFF I91 (store_1n[23], write_0a1d[23]);
  BUFF I92 (store_1n[24], write_0a1d[24]);
  BUFF I93 (store_1n[25], write_0a1d[25]);
  BUFF I94 (store_1n[26], write_0a1d[26]);
  BUFF I95 (store_1n[27], write_0a1d[27]);
  BUFF I96 (store_1n[28], write_0a1d[28]);
  BUFF I97 (store_1n[29], write_0a1d[29]);
  BUFF I98 (store_1n[30], write_0a1d[30]);
  BUFF I99 (store_1n[31], write_0a1d[31]);
  BUFF I100 (store_1n[32], write_0a1d[32]);
  BUFF I101 (store_1n[33], write_0a1d[33]);
  BUFF I102 (store_0n[0], write_0a0d[0]);
  BUFF I103 (store_0n[1], write_0a0d[1]);
  BUFF I104 (store_0n[2], write_0a0d[2]);
  BUFF I105 (store_0n[3], write_0a0d[3]);
  BUFF I106 (store_0n[4], write_0a0d[4]);
  BUFF I107 (store_0n[5], write_0a0d[5]);
  BUFF I108 (store_0n[6], write_0a0d[6]);
  BUFF I109 (store_0n[7], write_0a0d[7]);
  BUFF I110 (store_0n[8], write_0a0d[8]);
  BUFF I111 (store_0n[9], write_0a0d[9]);
  BUFF I112 (store_0n[10], write_0a0d[10]);
  BUFF I113 (store_0n[11], write_0a0d[11]);
  BUFF I114 (store_0n[12], write_0a0d[12]);
  BUFF I115 (store_0n[13], write_0a0d[13]);
  BUFF I116 (store_0n[14], write_0a0d[14]);
  BUFF I117 (store_0n[15], write_0a0d[15]);
  BUFF I118 (store_0n[16], write_0a0d[16]);
  BUFF I119 (store_0n[17], write_0a0d[17]);
  BUFF I120 (store_0n[18], write_0a0d[18]);
  BUFF I121 (store_0n[19], write_0a0d[19]);
  BUFF I122 (store_0n[20], write_0a0d[20]);
  BUFF I123 (store_0n[21], write_0a0d[21]);
  BUFF I124 (store_0n[22], write_0a0d[22]);
  BUFF I125 (store_0n[23], write_0a0d[23]);
  BUFF I126 (store_0n[24], write_0a0d[24]);
  BUFF I127 (store_0n[25], write_0a0d[25]);
  BUFF I128 (store_0n[26], write_0a0d[26]);
  BUFF I129 (store_0n[27], write_0a0d[27]);
  BUFF I130 (store_0n[28], write_0a0d[28]);
  BUFF I131 (store_0n[29], write_0a0d[29]);
  BUFF I132 (store_0n[30], write_0a0d[30]);
  BUFF I133 (store_0n[31], write_0a0d[31]);
  BUFF I134 (store_0n[32], write_0a0d[32]);
  BUFF I135 (store_0n[33], write_0a0d[33]);
  C2 I136 (trigger_0a, writeAck_0n, cd_0n);
  AND2 I137 (writeAck_0n, sigAck_0n, rReqOr_0n);
  NOR2 I138 (rReqOr_0n, readReq_0n, readReq_1n);
  BALSA_TELEM I139 (trigger_0r, sigAck_0n, signal_0r, signal_0a);
  C3 I140 (internal_0n[0], partCD_0n[0], partCD_0n[1], partCD_0n[2]);
  C3 I141 (internal_0n[1], partCD_0n[3], partCD_0n[4], partCD_0n[5]);
  C3 I142 (internal_0n[2], partCD_0n[6], partCD_0n[7], partCD_0n[8]);
  C3 I143 (internal_0n[3], partCD_0n[9], partCD_0n[10], partCD_0n[11]);
  C3 I144 (internal_0n[4], partCD_0n[12], partCD_0n[13], partCD_0n[14]);
  C3 I145 (internal_0n[5], partCD_0n[15], partCD_0n[16], partCD_0n[17]);
  C3 I146 (internal_0n[6], partCD_0n[18], partCD_0n[19], partCD_0n[20]);
  C3 I147 (internal_0n[7], partCD_0n[21], partCD_0n[22], partCD_0n[23]);
  C3 I148 (internal_0n[8], partCD_0n[24], partCD_0n[25], partCD_0n[26]);
  C3 I149 (internal_0n[9], partCD_0n[27], partCD_0n[28], partCD_0n[29]);
  C2 I150 (internal_0n[10], partCD_0n[30], partCD_0n[31]);
  C2 I151 (internal_0n[11], partCD_0n[32], partCD_0n[33]);
  C3 I152 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I153 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I154 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I155 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I156 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I157 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I158 (cd_0n, internal_0n[16], internal_0n[17]);
  OR2 I159 (partCD_0n[0], store_0n[0], store_1n[0]);
  OR2 I160 (partCD_0n[1], store_0n[1], store_1n[1]);
  OR2 I161 (partCD_0n[2], store_0n[2], store_1n[2]);
  OR2 I162 (partCD_0n[3], store_0n[3], store_1n[3]);
  OR2 I163 (partCD_0n[4], store_0n[4], store_1n[4]);
  OR2 I164 (partCD_0n[5], store_0n[5], store_1n[5]);
  OR2 I165 (partCD_0n[6], store_0n[6], store_1n[6]);
  OR2 I166 (partCD_0n[7], store_0n[7], store_1n[7]);
  OR2 I167 (partCD_0n[8], store_0n[8], store_1n[8]);
  OR2 I168 (partCD_0n[9], store_0n[9], store_1n[9]);
  OR2 I169 (partCD_0n[10], store_0n[10], store_1n[10]);
  OR2 I170 (partCD_0n[11], store_0n[11], store_1n[11]);
  OR2 I171 (partCD_0n[12], store_0n[12], store_1n[12]);
  OR2 I172 (partCD_0n[13], store_0n[13], store_1n[13]);
  OR2 I173 (partCD_0n[14], store_0n[14], store_1n[14]);
  OR2 I174 (partCD_0n[15], store_0n[15], store_1n[15]);
  OR2 I175 (partCD_0n[16], store_0n[16], store_1n[16]);
  OR2 I176 (partCD_0n[17], store_0n[17], store_1n[17]);
  OR2 I177 (partCD_0n[18], store_0n[18], store_1n[18]);
  OR2 I178 (partCD_0n[19], store_0n[19], store_1n[19]);
  OR2 I179 (partCD_0n[20], store_0n[20], store_1n[20]);
  OR2 I180 (partCD_0n[21], store_0n[21], store_1n[21]);
  OR2 I181 (partCD_0n[22], store_0n[22], store_1n[22]);
  OR2 I182 (partCD_0n[23], store_0n[23], store_1n[23]);
  OR2 I183 (partCD_0n[24], store_0n[24], store_1n[24]);
  OR2 I184 (partCD_0n[25], store_0n[25], store_1n[25]);
  OR2 I185 (partCD_0n[26], store_0n[26], store_1n[26]);
  OR2 I186 (partCD_0n[27], store_0n[27], store_1n[27]);
  OR2 I187 (partCD_0n[28], store_0n[28], store_1n[28]);
  OR2 I188 (partCD_0n[29], store_0n[29], store_1n[29]);
  OR2 I189 (partCD_0n[30], store_0n[30], store_1n[30]);
  OR2 I190 (partCD_0n[31], store_0n[31], store_1n[31]);
  OR2 I191 (partCD_0n[32], store_0n[32], store_1n[32]);
  OR2 I192 (partCD_0n[33], store_0n[33], store_1n[33]);
  BUFF I193 (write_0r, trigger_0r);
endmodule

module BrzActiveEagerFalseVariable_35_1_s0_ (
  trigger_0r, trigger_0a,
  write_0r, write_0a0d, write_0a1d,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d
);
  input trigger_0r;
  output trigger_0a;
  output write_0r;
  input [34:0] write_0a0d;
  input [34:0] write_0a1d;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output [34:0] read_0a0d;
  output [34:0] read_0a1d;
  wire [17:0] internal_0n;
  wire cd_0n;
  wire [34:0] partCD_0n;
  wire [34:0] store_0n;
  wire [34:0] store_1n;
  wire readReq_0n;
  wire writeAck_0n;
  wire sigAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I1 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I2 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I3 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I4 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I5 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I6 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I7 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I8 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I9 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I10 (read_0a1d[10], store_1n[10], readReq_0n);
  AND2 I11 (read_0a1d[11], store_1n[11], readReq_0n);
  AND2 I12 (read_0a1d[12], store_1n[12], readReq_0n);
  AND2 I13 (read_0a1d[13], store_1n[13], readReq_0n);
  AND2 I14 (read_0a1d[14], store_1n[14], readReq_0n);
  AND2 I15 (read_0a1d[15], store_1n[15], readReq_0n);
  AND2 I16 (read_0a1d[16], store_1n[16], readReq_0n);
  AND2 I17 (read_0a1d[17], store_1n[17], readReq_0n);
  AND2 I18 (read_0a1d[18], store_1n[18], readReq_0n);
  AND2 I19 (read_0a1d[19], store_1n[19], readReq_0n);
  AND2 I20 (read_0a1d[20], store_1n[20], readReq_0n);
  AND2 I21 (read_0a1d[21], store_1n[21], readReq_0n);
  AND2 I22 (read_0a1d[22], store_1n[22], readReq_0n);
  AND2 I23 (read_0a1d[23], store_1n[23], readReq_0n);
  AND2 I24 (read_0a1d[24], store_1n[24], readReq_0n);
  AND2 I25 (read_0a1d[25], store_1n[25], readReq_0n);
  AND2 I26 (read_0a1d[26], store_1n[26], readReq_0n);
  AND2 I27 (read_0a1d[27], store_1n[27], readReq_0n);
  AND2 I28 (read_0a1d[28], store_1n[28], readReq_0n);
  AND2 I29 (read_0a1d[29], store_1n[29], readReq_0n);
  AND2 I30 (read_0a1d[30], store_1n[30], readReq_0n);
  AND2 I31 (read_0a1d[31], store_1n[31], readReq_0n);
  AND2 I32 (read_0a1d[32], store_1n[32], readReq_0n);
  AND2 I33 (read_0a1d[33], store_1n[33], readReq_0n);
  AND2 I34 (read_0a1d[34], store_1n[34], readReq_0n);
  AND2 I35 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I36 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I37 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I38 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I39 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I40 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I41 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I42 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I43 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I44 (read_0a0d[9], store_0n[9], readReq_0n);
  AND2 I45 (read_0a0d[10], store_0n[10], readReq_0n);
  AND2 I46 (read_0a0d[11], store_0n[11], readReq_0n);
  AND2 I47 (read_0a0d[12], store_0n[12], readReq_0n);
  AND2 I48 (read_0a0d[13], store_0n[13], readReq_0n);
  AND2 I49 (read_0a0d[14], store_0n[14], readReq_0n);
  AND2 I50 (read_0a0d[15], store_0n[15], readReq_0n);
  AND2 I51 (read_0a0d[16], store_0n[16], readReq_0n);
  AND2 I52 (read_0a0d[17], store_0n[17], readReq_0n);
  AND2 I53 (read_0a0d[18], store_0n[18], readReq_0n);
  AND2 I54 (read_0a0d[19], store_0n[19], readReq_0n);
  AND2 I55 (read_0a0d[20], store_0n[20], readReq_0n);
  AND2 I56 (read_0a0d[21], store_0n[21], readReq_0n);
  AND2 I57 (read_0a0d[22], store_0n[22], readReq_0n);
  AND2 I58 (read_0a0d[23], store_0n[23], readReq_0n);
  AND2 I59 (read_0a0d[24], store_0n[24], readReq_0n);
  AND2 I60 (read_0a0d[25], store_0n[25], readReq_0n);
  AND2 I61 (read_0a0d[26], store_0n[26], readReq_0n);
  AND2 I62 (read_0a0d[27], store_0n[27], readReq_0n);
  AND2 I63 (read_0a0d[28], store_0n[28], readReq_0n);
  AND2 I64 (read_0a0d[29], store_0n[29], readReq_0n);
  AND2 I65 (read_0a0d[30], store_0n[30], readReq_0n);
  AND2 I66 (read_0a0d[31], store_0n[31], readReq_0n);
  AND2 I67 (read_0a0d[32], store_0n[32], readReq_0n);
  AND2 I68 (read_0a0d[33], store_0n[33], readReq_0n);
  AND2 I69 (read_0a0d[34], store_0n[34], readReq_0n);
  BUFF I70 (readReq_0n, read_0r);
  BUFF I71 (store_1n[0], write_0a1d[0]);
  BUFF I72 (store_1n[1], write_0a1d[1]);
  BUFF I73 (store_1n[2], write_0a1d[2]);
  BUFF I74 (store_1n[3], write_0a1d[3]);
  BUFF I75 (store_1n[4], write_0a1d[4]);
  BUFF I76 (store_1n[5], write_0a1d[5]);
  BUFF I77 (store_1n[6], write_0a1d[6]);
  BUFF I78 (store_1n[7], write_0a1d[7]);
  BUFF I79 (store_1n[8], write_0a1d[8]);
  BUFF I80 (store_1n[9], write_0a1d[9]);
  BUFF I81 (store_1n[10], write_0a1d[10]);
  BUFF I82 (store_1n[11], write_0a1d[11]);
  BUFF I83 (store_1n[12], write_0a1d[12]);
  BUFF I84 (store_1n[13], write_0a1d[13]);
  BUFF I85 (store_1n[14], write_0a1d[14]);
  BUFF I86 (store_1n[15], write_0a1d[15]);
  BUFF I87 (store_1n[16], write_0a1d[16]);
  BUFF I88 (store_1n[17], write_0a1d[17]);
  BUFF I89 (store_1n[18], write_0a1d[18]);
  BUFF I90 (store_1n[19], write_0a1d[19]);
  BUFF I91 (store_1n[20], write_0a1d[20]);
  BUFF I92 (store_1n[21], write_0a1d[21]);
  BUFF I93 (store_1n[22], write_0a1d[22]);
  BUFF I94 (store_1n[23], write_0a1d[23]);
  BUFF I95 (store_1n[24], write_0a1d[24]);
  BUFF I96 (store_1n[25], write_0a1d[25]);
  BUFF I97 (store_1n[26], write_0a1d[26]);
  BUFF I98 (store_1n[27], write_0a1d[27]);
  BUFF I99 (store_1n[28], write_0a1d[28]);
  BUFF I100 (store_1n[29], write_0a1d[29]);
  BUFF I101 (store_1n[30], write_0a1d[30]);
  BUFF I102 (store_1n[31], write_0a1d[31]);
  BUFF I103 (store_1n[32], write_0a1d[32]);
  BUFF I104 (store_1n[33], write_0a1d[33]);
  BUFF I105 (store_1n[34], write_0a1d[34]);
  BUFF I106 (store_0n[0], write_0a0d[0]);
  BUFF I107 (store_0n[1], write_0a0d[1]);
  BUFF I108 (store_0n[2], write_0a0d[2]);
  BUFF I109 (store_0n[3], write_0a0d[3]);
  BUFF I110 (store_0n[4], write_0a0d[4]);
  BUFF I111 (store_0n[5], write_0a0d[5]);
  BUFF I112 (store_0n[6], write_0a0d[6]);
  BUFF I113 (store_0n[7], write_0a0d[7]);
  BUFF I114 (store_0n[8], write_0a0d[8]);
  BUFF I115 (store_0n[9], write_0a0d[9]);
  BUFF I116 (store_0n[10], write_0a0d[10]);
  BUFF I117 (store_0n[11], write_0a0d[11]);
  BUFF I118 (store_0n[12], write_0a0d[12]);
  BUFF I119 (store_0n[13], write_0a0d[13]);
  BUFF I120 (store_0n[14], write_0a0d[14]);
  BUFF I121 (store_0n[15], write_0a0d[15]);
  BUFF I122 (store_0n[16], write_0a0d[16]);
  BUFF I123 (store_0n[17], write_0a0d[17]);
  BUFF I124 (store_0n[18], write_0a0d[18]);
  BUFF I125 (store_0n[19], write_0a0d[19]);
  BUFF I126 (store_0n[20], write_0a0d[20]);
  BUFF I127 (store_0n[21], write_0a0d[21]);
  BUFF I128 (store_0n[22], write_0a0d[22]);
  BUFF I129 (store_0n[23], write_0a0d[23]);
  BUFF I130 (store_0n[24], write_0a0d[24]);
  BUFF I131 (store_0n[25], write_0a0d[25]);
  BUFF I132 (store_0n[26], write_0a0d[26]);
  BUFF I133 (store_0n[27], write_0a0d[27]);
  BUFF I134 (store_0n[28], write_0a0d[28]);
  BUFF I135 (store_0n[29], write_0a0d[29]);
  BUFF I136 (store_0n[30], write_0a0d[30]);
  BUFF I137 (store_0n[31], write_0a0d[31]);
  BUFF I138 (store_0n[32], write_0a0d[32]);
  BUFF I139 (store_0n[33], write_0a0d[33]);
  BUFF I140 (store_0n[34], write_0a0d[34]);
  C2 I141 (trigger_0a, writeAck_0n, cd_0n);
  AND2 I142 (writeAck_0n, sigAck_0n, rReqOr_0n);
  INV I143 (rReqOr_0n, readReq_0n);
  BALSA_TELEM I144 (trigger_0r, sigAck_0n, signal_0r, signal_0a);
  C3 I145 (internal_0n[0], partCD_0n[0], partCD_0n[1], partCD_0n[2]);
  C3 I146 (internal_0n[1], partCD_0n[3], partCD_0n[4], partCD_0n[5]);
  C3 I147 (internal_0n[2], partCD_0n[6], partCD_0n[7], partCD_0n[8]);
  C3 I148 (internal_0n[3], partCD_0n[9], partCD_0n[10], partCD_0n[11]);
  C3 I149 (internal_0n[4], partCD_0n[12], partCD_0n[13], partCD_0n[14]);
  C3 I150 (internal_0n[5], partCD_0n[15], partCD_0n[16], partCD_0n[17]);
  C3 I151 (internal_0n[6], partCD_0n[18], partCD_0n[19], partCD_0n[20]);
  C3 I152 (internal_0n[7], partCD_0n[21], partCD_0n[22], partCD_0n[23]);
  C3 I153 (internal_0n[8], partCD_0n[24], partCD_0n[25], partCD_0n[26]);
  C3 I154 (internal_0n[9], partCD_0n[27], partCD_0n[28], partCD_0n[29]);
  C3 I155 (internal_0n[10], partCD_0n[30], partCD_0n[31], partCD_0n[32]);
  C2 I156 (internal_0n[11], partCD_0n[33], partCD_0n[34]);
  C3 I157 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I158 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I159 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I160 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I161 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I162 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I163 (cd_0n, internal_0n[16], internal_0n[17]);
  OR2 I164 (partCD_0n[0], store_0n[0], store_1n[0]);
  OR2 I165 (partCD_0n[1], store_0n[1], store_1n[1]);
  OR2 I166 (partCD_0n[2], store_0n[2], store_1n[2]);
  OR2 I167 (partCD_0n[3], store_0n[3], store_1n[3]);
  OR2 I168 (partCD_0n[4], store_0n[4], store_1n[4]);
  OR2 I169 (partCD_0n[5], store_0n[5], store_1n[5]);
  OR2 I170 (partCD_0n[6], store_0n[6], store_1n[6]);
  OR2 I171 (partCD_0n[7], store_0n[7], store_1n[7]);
  OR2 I172 (partCD_0n[8], store_0n[8], store_1n[8]);
  OR2 I173 (partCD_0n[9], store_0n[9], store_1n[9]);
  OR2 I174 (partCD_0n[10], store_0n[10], store_1n[10]);
  OR2 I175 (partCD_0n[11], store_0n[11], store_1n[11]);
  OR2 I176 (partCD_0n[12], store_0n[12], store_1n[12]);
  OR2 I177 (partCD_0n[13], store_0n[13], store_1n[13]);
  OR2 I178 (partCD_0n[14], store_0n[14], store_1n[14]);
  OR2 I179 (partCD_0n[15], store_0n[15], store_1n[15]);
  OR2 I180 (partCD_0n[16], store_0n[16], store_1n[16]);
  OR2 I181 (partCD_0n[17], store_0n[17], store_1n[17]);
  OR2 I182 (partCD_0n[18], store_0n[18], store_1n[18]);
  OR2 I183 (partCD_0n[19], store_0n[19], store_1n[19]);
  OR2 I184 (partCD_0n[20], store_0n[20], store_1n[20]);
  OR2 I185 (partCD_0n[21], store_0n[21], store_1n[21]);
  OR2 I186 (partCD_0n[22], store_0n[22], store_1n[22]);
  OR2 I187 (partCD_0n[23], store_0n[23], store_1n[23]);
  OR2 I188 (partCD_0n[24], store_0n[24], store_1n[24]);
  OR2 I189 (partCD_0n[25], store_0n[25], store_1n[25]);
  OR2 I190 (partCD_0n[26], store_0n[26], store_1n[26]);
  OR2 I191 (partCD_0n[27], store_0n[27], store_1n[27]);
  OR2 I192 (partCD_0n[28], store_0n[28], store_1n[28]);
  OR2 I193 (partCD_0n[29], store_0n[29], store_1n[29]);
  OR2 I194 (partCD_0n[30], store_0n[30], store_1n[30]);
  OR2 I195 (partCD_0n[31], store_0n[31], store_1n[31]);
  OR2 I196 (partCD_0n[32], store_0n[32], store_1n[32]);
  OR2 I197 (partCD_0n[33], store_0n[33], store_1n[33]);
  OR2 I198 (partCD_0n[34], store_0n[34], store_1n[34]);
  BUFF I199 (write_0r, trigger_0r);
endmodule

module BrzActiveEagerFalseVariable_35_2_s20_3_2e__m7m (
  trigger_0r, trigger_0a,
  write_0r, write_0a0d, write_0a1d,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d
);
  input trigger_0r;
  output trigger_0a;
  output write_0r;
  input [34:0] write_0a0d;
  input [34:0] write_0a1d;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output [31:0] read_0a0d;
  output [31:0] read_0a1d;
  input read_1r;
  output [2:0] read_1a0d;
  output [2:0] read_1a1d;
  wire [17:0] internal_0n;
  wire cd_0n;
  wire [34:0] partCD_0n;
  wire [34:0] store_0n;
  wire [34:0] store_1n;
  wire readReq_0n;
  wire readReq_1n;
  wire writeAck_0n;
  wire sigAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_1a1d[0], store_1n[0], readReq_1n);
  AND2 I1 (read_1a1d[1], store_1n[1], readReq_1n);
  AND2 I2 (read_1a1d[2], store_1n[2], readReq_1n);
  AND2 I3 (read_1a0d[0], store_0n[0], readReq_1n);
  AND2 I4 (read_1a0d[1], store_0n[1], readReq_1n);
  AND2 I5 (read_1a0d[2], store_0n[2], readReq_1n);
  AND2 I6 (read_0a1d[0], store_1n[3], readReq_0n);
  AND2 I7 (read_0a1d[1], store_1n[4], readReq_0n);
  AND2 I8 (read_0a1d[2], store_1n[5], readReq_0n);
  AND2 I9 (read_0a1d[3], store_1n[6], readReq_0n);
  AND2 I10 (read_0a1d[4], store_1n[7], readReq_0n);
  AND2 I11 (read_0a1d[5], store_1n[8], readReq_0n);
  AND2 I12 (read_0a1d[6], store_1n[9], readReq_0n);
  AND2 I13 (read_0a1d[7], store_1n[10], readReq_0n);
  AND2 I14 (read_0a1d[8], store_1n[11], readReq_0n);
  AND2 I15 (read_0a1d[9], store_1n[12], readReq_0n);
  AND2 I16 (read_0a1d[10], store_1n[13], readReq_0n);
  AND2 I17 (read_0a1d[11], store_1n[14], readReq_0n);
  AND2 I18 (read_0a1d[12], store_1n[15], readReq_0n);
  AND2 I19 (read_0a1d[13], store_1n[16], readReq_0n);
  AND2 I20 (read_0a1d[14], store_1n[17], readReq_0n);
  AND2 I21 (read_0a1d[15], store_1n[18], readReq_0n);
  AND2 I22 (read_0a1d[16], store_1n[19], readReq_0n);
  AND2 I23 (read_0a1d[17], store_1n[20], readReq_0n);
  AND2 I24 (read_0a1d[18], store_1n[21], readReq_0n);
  AND2 I25 (read_0a1d[19], store_1n[22], readReq_0n);
  AND2 I26 (read_0a1d[20], store_1n[23], readReq_0n);
  AND2 I27 (read_0a1d[21], store_1n[24], readReq_0n);
  AND2 I28 (read_0a1d[22], store_1n[25], readReq_0n);
  AND2 I29 (read_0a1d[23], store_1n[26], readReq_0n);
  AND2 I30 (read_0a1d[24], store_1n[27], readReq_0n);
  AND2 I31 (read_0a1d[25], store_1n[28], readReq_0n);
  AND2 I32 (read_0a1d[26], store_1n[29], readReq_0n);
  AND2 I33 (read_0a1d[27], store_1n[30], readReq_0n);
  AND2 I34 (read_0a1d[28], store_1n[31], readReq_0n);
  AND2 I35 (read_0a1d[29], store_1n[32], readReq_0n);
  AND2 I36 (read_0a1d[30], store_1n[33], readReq_0n);
  AND2 I37 (read_0a1d[31], store_1n[34], readReq_0n);
  AND2 I38 (read_0a0d[0], store_0n[3], readReq_0n);
  AND2 I39 (read_0a0d[1], store_0n[4], readReq_0n);
  AND2 I40 (read_0a0d[2], store_0n[5], readReq_0n);
  AND2 I41 (read_0a0d[3], store_0n[6], readReq_0n);
  AND2 I42 (read_0a0d[4], store_0n[7], readReq_0n);
  AND2 I43 (read_0a0d[5], store_0n[8], readReq_0n);
  AND2 I44 (read_0a0d[6], store_0n[9], readReq_0n);
  AND2 I45 (read_0a0d[7], store_0n[10], readReq_0n);
  AND2 I46 (read_0a0d[8], store_0n[11], readReq_0n);
  AND2 I47 (read_0a0d[9], store_0n[12], readReq_0n);
  AND2 I48 (read_0a0d[10], store_0n[13], readReq_0n);
  AND2 I49 (read_0a0d[11], store_0n[14], readReq_0n);
  AND2 I50 (read_0a0d[12], store_0n[15], readReq_0n);
  AND2 I51 (read_0a0d[13], store_0n[16], readReq_0n);
  AND2 I52 (read_0a0d[14], store_0n[17], readReq_0n);
  AND2 I53 (read_0a0d[15], store_0n[18], readReq_0n);
  AND2 I54 (read_0a0d[16], store_0n[19], readReq_0n);
  AND2 I55 (read_0a0d[17], store_0n[20], readReq_0n);
  AND2 I56 (read_0a0d[18], store_0n[21], readReq_0n);
  AND2 I57 (read_0a0d[19], store_0n[22], readReq_0n);
  AND2 I58 (read_0a0d[20], store_0n[23], readReq_0n);
  AND2 I59 (read_0a0d[21], store_0n[24], readReq_0n);
  AND2 I60 (read_0a0d[22], store_0n[25], readReq_0n);
  AND2 I61 (read_0a0d[23], store_0n[26], readReq_0n);
  AND2 I62 (read_0a0d[24], store_0n[27], readReq_0n);
  AND2 I63 (read_0a0d[25], store_0n[28], readReq_0n);
  AND2 I64 (read_0a0d[26], store_0n[29], readReq_0n);
  AND2 I65 (read_0a0d[27], store_0n[30], readReq_0n);
  AND2 I66 (read_0a0d[28], store_0n[31], readReq_0n);
  AND2 I67 (read_0a0d[29], store_0n[32], readReq_0n);
  AND2 I68 (read_0a0d[30], store_0n[33], readReq_0n);
  AND2 I69 (read_0a0d[31], store_0n[34], readReq_0n);
  BUFF I70 (readReq_0n, read_0r);
  BUFF I71 (readReq_1n, read_1r);
  BUFF I72 (store_1n[0], write_0a1d[0]);
  BUFF I73 (store_1n[1], write_0a1d[1]);
  BUFF I74 (store_1n[2], write_0a1d[2]);
  BUFF I75 (store_1n[3], write_0a1d[3]);
  BUFF I76 (store_1n[4], write_0a1d[4]);
  BUFF I77 (store_1n[5], write_0a1d[5]);
  BUFF I78 (store_1n[6], write_0a1d[6]);
  BUFF I79 (store_1n[7], write_0a1d[7]);
  BUFF I80 (store_1n[8], write_0a1d[8]);
  BUFF I81 (store_1n[9], write_0a1d[9]);
  BUFF I82 (store_1n[10], write_0a1d[10]);
  BUFF I83 (store_1n[11], write_0a1d[11]);
  BUFF I84 (store_1n[12], write_0a1d[12]);
  BUFF I85 (store_1n[13], write_0a1d[13]);
  BUFF I86 (store_1n[14], write_0a1d[14]);
  BUFF I87 (store_1n[15], write_0a1d[15]);
  BUFF I88 (store_1n[16], write_0a1d[16]);
  BUFF I89 (store_1n[17], write_0a1d[17]);
  BUFF I90 (store_1n[18], write_0a1d[18]);
  BUFF I91 (store_1n[19], write_0a1d[19]);
  BUFF I92 (store_1n[20], write_0a1d[20]);
  BUFF I93 (store_1n[21], write_0a1d[21]);
  BUFF I94 (store_1n[22], write_0a1d[22]);
  BUFF I95 (store_1n[23], write_0a1d[23]);
  BUFF I96 (store_1n[24], write_0a1d[24]);
  BUFF I97 (store_1n[25], write_0a1d[25]);
  BUFF I98 (store_1n[26], write_0a1d[26]);
  BUFF I99 (store_1n[27], write_0a1d[27]);
  BUFF I100 (store_1n[28], write_0a1d[28]);
  BUFF I101 (store_1n[29], write_0a1d[29]);
  BUFF I102 (store_1n[30], write_0a1d[30]);
  BUFF I103 (store_1n[31], write_0a1d[31]);
  BUFF I104 (store_1n[32], write_0a1d[32]);
  BUFF I105 (store_1n[33], write_0a1d[33]);
  BUFF I106 (store_1n[34], write_0a1d[34]);
  BUFF I107 (store_0n[0], write_0a0d[0]);
  BUFF I108 (store_0n[1], write_0a0d[1]);
  BUFF I109 (store_0n[2], write_0a0d[2]);
  BUFF I110 (store_0n[3], write_0a0d[3]);
  BUFF I111 (store_0n[4], write_0a0d[4]);
  BUFF I112 (store_0n[5], write_0a0d[5]);
  BUFF I113 (store_0n[6], write_0a0d[6]);
  BUFF I114 (store_0n[7], write_0a0d[7]);
  BUFF I115 (store_0n[8], write_0a0d[8]);
  BUFF I116 (store_0n[9], write_0a0d[9]);
  BUFF I117 (store_0n[10], write_0a0d[10]);
  BUFF I118 (store_0n[11], write_0a0d[11]);
  BUFF I119 (store_0n[12], write_0a0d[12]);
  BUFF I120 (store_0n[13], write_0a0d[13]);
  BUFF I121 (store_0n[14], write_0a0d[14]);
  BUFF I122 (store_0n[15], write_0a0d[15]);
  BUFF I123 (store_0n[16], write_0a0d[16]);
  BUFF I124 (store_0n[17], write_0a0d[17]);
  BUFF I125 (store_0n[18], write_0a0d[18]);
  BUFF I126 (store_0n[19], write_0a0d[19]);
  BUFF I127 (store_0n[20], write_0a0d[20]);
  BUFF I128 (store_0n[21], write_0a0d[21]);
  BUFF I129 (store_0n[22], write_0a0d[22]);
  BUFF I130 (store_0n[23], write_0a0d[23]);
  BUFF I131 (store_0n[24], write_0a0d[24]);
  BUFF I132 (store_0n[25], write_0a0d[25]);
  BUFF I133 (store_0n[26], write_0a0d[26]);
  BUFF I134 (store_0n[27], write_0a0d[27]);
  BUFF I135 (store_0n[28], write_0a0d[28]);
  BUFF I136 (store_0n[29], write_0a0d[29]);
  BUFF I137 (store_0n[30], write_0a0d[30]);
  BUFF I138 (store_0n[31], write_0a0d[31]);
  BUFF I139 (store_0n[32], write_0a0d[32]);
  BUFF I140 (store_0n[33], write_0a0d[33]);
  BUFF I141 (store_0n[34], write_0a0d[34]);
  C2 I142 (trigger_0a, writeAck_0n, cd_0n);
  AND2 I143 (writeAck_0n, sigAck_0n, rReqOr_0n);
  NOR2 I144 (rReqOr_0n, readReq_0n, readReq_1n);
  BALSA_TELEM I145 (trigger_0r, sigAck_0n, signal_0r, signal_0a);
  C3 I146 (internal_0n[0], partCD_0n[0], partCD_0n[1], partCD_0n[2]);
  C3 I147 (internal_0n[1], partCD_0n[3], partCD_0n[4], partCD_0n[5]);
  C3 I148 (internal_0n[2], partCD_0n[6], partCD_0n[7], partCD_0n[8]);
  C3 I149 (internal_0n[3], partCD_0n[9], partCD_0n[10], partCD_0n[11]);
  C3 I150 (internal_0n[4], partCD_0n[12], partCD_0n[13], partCD_0n[14]);
  C3 I151 (internal_0n[5], partCD_0n[15], partCD_0n[16], partCD_0n[17]);
  C3 I152 (internal_0n[6], partCD_0n[18], partCD_0n[19], partCD_0n[20]);
  C3 I153 (internal_0n[7], partCD_0n[21], partCD_0n[22], partCD_0n[23]);
  C3 I154 (internal_0n[8], partCD_0n[24], partCD_0n[25], partCD_0n[26]);
  C3 I155 (internal_0n[9], partCD_0n[27], partCD_0n[28], partCD_0n[29]);
  C3 I156 (internal_0n[10], partCD_0n[30], partCD_0n[31], partCD_0n[32]);
  C2 I157 (internal_0n[11], partCD_0n[33], partCD_0n[34]);
  C3 I158 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I159 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I160 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I161 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I162 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I163 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I164 (cd_0n, internal_0n[16], internal_0n[17]);
  OR2 I165 (partCD_0n[0], store_0n[0], store_1n[0]);
  OR2 I166 (partCD_0n[1], store_0n[1], store_1n[1]);
  OR2 I167 (partCD_0n[2], store_0n[2], store_1n[2]);
  OR2 I168 (partCD_0n[3], store_0n[3], store_1n[3]);
  OR2 I169 (partCD_0n[4], store_0n[4], store_1n[4]);
  OR2 I170 (partCD_0n[5], store_0n[5], store_1n[5]);
  OR2 I171 (partCD_0n[6], store_0n[6], store_1n[6]);
  OR2 I172 (partCD_0n[7], store_0n[7], store_1n[7]);
  OR2 I173 (partCD_0n[8], store_0n[8], store_1n[8]);
  OR2 I174 (partCD_0n[9], store_0n[9], store_1n[9]);
  OR2 I175 (partCD_0n[10], store_0n[10], store_1n[10]);
  OR2 I176 (partCD_0n[11], store_0n[11], store_1n[11]);
  OR2 I177 (partCD_0n[12], store_0n[12], store_1n[12]);
  OR2 I178 (partCD_0n[13], store_0n[13], store_1n[13]);
  OR2 I179 (partCD_0n[14], store_0n[14], store_1n[14]);
  OR2 I180 (partCD_0n[15], store_0n[15], store_1n[15]);
  OR2 I181 (partCD_0n[16], store_0n[16], store_1n[16]);
  OR2 I182 (partCD_0n[17], store_0n[17], store_1n[17]);
  OR2 I183 (partCD_0n[18], store_0n[18], store_1n[18]);
  OR2 I184 (partCD_0n[19], store_0n[19], store_1n[19]);
  OR2 I185 (partCD_0n[20], store_0n[20], store_1n[20]);
  OR2 I186 (partCD_0n[21], store_0n[21], store_1n[21]);
  OR2 I187 (partCD_0n[22], store_0n[22], store_1n[22]);
  OR2 I188 (partCD_0n[23], store_0n[23], store_1n[23]);
  OR2 I189 (partCD_0n[24], store_0n[24], store_1n[24]);
  OR2 I190 (partCD_0n[25], store_0n[25], store_1n[25]);
  OR2 I191 (partCD_0n[26], store_0n[26], store_1n[26]);
  OR2 I192 (partCD_0n[27], store_0n[27], store_1n[27]);
  OR2 I193 (partCD_0n[28], store_0n[28], store_1n[28]);
  OR2 I194 (partCD_0n[29], store_0n[29], store_1n[29]);
  OR2 I195 (partCD_0n[30], store_0n[30], store_1n[30]);
  OR2 I196 (partCD_0n[31], store_0n[31], store_1n[31]);
  OR2 I197 (partCD_0n[32], store_0n[32], store_1n[32]);
  OR2 I198 (partCD_0n[33], store_0n[33], store_1n[33]);
  OR2 I199 (partCD_0n[34], store_0n[34], store_1n[34]);
  BUFF I200 (write_0r, trigger_0r);
endmodule

module BrzActiveEagerFalseVariable_35_2_s11__3b0__m9m (
  trigger_0r, trigger_0a,
  write_0r, write_0a0d, write_0a1d,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d
);
  input trigger_0r;
  output trigger_0a;
  output write_0r;
  input [34:0] write_0a0d;
  input [34:0] write_0a1d;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output [34:0] read_0a0d;
  output [34:0] read_0a1d;
  input read_1r;
  output [1:0] read_1a0d;
  output [1:0] read_1a1d;
  wire [17:0] internal_0n;
  wire cd_0n;
  wire [34:0] partCD_0n;
  wire [34:0] store_0n;
  wire [34:0] store_1n;
  wire readReq_0n;
  wire readReq_1n;
  wire writeAck_0n;
  wire sigAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_1a1d[0], store_1n[0], readReq_1n);
  AND2 I1 (read_1a1d[1], store_1n[1], readReq_1n);
  AND2 I2 (read_1a0d[0], store_0n[0], readReq_1n);
  AND2 I3 (read_1a0d[1], store_0n[1], readReq_1n);
  AND2 I4 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I5 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I6 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I7 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I8 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I9 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I10 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I11 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I12 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I13 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I14 (read_0a1d[10], store_1n[10], readReq_0n);
  AND2 I15 (read_0a1d[11], store_1n[11], readReq_0n);
  AND2 I16 (read_0a1d[12], store_1n[12], readReq_0n);
  AND2 I17 (read_0a1d[13], store_1n[13], readReq_0n);
  AND2 I18 (read_0a1d[14], store_1n[14], readReq_0n);
  AND2 I19 (read_0a1d[15], store_1n[15], readReq_0n);
  AND2 I20 (read_0a1d[16], store_1n[16], readReq_0n);
  AND2 I21 (read_0a1d[17], store_1n[17], readReq_0n);
  AND2 I22 (read_0a1d[18], store_1n[18], readReq_0n);
  AND2 I23 (read_0a1d[19], store_1n[19], readReq_0n);
  AND2 I24 (read_0a1d[20], store_1n[20], readReq_0n);
  AND2 I25 (read_0a1d[21], store_1n[21], readReq_0n);
  AND2 I26 (read_0a1d[22], store_1n[22], readReq_0n);
  AND2 I27 (read_0a1d[23], store_1n[23], readReq_0n);
  AND2 I28 (read_0a1d[24], store_1n[24], readReq_0n);
  AND2 I29 (read_0a1d[25], store_1n[25], readReq_0n);
  AND2 I30 (read_0a1d[26], store_1n[26], readReq_0n);
  AND2 I31 (read_0a1d[27], store_1n[27], readReq_0n);
  AND2 I32 (read_0a1d[28], store_1n[28], readReq_0n);
  AND2 I33 (read_0a1d[29], store_1n[29], readReq_0n);
  AND2 I34 (read_0a1d[30], store_1n[30], readReq_0n);
  AND2 I35 (read_0a1d[31], store_1n[31], readReq_0n);
  AND2 I36 (read_0a1d[32], store_1n[32], readReq_0n);
  AND2 I37 (read_0a1d[33], store_1n[33], readReq_0n);
  AND2 I38 (read_0a1d[34], store_1n[34], readReq_0n);
  AND2 I39 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I40 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I41 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I42 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I43 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I44 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I45 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I46 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I47 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I48 (read_0a0d[9], store_0n[9], readReq_0n);
  AND2 I49 (read_0a0d[10], store_0n[10], readReq_0n);
  AND2 I50 (read_0a0d[11], store_0n[11], readReq_0n);
  AND2 I51 (read_0a0d[12], store_0n[12], readReq_0n);
  AND2 I52 (read_0a0d[13], store_0n[13], readReq_0n);
  AND2 I53 (read_0a0d[14], store_0n[14], readReq_0n);
  AND2 I54 (read_0a0d[15], store_0n[15], readReq_0n);
  AND2 I55 (read_0a0d[16], store_0n[16], readReq_0n);
  AND2 I56 (read_0a0d[17], store_0n[17], readReq_0n);
  AND2 I57 (read_0a0d[18], store_0n[18], readReq_0n);
  AND2 I58 (read_0a0d[19], store_0n[19], readReq_0n);
  AND2 I59 (read_0a0d[20], store_0n[20], readReq_0n);
  AND2 I60 (read_0a0d[21], store_0n[21], readReq_0n);
  AND2 I61 (read_0a0d[22], store_0n[22], readReq_0n);
  AND2 I62 (read_0a0d[23], store_0n[23], readReq_0n);
  AND2 I63 (read_0a0d[24], store_0n[24], readReq_0n);
  AND2 I64 (read_0a0d[25], store_0n[25], readReq_0n);
  AND2 I65 (read_0a0d[26], store_0n[26], readReq_0n);
  AND2 I66 (read_0a0d[27], store_0n[27], readReq_0n);
  AND2 I67 (read_0a0d[28], store_0n[28], readReq_0n);
  AND2 I68 (read_0a0d[29], store_0n[29], readReq_0n);
  AND2 I69 (read_0a0d[30], store_0n[30], readReq_0n);
  AND2 I70 (read_0a0d[31], store_0n[31], readReq_0n);
  AND2 I71 (read_0a0d[32], store_0n[32], readReq_0n);
  AND2 I72 (read_0a0d[33], store_0n[33], readReq_0n);
  AND2 I73 (read_0a0d[34], store_0n[34], readReq_0n);
  BUFF I74 (readReq_0n, read_0r);
  BUFF I75 (readReq_1n, read_1r);
  BUFF I76 (store_1n[0], write_0a1d[0]);
  BUFF I77 (store_1n[1], write_0a1d[1]);
  BUFF I78 (store_1n[2], write_0a1d[2]);
  BUFF I79 (store_1n[3], write_0a1d[3]);
  BUFF I80 (store_1n[4], write_0a1d[4]);
  BUFF I81 (store_1n[5], write_0a1d[5]);
  BUFF I82 (store_1n[6], write_0a1d[6]);
  BUFF I83 (store_1n[7], write_0a1d[7]);
  BUFF I84 (store_1n[8], write_0a1d[8]);
  BUFF I85 (store_1n[9], write_0a1d[9]);
  BUFF I86 (store_1n[10], write_0a1d[10]);
  BUFF I87 (store_1n[11], write_0a1d[11]);
  BUFF I88 (store_1n[12], write_0a1d[12]);
  BUFF I89 (store_1n[13], write_0a1d[13]);
  BUFF I90 (store_1n[14], write_0a1d[14]);
  BUFF I91 (store_1n[15], write_0a1d[15]);
  BUFF I92 (store_1n[16], write_0a1d[16]);
  BUFF I93 (store_1n[17], write_0a1d[17]);
  BUFF I94 (store_1n[18], write_0a1d[18]);
  BUFF I95 (store_1n[19], write_0a1d[19]);
  BUFF I96 (store_1n[20], write_0a1d[20]);
  BUFF I97 (store_1n[21], write_0a1d[21]);
  BUFF I98 (store_1n[22], write_0a1d[22]);
  BUFF I99 (store_1n[23], write_0a1d[23]);
  BUFF I100 (store_1n[24], write_0a1d[24]);
  BUFF I101 (store_1n[25], write_0a1d[25]);
  BUFF I102 (store_1n[26], write_0a1d[26]);
  BUFF I103 (store_1n[27], write_0a1d[27]);
  BUFF I104 (store_1n[28], write_0a1d[28]);
  BUFF I105 (store_1n[29], write_0a1d[29]);
  BUFF I106 (store_1n[30], write_0a1d[30]);
  BUFF I107 (store_1n[31], write_0a1d[31]);
  BUFF I108 (store_1n[32], write_0a1d[32]);
  BUFF I109 (store_1n[33], write_0a1d[33]);
  BUFF I110 (store_1n[34], write_0a1d[34]);
  BUFF I111 (store_0n[0], write_0a0d[0]);
  BUFF I112 (store_0n[1], write_0a0d[1]);
  BUFF I113 (store_0n[2], write_0a0d[2]);
  BUFF I114 (store_0n[3], write_0a0d[3]);
  BUFF I115 (store_0n[4], write_0a0d[4]);
  BUFF I116 (store_0n[5], write_0a0d[5]);
  BUFF I117 (store_0n[6], write_0a0d[6]);
  BUFF I118 (store_0n[7], write_0a0d[7]);
  BUFF I119 (store_0n[8], write_0a0d[8]);
  BUFF I120 (store_0n[9], write_0a0d[9]);
  BUFF I121 (store_0n[10], write_0a0d[10]);
  BUFF I122 (store_0n[11], write_0a0d[11]);
  BUFF I123 (store_0n[12], write_0a0d[12]);
  BUFF I124 (store_0n[13], write_0a0d[13]);
  BUFF I125 (store_0n[14], write_0a0d[14]);
  BUFF I126 (store_0n[15], write_0a0d[15]);
  BUFF I127 (store_0n[16], write_0a0d[16]);
  BUFF I128 (store_0n[17], write_0a0d[17]);
  BUFF I129 (store_0n[18], write_0a0d[18]);
  BUFF I130 (store_0n[19], write_0a0d[19]);
  BUFF I131 (store_0n[20], write_0a0d[20]);
  BUFF I132 (store_0n[21], write_0a0d[21]);
  BUFF I133 (store_0n[22], write_0a0d[22]);
  BUFF I134 (store_0n[23], write_0a0d[23]);
  BUFF I135 (store_0n[24], write_0a0d[24]);
  BUFF I136 (store_0n[25], write_0a0d[25]);
  BUFF I137 (store_0n[26], write_0a0d[26]);
  BUFF I138 (store_0n[27], write_0a0d[27]);
  BUFF I139 (store_0n[28], write_0a0d[28]);
  BUFF I140 (store_0n[29], write_0a0d[29]);
  BUFF I141 (store_0n[30], write_0a0d[30]);
  BUFF I142 (store_0n[31], write_0a0d[31]);
  BUFF I143 (store_0n[32], write_0a0d[32]);
  BUFF I144 (store_0n[33], write_0a0d[33]);
  BUFF I145 (store_0n[34], write_0a0d[34]);
  C2 I146 (trigger_0a, writeAck_0n, cd_0n);
  AND2 I147 (writeAck_0n, sigAck_0n, rReqOr_0n);
  NOR2 I148 (rReqOr_0n, readReq_0n, readReq_1n);
  BALSA_TELEM I149 (trigger_0r, sigAck_0n, signal_0r, signal_0a);
  C3 I150 (internal_0n[0], partCD_0n[0], partCD_0n[1], partCD_0n[2]);
  C3 I151 (internal_0n[1], partCD_0n[3], partCD_0n[4], partCD_0n[5]);
  C3 I152 (internal_0n[2], partCD_0n[6], partCD_0n[7], partCD_0n[8]);
  C3 I153 (internal_0n[3], partCD_0n[9], partCD_0n[10], partCD_0n[11]);
  C3 I154 (internal_0n[4], partCD_0n[12], partCD_0n[13], partCD_0n[14]);
  C3 I155 (internal_0n[5], partCD_0n[15], partCD_0n[16], partCD_0n[17]);
  C3 I156 (internal_0n[6], partCD_0n[18], partCD_0n[19], partCD_0n[20]);
  C3 I157 (internal_0n[7], partCD_0n[21], partCD_0n[22], partCD_0n[23]);
  C3 I158 (internal_0n[8], partCD_0n[24], partCD_0n[25], partCD_0n[26]);
  C3 I159 (internal_0n[9], partCD_0n[27], partCD_0n[28], partCD_0n[29]);
  C3 I160 (internal_0n[10], partCD_0n[30], partCD_0n[31], partCD_0n[32]);
  C2 I161 (internal_0n[11], partCD_0n[33], partCD_0n[34]);
  C3 I162 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I163 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I164 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I165 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I166 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I167 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I168 (cd_0n, internal_0n[16], internal_0n[17]);
  OR2 I169 (partCD_0n[0], store_0n[0], store_1n[0]);
  OR2 I170 (partCD_0n[1], store_0n[1], store_1n[1]);
  OR2 I171 (partCD_0n[2], store_0n[2], store_1n[2]);
  OR2 I172 (partCD_0n[3], store_0n[3], store_1n[3]);
  OR2 I173 (partCD_0n[4], store_0n[4], store_1n[4]);
  OR2 I174 (partCD_0n[5], store_0n[5], store_1n[5]);
  OR2 I175 (partCD_0n[6], store_0n[6], store_1n[6]);
  OR2 I176 (partCD_0n[7], store_0n[7], store_1n[7]);
  OR2 I177 (partCD_0n[8], store_0n[8], store_1n[8]);
  OR2 I178 (partCD_0n[9], store_0n[9], store_1n[9]);
  OR2 I179 (partCD_0n[10], store_0n[10], store_1n[10]);
  OR2 I180 (partCD_0n[11], store_0n[11], store_1n[11]);
  OR2 I181 (partCD_0n[12], store_0n[12], store_1n[12]);
  OR2 I182 (partCD_0n[13], store_0n[13], store_1n[13]);
  OR2 I183 (partCD_0n[14], store_0n[14], store_1n[14]);
  OR2 I184 (partCD_0n[15], store_0n[15], store_1n[15]);
  OR2 I185 (partCD_0n[16], store_0n[16], store_1n[16]);
  OR2 I186 (partCD_0n[17], store_0n[17], store_1n[17]);
  OR2 I187 (partCD_0n[18], store_0n[18], store_1n[18]);
  OR2 I188 (partCD_0n[19], store_0n[19], store_1n[19]);
  OR2 I189 (partCD_0n[20], store_0n[20], store_1n[20]);
  OR2 I190 (partCD_0n[21], store_0n[21], store_1n[21]);
  OR2 I191 (partCD_0n[22], store_0n[22], store_1n[22]);
  OR2 I192 (partCD_0n[23], store_0n[23], store_1n[23]);
  OR2 I193 (partCD_0n[24], store_0n[24], store_1n[24]);
  OR2 I194 (partCD_0n[25], store_0n[25], store_1n[25]);
  OR2 I195 (partCD_0n[26], store_0n[26], store_1n[26]);
  OR2 I196 (partCD_0n[27], store_0n[27], store_1n[27]);
  OR2 I197 (partCD_0n[28], store_0n[28], store_1n[28]);
  OR2 I198 (partCD_0n[29], store_0n[29], store_1n[29]);
  OR2 I199 (partCD_0n[30], store_0n[30], store_1n[30]);
  OR2 I200 (partCD_0n[31], store_0n[31], store_1n[31]);
  OR2 I201 (partCD_0n[32], store_0n[32], store_1n[32]);
  OR2 I202 (partCD_0n[33], store_0n[33], store_1n[33]);
  OR2 I203 (partCD_0n[34], store_0n[34], store_1n[34]);
  BUFF I204 (write_0r, trigger_0r);
endmodule

module BrzActiveEagerFalseVariable_35_3_s0_ (
  trigger_0r, trigger_0a,
  write_0r, write_0a0d, write_0a1d,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d,
  read_2r, read_2a0d, read_2a1d
);
  input trigger_0r;
  output trigger_0a;
  output write_0r;
  input [34:0] write_0a0d;
  input [34:0] write_0a1d;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output [34:0] read_0a0d;
  output [34:0] read_0a1d;
  input read_1r;
  output [34:0] read_1a0d;
  output [34:0] read_1a1d;
  input read_2r;
  output [34:0] read_2a0d;
  output [34:0] read_2a1d;
  wire [17:0] internal_0n;
  wire cd_0n;
  wire [34:0] partCD_0n;
  wire [34:0] store_0n;
  wire [34:0] store_1n;
  wire readReq_0n;
  wire readReq_1n;
  wire readReq_2n;
  wire writeAck_0n;
  wire sigAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_2a1d[0], store_1n[0], readReq_2n);
  AND2 I1 (read_2a1d[1], store_1n[1], readReq_2n);
  AND2 I2 (read_2a1d[2], store_1n[2], readReq_2n);
  AND2 I3 (read_2a1d[3], store_1n[3], readReq_2n);
  AND2 I4 (read_2a1d[4], store_1n[4], readReq_2n);
  AND2 I5 (read_2a1d[5], store_1n[5], readReq_2n);
  AND2 I6 (read_2a1d[6], store_1n[6], readReq_2n);
  AND2 I7 (read_2a1d[7], store_1n[7], readReq_2n);
  AND2 I8 (read_2a1d[8], store_1n[8], readReq_2n);
  AND2 I9 (read_2a1d[9], store_1n[9], readReq_2n);
  AND2 I10 (read_2a1d[10], store_1n[10], readReq_2n);
  AND2 I11 (read_2a1d[11], store_1n[11], readReq_2n);
  AND2 I12 (read_2a1d[12], store_1n[12], readReq_2n);
  AND2 I13 (read_2a1d[13], store_1n[13], readReq_2n);
  AND2 I14 (read_2a1d[14], store_1n[14], readReq_2n);
  AND2 I15 (read_2a1d[15], store_1n[15], readReq_2n);
  AND2 I16 (read_2a1d[16], store_1n[16], readReq_2n);
  AND2 I17 (read_2a1d[17], store_1n[17], readReq_2n);
  AND2 I18 (read_2a1d[18], store_1n[18], readReq_2n);
  AND2 I19 (read_2a1d[19], store_1n[19], readReq_2n);
  AND2 I20 (read_2a1d[20], store_1n[20], readReq_2n);
  AND2 I21 (read_2a1d[21], store_1n[21], readReq_2n);
  AND2 I22 (read_2a1d[22], store_1n[22], readReq_2n);
  AND2 I23 (read_2a1d[23], store_1n[23], readReq_2n);
  AND2 I24 (read_2a1d[24], store_1n[24], readReq_2n);
  AND2 I25 (read_2a1d[25], store_1n[25], readReq_2n);
  AND2 I26 (read_2a1d[26], store_1n[26], readReq_2n);
  AND2 I27 (read_2a1d[27], store_1n[27], readReq_2n);
  AND2 I28 (read_2a1d[28], store_1n[28], readReq_2n);
  AND2 I29 (read_2a1d[29], store_1n[29], readReq_2n);
  AND2 I30 (read_2a1d[30], store_1n[30], readReq_2n);
  AND2 I31 (read_2a1d[31], store_1n[31], readReq_2n);
  AND2 I32 (read_2a1d[32], store_1n[32], readReq_2n);
  AND2 I33 (read_2a1d[33], store_1n[33], readReq_2n);
  AND2 I34 (read_2a1d[34], store_1n[34], readReq_2n);
  AND2 I35 (read_2a0d[0], store_0n[0], readReq_2n);
  AND2 I36 (read_2a0d[1], store_0n[1], readReq_2n);
  AND2 I37 (read_2a0d[2], store_0n[2], readReq_2n);
  AND2 I38 (read_2a0d[3], store_0n[3], readReq_2n);
  AND2 I39 (read_2a0d[4], store_0n[4], readReq_2n);
  AND2 I40 (read_2a0d[5], store_0n[5], readReq_2n);
  AND2 I41 (read_2a0d[6], store_0n[6], readReq_2n);
  AND2 I42 (read_2a0d[7], store_0n[7], readReq_2n);
  AND2 I43 (read_2a0d[8], store_0n[8], readReq_2n);
  AND2 I44 (read_2a0d[9], store_0n[9], readReq_2n);
  AND2 I45 (read_2a0d[10], store_0n[10], readReq_2n);
  AND2 I46 (read_2a0d[11], store_0n[11], readReq_2n);
  AND2 I47 (read_2a0d[12], store_0n[12], readReq_2n);
  AND2 I48 (read_2a0d[13], store_0n[13], readReq_2n);
  AND2 I49 (read_2a0d[14], store_0n[14], readReq_2n);
  AND2 I50 (read_2a0d[15], store_0n[15], readReq_2n);
  AND2 I51 (read_2a0d[16], store_0n[16], readReq_2n);
  AND2 I52 (read_2a0d[17], store_0n[17], readReq_2n);
  AND2 I53 (read_2a0d[18], store_0n[18], readReq_2n);
  AND2 I54 (read_2a0d[19], store_0n[19], readReq_2n);
  AND2 I55 (read_2a0d[20], store_0n[20], readReq_2n);
  AND2 I56 (read_2a0d[21], store_0n[21], readReq_2n);
  AND2 I57 (read_2a0d[22], store_0n[22], readReq_2n);
  AND2 I58 (read_2a0d[23], store_0n[23], readReq_2n);
  AND2 I59 (read_2a0d[24], store_0n[24], readReq_2n);
  AND2 I60 (read_2a0d[25], store_0n[25], readReq_2n);
  AND2 I61 (read_2a0d[26], store_0n[26], readReq_2n);
  AND2 I62 (read_2a0d[27], store_0n[27], readReq_2n);
  AND2 I63 (read_2a0d[28], store_0n[28], readReq_2n);
  AND2 I64 (read_2a0d[29], store_0n[29], readReq_2n);
  AND2 I65 (read_2a0d[30], store_0n[30], readReq_2n);
  AND2 I66 (read_2a0d[31], store_0n[31], readReq_2n);
  AND2 I67 (read_2a0d[32], store_0n[32], readReq_2n);
  AND2 I68 (read_2a0d[33], store_0n[33], readReq_2n);
  AND2 I69 (read_2a0d[34], store_0n[34], readReq_2n);
  AND2 I70 (read_1a1d[0], store_1n[0], readReq_1n);
  AND2 I71 (read_1a1d[1], store_1n[1], readReq_1n);
  AND2 I72 (read_1a1d[2], store_1n[2], readReq_1n);
  AND2 I73 (read_1a1d[3], store_1n[3], readReq_1n);
  AND2 I74 (read_1a1d[4], store_1n[4], readReq_1n);
  AND2 I75 (read_1a1d[5], store_1n[5], readReq_1n);
  AND2 I76 (read_1a1d[6], store_1n[6], readReq_1n);
  AND2 I77 (read_1a1d[7], store_1n[7], readReq_1n);
  AND2 I78 (read_1a1d[8], store_1n[8], readReq_1n);
  AND2 I79 (read_1a1d[9], store_1n[9], readReq_1n);
  AND2 I80 (read_1a1d[10], store_1n[10], readReq_1n);
  AND2 I81 (read_1a1d[11], store_1n[11], readReq_1n);
  AND2 I82 (read_1a1d[12], store_1n[12], readReq_1n);
  AND2 I83 (read_1a1d[13], store_1n[13], readReq_1n);
  AND2 I84 (read_1a1d[14], store_1n[14], readReq_1n);
  AND2 I85 (read_1a1d[15], store_1n[15], readReq_1n);
  AND2 I86 (read_1a1d[16], store_1n[16], readReq_1n);
  AND2 I87 (read_1a1d[17], store_1n[17], readReq_1n);
  AND2 I88 (read_1a1d[18], store_1n[18], readReq_1n);
  AND2 I89 (read_1a1d[19], store_1n[19], readReq_1n);
  AND2 I90 (read_1a1d[20], store_1n[20], readReq_1n);
  AND2 I91 (read_1a1d[21], store_1n[21], readReq_1n);
  AND2 I92 (read_1a1d[22], store_1n[22], readReq_1n);
  AND2 I93 (read_1a1d[23], store_1n[23], readReq_1n);
  AND2 I94 (read_1a1d[24], store_1n[24], readReq_1n);
  AND2 I95 (read_1a1d[25], store_1n[25], readReq_1n);
  AND2 I96 (read_1a1d[26], store_1n[26], readReq_1n);
  AND2 I97 (read_1a1d[27], store_1n[27], readReq_1n);
  AND2 I98 (read_1a1d[28], store_1n[28], readReq_1n);
  AND2 I99 (read_1a1d[29], store_1n[29], readReq_1n);
  AND2 I100 (read_1a1d[30], store_1n[30], readReq_1n);
  AND2 I101 (read_1a1d[31], store_1n[31], readReq_1n);
  AND2 I102 (read_1a1d[32], store_1n[32], readReq_1n);
  AND2 I103 (read_1a1d[33], store_1n[33], readReq_1n);
  AND2 I104 (read_1a1d[34], store_1n[34], readReq_1n);
  AND2 I105 (read_1a0d[0], store_0n[0], readReq_1n);
  AND2 I106 (read_1a0d[1], store_0n[1], readReq_1n);
  AND2 I107 (read_1a0d[2], store_0n[2], readReq_1n);
  AND2 I108 (read_1a0d[3], store_0n[3], readReq_1n);
  AND2 I109 (read_1a0d[4], store_0n[4], readReq_1n);
  AND2 I110 (read_1a0d[5], store_0n[5], readReq_1n);
  AND2 I111 (read_1a0d[6], store_0n[6], readReq_1n);
  AND2 I112 (read_1a0d[7], store_0n[7], readReq_1n);
  AND2 I113 (read_1a0d[8], store_0n[8], readReq_1n);
  AND2 I114 (read_1a0d[9], store_0n[9], readReq_1n);
  AND2 I115 (read_1a0d[10], store_0n[10], readReq_1n);
  AND2 I116 (read_1a0d[11], store_0n[11], readReq_1n);
  AND2 I117 (read_1a0d[12], store_0n[12], readReq_1n);
  AND2 I118 (read_1a0d[13], store_0n[13], readReq_1n);
  AND2 I119 (read_1a0d[14], store_0n[14], readReq_1n);
  AND2 I120 (read_1a0d[15], store_0n[15], readReq_1n);
  AND2 I121 (read_1a0d[16], store_0n[16], readReq_1n);
  AND2 I122 (read_1a0d[17], store_0n[17], readReq_1n);
  AND2 I123 (read_1a0d[18], store_0n[18], readReq_1n);
  AND2 I124 (read_1a0d[19], store_0n[19], readReq_1n);
  AND2 I125 (read_1a0d[20], store_0n[20], readReq_1n);
  AND2 I126 (read_1a0d[21], store_0n[21], readReq_1n);
  AND2 I127 (read_1a0d[22], store_0n[22], readReq_1n);
  AND2 I128 (read_1a0d[23], store_0n[23], readReq_1n);
  AND2 I129 (read_1a0d[24], store_0n[24], readReq_1n);
  AND2 I130 (read_1a0d[25], store_0n[25], readReq_1n);
  AND2 I131 (read_1a0d[26], store_0n[26], readReq_1n);
  AND2 I132 (read_1a0d[27], store_0n[27], readReq_1n);
  AND2 I133 (read_1a0d[28], store_0n[28], readReq_1n);
  AND2 I134 (read_1a0d[29], store_0n[29], readReq_1n);
  AND2 I135 (read_1a0d[30], store_0n[30], readReq_1n);
  AND2 I136 (read_1a0d[31], store_0n[31], readReq_1n);
  AND2 I137 (read_1a0d[32], store_0n[32], readReq_1n);
  AND2 I138 (read_1a0d[33], store_0n[33], readReq_1n);
  AND2 I139 (read_1a0d[34], store_0n[34], readReq_1n);
  AND2 I140 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I141 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I142 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I143 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I144 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I145 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I146 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I147 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I148 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I149 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I150 (read_0a1d[10], store_1n[10], readReq_0n);
  AND2 I151 (read_0a1d[11], store_1n[11], readReq_0n);
  AND2 I152 (read_0a1d[12], store_1n[12], readReq_0n);
  AND2 I153 (read_0a1d[13], store_1n[13], readReq_0n);
  AND2 I154 (read_0a1d[14], store_1n[14], readReq_0n);
  AND2 I155 (read_0a1d[15], store_1n[15], readReq_0n);
  AND2 I156 (read_0a1d[16], store_1n[16], readReq_0n);
  AND2 I157 (read_0a1d[17], store_1n[17], readReq_0n);
  AND2 I158 (read_0a1d[18], store_1n[18], readReq_0n);
  AND2 I159 (read_0a1d[19], store_1n[19], readReq_0n);
  AND2 I160 (read_0a1d[20], store_1n[20], readReq_0n);
  AND2 I161 (read_0a1d[21], store_1n[21], readReq_0n);
  AND2 I162 (read_0a1d[22], store_1n[22], readReq_0n);
  AND2 I163 (read_0a1d[23], store_1n[23], readReq_0n);
  AND2 I164 (read_0a1d[24], store_1n[24], readReq_0n);
  AND2 I165 (read_0a1d[25], store_1n[25], readReq_0n);
  AND2 I166 (read_0a1d[26], store_1n[26], readReq_0n);
  AND2 I167 (read_0a1d[27], store_1n[27], readReq_0n);
  AND2 I168 (read_0a1d[28], store_1n[28], readReq_0n);
  AND2 I169 (read_0a1d[29], store_1n[29], readReq_0n);
  AND2 I170 (read_0a1d[30], store_1n[30], readReq_0n);
  AND2 I171 (read_0a1d[31], store_1n[31], readReq_0n);
  AND2 I172 (read_0a1d[32], store_1n[32], readReq_0n);
  AND2 I173 (read_0a1d[33], store_1n[33], readReq_0n);
  AND2 I174 (read_0a1d[34], store_1n[34], readReq_0n);
  AND2 I175 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I176 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I177 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I178 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I179 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I180 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I181 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I182 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I183 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I184 (read_0a0d[9], store_0n[9], readReq_0n);
  AND2 I185 (read_0a0d[10], store_0n[10], readReq_0n);
  AND2 I186 (read_0a0d[11], store_0n[11], readReq_0n);
  AND2 I187 (read_0a0d[12], store_0n[12], readReq_0n);
  AND2 I188 (read_0a0d[13], store_0n[13], readReq_0n);
  AND2 I189 (read_0a0d[14], store_0n[14], readReq_0n);
  AND2 I190 (read_0a0d[15], store_0n[15], readReq_0n);
  AND2 I191 (read_0a0d[16], store_0n[16], readReq_0n);
  AND2 I192 (read_0a0d[17], store_0n[17], readReq_0n);
  AND2 I193 (read_0a0d[18], store_0n[18], readReq_0n);
  AND2 I194 (read_0a0d[19], store_0n[19], readReq_0n);
  AND2 I195 (read_0a0d[20], store_0n[20], readReq_0n);
  AND2 I196 (read_0a0d[21], store_0n[21], readReq_0n);
  AND2 I197 (read_0a0d[22], store_0n[22], readReq_0n);
  AND2 I198 (read_0a0d[23], store_0n[23], readReq_0n);
  AND2 I199 (read_0a0d[24], store_0n[24], readReq_0n);
  AND2 I200 (read_0a0d[25], store_0n[25], readReq_0n);
  AND2 I201 (read_0a0d[26], store_0n[26], readReq_0n);
  AND2 I202 (read_0a0d[27], store_0n[27], readReq_0n);
  AND2 I203 (read_0a0d[28], store_0n[28], readReq_0n);
  AND2 I204 (read_0a0d[29], store_0n[29], readReq_0n);
  AND2 I205 (read_0a0d[30], store_0n[30], readReq_0n);
  AND2 I206 (read_0a0d[31], store_0n[31], readReq_0n);
  AND2 I207 (read_0a0d[32], store_0n[32], readReq_0n);
  AND2 I208 (read_0a0d[33], store_0n[33], readReq_0n);
  AND2 I209 (read_0a0d[34], store_0n[34], readReq_0n);
  BUFF I210 (readReq_0n, read_0r);
  BUFF I211 (readReq_1n, read_1r);
  BUFF I212 (readReq_2n, read_2r);
  BUFF I213 (store_1n[0], write_0a1d[0]);
  BUFF I214 (store_1n[1], write_0a1d[1]);
  BUFF I215 (store_1n[2], write_0a1d[2]);
  BUFF I216 (store_1n[3], write_0a1d[3]);
  BUFF I217 (store_1n[4], write_0a1d[4]);
  BUFF I218 (store_1n[5], write_0a1d[5]);
  BUFF I219 (store_1n[6], write_0a1d[6]);
  BUFF I220 (store_1n[7], write_0a1d[7]);
  BUFF I221 (store_1n[8], write_0a1d[8]);
  BUFF I222 (store_1n[9], write_0a1d[9]);
  BUFF I223 (store_1n[10], write_0a1d[10]);
  BUFF I224 (store_1n[11], write_0a1d[11]);
  BUFF I225 (store_1n[12], write_0a1d[12]);
  BUFF I226 (store_1n[13], write_0a1d[13]);
  BUFF I227 (store_1n[14], write_0a1d[14]);
  BUFF I228 (store_1n[15], write_0a1d[15]);
  BUFF I229 (store_1n[16], write_0a1d[16]);
  BUFF I230 (store_1n[17], write_0a1d[17]);
  BUFF I231 (store_1n[18], write_0a1d[18]);
  BUFF I232 (store_1n[19], write_0a1d[19]);
  BUFF I233 (store_1n[20], write_0a1d[20]);
  BUFF I234 (store_1n[21], write_0a1d[21]);
  BUFF I235 (store_1n[22], write_0a1d[22]);
  BUFF I236 (store_1n[23], write_0a1d[23]);
  BUFF I237 (store_1n[24], write_0a1d[24]);
  BUFF I238 (store_1n[25], write_0a1d[25]);
  BUFF I239 (store_1n[26], write_0a1d[26]);
  BUFF I240 (store_1n[27], write_0a1d[27]);
  BUFF I241 (store_1n[28], write_0a1d[28]);
  BUFF I242 (store_1n[29], write_0a1d[29]);
  BUFF I243 (store_1n[30], write_0a1d[30]);
  BUFF I244 (store_1n[31], write_0a1d[31]);
  BUFF I245 (store_1n[32], write_0a1d[32]);
  BUFF I246 (store_1n[33], write_0a1d[33]);
  BUFF I247 (store_1n[34], write_0a1d[34]);
  BUFF I248 (store_0n[0], write_0a0d[0]);
  BUFF I249 (store_0n[1], write_0a0d[1]);
  BUFF I250 (store_0n[2], write_0a0d[2]);
  BUFF I251 (store_0n[3], write_0a0d[3]);
  BUFF I252 (store_0n[4], write_0a0d[4]);
  BUFF I253 (store_0n[5], write_0a0d[5]);
  BUFF I254 (store_0n[6], write_0a0d[6]);
  BUFF I255 (store_0n[7], write_0a0d[7]);
  BUFF I256 (store_0n[8], write_0a0d[8]);
  BUFF I257 (store_0n[9], write_0a0d[9]);
  BUFF I258 (store_0n[10], write_0a0d[10]);
  BUFF I259 (store_0n[11], write_0a0d[11]);
  BUFF I260 (store_0n[12], write_0a0d[12]);
  BUFF I261 (store_0n[13], write_0a0d[13]);
  BUFF I262 (store_0n[14], write_0a0d[14]);
  BUFF I263 (store_0n[15], write_0a0d[15]);
  BUFF I264 (store_0n[16], write_0a0d[16]);
  BUFF I265 (store_0n[17], write_0a0d[17]);
  BUFF I266 (store_0n[18], write_0a0d[18]);
  BUFF I267 (store_0n[19], write_0a0d[19]);
  BUFF I268 (store_0n[20], write_0a0d[20]);
  BUFF I269 (store_0n[21], write_0a0d[21]);
  BUFF I270 (store_0n[22], write_0a0d[22]);
  BUFF I271 (store_0n[23], write_0a0d[23]);
  BUFF I272 (store_0n[24], write_0a0d[24]);
  BUFF I273 (store_0n[25], write_0a0d[25]);
  BUFF I274 (store_0n[26], write_0a0d[26]);
  BUFF I275 (store_0n[27], write_0a0d[27]);
  BUFF I276 (store_0n[28], write_0a0d[28]);
  BUFF I277 (store_0n[29], write_0a0d[29]);
  BUFF I278 (store_0n[30], write_0a0d[30]);
  BUFF I279 (store_0n[31], write_0a0d[31]);
  BUFF I280 (store_0n[32], write_0a0d[32]);
  BUFF I281 (store_0n[33], write_0a0d[33]);
  BUFF I282 (store_0n[34], write_0a0d[34]);
  C2 I283 (trigger_0a, writeAck_0n, cd_0n);
  AND2 I284 (writeAck_0n, sigAck_0n, rReqOr_0n);
  NOR3 I285 (rReqOr_0n, readReq_0n, readReq_1n, readReq_2n);
  BALSA_TELEM I286 (trigger_0r, sigAck_0n, signal_0r, signal_0a);
  C3 I287 (internal_0n[0], partCD_0n[0], partCD_0n[1], partCD_0n[2]);
  C3 I288 (internal_0n[1], partCD_0n[3], partCD_0n[4], partCD_0n[5]);
  C3 I289 (internal_0n[2], partCD_0n[6], partCD_0n[7], partCD_0n[8]);
  C3 I290 (internal_0n[3], partCD_0n[9], partCD_0n[10], partCD_0n[11]);
  C3 I291 (internal_0n[4], partCD_0n[12], partCD_0n[13], partCD_0n[14]);
  C3 I292 (internal_0n[5], partCD_0n[15], partCD_0n[16], partCD_0n[17]);
  C3 I293 (internal_0n[6], partCD_0n[18], partCD_0n[19], partCD_0n[20]);
  C3 I294 (internal_0n[7], partCD_0n[21], partCD_0n[22], partCD_0n[23]);
  C3 I295 (internal_0n[8], partCD_0n[24], partCD_0n[25], partCD_0n[26]);
  C3 I296 (internal_0n[9], partCD_0n[27], partCD_0n[28], partCD_0n[29]);
  C3 I297 (internal_0n[10], partCD_0n[30], partCD_0n[31], partCD_0n[32]);
  C2 I298 (internal_0n[11], partCD_0n[33], partCD_0n[34]);
  C3 I299 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I300 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I301 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I302 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I303 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I304 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I305 (cd_0n, internal_0n[16], internal_0n[17]);
  OR2 I306 (partCD_0n[0], store_0n[0], store_1n[0]);
  OR2 I307 (partCD_0n[1], store_0n[1], store_1n[1]);
  OR2 I308 (partCD_0n[2], store_0n[2], store_1n[2]);
  OR2 I309 (partCD_0n[3], store_0n[3], store_1n[3]);
  OR2 I310 (partCD_0n[4], store_0n[4], store_1n[4]);
  OR2 I311 (partCD_0n[5], store_0n[5], store_1n[5]);
  OR2 I312 (partCD_0n[6], store_0n[6], store_1n[6]);
  OR2 I313 (partCD_0n[7], store_0n[7], store_1n[7]);
  OR2 I314 (partCD_0n[8], store_0n[8], store_1n[8]);
  OR2 I315 (partCD_0n[9], store_0n[9], store_1n[9]);
  OR2 I316 (partCD_0n[10], store_0n[10], store_1n[10]);
  OR2 I317 (partCD_0n[11], store_0n[11], store_1n[11]);
  OR2 I318 (partCD_0n[12], store_0n[12], store_1n[12]);
  OR2 I319 (partCD_0n[13], store_0n[13], store_1n[13]);
  OR2 I320 (partCD_0n[14], store_0n[14], store_1n[14]);
  OR2 I321 (partCD_0n[15], store_0n[15], store_1n[15]);
  OR2 I322 (partCD_0n[16], store_0n[16], store_1n[16]);
  OR2 I323 (partCD_0n[17], store_0n[17], store_1n[17]);
  OR2 I324 (partCD_0n[18], store_0n[18], store_1n[18]);
  OR2 I325 (partCD_0n[19], store_0n[19], store_1n[19]);
  OR2 I326 (partCD_0n[20], store_0n[20], store_1n[20]);
  OR2 I327 (partCD_0n[21], store_0n[21], store_1n[21]);
  OR2 I328 (partCD_0n[22], store_0n[22], store_1n[22]);
  OR2 I329 (partCD_0n[23], store_0n[23], store_1n[23]);
  OR2 I330 (partCD_0n[24], store_0n[24], store_1n[24]);
  OR2 I331 (partCD_0n[25], store_0n[25], store_1n[25]);
  OR2 I332 (partCD_0n[26], store_0n[26], store_1n[26]);
  OR2 I333 (partCD_0n[27], store_0n[27], store_1n[27]);
  OR2 I334 (partCD_0n[28], store_0n[28], store_1n[28]);
  OR2 I335 (partCD_0n[29], store_0n[29], store_1n[29]);
  OR2 I336 (partCD_0n[30], store_0n[30], store_1n[30]);
  OR2 I337 (partCD_0n[31], store_0n[31], store_1n[31]);
  OR2 I338 (partCD_0n[32], store_0n[32], store_1n[32]);
  OR2 I339 (partCD_0n[33], store_0n[33], store_1n[33]);
  OR2 I340 (partCD_0n[34], store_0n[34], store_1n[34]);
  BUFF I341 (write_0r, trigger_0r);
endmodule

module BrzActiveEagerFalseVariable_35_7_s63__3b0__m11m (
  trigger_0r, trigger_0a,
  write_0r, write_0a0d, write_0a1d,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d,
  read_2r, read_2a0d, read_2a1d,
  read_3r, read_3a0d, read_3a1d,
  read_4r, read_4a0d, read_4a1d,
  read_5r, read_5a0d, read_5a1d,
  read_6r, read_6a0d, read_6a1d
);
  input trigger_0r;
  output trigger_0a;
  output write_0r;
  input [34:0] write_0a0d;
  input [34:0] write_0a1d;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output [34:0] read_0a0d;
  output [34:0] read_0a1d;
  input read_1r;
  output [33:0] read_1a0d;
  output [33:0] read_1a1d;
  input read_2r;
  output [32:0] read_2a0d;
  output [32:0] read_2a1d;
  input read_3r;
  output [31:0] read_3a0d;
  output [31:0] read_3a1d;
  input read_4r;
  output [34:0] read_4a0d;
  output [34:0] read_4a1d;
  input read_5r;
  output read_5a0d;
  output read_5a1d;
  input read_6r;
  output read_6a0d;
  output read_6a1d;
  wire [20:0] internal_0n;
  wire cd_0n;
  wire [34:0] partCD_0n;
  wire [34:0] store_0n;
  wire [34:0] store_1n;
  wire readReq_0n;
  wire readReq_1n;
  wire readReq_2n;
  wire readReq_3n;
  wire readReq_4n;
  wire readReq_5n;
  wire readReq_6n;
  wire writeAck_0n;
  wire sigAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_6a1d, store_1n[32], readReq_6n);
  AND2 I1 (read_6a0d, store_0n[32], readReq_6n);
  AND2 I2 (read_5a1d, store_1n[0], readReq_5n);
  AND2 I3 (read_5a0d, store_0n[0], readReq_5n);
  AND2 I4 (read_4a1d[0], store_1n[0], readReq_4n);
  AND2 I5 (read_4a1d[1], store_1n[1], readReq_4n);
  AND2 I6 (read_4a1d[2], store_1n[2], readReq_4n);
  AND2 I7 (read_4a1d[3], store_1n[3], readReq_4n);
  AND2 I8 (read_4a1d[4], store_1n[4], readReq_4n);
  AND2 I9 (read_4a1d[5], store_1n[5], readReq_4n);
  AND2 I10 (read_4a1d[6], store_1n[6], readReq_4n);
  AND2 I11 (read_4a1d[7], store_1n[7], readReq_4n);
  AND2 I12 (read_4a1d[8], store_1n[8], readReq_4n);
  AND2 I13 (read_4a1d[9], store_1n[9], readReq_4n);
  AND2 I14 (read_4a1d[10], store_1n[10], readReq_4n);
  AND2 I15 (read_4a1d[11], store_1n[11], readReq_4n);
  AND2 I16 (read_4a1d[12], store_1n[12], readReq_4n);
  AND2 I17 (read_4a1d[13], store_1n[13], readReq_4n);
  AND2 I18 (read_4a1d[14], store_1n[14], readReq_4n);
  AND2 I19 (read_4a1d[15], store_1n[15], readReq_4n);
  AND2 I20 (read_4a1d[16], store_1n[16], readReq_4n);
  AND2 I21 (read_4a1d[17], store_1n[17], readReq_4n);
  AND2 I22 (read_4a1d[18], store_1n[18], readReq_4n);
  AND2 I23 (read_4a1d[19], store_1n[19], readReq_4n);
  AND2 I24 (read_4a1d[20], store_1n[20], readReq_4n);
  AND2 I25 (read_4a1d[21], store_1n[21], readReq_4n);
  AND2 I26 (read_4a1d[22], store_1n[22], readReq_4n);
  AND2 I27 (read_4a1d[23], store_1n[23], readReq_4n);
  AND2 I28 (read_4a1d[24], store_1n[24], readReq_4n);
  AND2 I29 (read_4a1d[25], store_1n[25], readReq_4n);
  AND2 I30 (read_4a1d[26], store_1n[26], readReq_4n);
  AND2 I31 (read_4a1d[27], store_1n[27], readReq_4n);
  AND2 I32 (read_4a1d[28], store_1n[28], readReq_4n);
  AND2 I33 (read_4a1d[29], store_1n[29], readReq_4n);
  AND2 I34 (read_4a1d[30], store_1n[30], readReq_4n);
  AND2 I35 (read_4a1d[31], store_1n[31], readReq_4n);
  AND2 I36 (read_4a1d[32], store_1n[32], readReq_4n);
  AND2 I37 (read_4a1d[33], store_1n[33], readReq_4n);
  AND2 I38 (read_4a1d[34], store_1n[34], readReq_4n);
  AND2 I39 (read_4a0d[0], store_0n[0], readReq_4n);
  AND2 I40 (read_4a0d[1], store_0n[1], readReq_4n);
  AND2 I41 (read_4a0d[2], store_0n[2], readReq_4n);
  AND2 I42 (read_4a0d[3], store_0n[3], readReq_4n);
  AND2 I43 (read_4a0d[4], store_0n[4], readReq_4n);
  AND2 I44 (read_4a0d[5], store_0n[5], readReq_4n);
  AND2 I45 (read_4a0d[6], store_0n[6], readReq_4n);
  AND2 I46 (read_4a0d[7], store_0n[7], readReq_4n);
  AND2 I47 (read_4a0d[8], store_0n[8], readReq_4n);
  AND2 I48 (read_4a0d[9], store_0n[9], readReq_4n);
  AND2 I49 (read_4a0d[10], store_0n[10], readReq_4n);
  AND2 I50 (read_4a0d[11], store_0n[11], readReq_4n);
  AND2 I51 (read_4a0d[12], store_0n[12], readReq_4n);
  AND2 I52 (read_4a0d[13], store_0n[13], readReq_4n);
  AND2 I53 (read_4a0d[14], store_0n[14], readReq_4n);
  AND2 I54 (read_4a0d[15], store_0n[15], readReq_4n);
  AND2 I55 (read_4a0d[16], store_0n[16], readReq_4n);
  AND2 I56 (read_4a0d[17], store_0n[17], readReq_4n);
  AND2 I57 (read_4a0d[18], store_0n[18], readReq_4n);
  AND2 I58 (read_4a0d[19], store_0n[19], readReq_4n);
  AND2 I59 (read_4a0d[20], store_0n[20], readReq_4n);
  AND2 I60 (read_4a0d[21], store_0n[21], readReq_4n);
  AND2 I61 (read_4a0d[22], store_0n[22], readReq_4n);
  AND2 I62 (read_4a0d[23], store_0n[23], readReq_4n);
  AND2 I63 (read_4a0d[24], store_0n[24], readReq_4n);
  AND2 I64 (read_4a0d[25], store_0n[25], readReq_4n);
  AND2 I65 (read_4a0d[26], store_0n[26], readReq_4n);
  AND2 I66 (read_4a0d[27], store_0n[27], readReq_4n);
  AND2 I67 (read_4a0d[28], store_0n[28], readReq_4n);
  AND2 I68 (read_4a0d[29], store_0n[29], readReq_4n);
  AND2 I69 (read_4a0d[30], store_0n[30], readReq_4n);
  AND2 I70 (read_4a0d[31], store_0n[31], readReq_4n);
  AND2 I71 (read_4a0d[32], store_0n[32], readReq_4n);
  AND2 I72 (read_4a0d[33], store_0n[33], readReq_4n);
  AND2 I73 (read_4a0d[34], store_0n[34], readReq_4n);
  AND2 I74 (read_3a1d[0], store_1n[1], readReq_3n);
  AND2 I75 (read_3a1d[1], store_1n[2], readReq_3n);
  AND2 I76 (read_3a1d[2], store_1n[3], readReq_3n);
  AND2 I77 (read_3a1d[3], store_1n[4], readReq_3n);
  AND2 I78 (read_3a1d[4], store_1n[5], readReq_3n);
  AND2 I79 (read_3a1d[5], store_1n[6], readReq_3n);
  AND2 I80 (read_3a1d[6], store_1n[7], readReq_3n);
  AND2 I81 (read_3a1d[7], store_1n[8], readReq_3n);
  AND2 I82 (read_3a1d[8], store_1n[9], readReq_3n);
  AND2 I83 (read_3a1d[9], store_1n[10], readReq_3n);
  AND2 I84 (read_3a1d[10], store_1n[11], readReq_3n);
  AND2 I85 (read_3a1d[11], store_1n[12], readReq_3n);
  AND2 I86 (read_3a1d[12], store_1n[13], readReq_3n);
  AND2 I87 (read_3a1d[13], store_1n[14], readReq_3n);
  AND2 I88 (read_3a1d[14], store_1n[15], readReq_3n);
  AND2 I89 (read_3a1d[15], store_1n[16], readReq_3n);
  AND2 I90 (read_3a1d[16], store_1n[17], readReq_3n);
  AND2 I91 (read_3a1d[17], store_1n[18], readReq_3n);
  AND2 I92 (read_3a1d[18], store_1n[19], readReq_3n);
  AND2 I93 (read_3a1d[19], store_1n[20], readReq_3n);
  AND2 I94 (read_3a1d[20], store_1n[21], readReq_3n);
  AND2 I95 (read_3a1d[21], store_1n[22], readReq_3n);
  AND2 I96 (read_3a1d[22], store_1n[23], readReq_3n);
  AND2 I97 (read_3a1d[23], store_1n[24], readReq_3n);
  AND2 I98 (read_3a1d[24], store_1n[25], readReq_3n);
  AND2 I99 (read_3a1d[25], store_1n[26], readReq_3n);
  AND2 I100 (read_3a1d[26], store_1n[27], readReq_3n);
  AND2 I101 (read_3a1d[27], store_1n[28], readReq_3n);
  AND2 I102 (read_3a1d[28], store_1n[29], readReq_3n);
  AND2 I103 (read_3a1d[29], store_1n[30], readReq_3n);
  AND2 I104 (read_3a1d[30], store_1n[31], readReq_3n);
  AND2 I105 (read_3a1d[31], store_1n[32], readReq_3n);
  AND2 I106 (read_3a0d[0], store_0n[1], readReq_3n);
  AND2 I107 (read_3a0d[1], store_0n[2], readReq_3n);
  AND2 I108 (read_3a0d[2], store_0n[3], readReq_3n);
  AND2 I109 (read_3a0d[3], store_0n[4], readReq_3n);
  AND2 I110 (read_3a0d[4], store_0n[5], readReq_3n);
  AND2 I111 (read_3a0d[5], store_0n[6], readReq_3n);
  AND2 I112 (read_3a0d[6], store_0n[7], readReq_3n);
  AND2 I113 (read_3a0d[7], store_0n[8], readReq_3n);
  AND2 I114 (read_3a0d[8], store_0n[9], readReq_3n);
  AND2 I115 (read_3a0d[9], store_0n[10], readReq_3n);
  AND2 I116 (read_3a0d[10], store_0n[11], readReq_3n);
  AND2 I117 (read_3a0d[11], store_0n[12], readReq_3n);
  AND2 I118 (read_3a0d[12], store_0n[13], readReq_3n);
  AND2 I119 (read_3a0d[13], store_0n[14], readReq_3n);
  AND2 I120 (read_3a0d[14], store_0n[15], readReq_3n);
  AND2 I121 (read_3a0d[15], store_0n[16], readReq_3n);
  AND2 I122 (read_3a0d[16], store_0n[17], readReq_3n);
  AND2 I123 (read_3a0d[17], store_0n[18], readReq_3n);
  AND2 I124 (read_3a0d[18], store_0n[19], readReq_3n);
  AND2 I125 (read_3a0d[19], store_0n[20], readReq_3n);
  AND2 I126 (read_3a0d[20], store_0n[21], readReq_3n);
  AND2 I127 (read_3a0d[21], store_0n[22], readReq_3n);
  AND2 I128 (read_3a0d[22], store_0n[23], readReq_3n);
  AND2 I129 (read_3a0d[23], store_0n[24], readReq_3n);
  AND2 I130 (read_3a0d[24], store_0n[25], readReq_3n);
  AND2 I131 (read_3a0d[25], store_0n[26], readReq_3n);
  AND2 I132 (read_3a0d[26], store_0n[27], readReq_3n);
  AND2 I133 (read_3a0d[27], store_0n[28], readReq_3n);
  AND2 I134 (read_3a0d[28], store_0n[29], readReq_3n);
  AND2 I135 (read_3a0d[29], store_0n[30], readReq_3n);
  AND2 I136 (read_3a0d[30], store_0n[31], readReq_3n);
  AND2 I137 (read_3a0d[31], store_0n[32], readReq_3n);
  AND2 I138 (read_2a1d[0], store_1n[0], readReq_2n);
  AND2 I139 (read_2a1d[1], store_1n[1], readReq_2n);
  AND2 I140 (read_2a1d[2], store_1n[2], readReq_2n);
  AND2 I141 (read_2a1d[3], store_1n[3], readReq_2n);
  AND2 I142 (read_2a1d[4], store_1n[4], readReq_2n);
  AND2 I143 (read_2a1d[5], store_1n[5], readReq_2n);
  AND2 I144 (read_2a1d[6], store_1n[6], readReq_2n);
  AND2 I145 (read_2a1d[7], store_1n[7], readReq_2n);
  AND2 I146 (read_2a1d[8], store_1n[8], readReq_2n);
  AND2 I147 (read_2a1d[9], store_1n[9], readReq_2n);
  AND2 I148 (read_2a1d[10], store_1n[10], readReq_2n);
  AND2 I149 (read_2a1d[11], store_1n[11], readReq_2n);
  AND2 I150 (read_2a1d[12], store_1n[12], readReq_2n);
  AND2 I151 (read_2a1d[13], store_1n[13], readReq_2n);
  AND2 I152 (read_2a1d[14], store_1n[14], readReq_2n);
  AND2 I153 (read_2a1d[15], store_1n[15], readReq_2n);
  AND2 I154 (read_2a1d[16], store_1n[16], readReq_2n);
  AND2 I155 (read_2a1d[17], store_1n[17], readReq_2n);
  AND2 I156 (read_2a1d[18], store_1n[18], readReq_2n);
  AND2 I157 (read_2a1d[19], store_1n[19], readReq_2n);
  AND2 I158 (read_2a1d[20], store_1n[20], readReq_2n);
  AND2 I159 (read_2a1d[21], store_1n[21], readReq_2n);
  AND2 I160 (read_2a1d[22], store_1n[22], readReq_2n);
  AND2 I161 (read_2a1d[23], store_1n[23], readReq_2n);
  AND2 I162 (read_2a1d[24], store_1n[24], readReq_2n);
  AND2 I163 (read_2a1d[25], store_1n[25], readReq_2n);
  AND2 I164 (read_2a1d[26], store_1n[26], readReq_2n);
  AND2 I165 (read_2a1d[27], store_1n[27], readReq_2n);
  AND2 I166 (read_2a1d[28], store_1n[28], readReq_2n);
  AND2 I167 (read_2a1d[29], store_1n[29], readReq_2n);
  AND2 I168 (read_2a1d[30], store_1n[30], readReq_2n);
  AND2 I169 (read_2a1d[31], store_1n[31], readReq_2n);
  AND2 I170 (read_2a1d[32], store_1n[32], readReq_2n);
  AND2 I171 (read_2a0d[0], store_0n[0], readReq_2n);
  AND2 I172 (read_2a0d[1], store_0n[1], readReq_2n);
  AND2 I173 (read_2a0d[2], store_0n[2], readReq_2n);
  AND2 I174 (read_2a0d[3], store_0n[3], readReq_2n);
  AND2 I175 (read_2a0d[4], store_0n[4], readReq_2n);
  AND2 I176 (read_2a0d[5], store_0n[5], readReq_2n);
  AND2 I177 (read_2a0d[6], store_0n[6], readReq_2n);
  AND2 I178 (read_2a0d[7], store_0n[7], readReq_2n);
  AND2 I179 (read_2a0d[8], store_0n[8], readReq_2n);
  AND2 I180 (read_2a0d[9], store_0n[9], readReq_2n);
  AND2 I181 (read_2a0d[10], store_0n[10], readReq_2n);
  AND2 I182 (read_2a0d[11], store_0n[11], readReq_2n);
  AND2 I183 (read_2a0d[12], store_0n[12], readReq_2n);
  AND2 I184 (read_2a0d[13], store_0n[13], readReq_2n);
  AND2 I185 (read_2a0d[14], store_0n[14], readReq_2n);
  AND2 I186 (read_2a0d[15], store_0n[15], readReq_2n);
  AND2 I187 (read_2a0d[16], store_0n[16], readReq_2n);
  AND2 I188 (read_2a0d[17], store_0n[17], readReq_2n);
  AND2 I189 (read_2a0d[18], store_0n[18], readReq_2n);
  AND2 I190 (read_2a0d[19], store_0n[19], readReq_2n);
  AND2 I191 (read_2a0d[20], store_0n[20], readReq_2n);
  AND2 I192 (read_2a0d[21], store_0n[21], readReq_2n);
  AND2 I193 (read_2a0d[22], store_0n[22], readReq_2n);
  AND2 I194 (read_2a0d[23], store_0n[23], readReq_2n);
  AND2 I195 (read_2a0d[24], store_0n[24], readReq_2n);
  AND2 I196 (read_2a0d[25], store_0n[25], readReq_2n);
  AND2 I197 (read_2a0d[26], store_0n[26], readReq_2n);
  AND2 I198 (read_2a0d[27], store_0n[27], readReq_2n);
  AND2 I199 (read_2a0d[28], store_0n[28], readReq_2n);
  AND2 I200 (read_2a0d[29], store_0n[29], readReq_2n);
  AND2 I201 (read_2a0d[30], store_0n[30], readReq_2n);
  AND2 I202 (read_2a0d[31], store_0n[31], readReq_2n);
  AND2 I203 (read_2a0d[32], store_0n[32], readReq_2n);
  AND2 I204 (read_1a1d[0], store_1n[0], readReq_1n);
  AND2 I205 (read_1a1d[1], store_1n[1], readReq_1n);
  AND2 I206 (read_1a1d[2], store_1n[2], readReq_1n);
  AND2 I207 (read_1a1d[3], store_1n[3], readReq_1n);
  AND2 I208 (read_1a1d[4], store_1n[4], readReq_1n);
  AND2 I209 (read_1a1d[5], store_1n[5], readReq_1n);
  AND2 I210 (read_1a1d[6], store_1n[6], readReq_1n);
  AND2 I211 (read_1a1d[7], store_1n[7], readReq_1n);
  AND2 I212 (read_1a1d[8], store_1n[8], readReq_1n);
  AND2 I213 (read_1a1d[9], store_1n[9], readReq_1n);
  AND2 I214 (read_1a1d[10], store_1n[10], readReq_1n);
  AND2 I215 (read_1a1d[11], store_1n[11], readReq_1n);
  AND2 I216 (read_1a1d[12], store_1n[12], readReq_1n);
  AND2 I217 (read_1a1d[13], store_1n[13], readReq_1n);
  AND2 I218 (read_1a1d[14], store_1n[14], readReq_1n);
  AND2 I219 (read_1a1d[15], store_1n[15], readReq_1n);
  AND2 I220 (read_1a1d[16], store_1n[16], readReq_1n);
  AND2 I221 (read_1a1d[17], store_1n[17], readReq_1n);
  AND2 I222 (read_1a1d[18], store_1n[18], readReq_1n);
  AND2 I223 (read_1a1d[19], store_1n[19], readReq_1n);
  AND2 I224 (read_1a1d[20], store_1n[20], readReq_1n);
  AND2 I225 (read_1a1d[21], store_1n[21], readReq_1n);
  AND2 I226 (read_1a1d[22], store_1n[22], readReq_1n);
  AND2 I227 (read_1a1d[23], store_1n[23], readReq_1n);
  AND2 I228 (read_1a1d[24], store_1n[24], readReq_1n);
  AND2 I229 (read_1a1d[25], store_1n[25], readReq_1n);
  AND2 I230 (read_1a1d[26], store_1n[26], readReq_1n);
  AND2 I231 (read_1a1d[27], store_1n[27], readReq_1n);
  AND2 I232 (read_1a1d[28], store_1n[28], readReq_1n);
  AND2 I233 (read_1a1d[29], store_1n[29], readReq_1n);
  AND2 I234 (read_1a1d[30], store_1n[30], readReq_1n);
  AND2 I235 (read_1a1d[31], store_1n[31], readReq_1n);
  AND2 I236 (read_1a1d[32], store_1n[32], readReq_1n);
  AND2 I237 (read_1a1d[33], store_1n[33], readReq_1n);
  AND2 I238 (read_1a0d[0], store_0n[0], readReq_1n);
  AND2 I239 (read_1a0d[1], store_0n[1], readReq_1n);
  AND2 I240 (read_1a0d[2], store_0n[2], readReq_1n);
  AND2 I241 (read_1a0d[3], store_0n[3], readReq_1n);
  AND2 I242 (read_1a0d[4], store_0n[4], readReq_1n);
  AND2 I243 (read_1a0d[5], store_0n[5], readReq_1n);
  AND2 I244 (read_1a0d[6], store_0n[6], readReq_1n);
  AND2 I245 (read_1a0d[7], store_0n[7], readReq_1n);
  AND2 I246 (read_1a0d[8], store_0n[8], readReq_1n);
  AND2 I247 (read_1a0d[9], store_0n[9], readReq_1n);
  AND2 I248 (read_1a0d[10], store_0n[10], readReq_1n);
  AND2 I249 (read_1a0d[11], store_0n[11], readReq_1n);
  AND2 I250 (read_1a0d[12], store_0n[12], readReq_1n);
  AND2 I251 (read_1a0d[13], store_0n[13], readReq_1n);
  AND2 I252 (read_1a0d[14], store_0n[14], readReq_1n);
  AND2 I253 (read_1a0d[15], store_0n[15], readReq_1n);
  AND2 I254 (read_1a0d[16], store_0n[16], readReq_1n);
  AND2 I255 (read_1a0d[17], store_0n[17], readReq_1n);
  AND2 I256 (read_1a0d[18], store_0n[18], readReq_1n);
  AND2 I257 (read_1a0d[19], store_0n[19], readReq_1n);
  AND2 I258 (read_1a0d[20], store_0n[20], readReq_1n);
  AND2 I259 (read_1a0d[21], store_0n[21], readReq_1n);
  AND2 I260 (read_1a0d[22], store_0n[22], readReq_1n);
  AND2 I261 (read_1a0d[23], store_0n[23], readReq_1n);
  AND2 I262 (read_1a0d[24], store_0n[24], readReq_1n);
  AND2 I263 (read_1a0d[25], store_0n[25], readReq_1n);
  AND2 I264 (read_1a0d[26], store_0n[26], readReq_1n);
  AND2 I265 (read_1a0d[27], store_0n[27], readReq_1n);
  AND2 I266 (read_1a0d[28], store_0n[28], readReq_1n);
  AND2 I267 (read_1a0d[29], store_0n[29], readReq_1n);
  AND2 I268 (read_1a0d[30], store_0n[30], readReq_1n);
  AND2 I269 (read_1a0d[31], store_0n[31], readReq_1n);
  AND2 I270 (read_1a0d[32], store_0n[32], readReq_1n);
  AND2 I271 (read_1a0d[33], store_0n[33], readReq_1n);
  AND2 I272 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I273 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I274 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I275 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I276 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I277 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I278 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I279 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I280 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I281 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I282 (read_0a1d[10], store_1n[10], readReq_0n);
  AND2 I283 (read_0a1d[11], store_1n[11], readReq_0n);
  AND2 I284 (read_0a1d[12], store_1n[12], readReq_0n);
  AND2 I285 (read_0a1d[13], store_1n[13], readReq_0n);
  AND2 I286 (read_0a1d[14], store_1n[14], readReq_0n);
  AND2 I287 (read_0a1d[15], store_1n[15], readReq_0n);
  AND2 I288 (read_0a1d[16], store_1n[16], readReq_0n);
  AND2 I289 (read_0a1d[17], store_1n[17], readReq_0n);
  AND2 I290 (read_0a1d[18], store_1n[18], readReq_0n);
  AND2 I291 (read_0a1d[19], store_1n[19], readReq_0n);
  AND2 I292 (read_0a1d[20], store_1n[20], readReq_0n);
  AND2 I293 (read_0a1d[21], store_1n[21], readReq_0n);
  AND2 I294 (read_0a1d[22], store_1n[22], readReq_0n);
  AND2 I295 (read_0a1d[23], store_1n[23], readReq_0n);
  AND2 I296 (read_0a1d[24], store_1n[24], readReq_0n);
  AND2 I297 (read_0a1d[25], store_1n[25], readReq_0n);
  AND2 I298 (read_0a1d[26], store_1n[26], readReq_0n);
  AND2 I299 (read_0a1d[27], store_1n[27], readReq_0n);
  AND2 I300 (read_0a1d[28], store_1n[28], readReq_0n);
  AND2 I301 (read_0a1d[29], store_1n[29], readReq_0n);
  AND2 I302 (read_0a1d[30], store_1n[30], readReq_0n);
  AND2 I303 (read_0a1d[31], store_1n[31], readReq_0n);
  AND2 I304 (read_0a1d[32], store_1n[32], readReq_0n);
  AND2 I305 (read_0a1d[33], store_1n[33], readReq_0n);
  AND2 I306 (read_0a1d[34], store_1n[34], readReq_0n);
  AND2 I307 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I308 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I309 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I310 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I311 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I312 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I313 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I314 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I315 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I316 (read_0a0d[9], store_0n[9], readReq_0n);
  AND2 I317 (read_0a0d[10], store_0n[10], readReq_0n);
  AND2 I318 (read_0a0d[11], store_0n[11], readReq_0n);
  AND2 I319 (read_0a0d[12], store_0n[12], readReq_0n);
  AND2 I320 (read_0a0d[13], store_0n[13], readReq_0n);
  AND2 I321 (read_0a0d[14], store_0n[14], readReq_0n);
  AND2 I322 (read_0a0d[15], store_0n[15], readReq_0n);
  AND2 I323 (read_0a0d[16], store_0n[16], readReq_0n);
  AND2 I324 (read_0a0d[17], store_0n[17], readReq_0n);
  AND2 I325 (read_0a0d[18], store_0n[18], readReq_0n);
  AND2 I326 (read_0a0d[19], store_0n[19], readReq_0n);
  AND2 I327 (read_0a0d[20], store_0n[20], readReq_0n);
  AND2 I328 (read_0a0d[21], store_0n[21], readReq_0n);
  AND2 I329 (read_0a0d[22], store_0n[22], readReq_0n);
  AND2 I330 (read_0a0d[23], store_0n[23], readReq_0n);
  AND2 I331 (read_0a0d[24], store_0n[24], readReq_0n);
  AND2 I332 (read_0a0d[25], store_0n[25], readReq_0n);
  AND2 I333 (read_0a0d[26], store_0n[26], readReq_0n);
  AND2 I334 (read_0a0d[27], store_0n[27], readReq_0n);
  AND2 I335 (read_0a0d[28], store_0n[28], readReq_0n);
  AND2 I336 (read_0a0d[29], store_0n[29], readReq_0n);
  AND2 I337 (read_0a0d[30], store_0n[30], readReq_0n);
  AND2 I338 (read_0a0d[31], store_0n[31], readReq_0n);
  AND2 I339 (read_0a0d[32], store_0n[32], readReq_0n);
  AND2 I340 (read_0a0d[33], store_0n[33], readReq_0n);
  AND2 I341 (read_0a0d[34], store_0n[34], readReq_0n);
  BUFF I342 (readReq_0n, read_0r);
  BUFF I343 (readReq_1n, read_1r);
  BUFF I344 (readReq_2n, read_2r);
  BUFF I345 (readReq_3n, read_3r);
  BUFF I346 (readReq_4n, read_4r);
  BUFF I347 (readReq_5n, read_5r);
  BUFF I348 (readReq_6n, read_6r);
  BUFF I349 (store_1n[0], write_0a1d[0]);
  BUFF I350 (store_1n[1], write_0a1d[1]);
  BUFF I351 (store_1n[2], write_0a1d[2]);
  BUFF I352 (store_1n[3], write_0a1d[3]);
  BUFF I353 (store_1n[4], write_0a1d[4]);
  BUFF I354 (store_1n[5], write_0a1d[5]);
  BUFF I355 (store_1n[6], write_0a1d[6]);
  BUFF I356 (store_1n[7], write_0a1d[7]);
  BUFF I357 (store_1n[8], write_0a1d[8]);
  BUFF I358 (store_1n[9], write_0a1d[9]);
  BUFF I359 (store_1n[10], write_0a1d[10]);
  BUFF I360 (store_1n[11], write_0a1d[11]);
  BUFF I361 (store_1n[12], write_0a1d[12]);
  BUFF I362 (store_1n[13], write_0a1d[13]);
  BUFF I363 (store_1n[14], write_0a1d[14]);
  BUFF I364 (store_1n[15], write_0a1d[15]);
  BUFF I365 (store_1n[16], write_0a1d[16]);
  BUFF I366 (store_1n[17], write_0a1d[17]);
  BUFF I367 (store_1n[18], write_0a1d[18]);
  BUFF I368 (store_1n[19], write_0a1d[19]);
  BUFF I369 (store_1n[20], write_0a1d[20]);
  BUFF I370 (store_1n[21], write_0a1d[21]);
  BUFF I371 (store_1n[22], write_0a1d[22]);
  BUFF I372 (store_1n[23], write_0a1d[23]);
  BUFF I373 (store_1n[24], write_0a1d[24]);
  BUFF I374 (store_1n[25], write_0a1d[25]);
  BUFF I375 (store_1n[26], write_0a1d[26]);
  BUFF I376 (store_1n[27], write_0a1d[27]);
  BUFF I377 (store_1n[28], write_0a1d[28]);
  BUFF I378 (store_1n[29], write_0a1d[29]);
  BUFF I379 (store_1n[30], write_0a1d[30]);
  BUFF I380 (store_1n[31], write_0a1d[31]);
  BUFF I381 (store_1n[32], write_0a1d[32]);
  BUFF I382 (store_1n[33], write_0a1d[33]);
  BUFF I383 (store_1n[34], write_0a1d[34]);
  BUFF I384 (store_0n[0], write_0a0d[0]);
  BUFF I385 (store_0n[1], write_0a0d[1]);
  BUFF I386 (store_0n[2], write_0a0d[2]);
  BUFF I387 (store_0n[3], write_0a0d[3]);
  BUFF I388 (store_0n[4], write_0a0d[4]);
  BUFF I389 (store_0n[5], write_0a0d[5]);
  BUFF I390 (store_0n[6], write_0a0d[6]);
  BUFF I391 (store_0n[7], write_0a0d[7]);
  BUFF I392 (store_0n[8], write_0a0d[8]);
  BUFF I393 (store_0n[9], write_0a0d[9]);
  BUFF I394 (store_0n[10], write_0a0d[10]);
  BUFF I395 (store_0n[11], write_0a0d[11]);
  BUFF I396 (store_0n[12], write_0a0d[12]);
  BUFF I397 (store_0n[13], write_0a0d[13]);
  BUFF I398 (store_0n[14], write_0a0d[14]);
  BUFF I399 (store_0n[15], write_0a0d[15]);
  BUFF I400 (store_0n[16], write_0a0d[16]);
  BUFF I401 (store_0n[17], write_0a0d[17]);
  BUFF I402 (store_0n[18], write_0a0d[18]);
  BUFF I403 (store_0n[19], write_0a0d[19]);
  BUFF I404 (store_0n[20], write_0a0d[20]);
  BUFF I405 (store_0n[21], write_0a0d[21]);
  BUFF I406 (store_0n[22], write_0a0d[22]);
  BUFF I407 (store_0n[23], write_0a0d[23]);
  BUFF I408 (store_0n[24], write_0a0d[24]);
  BUFF I409 (store_0n[25], write_0a0d[25]);
  BUFF I410 (store_0n[26], write_0a0d[26]);
  BUFF I411 (store_0n[27], write_0a0d[27]);
  BUFF I412 (store_0n[28], write_0a0d[28]);
  BUFF I413 (store_0n[29], write_0a0d[29]);
  BUFF I414 (store_0n[30], write_0a0d[30]);
  BUFF I415 (store_0n[31], write_0a0d[31]);
  BUFF I416 (store_0n[32], write_0a0d[32]);
  BUFF I417 (store_0n[33], write_0a0d[33]);
  BUFF I418 (store_0n[34], write_0a0d[34]);
  C2 I419 (trigger_0a, writeAck_0n, cd_0n);
  AND2 I420 (writeAck_0n, sigAck_0n, rReqOr_0n);
  NOR3 I421 (internal_0n[0], readReq_0n, readReq_1n, readReq_2n);
  NOR2 I422 (internal_0n[1], readReq_3n, readReq_4n);
  NOR2 I423 (internal_0n[2], readReq_5n, readReq_6n);
  AND3 I424 (rReqOr_0n, internal_0n[0], internal_0n[1], internal_0n[2]);
  BALSA_TELEM I425 (trigger_0r, sigAck_0n, signal_0r, signal_0a);
  C3 I426 (internal_0n[3], partCD_0n[0], partCD_0n[1], partCD_0n[2]);
  C3 I427 (internal_0n[4], partCD_0n[3], partCD_0n[4], partCD_0n[5]);
  C3 I428 (internal_0n[5], partCD_0n[6], partCD_0n[7], partCD_0n[8]);
  C3 I429 (internal_0n[6], partCD_0n[9], partCD_0n[10], partCD_0n[11]);
  C3 I430 (internal_0n[7], partCD_0n[12], partCD_0n[13], partCD_0n[14]);
  C3 I431 (internal_0n[8], partCD_0n[15], partCD_0n[16], partCD_0n[17]);
  C3 I432 (internal_0n[9], partCD_0n[18], partCD_0n[19], partCD_0n[20]);
  C3 I433 (internal_0n[10], partCD_0n[21], partCD_0n[22], partCD_0n[23]);
  C3 I434 (internal_0n[11], partCD_0n[24], partCD_0n[25], partCD_0n[26]);
  C3 I435 (internal_0n[12], partCD_0n[27], partCD_0n[28], partCD_0n[29]);
  C3 I436 (internal_0n[13], partCD_0n[30], partCD_0n[31], partCD_0n[32]);
  C2 I437 (internal_0n[14], partCD_0n[33], partCD_0n[34]);
  C3 I438 (internal_0n[15], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I439 (internal_0n[16], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I440 (internal_0n[17], internal_0n[9], internal_0n[10], internal_0n[11]);
  C3 I441 (internal_0n[18], internal_0n[12], internal_0n[13], internal_0n[14]);
  C2 I442 (internal_0n[19], internal_0n[15], internal_0n[16]);
  C2 I443 (internal_0n[20], internal_0n[17], internal_0n[18]);
  C2 I444 (cd_0n, internal_0n[19], internal_0n[20]);
  OR2 I445 (partCD_0n[0], store_0n[0], store_1n[0]);
  OR2 I446 (partCD_0n[1], store_0n[1], store_1n[1]);
  OR2 I447 (partCD_0n[2], store_0n[2], store_1n[2]);
  OR2 I448 (partCD_0n[3], store_0n[3], store_1n[3]);
  OR2 I449 (partCD_0n[4], store_0n[4], store_1n[4]);
  OR2 I450 (partCD_0n[5], store_0n[5], store_1n[5]);
  OR2 I451 (partCD_0n[6], store_0n[6], store_1n[6]);
  OR2 I452 (partCD_0n[7], store_0n[7], store_1n[7]);
  OR2 I453 (partCD_0n[8], store_0n[8], store_1n[8]);
  OR2 I454 (partCD_0n[9], store_0n[9], store_1n[9]);
  OR2 I455 (partCD_0n[10], store_0n[10], store_1n[10]);
  OR2 I456 (partCD_0n[11], store_0n[11], store_1n[11]);
  OR2 I457 (partCD_0n[12], store_0n[12], store_1n[12]);
  OR2 I458 (partCD_0n[13], store_0n[13], store_1n[13]);
  OR2 I459 (partCD_0n[14], store_0n[14], store_1n[14]);
  OR2 I460 (partCD_0n[15], store_0n[15], store_1n[15]);
  OR2 I461 (partCD_0n[16], store_0n[16], store_1n[16]);
  OR2 I462 (partCD_0n[17], store_0n[17], store_1n[17]);
  OR2 I463 (partCD_0n[18], store_0n[18], store_1n[18]);
  OR2 I464 (partCD_0n[19], store_0n[19], store_1n[19]);
  OR2 I465 (partCD_0n[20], store_0n[20], store_1n[20]);
  OR2 I466 (partCD_0n[21], store_0n[21], store_1n[21]);
  OR2 I467 (partCD_0n[22], store_0n[22], store_1n[22]);
  OR2 I468 (partCD_0n[23], store_0n[23], store_1n[23]);
  OR2 I469 (partCD_0n[24], store_0n[24], store_1n[24]);
  OR2 I470 (partCD_0n[25], store_0n[25], store_1n[25]);
  OR2 I471 (partCD_0n[26], store_0n[26], store_1n[26]);
  OR2 I472 (partCD_0n[27], store_0n[27], store_1n[27]);
  OR2 I473 (partCD_0n[28], store_0n[28], store_1n[28]);
  OR2 I474 (partCD_0n[29], store_0n[29], store_1n[29]);
  OR2 I475 (partCD_0n[30], store_0n[30], store_1n[30]);
  OR2 I476 (partCD_0n[31], store_0n[31], store_1n[31]);
  OR2 I477 (partCD_0n[32], store_0n[32], store_1n[32]);
  OR2 I478 (partCD_0n[33], store_0n[33], store_1n[33]);
  OR2 I479 (partCD_0n[34], store_0n[34], store_1n[34]);
  BUFF I480 (write_0r, trigger_0r);
endmodule

module BrzActiveEagerFalseVariable_36_2_s11__3b0__m13m (
  trigger_0r, trigger_0a,
  write_0r, write_0a0d, write_0a1d,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d
);
  input trigger_0r;
  output trigger_0a;
  output write_0r;
  input [35:0] write_0a0d;
  input [35:0] write_0a1d;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output [35:0] read_0a0d;
  output [35:0] read_0a1d;
  input read_1r;
  output [3:0] read_1a0d;
  output [3:0] read_1a1d;
  wire [17:0] internal_0n;
  wire cd_0n;
  wire [35:0] partCD_0n;
  wire [35:0] store_0n;
  wire [35:0] store_1n;
  wire readReq_0n;
  wire readReq_1n;
  wire writeAck_0n;
  wire sigAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_1a1d[0], store_1n[0], readReq_1n);
  AND2 I1 (read_1a1d[1], store_1n[1], readReq_1n);
  AND2 I2 (read_1a1d[2], store_1n[2], readReq_1n);
  AND2 I3 (read_1a1d[3], store_1n[3], readReq_1n);
  AND2 I4 (read_1a0d[0], store_0n[0], readReq_1n);
  AND2 I5 (read_1a0d[1], store_0n[1], readReq_1n);
  AND2 I6 (read_1a0d[2], store_0n[2], readReq_1n);
  AND2 I7 (read_1a0d[3], store_0n[3], readReq_1n);
  AND2 I8 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I9 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I10 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I11 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I12 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I13 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I14 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I15 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I16 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I17 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I18 (read_0a1d[10], store_1n[10], readReq_0n);
  AND2 I19 (read_0a1d[11], store_1n[11], readReq_0n);
  AND2 I20 (read_0a1d[12], store_1n[12], readReq_0n);
  AND2 I21 (read_0a1d[13], store_1n[13], readReq_0n);
  AND2 I22 (read_0a1d[14], store_1n[14], readReq_0n);
  AND2 I23 (read_0a1d[15], store_1n[15], readReq_0n);
  AND2 I24 (read_0a1d[16], store_1n[16], readReq_0n);
  AND2 I25 (read_0a1d[17], store_1n[17], readReq_0n);
  AND2 I26 (read_0a1d[18], store_1n[18], readReq_0n);
  AND2 I27 (read_0a1d[19], store_1n[19], readReq_0n);
  AND2 I28 (read_0a1d[20], store_1n[20], readReq_0n);
  AND2 I29 (read_0a1d[21], store_1n[21], readReq_0n);
  AND2 I30 (read_0a1d[22], store_1n[22], readReq_0n);
  AND2 I31 (read_0a1d[23], store_1n[23], readReq_0n);
  AND2 I32 (read_0a1d[24], store_1n[24], readReq_0n);
  AND2 I33 (read_0a1d[25], store_1n[25], readReq_0n);
  AND2 I34 (read_0a1d[26], store_1n[26], readReq_0n);
  AND2 I35 (read_0a1d[27], store_1n[27], readReq_0n);
  AND2 I36 (read_0a1d[28], store_1n[28], readReq_0n);
  AND2 I37 (read_0a1d[29], store_1n[29], readReq_0n);
  AND2 I38 (read_0a1d[30], store_1n[30], readReq_0n);
  AND2 I39 (read_0a1d[31], store_1n[31], readReq_0n);
  AND2 I40 (read_0a1d[32], store_1n[32], readReq_0n);
  AND2 I41 (read_0a1d[33], store_1n[33], readReq_0n);
  AND2 I42 (read_0a1d[34], store_1n[34], readReq_0n);
  AND2 I43 (read_0a1d[35], store_1n[35], readReq_0n);
  AND2 I44 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I45 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I46 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I47 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I48 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I49 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I50 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I51 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I52 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I53 (read_0a0d[9], store_0n[9], readReq_0n);
  AND2 I54 (read_0a0d[10], store_0n[10], readReq_0n);
  AND2 I55 (read_0a0d[11], store_0n[11], readReq_0n);
  AND2 I56 (read_0a0d[12], store_0n[12], readReq_0n);
  AND2 I57 (read_0a0d[13], store_0n[13], readReq_0n);
  AND2 I58 (read_0a0d[14], store_0n[14], readReq_0n);
  AND2 I59 (read_0a0d[15], store_0n[15], readReq_0n);
  AND2 I60 (read_0a0d[16], store_0n[16], readReq_0n);
  AND2 I61 (read_0a0d[17], store_0n[17], readReq_0n);
  AND2 I62 (read_0a0d[18], store_0n[18], readReq_0n);
  AND2 I63 (read_0a0d[19], store_0n[19], readReq_0n);
  AND2 I64 (read_0a0d[20], store_0n[20], readReq_0n);
  AND2 I65 (read_0a0d[21], store_0n[21], readReq_0n);
  AND2 I66 (read_0a0d[22], store_0n[22], readReq_0n);
  AND2 I67 (read_0a0d[23], store_0n[23], readReq_0n);
  AND2 I68 (read_0a0d[24], store_0n[24], readReq_0n);
  AND2 I69 (read_0a0d[25], store_0n[25], readReq_0n);
  AND2 I70 (read_0a0d[26], store_0n[26], readReq_0n);
  AND2 I71 (read_0a0d[27], store_0n[27], readReq_0n);
  AND2 I72 (read_0a0d[28], store_0n[28], readReq_0n);
  AND2 I73 (read_0a0d[29], store_0n[29], readReq_0n);
  AND2 I74 (read_0a0d[30], store_0n[30], readReq_0n);
  AND2 I75 (read_0a0d[31], store_0n[31], readReq_0n);
  AND2 I76 (read_0a0d[32], store_0n[32], readReq_0n);
  AND2 I77 (read_0a0d[33], store_0n[33], readReq_0n);
  AND2 I78 (read_0a0d[34], store_0n[34], readReq_0n);
  AND2 I79 (read_0a0d[35], store_0n[35], readReq_0n);
  BUFF I80 (readReq_0n, read_0r);
  BUFF I81 (readReq_1n, read_1r);
  BUFF I82 (store_1n[0], write_0a1d[0]);
  BUFF I83 (store_1n[1], write_0a1d[1]);
  BUFF I84 (store_1n[2], write_0a1d[2]);
  BUFF I85 (store_1n[3], write_0a1d[3]);
  BUFF I86 (store_1n[4], write_0a1d[4]);
  BUFF I87 (store_1n[5], write_0a1d[5]);
  BUFF I88 (store_1n[6], write_0a1d[6]);
  BUFF I89 (store_1n[7], write_0a1d[7]);
  BUFF I90 (store_1n[8], write_0a1d[8]);
  BUFF I91 (store_1n[9], write_0a1d[9]);
  BUFF I92 (store_1n[10], write_0a1d[10]);
  BUFF I93 (store_1n[11], write_0a1d[11]);
  BUFF I94 (store_1n[12], write_0a1d[12]);
  BUFF I95 (store_1n[13], write_0a1d[13]);
  BUFF I96 (store_1n[14], write_0a1d[14]);
  BUFF I97 (store_1n[15], write_0a1d[15]);
  BUFF I98 (store_1n[16], write_0a1d[16]);
  BUFF I99 (store_1n[17], write_0a1d[17]);
  BUFF I100 (store_1n[18], write_0a1d[18]);
  BUFF I101 (store_1n[19], write_0a1d[19]);
  BUFF I102 (store_1n[20], write_0a1d[20]);
  BUFF I103 (store_1n[21], write_0a1d[21]);
  BUFF I104 (store_1n[22], write_0a1d[22]);
  BUFF I105 (store_1n[23], write_0a1d[23]);
  BUFF I106 (store_1n[24], write_0a1d[24]);
  BUFF I107 (store_1n[25], write_0a1d[25]);
  BUFF I108 (store_1n[26], write_0a1d[26]);
  BUFF I109 (store_1n[27], write_0a1d[27]);
  BUFF I110 (store_1n[28], write_0a1d[28]);
  BUFF I111 (store_1n[29], write_0a1d[29]);
  BUFF I112 (store_1n[30], write_0a1d[30]);
  BUFF I113 (store_1n[31], write_0a1d[31]);
  BUFF I114 (store_1n[32], write_0a1d[32]);
  BUFF I115 (store_1n[33], write_0a1d[33]);
  BUFF I116 (store_1n[34], write_0a1d[34]);
  BUFF I117 (store_1n[35], write_0a1d[35]);
  BUFF I118 (store_0n[0], write_0a0d[0]);
  BUFF I119 (store_0n[1], write_0a0d[1]);
  BUFF I120 (store_0n[2], write_0a0d[2]);
  BUFF I121 (store_0n[3], write_0a0d[3]);
  BUFF I122 (store_0n[4], write_0a0d[4]);
  BUFF I123 (store_0n[5], write_0a0d[5]);
  BUFF I124 (store_0n[6], write_0a0d[6]);
  BUFF I125 (store_0n[7], write_0a0d[7]);
  BUFF I126 (store_0n[8], write_0a0d[8]);
  BUFF I127 (store_0n[9], write_0a0d[9]);
  BUFF I128 (store_0n[10], write_0a0d[10]);
  BUFF I129 (store_0n[11], write_0a0d[11]);
  BUFF I130 (store_0n[12], write_0a0d[12]);
  BUFF I131 (store_0n[13], write_0a0d[13]);
  BUFF I132 (store_0n[14], write_0a0d[14]);
  BUFF I133 (store_0n[15], write_0a0d[15]);
  BUFF I134 (store_0n[16], write_0a0d[16]);
  BUFF I135 (store_0n[17], write_0a0d[17]);
  BUFF I136 (store_0n[18], write_0a0d[18]);
  BUFF I137 (store_0n[19], write_0a0d[19]);
  BUFF I138 (store_0n[20], write_0a0d[20]);
  BUFF I139 (store_0n[21], write_0a0d[21]);
  BUFF I140 (store_0n[22], write_0a0d[22]);
  BUFF I141 (store_0n[23], write_0a0d[23]);
  BUFF I142 (store_0n[24], write_0a0d[24]);
  BUFF I143 (store_0n[25], write_0a0d[25]);
  BUFF I144 (store_0n[26], write_0a0d[26]);
  BUFF I145 (store_0n[27], write_0a0d[27]);
  BUFF I146 (store_0n[28], write_0a0d[28]);
  BUFF I147 (store_0n[29], write_0a0d[29]);
  BUFF I148 (store_0n[30], write_0a0d[30]);
  BUFF I149 (store_0n[31], write_0a0d[31]);
  BUFF I150 (store_0n[32], write_0a0d[32]);
  BUFF I151 (store_0n[33], write_0a0d[33]);
  BUFF I152 (store_0n[34], write_0a0d[34]);
  BUFF I153 (store_0n[35], write_0a0d[35]);
  C2 I154 (trigger_0a, writeAck_0n, cd_0n);
  AND2 I155 (writeAck_0n, sigAck_0n, rReqOr_0n);
  NOR2 I156 (rReqOr_0n, readReq_0n, readReq_1n);
  BALSA_TELEM I157 (trigger_0r, sigAck_0n, signal_0r, signal_0a);
  C3 I158 (internal_0n[0], partCD_0n[0], partCD_0n[1], partCD_0n[2]);
  C3 I159 (internal_0n[1], partCD_0n[3], partCD_0n[4], partCD_0n[5]);
  C3 I160 (internal_0n[2], partCD_0n[6], partCD_0n[7], partCD_0n[8]);
  C3 I161 (internal_0n[3], partCD_0n[9], partCD_0n[10], partCD_0n[11]);
  C3 I162 (internal_0n[4], partCD_0n[12], partCD_0n[13], partCD_0n[14]);
  C3 I163 (internal_0n[5], partCD_0n[15], partCD_0n[16], partCD_0n[17]);
  C3 I164 (internal_0n[6], partCD_0n[18], partCD_0n[19], partCD_0n[20]);
  C3 I165 (internal_0n[7], partCD_0n[21], partCD_0n[22], partCD_0n[23]);
  C3 I166 (internal_0n[8], partCD_0n[24], partCD_0n[25], partCD_0n[26]);
  C3 I167 (internal_0n[9], partCD_0n[27], partCD_0n[28], partCD_0n[29]);
  C3 I168 (internal_0n[10], partCD_0n[30], partCD_0n[31], partCD_0n[32]);
  C3 I169 (internal_0n[11], partCD_0n[33], partCD_0n[34], partCD_0n[35]);
  C3 I170 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I171 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I172 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I173 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I174 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I175 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I176 (cd_0n, internal_0n[16], internal_0n[17]);
  OR2 I177 (partCD_0n[0], store_0n[0], store_1n[0]);
  OR2 I178 (partCD_0n[1], store_0n[1], store_1n[1]);
  OR2 I179 (partCD_0n[2], store_0n[2], store_1n[2]);
  OR2 I180 (partCD_0n[3], store_0n[3], store_1n[3]);
  OR2 I181 (partCD_0n[4], store_0n[4], store_1n[4]);
  OR2 I182 (partCD_0n[5], store_0n[5], store_1n[5]);
  OR2 I183 (partCD_0n[6], store_0n[6], store_1n[6]);
  OR2 I184 (partCD_0n[7], store_0n[7], store_1n[7]);
  OR2 I185 (partCD_0n[8], store_0n[8], store_1n[8]);
  OR2 I186 (partCD_0n[9], store_0n[9], store_1n[9]);
  OR2 I187 (partCD_0n[10], store_0n[10], store_1n[10]);
  OR2 I188 (partCD_0n[11], store_0n[11], store_1n[11]);
  OR2 I189 (partCD_0n[12], store_0n[12], store_1n[12]);
  OR2 I190 (partCD_0n[13], store_0n[13], store_1n[13]);
  OR2 I191 (partCD_0n[14], store_0n[14], store_1n[14]);
  OR2 I192 (partCD_0n[15], store_0n[15], store_1n[15]);
  OR2 I193 (partCD_0n[16], store_0n[16], store_1n[16]);
  OR2 I194 (partCD_0n[17], store_0n[17], store_1n[17]);
  OR2 I195 (partCD_0n[18], store_0n[18], store_1n[18]);
  OR2 I196 (partCD_0n[19], store_0n[19], store_1n[19]);
  OR2 I197 (partCD_0n[20], store_0n[20], store_1n[20]);
  OR2 I198 (partCD_0n[21], store_0n[21], store_1n[21]);
  OR2 I199 (partCD_0n[22], store_0n[22], store_1n[22]);
  OR2 I200 (partCD_0n[23], store_0n[23], store_1n[23]);
  OR2 I201 (partCD_0n[24], store_0n[24], store_1n[24]);
  OR2 I202 (partCD_0n[25], store_0n[25], store_1n[25]);
  OR2 I203 (partCD_0n[26], store_0n[26], store_1n[26]);
  OR2 I204 (partCD_0n[27], store_0n[27], store_1n[27]);
  OR2 I205 (partCD_0n[28], store_0n[28], store_1n[28]);
  OR2 I206 (partCD_0n[29], store_0n[29], store_1n[29]);
  OR2 I207 (partCD_0n[30], store_0n[30], store_1n[30]);
  OR2 I208 (partCD_0n[31], store_0n[31], store_1n[31]);
  OR2 I209 (partCD_0n[32], store_0n[32], store_1n[32]);
  OR2 I210 (partCD_0n[33], store_0n[33], store_1n[33]);
  OR2 I211 (partCD_0n[34], store_0n[34], store_1n[34]);
  OR2 I212 (partCD_0n[35], store_0n[35], store_1n[35]);
  BUFF I213 (write_0r, trigger_0r);
endmodule

module BrzActiveEagerNullAdapt_1 (
  trigger_0r, trigger_0a,
  inp_0r, inp_0a0d, inp_0a1d,
  signal_0r, signal_0a
);
  input trigger_0r;
  output trigger_0a;
  output inp_0r;
  input inp_0a0d;
  input inp_0a1d;
  output signal_0r;
  input signal_0a;
  wire partCD_0n;
  wire cd_0n;
  wire writeAck_0n;
  C2 I0 (trigger_0a, writeAck_0n, cd_0n);
  BALSA_TELEM I1 (trigger_0r, writeAck_0n, signal_0r, signal_0a);
  BUFF I2 (cd_0n, partCD_0n);
  OR2 I3 (partCD_0n, inp_0a0d, inp_0a1d);
  BUFF I4 (inp_0r, trigger_0r);
endmodule

module BrzActiveEagerNullAdapt_32 (
  trigger_0r, trigger_0a,
  inp_0r, inp_0a0d, inp_0a1d,
  signal_0r, signal_0a
);
  input trigger_0r;
  output trigger_0a;
  output inp_0r;
  input [31:0] inp_0a0d;
  input [31:0] inp_0a1d;
  output signal_0r;
  input signal_0a;
  wire [16:0] internal_0n;
  wire [31:0] partCD_0n;
  wire cd_0n;
  wire writeAck_0n;
  C2 I0 (trigger_0a, writeAck_0n, cd_0n);
  BALSA_TELEM I1 (trigger_0r, writeAck_0n, signal_0r, signal_0a);
  C3 I2 (internal_0n[0], partCD_0n[0], partCD_0n[1], partCD_0n[2]);
  C3 I3 (internal_0n[1], partCD_0n[3], partCD_0n[4], partCD_0n[5]);
  C3 I4 (internal_0n[2], partCD_0n[6], partCD_0n[7], partCD_0n[8]);
  C3 I5 (internal_0n[3], partCD_0n[9], partCD_0n[10], partCD_0n[11]);
  C3 I6 (internal_0n[4], partCD_0n[12], partCD_0n[13], partCD_0n[14]);
  C3 I7 (internal_0n[5], partCD_0n[15], partCD_0n[16], partCD_0n[17]);
  C3 I8 (internal_0n[6], partCD_0n[18], partCD_0n[19], partCD_0n[20]);
  C3 I9 (internal_0n[7], partCD_0n[21], partCD_0n[22], partCD_0n[23]);
  C3 I10 (internal_0n[8], partCD_0n[24], partCD_0n[25], partCD_0n[26]);
  C3 I11 (internal_0n[9], partCD_0n[27], partCD_0n[28], partCD_0n[29]);
  C2 I12 (internal_0n[10], partCD_0n[30], partCD_0n[31]);
  C3 I13 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I14 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I15 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I16 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I17 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I18 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I19 (cd_0n, internal_0n[15], internal_0n[16]);
  OR2 I20 (partCD_0n[0], inp_0a0d[0], inp_0a1d[0]);
  OR2 I21 (partCD_0n[1], inp_0a0d[1], inp_0a1d[1]);
  OR2 I22 (partCD_0n[2], inp_0a0d[2], inp_0a1d[2]);
  OR2 I23 (partCD_0n[3], inp_0a0d[3], inp_0a1d[3]);
  OR2 I24 (partCD_0n[4], inp_0a0d[4], inp_0a1d[4]);
  OR2 I25 (partCD_0n[5], inp_0a0d[5], inp_0a1d[5]);
  OR2 I26 (partCD_0n[6], inp_0a0d[6], inp_0a1d[6]);
  OR2 I27 (partCD_0n[7], inp_0a0d[7], inp_0a1d[7]);
  OR2 I28 (partCD_0n[8], inp_0a0d[8], inp_0a1d[8]);
  OR2 I29 (partCD_0n[9], inp_0a0d[9], inp_0a1d[9]);
  OR2 I30 (partCD_0n[10], inp_0a0d[10], inp_0a1d[10]);
  OR2 I31 (partCD_0n[11], inp_0a0d[11], inp_0a1d[11]);
  OR2 I32 (partCD_0n[12], inp_0a0d[12], inp_0a1d[12]);
  OR2 I33 (partCD_0n[13], inp_0a0d[13], inp_0a1d[13]);
  OR2 I34 (partCD_0n[14], inp_0a0d[14], inp_0a1d[14]);
  OR2 I35 (partCD_0n[15], inp_0a0d[15], inp_0a1d[15]);
  OR2 I36 (partCD_0n[16], inp_0a0d[16], inp_0a1d[16]);
  OR2 I37 (partCD_0n[17], inp_0a0d[17], inp_0a1d[17]);
  OR2 I38 (partCD_0n[18], inp_0a0d[18], inp_0a1d[18]);
  OR2 I39 (partCD_0n[19], inp_0a0d[19], inp_0a1d[19]);
  OR2 I40 (partCD_0n[20], inp_0a0d[20], inp_0a1d[20]);
  OR2 I41 (partCD_0n[21], inp_0a0d[21], inp_0a1d[21]);
  OR2 I42 (partCD_0n[22], inp_0a0d[22], inp_0a1d[22]);
  OR2 I43 (partCD_0n[23], inp_0a0d[23], inp_0a1d[23]);
  OR2 I44 (partCD_0n[24], inp_0a0d[24], inp_0a1d[24]);
  OR2 I45 (partCD_0n[25], inp_0a0d[25], inp_0a1d[25]);
  OR2 I46 (partCD_0n[26], inp_0a0d[26], inp_0a1d[26]);
  OR2 I47 (partCD_0n[27], inp_0a0d[27], inp_0a1d[27]);
  OR2 I48 (partCD_0n[28], inp_0a0d[28], inp_0a1d[28]);
  OR2 I49 (partCD_0n[29], inp_0a0d[29], inp_0a1d[29]);
  OR2 I50 (partCD_0n[30], inp_0a0d[30], inp_0a1d[30]);
  OR2 I51 (partCD_0n[31], inp_0a0d[31], inp_0a1d[31]);
  BUFF I52 (inp_0r, trigger_0r);
endmodule

module BrzAdapt_10_9_s5_false_s5_false (
  out_0r, out_0a0d, out_0a1d,
  inp_0r, inp_0a0d, inp_0a1d
);
  input out_0r;
  output [9:0] out_0a0d;
  output [9:0] out_0a1d;
  output inp_0r;
  input [8:0] inp_0a0d;
  input [8:0] inp_0a1d;
  wire extendf_0n;
  wire extendt_0n;
  supply0 gnd;
  BUFF I0 (out_0a1d[9], gnd);
  BUFF I1 (out_0a0d[9], out_0r);
  BUFF I2 (out_0a1d[0], inp_0a1d[0]);
  BUFF I3 (out_0a1d[1], inp_0a1d[1]);
  BUFF I4 (out_0a1d[2], inp_0a1d[2]);
  BUFF I5 (out_0a1d[3], inp_0a1d[3]);
  BUFF I6 (out_0a1d[4], inp_0a1d[4]);
  BUFF I7 (out_0a1d[5], inp_0a1d[5]);
  BUFF I8 (out_0a1d[6], inp_0a1d[6]);
  BUFF I9 (out_0a1d[7], inp_0a1d[7]);
  BUFF I10 (out_0a1d[8], inp_0a1d[8]);
  BUFF I11 (out_0a0d[0], inp_0a0d[0]);
  BUFF I12 (out_0a0d[1], inp_0a0d[1]);
  BUFF I13 (out_0a0d[2], inp_0a0d[2]);
  BUFF I14 (out_0a0d[3], inp_0a0d[3]);
  BUFF I15 (out_0a0d[4], inp_0a0d[4]);
  BUFF I16 (out_0a0d[5], inp_0a0d[5]);
  BUFF I17 (out_0a0d[6], inp_0a0d[6]);
  BUFF I18 (out_0a0d[7], inp_0a0d[7]);
  BUFF I19 (out_0a0d[8], inp_0a0d[8]);
  BUFF I20 (inp_0r, out_0r);
endmodule

module BrzAdapt_32_35_s5_false_s5_false (
  out_0r, out_0a0d, out_0a1d,
  inp_0r, inp_0a0d, inp_0a1d
);
  input out_0r;
  output [31:0] out_0a0d;
  output [31:0] out_0a1d;
  output inp_0r;
  input [34:0] inp_0a0d;
  input [34:0] inp_0a1d;
  wire extendf_0n;
  wire extendt_0n;
  BUFF I0 (out_0a1d[0], inp_0a1d[0]);
  BUFF I1 (out_0a1d[1], inp_0a1d[1]);
  BUFF I2 (out_0a1d[2], inp_0a1d[2]);
  BUFF I3 (out_0a1d[3], inp_0a1d[3]);
  BUFF I4 (out_0a1d[4], inp_0a1d[4]);
  BUFF I5 (out_0a1d[5], inp_0a1d[5]);
  BUFF I6 (out_0a1d[6], inp_0a1d[6]);
  BUFF I7 (out_0a1d[7], inp_0a1d[7]);
  BUFF I8 (out_0a1d[8], inp_0a1d[8]);
  BUFF I9 (out_0a1d[9], inp_0a1d[9]);
  BUFF I10 (out_0a1d[10], inp_0a1d[10]);
  BUFF I11 (out_0a1d[11], inp_0a1d[11]);
  BUFF I12 (out_0a1d[12], inp_0a1d[12]);
  BUFF I13 (out_0a1d[13], inp_0a1d[13]);
  BUFF I14 (out_0a1d[14], inp_0a1d[14]);
  BUFF I15 (out_0a1d[15], inp_0a1d[15]);
  BUFF I16 (out_0a1d[16], inp_0a1d[16]);
  BUFF I17 (out_0a1d[17], inp_0a1d[17]);
  BUFF I18 (out_0a1d[18], inp_0a1d[18]);
  BUFF I19 (out_0a1d[19], inp_0a1d[19]);
  BUFF I20 (out_0a1d[20], inp_0a1d[20]);
  BUFF I21 (out_0a1d[21], inp_0a1d[21]);
  BUFF I22 (out_0a1d[22], inp_0a1d[22]);
  BUFF I23 (out_0a1d[23], inp_0a1d[23]);
  BUFF I24 (out_0a1d[24], inp_0a1d[24]);
  BUFF I25 (out_0a1d[25], inp_0a1d[25]);
  BUFF I26 (out_0a1d[26], inp_0a1d[26]);
  BUFF I27 (out_0a1d[27], inp_0a1d[27]);
  BUFF I28 (out_0a1d[28], inp_0a1d[28]);
  BUFF I29 (out_0a1d[29], inp_0a1d[29]);
  BUFF I30 (out_0a1d[30], inp_0a1d[30]);
  BUFF I31 (out_0a1d[31], inp_0a1d[31]);
  BUFF I32 (out_0a0d[0], inp_0a0d[0]);
  BUFF I33 (out_0a0d[1], inp_0a0d[1]);
  BUFF I34 (out_0a0d[2], inp_0a0d[2]);
  BUFF I35 (out_0a0d[3], inp_0a0d[3]);
  BUFF I36 (out_0a0d[4], inp_0a0d[4]);
  BUFF I37 (out_0a0d[5], inp_0a0d[5]);
  BUFF I38 (out_0a0d[6], inp_0a0d[6]);
  BUFF I39 (out_0a0d[7], inp_0a0d[7]);
  BUFF I40 (out_0a0d[8], inp_0a0d[8]);
  BUFF I41 (out_0a0d[9], inp_0a0d[9]);
  BUFF I42 (out_0a0d[10], inp_0a0d[10]);
  BUFF I43 (out_0a0d[11], inp_0a0d[11]);
  BUFF I44 (out_0a0d[12], inp_0a0d[12]);
  BUFF I45 (out_0a0d[13], inp_0a0d[13]);
  BUFF I46 (out_0a0d[14], inp_0a0d[14]);
  BUFF I47 (out_0a0d[15], inp_0a0d[15]);
  BUFF I48 (out_0a0d[16], inp_0a0d[16]);
  BUFF I49 (out_0a0d[17], inp_0a0d[17]);
  BUFF I50 (out_0a0d[18], inp_0a0d[18]);
  BUFF I51 (out_0a0d[19], inp_0a0d[19]);
  BUFF I52 (out_0a0d[20], inp_0a0d[20]);
  BUFF I53 (out_0a0d[21], inp_0a0d[21]);
  BUFF I54 (out_0a0d[22], inp_0a0d[22]);
  BUFF I55 (out_0a0d[23], inp_0a0d[23]);
  BUFF I56 (out_0a0d[24], inp_0a0d[24]);
  BUFF I57 (out_0a0d[25], inp_0a0d[25]);
  BUFF I58 (out_0a0d[26], inp_0a0d[26]);
  BUFF I59 (out_0a0d[27], inp_0a0d[27]);
  BUFF I60 (out_0a0d[28], inp_0a0d[28]);
  BUFF I61 (out_0a0d[29], inp_0a0d[29]);
  BUFF I62 (out_0a0d[30], inp_0a0d[30]);
  BUFF I63 (out_0a0d[31], inp_0a0d[31]);
  BUFF I64 (inp_0r, out_0r);
endmodule

module BrzAdapt_35_4_s4_true_s4_true (
  out_0r, out_0a0d, out_0a1d,
  inp_0r, inp_0a0d, inp_0a1d
);
  input out_0r;
  output [34:0] out_0a0d;
  output [34:0] out_0a1d;
  output inp_0r;
  input [3:0] inp_0a0d;
  input [3:0] inp_0a1d;
  wire extendf_0n;
  wire extendt_0n;
  BUFF I0 (out_0a1d[4], extendt_0n);
  BUFF I1 (out_0a1d[5], extendt_0n);
  BUFF I2 (out_0a1d[6], extendt_0n);
  BUFF I3 (out_0a1d[7], extendt_0n);
  BUFF I4 (out_0a1d[8], extendt_0n);
  BUFF I5 (out_0a1d[9], extendt_0n);
  BUFF I6 (out_0a1d[10], extendt_0n);
  BUFF I7 (out_0a1d[11], extendt_0n);
  BUFF I8 (out_0a1d[12], extendt_0n);
  BUFF I9 (out_0a1d[13], extendt_0n);
  BUFF I10 (out_0a1d[14], extendt_0n);
  BUFF I11 (out_0a1d[15], extendt_0n);
  BUFF I12 (out_0a1d[16], extendt_0n);
  BUFF I13 (out_0a1d[17], extendt_0n);
  BUFF I14 (out_0a1d[18], extendt_0n);
  BUFF I15 (out_0a1d[19], extendt_0n);
  BUFF I16 (out_0a1d[20], extendt_0n);
  BUFF I17 (out_0a1d[21], extendt_0n);
  BUFF I18 (out_0a1d[22], extendt_0n);
  BUFF I19 (out_0a1d[23], extendt_0n);
  BUFF I20 (out_0a1d[24], extendt_0n);
  BUFF I21 (out_0a1d[25], extendt_0n);
  BUFF I22 (out_0a1d[26], extendt_0n);
  BUFF I23 (out_0a1d[27], extendt_0n);
  BUFF I24 (out_0a1d[28], extendt_0n);
  BUFF I25 (out_0a1d[29], extendt_0n);
  BUFF I26 (out_0a1d[30], extendt_0n);
  BUFF I27 (out_0a1d[31], extendt_0n);
  BUFF I28 (out_0a1d[32], extendt_0n);
  BUFF I29 (out_0a1d[33], extendt_0n);
  BUFF I30 (out_0a1d[34], extendt_0n);
  BUFF I31 (out_0a0d[4], extendf_0n);
  BUFF I32 (out_0a0d[5], extendf_0n);
  BUFF I33 (out_0a0d[6], extendf_0n);
  BUFF I34 (out_0a0d[7], extendf_0n);
  BUFF I35 (out_0a0d[8], extendf_0n);
  BUFF I36 (out_0a0d[9], extendf_0n);
  BUFF I37 (out_0a0d[10], extendf_0n);
  BUFF I38 (out_0a0d[11], extendf_0n);
  BUFF I39 (out_0a0d[12], extendf_0n);
  BUFF I40 (out_0a0d[13], extendf_0n);
  BUFF I41 (out_0a0d[14], extendf_0n);
  BUFF I42 (out_0a0d[15], extendf_0n);
  BUFF I43 (out_0a0d[16], extendf_0n);
  BUFF I44 (out_0a0d[17], extendf_0n);
  BUFF I45 (out_0a0d[18], extendf_0n);
  BUFF I46 (out_0a0d[19], extendf_0n);
  BUFF I47 (out_0a0d[20], extendf_0n);
  BUFF I48 (out_0a0d[21], extendf_0n);
  BUFF I49 (out_0a0d[22], extendf_0n);
  BUFF I50 (out_0a0d[23], extendf_0n);
  BUFF I51 (out_0a0d[24], extendf_0n);
  BUFF I52 (out_0a0d[25], extendf_0n);
  BUFF I53 (out_0a0d[26], extendf_0n);
  BUFF I54 (out_0a0d[27], extendf_0n);
  BUFF I55 (out_0a0d[28], extendf_0n);
  BUFF I56 (out_0a0d[29], extendf_0n);
  BUFF I57 (out_0a0d[30], extendf_0n);
  BUFF I58 (out_0a0d[31], extendf_0n);
  BUFF I59 (out_0a0d[32], extendf_0n);
  BUFF I60 (out_0a0d[33], extendf_0n);
  BUFF I61 (out_0a0d[34], extendf_0n);
  BUFF I62 (extendt_0n, inp_0a1d[3]);
  BUFF I63 (extendf_0n, inp_0a0d[3]);
  BUFF I64 (out_0a1d[0], inp_0a1d[0]);
  BUFF I65 (out_0a1d[1], inp_0a1d[1]);
  BUFF I66 (out_0a1d[2], inp_0a1d[2]);
  BUFF I67 (out_0a1d[3], inp_0a1d[3]);
  BUFF I68 (out_0a0d[0], inp_0a0d[0]);
  BUFF I69 (out_0a0d[1], inp_0a0d[1]);
  BUFF I70 (out_0a0d[2], inp_0a0d[2]);
  BUFF I71 (out_0a0d[3], inp_0a0d[3]);
  BUFF I72 (inp_0r, out_0r);
endmodule

module BrzAdapt_35_32_s5_false_s5_false (
  out_0r, out_0a0d, out_0a1d,
  inp_0r, inp_0a0d, inp_0a1d
);
  input out_0r;
  output [34:0] out_0a0d;
  output [34:0] out_0a1d;
  output inp_0r;
  input [31:0] inp_0a0d;
  input [31:0] inp_0a1d;
  wire extendf_0n;
  wire extendt_0n;
  supply0 gnd;
  BUFF I0 (out_0a1d[32], gnd);
  BUFF I1 (out_0a1d[33], gnd);
  BUFF I2 (out_0a1d[34], gnd);
  BUFF I3 (out_0a0d[32], out_0r);
  BUFF I4 (out_0a0d[33], out_0r);
  BUFF I5 (out_0a0d[34], out_0r);
  BUFF I6 (out_0a1d[0], inp_0a1d[0]);
  BUFF I7 (out_0a1d[1], inp_0a1d[1]);
  BUFF I8 (out_0a1d[2], inp_0a1d[2]);
  BUFF I9 (out_0a1d[3], inp_0a1d[3]);
  BUFF I10 (out_0a1d[4], inp_0a1d[4]);
  BUFF I11 (out_0a1d[5], inp_0a1d[5]);
  BUFF I12 (out_0a1d[6], inp_0a1d[6]);
  BUFF I13 (out_0a1d[7], inp_0a1d[7]);
  BUFF I14 (out_0a1d[8], inp_0a1d[8]);
  BUFF I15 (out_0a1d[9], inp_0a1d[9]);
  BUFF I16 (out_0a1d[10], inp_0a1d[10]);
  BUFF I17 (out_0a1d[11], inp_0a1d[11]);
  BUFF I18 (out_0a1d[12], inp_0a1d[12]);
  BUFF I19 (out_0a1d[13], inp_0a1d[13]);
  BUFF I20 (out_0a1d[14], inp_0a1d[14]);
  BUFF I21 (out_0a1d[15], inp_0a1d[15]);
  BUFF I22 (out_0a1d[16], inp_0a1d[16]);
  BUFF I23 (out_0a1d[17], inp_0a1d[17]);
  BUFF I24 (out_0a1d[18], inp_0a1d[18]);
  BUFF I25 (out_0a1d[19], inp_0a1d[19]);
  BUFF I26 (out_0a1d[20], inp_0a1d[20]);
  BUFF I27 (out_0a1d[21], inp_0a1d[21]);
  BUFF I28 (out_0a1d[22], inp_0a1d[22]);
  BUFF I29 (out_0a1d[23], inp_0a1d[23]);
  BUFF I30 (out_0a1d[24], inp_0a1d[24]);
  BUFF I31 (out_0a1d[25], inp_0a1d[25]);
  BUFF I32 (out_0a1d[26], inp_0a1d[26]);
  BUFF I33 (out_0a1d[27], inp_0a1d[27]);
  BUFF I34 (out_0a1d[28], inp_0a1d[28]);
  BUFF I35 (out_0a1d[29], inp_0a1d[29]);
  BUFF I36 (out_0a1d[30], inp_0a1d[30]);
  BUFF I37 (out_0a1d[31], inp_0a1d[31]);
  BUFF I38 (out_0a0d[0], inp_0a0d[0]);
  BUFF I39 (out_0a0d[1], inp_0a0d[1]);
  BUFF I40 (out_0a0d[2], inp_0a0d[2]);
  BUFF I41 (out_0a0d[3], inp_0a0d[3]);
  BUFF I42 (out_0a0d[4], inp_0a0d[4]);
  BUFF I43 (out_0a0d[5], inp_0a0d[5]);
  BUFF I44 (out_0a0d[6], inp_0a0d[6]);
  BUFF I45 (out_0a0d[7], inp_0a0d[7]);
  BUFF I46 (out_0a0d[8], inp_0a0d[8]);
  BUFF I47 (out_0a0d[9], inp_0a0d[9]);
  BUFF I48 (out_0a0d[10], inp_0a0d[10]);
  BUFF I49 (out_0a0d[11], inp_0a0d[11]);
  BUFF I50 (out_0a0d[12], inp_0a0d[12]);
  BUFF I51 (out_0a0d[13], inp_0a0d[13]);
  BUFF I52 (out_0a0d[14], inp_0a0d[14]);
  BUFF I53 (out_0a0d[15], inp_0a0d[15]);
  BUFF I54 (out_0a0d[16], inp_0a0d[16]);
  BUFF I55 (out_0a0d[17], inp_0a0d[17]);
  BUFF I56 (out_0a0d[18], inp_0a0d[18]);
  BUFF I57 (out_0a0d[19], inp_0a0d[19]);
  BUFF I58 (out_0a0d[20], inp_0a0d[20]);
  BUFF I59 (out_0a0d[21], inp_0a0d[21]);
  BUFF I60 (out_0a0d[22], inp_0a0d[22]);
  BUFF I61 (out_0a0d[23], inp_0a0d[23]);
  BUFF I62 (out_0a0d[24], inp_0a0d[24]);
  BUFF I63 (out_0a0d[25], inp_0a0d[25]);
  BUFF I64 (out_0a0d[26], inp_0a0d[26]);
  BUFF I65 (out_0a0d[27], inp_0a0d[27]);
  BUFF I66 (out_0a0d[28], inp_0a0d[28]);
  BUFF I67 (out_0a0d[29], inp_0a0d[29]);
  BUFF I68 (out_0a0d[30], inp_0a0d[30]);
  BUFF I69 (out_0a0d[31], inp_0a0d[31]);
  BUFF I70 (inp_0r, out_0r);
endmodule

module BrzAdapt_35_32_s4_true_s4_true (
  out_0r, out_0a0d, out_0a1d,
  inp_0r, inp_0a0d, inp_0a1d
);
  input out_0r;
  output [34:0] out_0a0d;
  output [34:0] out_0a1d;
  output inp_0r;
  input [31:0] inp_0a0d;
  input [31:0] inp_0a1d;
  wire extendf_0n;
  wire extendt_0n;
  BUFF I0 (out_0a1d[32], extendt_0n);
  BUFF I1 (out_0a1d[33], extendt_0n);
  BUFF I2 (out_0a1d[34], extendt_0n);
  BUFF I3 (out_0a0d[32], extendf_0n);
  BUFF I4 (out_0a0d[33], extendf_0n);
  BUFF I5 (out_0a0d[34], extendf_0n);
  BUFF I6 (extendt_0n, inp_0a1d[31]);
  BUFF I7 (extendf_0n, inp_0a0d[31]);
  BUFF I8 (out_0a1d[0], inp_0a1d[0]);
  BUFF I9 (out_0a1d[1], inp_0a1d[1]);
  BUFF I10 (out_0a1d[2], inp_0a1d[2]);
  BUFF I11 (out_0a1d[3], inp_0a1d[3]);
  BUFF I12 (out_0a1d[4], inp_0a1d[4]);
  BUFF I13 (out_0a1d[5], inp_0a1d[5]);
  BUFF I14 (out_0a1d[6], inp_0a1d[6]);
  BUFF I15 (out_0a1d[7], inp_0a1d[7]);
  BUFF I16 (out_0a1d[8], inp_0a1d[8]);
  BUFF I17 (out_0a1d[9], inp_0a1d[9]);
  BUFF I18 (out_0a1d[10], inp_0a1d[10]);
  BUFF I19 (out_0a1d[11], inp_0a1d[11]);
  BUFF I20 (out_0a1d[12], inp_0a1d[12]);
  BUFF I21 (out_0a1d[13], inp_0a1d[13]);
  BUFF I22 (out_0a1d[14], inp_0a1d[14]);
  BUFF I23 (out_0a1d[15], inp_0a1d[15]);
  BUFF I24 (out_0a1d[16], inp_0a1d[16]);
  BUFF I25 (out_0a1d[17], inp_0a1d[17]);
  BUFF I26 (out_0a1d[18], inp_0a1d[18]);
  BUFF I27 (out_0a1d[19], inp_0a1d[19]);
  BUFF I28 (out_0a1d[20], inp_0a1d[20]);
  BUFF I29 (out_0a1d[21], inp_0a1d[21]);
  BUFF I30 (out_0a1d[22], inp_0a1d[22]);
  BUFF I31 (out_0a1d[23], inp_0a1d[23]);
  BUFF I32 (out_0a1d[24], inp_0a1d[24]);
  BUFF I33 (out_0a1d[25], inp_0a1d[25]);
  BUFF I34 (out_0a1d[26], inp_0a1d[26]);
  BUFF I35 (out_0a1d[27], inp_0a1d[27]);
  BUFF I36 (out_0a1d[28], inp_0a1d[28]);
  BUFF I37 (out_0a1d[29], inp_0a1d[29]);
  BUFF I38 (out_0a1d[30], inp_0a1d[30]);
  BUFF I39 (out_0a1d[31], inp_0a1d[31]);
  BUFF I40 (out_0a0d[0], inp_0a0d[0]);
  BUFF I41 (out_0a0d[1], inp_0a0d[1]);
  BUFF I42 (out_0a0d[2], inp_0a0d[2]);
  BUFF I43 (out_0a0d[3], inp_0a0d[3]);
  BUFF I44 (out_0a0d[4], inp_0a0d[4]);
  BUFF I45 (out_0a0d[5], inp_0a0d[5]);
  BUFF I46 (out_0a0d[6], inp_0a0d[6]);
  BUFF I47 (out_0a0d[7], inp_0a0d[7]);
  BUFF I48 (out_0a0d[8], inp_0a0d[8]);
  BUFF I49 (out_0a0d[9], inp_0a0d[9]);
  BUFF I50 (out_0a0d[10], inp_0a0d[10]);
  BUFF I51 (out_0a0d[11], inp_0a0d[11]);
  BUFF I52 (out_0a0d[12], inp_0a0d[12]);
  BUFF I53 (out_0a0d[13], inp_0a0d[13]);
  BUFF I54 (out_0a0d[14], inp_0a0d[14]);
  BUFF I55 (out_0a0d[15], inp_0a0d[15]);
  BUFF I56 (out_0a0d[16], inp_0a0d[16]);
  BUFF I57 (out_0a0d[17], inp_0a0d[17]);
  BUFF I58 (out_0a0d[18], inp_0a0d[18]);
  BUFF I59 (out_0a0d[19], inp_0a0d[19]);
  BUFF I60 (out_0a0d[20], inp_0a0d[20]);
  BUFF I61 (out_0a0d[21], inp_0a0d[21]);
  BUFF I62 (out_0a0d[22], inp_0a0d[22]);
  BUFF I63 (out_0a0d[23], inp_0a0d[23]);
  BUFF I64 (out_0a0d[24], inp_0a0d[24]);
  BUFF I65 (out_0a0d[25], inp_0a0d[25]);
  BUFF I66 (out_0a0d[26], inp_0a0d[26]);
  BUFF I67 (out_0a0d[27], inp_0a0d[27]);
  BUFF I68 (out_0a0d[28], inp_0a0d[28]);
  BUFF I69 (out_0a0d[29], inp_0a0d[29]);
  BUFF I70 (out_0a0d[30], inp_0a0d[30]);
  BUFF I71 (out_0a0d[31], inp_0a0d[31]);
  BUFF I72 (inp_0r, out_0r);
endmodule

module BrzAdapt_36_33_s5_false_s5_false (
  out_0r, out_0a0d, out_0a1d,
  inp_0r, inp_0a0d, inp_0a1d
);
  input out_0r;
  output [35:0] out_0a0d;
  output [35:0] out_0a1d;
  output inp_0r;
  input [32:0] inp_0a0d;
  input [32:0] inp_0a1d;
  wire extendf_0n;
  wire extendt_0n;
  supply0 gnd;
  BUFF I0 (out_0a1d[33], gnd);
  BUFF I1 (out_0a1d[34], gnd);
  BUFF I2 (out_0a1d[35], gnd);
  BUFF I3 (out_0a0d[33], out_0r);
  BUFF I4 (out_0a0d[34], out_0r);
  BUFF I5 (out_0a0d[35], out_0r);
  BUFF I6 (out_0a1d[0], inp_0a1d[0]);
  BUFF I7 (out_0a1d[1], inp_0a1d[1]);
  BUFF I8 (out_0a1d[2], inp_0a1d[2]);
  BUFF I9 (out_0a1d[3], inp_0a1d[3]);
  BUFF I10 (out_0a1d[4], inp_0a1d[4]);
  BUFF I11 (out_0a1d[5], inp_0a1d[5]);
  BUFF I12 (out_0a1d[6], inp_0a1d[6]);
  BUFF I13 (out_0a1d[7], inp_0a1d[7]);
  BUFF I14 (out_0a1d[8], inp_0a1d[8]);
  BUFF I15 (out_0a1d[9], inp_0a1d[9]);
  BUFF I16 (out_0a1d[10], inp_0a1d[10]);
  BUFF I17 (out_0a1d[11], inp_0a1d[11]);
  BUFF I18 (out_0a1d[12], inp_0a1d[12]);
  BUFF I19 (out_0a1d[13], inp_0a1d[13]);
  BUFF I20 (out_0a1d[14], inp_0a1d[14]);
  BUFF I21 (out_0a1d[15], inp_0a1d[15]);
  BUFF I22 (out_0a1d[16], inp_0a1d[16]);
  BUFF I23 (out_0a1d[17], inp_0a1d[17]);
  BUFF I24 (out_0a1d[18], inp_0a1d[18]);
  BUFF I25 (out_0a1d[19], inp_0a1d[19]);
  BUFF I26 (out_0a1d[20], inp_0a1d[20]);
  BUFF I27 (out_0a1d[21], inp_0a1d[21]);
  BUFF I28 (out_0a1d[22], inp_0a1d[22]);
  BUFF I29 (out_0a1d[23], inp_0a1d[23]);
  BUFF I30 (out_0a1d[24], inp_0a1d[24]);
  BUFF I31 (out_0a1d[25], inp_0a1d[25]);
  BUFF I32 (out_0a1d[26], inp_0a1d[26]);
  BUFF I33 (out_0a1d[27], inp_0a1d[27]);
  BUFF I34 (out_0a1d[28], inp_0a1d[28]);
  BUFF I35 (out_0a1d[29], inp_0a1d[29]);
  BUFF I36 (out_0a1d[30], inp_0a1d[30]);
  BUFF I37 (out_0a1d[31], inp_0a1d[31]);
  BUFF I38 (out_0a1d[32], inp_0a1d[32]);
  BUFF I39 (out_0a0d[0], inp_0a0d[0]);
  BUFF I40 (out_0a0d[1], inp_0a0d[1]);
  BUFF I41 (out_0a0d[2], inp_0a0d[2]);
  BUFF I42 (out_0a0d[3], inp_0a0d[3]);
  BUFF I43 (out_0a0d[4], inp_0a0d[4]);
  BUFF I44 (out_0a0d[5], inp_0a0d[5]);
  BUFF I45 (out_0a0d[6], inp_0a0d[6]);
  BUFF I46 (out_0a0d[7], inp_0a0d[7]);
  BUFF I47 (out_0a0d[8], inp_0a0d[8]);
  BUFF I48 (out_0a0d[9], inp_0a0d[9]);
  BUFF I49 (out_0a0d[10], inp_0a0d[10]);
  BUFF I50 (out_0a0d[11], inp_0a0d[11]);
  BUFF I51 (out_0a0d[12], inp_0a0d[12]);
  BUFF I52 (out_0a0d[13], inp_0a0d[13]);
  BUFF I53 (out_0a0d[14], inp_0a0d[14]);
  BUFF I54 (out_0a0d[15], inp_0a0d[15]);
  BUFF I55 (out_0a0d[16], inp_0a0d[16]);
  BUFF I56 (out_0a0d[17], inp_0a0d[17]);
  BUFF I57 (out_0a0d[18], inp_0a0d[18]);
  BUFF I58 (out_0a0d[19], inp_0a0d[19]);
  BUFF I59 (out_0a0d[20], inp_0a0d[20]);
  BUFF I60 (out_0a0d[21], inp_0a0d[21]);
  BUFF I61 (out_0a0d[22], inp_0a0d[22]);
  BUFF I62 (out_0a0d[23], inp_0a0d[23]);
  BUFF I63 (out_0a0d[24], inp_0a0d[24]);
  BUFF I64 (out_0a0d[25], inp_0a0d[25]);
  BUFF I65 (out_0a0d[26], inp_0a0d[26]);
  BUFF I66 (out_0a0d[27], inp_0a0d[27]);
  BUFF I67 (out_0a0d[28], inp_0a0d[28]);
  BUFF I68 (out_0a0d[29], inp_0a0d[29]);
  BUFF I69 (out_0a0d[30], inp_0a0d[30]);
  BUFF I70 (out_0a0d[31], inp_0a0d[31]);
  BUFF I71 (out_0a0d[32], inp_0a0d[32]);
  BUFF I72 (inp_0r, out_0r);
endmodule

module BrzAdapt_36_33_s4_true_s4_true (
  out_0r, out_0a0d, out_0a1d,
  inp_0r, inp_0a0d, inp_0a1d
);
  input out_0r;
  output [35:0] out_0a0d;
  output [35:0] out_0a1d;
  output inp_0r;
  input [32:0] inp_0a0d;
  input [32:0] inp_0a1d;
  wire extendf_0n;
  wire extendt_0n;
  BUFF I0 (out_0a1d[33], extendt_0n);
  BUFF I1 (out_0a1d[34], extendt_0n);
  BUFF I2 (out_0a1d[35], extendt_0n);
  BUFF I3 (out_0a0d[33], extendf_0n);
  BUFF I4 (out_0a0d[34], extendf_0n);
  BUFF I5 (out_0a0d[35], extendf_0n);
  BUFF I6 (extendt_0n, inp_0a1d[32]);
  BUFF I7 (extendf_0n, inp_0a0d[32]);
  BUFF I8 (out_0a1d[0], inp_0a1d[0]);
  BUFF I9 (out_0a1d[1], inp_0a1d[1]);
  BUFF I10 (out_0a1d[2], inp_0a1d[2]);
  BUFF I11 (out_0a1d[3], inp_0a1d[3]);
  BUFF I12 (out_0a1d[4], inp_0a1d[4]);
  BUFF I13 (out_0a1d[5], inp_0a1d[5]);
  BUFF I14 (out_0a1d[6], inp_0a1d[6]);
  BUFF I15 (out_0a1d[7], inp_0a1d[7]);
  BUFF I16 (out_0a1d[8], inp_0a1d[8]);
  BUFF I17 (out_0a1d[9], inp_0a1d[9]);
  BUFF I18 (out_0a1d[10], inp_0a1d[10]);
  BUFF I19 (out_0a1d[11], inp_0a1d[11]);
  BUFF I20 (out_0a1d[12], inp_0a1d[12]);
  BUFF I21 (out_0a1d[13], inp_0a1d[13]);
  BUFF I22 (out_0a1d[14], inp_0a1d[14]);
  BUFF I23 (out_0a1d[15], inp_0a1d[15]);
  BUFF I24 (out_0a1d[16], inp_0a1d[16]);
  BUFF I25 (out_0a1d[17], inp_0a1d[17]);
  BUFF I26 (out_0a1d[18], inp_0a1d[18]);
  BUFF I27 (out_0a1d[19], inp_0a1d[19]);
  BUFF I28 (out_0a1d[20], inp_0a1d[20]);
  BUFF I29 (out_0a1d[21], inp_0a1d[21]);
  BUFF I30 (out_0a1d[22], inp_0a1d[22]);
  BUFF I31 (out_0a1d[23], inp_0a1d[23]);
  BUFF I32 (out_0a1d[24], inp_0a1d[24]);
  BUFF I33 (out_0a1d[25], inp_0a1d[25]);
  BUFF I34 (out_0a1d[26], inp_0a1d[26]);
  BUFF I35 (out_0a1d[27], inp_0a1d[27]);
  BUFF I36 (out_0a1d[28], inp_0a1d[28]);
  BUFF I37 (out_0a1d[29], inp_0a1d[29]);
  BUFF I38 (out_0a1d[30], inp_0a1d[30]);
  BUFF I39 (out_0a1d[31], inp_0a1d[31]);
  BUFF I40 (out_0a1d[32], inp_0a1d[32]);
  BUFF I41 (out_0a0d[0], inp_0a0d[0]);
  BUFF I42 (out_0a0d[1], inp_0a0d[1]);
  BUFF I43 (out_0a0d[2], inp_0a0d[2]);
  BUFF I44 (out_0a0d[3], inp_0a0d[3]);
  BUFF I45 (out_0a0d[4], inp_0a0d[4]);
  BUFF I46 (out_0a0d[5], inp_0a0d[5]);
  BUFF I47 (out_0a0d[6], inp_0a0d[6]);
  BUFF I48 (out_0a0d[7], inp_0a0d[7]);
  BUFF I49 (out_0a0d[8], inp_0a0d[8]);
  BUFF I50 (out_0a0d[9], inp_0a0d[9]);
  BUFF I51 (out_0a0d[10], inp_0a0d[10]);
  BUFF I52 (out_0a0d[11], inp_0a0d[11]);
  BUFF I53 (out_0a0d[12], inp_0a0d[12]);
  BUFF I54 (out_0a0d[13], inp_0a0d[13]);
  BUFF I55 (out_0a0d[14], inp_0a0d[14]);
  BUFF I56 (out_0a0d[15], inp_0a0d[15]);
  BUFF I57 (out_0a0d[16], inp_0a0d[16]);
  BUFF I58 (out_0a0d[17], inp_0a0d[17]);
  BUFF I59 (out_0a0d[18], inp_0a0d[18]);
  BUFF I60 (out_0a0d[19], inp_0a0d[19]);
  BUFF I61 (out_0a0d[20], inp_0a0d[20]);
  BUFF I62 (out_0a0d[21], inp_0a0d[21]);
  BUFF I63 (out_0a0d[22], inp_0a0d[22]);
  BUFF I64 (out_0a0d[23], inp_0a0d[23]);
  BUFF I65 (out_0a0d[24], inp_0a0d[24]);
  BUFF I66 (out_0a0d[25], inp_0a0d[25]);
  BUFF I67 (out_0a0d[26], inp_0a0d[26]);
  BUFF I68 (out_0a0d[27], inp_0a0d[27]);
  BUFF I69 (out_0a0d[28], inp_0a0d[28]);
  BUFF I70 (out_0a0d[29], inp_0a0d[29]);
  BUFF I71 (out_0a0d[30], inp_0a0d[30]);
  BUFF I72 (out_0a0d[31], inp_0a0d[31]);
  BUFF I73 (out_0a0d[32], inp_0a0d[32]);
  BUFF I74 (inp_0r, out_0r);
endmodule

module BrzAdapt_36_35_s5_false_s5_false (
  out_0r, out_0a0d, out_0a1d,
  inp_0r, inp_0a0d, inp_0a1d
);
  input out_0r;
  output [35:0] out_0a0d;
  output [35:0] out_0a1d;
  output inp_0r;
  input [34:0] inp_0a0d;
  input [34:0] inp_0a1d;
  wire extendf_0n;
  wire extendt_0n;
  supply0 gnd;
  BUFF I0 (out_0a1d[35], gnd);
  BUFF I1 (out_0a0d[35], out_0r);
  BUFF I2 (out_0a1d[0], inp_0a1d[0]);
  BUFF I3 (out_0a1d[1], inp_0a1d[1]);
  BUFF I4 (out_0a1d[2], inp_0a1d[2]);
  BUFF I5 (out_0a1d[3], inp_0a1d[3]);
  BUFF I6 (out_0a1d[4], inp_0a1d[4]);
  BUFF I7 (out_0a1d[5], inp_0a1d[5]);
  BUFF I8 (out_0a1d[6], inp_0a1d[6]);
  BUFF I9 (out_0a1d[7], inp_0a1d[7]);
  BUFF I10 (out_0a1d[8], inp_0a1d[8]);
  BUFF I11 (out_0a1d[9], inp_0a1d[9]);
  BUFF I12 (out_0a1d[10], inp_0a1d[10]);
  BUFF I13 (out_0a1d[11], inp_0a1d[11]);
  BUFF I14 (out_0a1d[12], inp_0a1d[12]);
  BUFF I15 (out_0a1d[13], inp_0a1d[13]);
  BUFF I16 (out_0a1d[14], inp_0a1d[14]);
  BUFF I17 (out_0a1d[15], inp_0a1d[15]);
  BUFF I18 (out_0a1d[16], inp_0a1d[16]);
  BUFF I19 (out_0a1d[17], inp_0a1d[17]);
  BUFF I20 (out_0a1d[18], inp_0a1d[18]);
  BUFF I21 (out_0a1d[19], inp_0a1d[19]);
  BUFF I22 (out_0a1d[20], inp_0a1d[20]);
  BUFF I23 (out_0a1d[21], inp_0a1d[21]);
  BUFF I24 (out_0a1d[22], inp_0a1d[22]);
  BUFF I25 (out_0a1d[23], inp_0a1d[23]);
  BUFF I26 (out_0a1d[24], inp_0a1d[24]);
  BUFF I27 (out_0a1d[25], inp_0a1d[25]);
  BUFF I28 (out_0a1d[26], inp_0a1d[26]);
  BUFF I29 (out_0a1d[27], inp_0a1d[27]);
  BUFF I30 (out_0a1d[28], inp_0a1d[28]);
  BUFF I31 (out_0a1d[29], inp_0a1d[29]);
  BUFF I32 (out_0a1d[30], inp_0a1d[30]);
  BUFF I33 (out_0a1d[31], inp_0a1d[31]);
  BUFF I34 (out_0a1d[32], inp_0a1d[32]);
  BUFF I35 (out_0a1d[33], inp_0a1d[33]);
  BUFF I36 (out_0a1d[34], inp_0a1d[34]);
  BUFF I37 (out_0a0d[0], inp_0a0d[0]);
  BUFF I38 (out_0a0d[1], inp_0a0d[1]);
  BUFF I39 (out_0a0d[2], inp_0a0d[2]);
  BUFF I40 (out_0a0d[3], inp_0a0d[3]);
  BUFF I41 (out_0a0d[4], inp_0a0d[4]);
  BUFF I42 (out_0a0d[5], inp_0a0d[5]);
  BUFF I43 (out_0a0d[6], inp_0a0d[6]);
  BUFF I44 (out_0a0d[7], inp_0a0d[7]);
  BUFF I45 (out_0a0d[8], inp_0a0d[8]);
  BUFF I46 (out_0a0d[9], inp_0a0d[9]);
  BUFF I47 (out_0a0d[10], inp_0a0d[10]);
  BUFF I48 (out_0a0d[11], inp_0a0d[11]);
  BUFF I49 (out_0a0d[12], inp_0a0d[12]);
  BUFF I50 (out_0a0d[13], inp_0a0d[13]);
  BUFF I51 (out_0a0d[14], inp_0a0d[14]);
  BUFF I52 (out_0a0d[15], inp_0a0d[15]);
  BUFF I53 (out_0a0d[16], inp_0a0d[16]);
  BUFF I54 (out_0a0d[17], inp_0a0d[17]);
  BUFF I55 (out_0a0d[18], inp_0a0d[18]);
  BUFF I56 (out_0a0d[19], inp_0a0d[19]);
  BUFF I57 (out_0a0d[20], inp_0a0d[20]);
  BUFF I58 (out_0a0d[21], inp_0a0d[21]);
  BUFF I59 (out_0a0d[22], inp_0a0d[22]);
  BUFF I60 (out_0a0d[23], inp_0a0d[23]);
  BUFF I61 (out_0a0d[24], inp_0a0d[24]);
  BUFF I62 (out_0a0d[25], inp_0a0d[25]);
  BUFF I63 (out_0a0d[26], inp_0a0d[26]);
  BUFF I64 (out_0a0d[27], inp_0a0d[27]);
  BUFF I65 (out_0a0d[28], inp_0a0d[28]);
  BUFF I66 (out_0a0d[29], inp_0a0d[29]);
  BUFF I67 (out_0a0d[30], inp_0a0d[30]);
  BUFF I68 (out_0a0d[31], inp_0a0d[31]);
  BUFF I69 (out_0a0d[32], inp_0a0d[32]);
  BUFF I70 (out_0a0d[33], inp_0a0d[33]);
  BUFF I71 (out_0a0d[34], inp_0a0d[34]);
  BUFF I72 (inp_0r, out_0r);
endmodule

module DRAND2 (
  i0_0,
  i0_1,
  i1_0,
  i1_1,
  q_0,
  q_1
);
  input i0_0;
  input i0_1;
  input i1_0;
  input i1_1;
  output q_0;
  output q_1;
  wire n0_0n;
  wire n1_0n;
  wire n2_0n;
  OR3 I0 (q_0, n0_0n, n1_0n, n2_0n);
  C2 I1 (n0_0n, i0_0, i1_0);
  C2 I2 (n1_0n, i0_0, i1_1);
  C2 I3 (n2_0n, i0_1, i1_0);
  C2 I4 (q_1, i0_1, i1_1);
endmodule

module BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m15m (
  out_0r, out_0a0d, out_0a1d,
  inpA_0r, inpA_0a0d, inpA_0a1d,
  inpB_0r, inpB_0a0d, inpB_0a1d
);
  input out_0r;
  output out_0a0d;
  output out_0a1d;
  output inpA_0r;
  input inpA_0a0d;
  input inpA_0a1d;
  output inpB_0r;
  input inpB_0a0d;
  input inpB_0a1d;
  wire n1_0n;
  wire n0_0n;
  wire w1_0n;
  wire w0_0n;
  DRAND2 I0 (n0_0n, n1_0n, w0_0n, w1_0n, out_0a0d, out_0a1d);
  BUFF I1 (n0_0n, inpB_0a0d);
  BUFF I2 (n1_0n, inpB_0a1d);
  BUFF I3 (w0_0n, inpA_0a0d);
  BUFF I4 (w1_0n, inpA_0a1d);
  BUFF I5 (inpA_0r, out_0r);
  BUFF I6 (inpB_0r, out_0r);
endmodule

module AO222 (
  q,
  i0,
  i1,
  i2,
  i3,
  i4,
  i5
);
  output q;
  input i0;
  input i1;
  input i2;
  input i3;
  input i4;
  input i5;
  wire [2:0] int_0n;
  OR3 I0 (q, int_0n[0], int_0n[1], int_0n[2]);
  AND2 I1 (int_0n[2], i4, i5);
  AND2 I2 (int_0n[1], i2, i3);
  AND2 I3 (int_0n[0], i0, i1);
endmodule

module DRFA (
  a0,
  a1,
  b0,
  b1,
  ci0,
  ci1,
  co0,
  co1,
  sum0,
  sum1
);
  input a0;
  input a1;
  input b0;
  input b1;
  input ci0;
  input ci1;
  output co0;
  output co1;
  output sum0;
  output sum1;
  wire [7:0] internal_0n;
  wire [7:0] minterm_0n;
  AO222 I0 (co0, a0, b0, a0, ci0, b0, ci0);
  AO222 I1 (co1, a1, b1, a1, ci1, b1, ci1);
  NAND2 I2 (sum0, internal_0n[4], internal_0n[5]);
  NOR2 I3 (internal_0n[5], minterm_0n[5], minterm_0n[6]);
  NOR2 I4 (internal_0n[4], minterm_0n[0], minterm_0n[3]);
  NAND2 I5 (sum1, internal_0n[6], internal_0n[7]);
  NOR2 I6 (internal_0n[7], minterm_0n[4], minterm_0n[7]);
  NOR2 I7 (internal_0n[6], minterm_0n[1], minterm_0n[2]);
  C3 I8 (minterm_0n[7], a1, b1, ci1);
  C3 I9 (minterm_0n[6], a1, b1, ci0);
  C3 I10 (minterm_0n[5], a1, b0, ci1);
  C3 I11 (minterm_0n[4], a1, b0, ci0);
  C3 I12 (minterm_0n[3], a0, b1, ci1);
  C3 I13 (minterm_0n[2], a0, b1, ci0);
  C3 I14 (minterm_0n[1], a0, b0, ci1);
  C3 I15 (minterm_0n[0], a0, b0, ci0);
endmodule

module BrzBinaryFunc_34_33_33_s3_Add_s5_false_s5__m17m (
  out_0r, out_0a0d, out_0a1d,
  inpA_0r, inpA_0a0d, inpA_0a1d,
  inpB_0r, inpB_0a0d, inpB_0a1d
);
  input out_0r;
  output [33:0] out_0a0d;
  output [33:0] out_0a1d;
  output inpA_0r;
  input [32:0] inpA_0a0d;
  input [32:0] inpA_0a1d;
  output inpB_0r;
  input [32:0] inpB_0a0d;
  input [32:0] inpB_0a1d;
  wire [32:0] n1_0n;
  wire [32:0] n0_0n;
  wire [32:0] w1_0n;
  wire [32:0] w0_0n;
  wire [33:0] c1_0n;
  wire [33:0] c0_0n;
  supply0 gnd;
  BUFF I0 (out_0a0d[33], c0_0n[33]);
  BUFF I1 (out_0a1d[33], c1_0n[33]);
  BUFF I2 (c0_0n[0], out_0r);
  BUFF I3 (c1_0n[0], gnd);
  DRFA I4 (n0_0n[32], n1_0n[32], w0_0n[32], w1_0n[32], c0_0n[32], c1_0n[32], c0_0n[33], c1_0n[33], out_0a0d[32], out_0a1d[32]);
  DRFA I5 (n0_0n[0], n1_0n[0], w0_0n[0], w1_0n[0], c0_0n[0], c1_0n[0], c0_0n[1], c1_0n[1], out_0a0d[0], out_0a1d[0]);
  DRFA I6 (n0_0n[1], n1_0n[1], w0_0n[1], w1_0n[1], c0_0n[1], c1_0n[1], c0_0n[2], c1_0n[2], out_0a0d[1], out_0a1d[1]);
  DRFA I7 (n0_0n[2], n1_0n[2], w0_0n[2], w1_0n[2], c0_0n[2], c1_0n[2], c0_0n[3], c1_0n[3], out_0a0d[2], out_0a1d[2]);
  DRFA I8 (n0_0n[3], n1_0n[3], w0_0n[3], w1_0n[3], c0_0n[3], c1_0n[3], c0_0n[4], c1_0n[4], out_0a0d[3], out_0a1d[3]);
  DRFA I9 (n0_0n[4], n1_0n[4], w0_0n[4], w1_0n[4], c0_0n[4], c1_0n[4], c0_0n[5], c1_0n[5], out_0a0d[4], out_0a1d[4]);
  DRFA I10 (n0_0n[5], n1_0n[5], w0_0n[5], w1_0n[5], c0_0n[5], c1_0n[5], c0_0n[6], c1_0n[6], out_0a0d[5], out_0a1d[5]);
  DRFA I11 (n0_0n[6], n1_0n[6], w0_0n[6], w1_0n[6], c0_0n[6], c1_0n[6], c0_0n[7], c1_0n[7], out_0a0d[6], out_0a1d[6]);
  DRFA I12 (n0_0n[7], n1_0n[7], w0_0n[7], w1_0n[7], c0_0n[7], c1_0n[7], c0_0n[8], c1_0n[8], out_0a0d[7], out_0a1d[7]);
  DRFA I13 (n0_0n[8], n1_0n[8], w0_0n[8], w1_0n[8], c0_0n[8], c1_0n[8], c0_0n[9], c1_0n[9], out_0a0d[8], out_0a1d[8]);
  DRFA I14 (n0_0n[9], n1_0n[9], w0_0n[9], w1_0n[9], c0_0n[9], c1_0n[9], c0_0n[10], c1_0n[10], out_0a0d[9], out_0a1d[9]);
  DRFA I15 (n0_0n[10], n1_0n[10], w0_0n[10], w1_0n[10], c0_0n[10], c1_0n[10], c0_0n[11], c1_0n[11], out_0a0d[10], out_0a1d[10]);
  DRFA I16 (n0_0n[11], n1_0n[11], w0_0n[11], w1_0n[11], c0_0n[11], c1_0n[11], c0_0n[12], c1_0n[12], out_0a0d[11], out_0a1d[11]);
  DRFA I17 (n0_0n[12], n1_0n[12], w0_0n[12], w1_0n[12], c0_0n[12], c1_0n[12], c0_0n[13], c1_0n[13], out_0a0d[12], out_0a1d[12]);
  DRFA I18 (n0_0n[13], n1_0n[13], w0_0n[13], w1_0n[13], c0_0n[13], c1_0n[13], c0_0n[14], c1_0n[14], out_0a0d[13], out_0a1d[13]);
  DRFA I19 (n0_0n[14], n1_0n[14], w0_0n[14], w1_0n[14], c0_0n[14], c1_0n[14], c0_0n[15], c1_0n[15], out_0a0d[14], out_0a1d[14]);
  DRFA I20 (n0_0n[15], n1_0n[15], w0_0n[15], w1_0n[15], c0_0n[15], c1_0n[15], c0_0n[16], c1_0n[16], out_0a0d[15], out_0a1d[15]);
  DRFA I21 (n0_0n[16], n1_0n[16], w0_0n[16], w1_0n[16], c0_0n[16], c1_0n[16], c0_0n[17], c1_0n[17], out_0a0d[16], out_0a1d[16]);
  DRFA I22 (n0_0n[17], n1_0n[17], w0_0n[17], w1_0n[17], c0_0n[17], c1_0n[17], c0_0n[18], c1_0n[18], out_0a0d[17], out_0a1d[17]);
  DRFA I23 (n0_0n[18], n1_0n[18], w0_0n[18], w1_0n[18], c0_0n[18], c1_0n[18], c0_0n[19], c1_0n[19], out_0a0d[18], out_0a1d[18]);
  DRFA I24 (n0_0n[19], n1_0n[19], w0_0n[19], w1_0n[19], c0_0n[19], c1_0n[19], c0_0n[20], c1_0n[20], out_0a0d[19], out_0a1d[19]);
  DRFA I25 (n0_0n[20], n1_0n[20], w0_0n[20], w1_0n[20], c0_0n[20], c1_0n[20], c0_0n[21], c1_0n[21], out_0a0d[20], out_0a1d[20]);
  DRFA I26 (n0_0n[21], n1_0n[21], w0_0n[21], w1_0n[21], c0_0n[21], c1_0n[21], c0_0n[22], c1_0n[22], out_0a0d[21], out_0a1d[21]);
  DRFA I27 (n0_0n[22], n1_0n[22], w0_0n[22], w1_0n[22], c0_0n[22], c1_0n[22], c0_0n[23], c1_0n[23], out_0a0d[22], out_0a1d[22]);
  DRFA I28 (n0_0n[23], n1_0n[23], w0_0n[23], w1_0n[23], c0_0n[23], c1_0n[23], c0_0n[24], c1_0n[24], out_0a0d[23], out_0a1d[23]);
  DRFA I29 (n0_0n[24], n1_0n[24], w0_0n[24], w1_0n[24], c0_0n[24], c1_0n[24], c0_0n[25], c1_0n[25], out_0a0d[24], out_0a1d[24]);
  DRFA I30 (n0_0n[25], n1_0n[25], w0_0n[25], w1_0n[25], c0_0n[25], c1_0n[25], c0_0n[26], c1_0n[26], out_0a0d[25], out_0a1d[25]);
  DRFA I31 (n0_0n[26], n1_0n[26], w0_0n[26], w1_0n[26], c0_0n[26], c1_0n[26], c0_0n[27], c1_0n[27], out_0a0d[26], out_0a1d[26]);
  DRFA I32 (n0_0n[27], n1_0n[27], w0_0n[27], w1_0n[27], c0_0n[27], c1_0n[27], c0_0n[28], c1_0n[28], out_0a0d[27], out_0a1d[27]);
  DRFA I33 (n0_0n[28], n1_0n[28], w0_0n[28], w1_0n[28], c0_0n[28], c1_0n[28], c0_0n[29], c1_0n[29], out_0a0d[28], out_0a1d[28]);
  DRFA I34 (n0_0n[29], n1_0n[29], w0_0n[29], w1_0n[29], c0_0n[29], c1_0n[29], c0_0n[30], c1_0n[30], out_0a0d[29], out_0a1d[29]);
  DRFA I35 (n0_0n[30], n1_0n[30], w0_0n[30], w1_0n[30], c0_0n[30], c1_0n[30], c0_0n[31], c1_0n[31], out_0a0d[30], out_0a1d[30]);
  DRFA I36 (n0_0n[31], n1_0n[31], w0_0n[31], w1_0n[31], c0_0n[31], c1_0n[31], c0_0n[32], c1_0n[32], out_0a0d[31], out_0a1d[31]);
  BUFF I37 (n0_0n[0], inpB_0a0d[0]);
  BUFF I38 (n0_0n[1], inpB_0a0d[1]);
  BUFF I39 (n0_0n[2], inpB_0a0d[2]);
  BUFF I40 (n0_0n[3], inpB_0a0d[3]);
  BUFF I41 (n0_0n[4], inpB_0a0d[4]);
  BUFF I42 (n0_0n[5], inpB_0a0d[5]);
  BUFF I43 (n0_0n[6], inpB_0a0d[6]);
  BUFF I44 (n0_0n[7], inpB_0a0d[7]);
  BUFF I45 (n0_0n[8], inpB_0a0d[8]);
  BUFF I46 (n0_0n[9], inpB_0a0d[9]);
  BUFF I47 (n0_0n[10], inpB_0a0d[10]);
  BUFF I48 (n0_0n[11], inpB_0a0d[11]);
  BUFF I49 (n0_0n[12], inpB_0a0d[12]);
  BUFF I50 (n0_0n[13], inpB_0a0d[13]);
  BUFF I51 (n0_0n[14], inpB_0a0d[14]);
  BUFF I52 (n0_0n[15], inpB_0a0d[15]);
  BUFF I53 (n0_0n[16], inpB_0a0d[16]);
  BUFF I54 (n0_0n[17], inpB_0a0d[17]);
  BUFF I55 (n0_0n[18], inpB_0a0d[18]);
  BUFF I56 (n0_0n[19], inpB_0a0d[19]);
  BUFF I57 (n0_0n[20], inpB_0a0d[20]);
  BUFF I58 (n0_0n[21], inpB_0a0d[21]);
  BUFF I59 (n0_0n[22], inpB_0a0d[22]);
  BUFF I60 (n0_0n[23], inpB_0a0d[23]);
  BUFF I61 (n0_0n[24], inpB_0a0d[24]);
  BUFF I62 (n0_0n[25], inpB_0a0d[25]);
  BUFF I63 (n0_0n[26], inpB_0a0d[26]);
  BUFF I64 (n0_0n[27], inpB_0a0d[27]);
  BUFF I65 (n0_0n[28], inpB_0a0d[28]);
  BUFF I66 (n0_0n[29], inpB_0a0d[29]);
  BUFF I67 (n0_0n[30], inpB_0a0d[30]);
  BUFF I68 (n0_0n[31], inpB_0a0d[31]);
  BUFF I69 (n0_0n[32], inpB_0a0d[32]);
  BUFF I70 (n1_0n[0], inpB_0a1d[0]);
  BUFF I71 (n1_0n[1], inpB_0a1d[1]);
  BUFF I72 (n1_0n[2], inpB_0a1d[2]);
  BUFF I73 (n1_0n[3], inpB_0a1d[3]);
  BUFF I74 (n1_0n[4], inpB_0a1d[4]);
  BUFF I75 (n1_0n[5], inpB_0a1d[5]);
  BUFF I76 (n1_0n[6], inpB_0a1d[6]);
  BUFF I77 (n1_0n[7], inpB_0a1d[7]);
  BUFF I78 (n1_0n[8], inpB_0a1d[8]);
  BUFF I79 (n1_0n[9], inpB_0a1d[9]);
  BUFF I80 (n1_0n[10], inpB_0a1d[10]);
  BUFF I81 (n1_0n[11], inpB_0a1d[11]);
  BUFF I82 (n1_0n[12], inpB_0a1d[12]);
  BUFF I83 (n1_0n[13], inpB_0a1d[13]);
  BUFF I84 (n1_0n[14], inpB_0a1d[14]);
  BUFF I85 (n1_0n[15], inpB_0a1d[15]);
  BUFF I86 (n1_0n[16], inpB_0a1d[16]);
  BUFF I87 (n1_0n[17], inpB_0a1d[17]);
  BUFF I88 (n1_0n[18], inpB_0a1d[18]);
  BUFF I89 (n1_0n[19], inpB_0a1d[19]);
  BUFF I90 (n1_0n[20], inpB_0a1d[20]);
  BUFF I91 (n1_0n[21], inpB_0a1d[21]);
  BUFF I92 (n1_0n[22], inpB_0a1d[22]);
  BUFF I93 (n1_0n[23], inpB_0a1d[23]);
  BUFF I94 (n1_0n[24], inpB_0a1d[24]);
  BUFF I95 (n1_0n[25], inpB_0a1d[25]);
  BUFF I96 (n1_0n[26], inpB_0a1d[26]);
  BUFF I97 (n1_0n[27], inpB_0a1d[27]);
  BUFF I98 (n1_0n[28], inpB_0a1d[28]);
  BUFF I99 (n1_0n[29], inpB_0a1d[29]);
  BUFF I100 (n1_0n[30], inpB_0a1d[30]);
  BUFF I101 (n1_0n[31], inpB_0a1d[31]);
  BUFF I102 (n1_0n[32], inpB_0a1d[32]);
  BUFF I103 (w0_0n[0], inpA_0a0d[0]);
  BUFF I104 (w0_0n[1], inpA_0a0d[1]);
  BUFF I105 (w0_0n[2], inpA_0a0d[2]);
  BUFF I106 (w0_0n[3], inpA_0a0d[3]);
  BUFF I107 (w0_0n[4], inpA_0a0d[4]);
  BUFF I108 (w0_0n[5], inpA_0a0d[5]);
  BUFF I109 (w0_0n[6], inpA_0a0d[6]);
  BUFF I110 (w0_0n[7], inpA_0a0d[7]);
  BUFF I111 (w0_0n[8], inpA_0a0d[8]);
  BUFF I112 (w0_0n[9], inpA_0a0d[9]);
  BUFF I113 (w0_0n[10], inpA_0a0d[10]);
  BUFF I114 (w0_0n[11], inpA_0a0d[11]);
  BUFF I115 (w0_0n[12], inpA_0a0d[12]);
  BUFF I116 (w0_0n[13], inpA_0a0d[13]);
  BUFF I117 (w0_0n[14], inpA_0a0d[14]);
  BUFF I118 (w0_0n[15], inpA_0a0d[15]);
  BUFF I119 (w0_0n[16], inpA_0a0d[16]);
  BUFF I120 (w0_0n[17], inpA_0a0d[17]);
  BUFF I121 (w0_0n[18], inpA_0a0d[18]);
  BUFF I122 (w0_0n[19], inpA_0a0d[19]);
  BUFF I123 (w0_0n[20], inpA_0a0d[20]);
  BUFF I124 (w0_0n[21], inpA_0a0d[21]);
  BUFF I125 (w0_0n[22], inpA_0a0d[22]);
  BUFF I126 (w0_0n[23], inpA_0a0d[23]);
  BUFF I127 (w0_0n[24], inpA_0a0d[24]);
  BUFF I128 (w0_0n[25], inpA_0a0d[25]);
  BUFF I129 (w0_0n[26], inpA_0a0d[26]);
  BUFF I130 (w0_0n[27], inpA_0a0d[27]);
  BUFF I131 (w0_0n[28], inpA_0a0d[28]);
  BUFF I132 (w0_0n[29], inpA_0a0d[29]);
  BUFF I133 (w0_0n[30], inpA_0a0d[30]);
  BUFF I134 (w0_0n[31], inpA_0a0d[31]);
  BUFF I135 (w0_0n[32], inpA_0a0d[32]);
  BUFF I136 (w1_0n[0], inpA_0a1d[0]);
  BUFF I137 (w1_0n[1], inpA_0a1d[1]);
  BUFF I138 (w1_0n[2], inpA_0a1d[2]);
  BUFF I139 (w1_0n[3], inpA_0a1d[3]);
  BUFF I140 (w1_0n[4], inpA_0a1d[4]);
  BUFF I141 (w1_0n[5], inpA_0a1d[5]);
  BUFF I142 (w1_0n[6], inpA_0a1d[6]);
  BUFF I143 (w1_0n[7], inpA_0a1d[7]);
  BUFF I144 (w1_0n[8], inpA_0a1d[8]);
  BUFF I145 (w1_0n[9], inpA_0a1d[9]);
  BUFF I146 (w1_0n[10], inpA_0a1d[10]);
  BUFF I147 (w1_0n[11], inpA_0a1d[11]);
  BUFF I148 (w1_0n[12], inpA_0a1d[12]);
  BUFF I149 (w1_0n[13], inpA_0a1d[13]);
  BUFF I150 (w1_0n[14], inpA_0a1d[14]);
  BUFF I151 (w1_0n[15], inpA_0a1d[15]);
  BUFF I152 (w1_0n[16], inpA_0a1d[16]);
  BUFF I153 (w1_0n[17], inpA_0a1d[17]);
  BUFF I154 (w1_0n[18], inpA_0a1d[18]);
  BUFF I155 (w1_0n[19], inpA_0a1d[19]);
  BUFF I156 (w1_0n[20], inpA_0a1d[20]);
  BUFF I157 (w1_0n[21], inpA_0a1d[21]);
  BUFF I158 (w1_0n[22], inpA_0a1d[22]);
  BUFF I159 (w1_0n[23], inpA_0a1d[23]);
  BUFF I160 (w1_0n[24], inpA_0a1d[24]);
  BUFF I161 (w1_0n[25], inpA_0a1d[25]);
  BUFF I162 (w1_0n[26], inpA_0a1d[26]);
  BUFF I163 (w1_0n[27], inpA_0a1d[27]);
  BUFF I164 (w1_0n[28], inpA_0a1d[28]);
  BUFF I165 (w1_0n[29], inpA_0a1d[29]);
  BUFF I166 (w1_0n[30], inpA_0a1d[30]);
  BUFF I167 (w1_0n[31], inpA_0a1d[31]);
  BUFF I168 (w1_0n[32], inpA_0a1d[32]);
  BUFF I169 (inpA_0r, out_0r);
  BUFF I170 (inpB_0r, out_0r);
endmodule

module BrzBinaryFunc_35_35_35_s3_And_s5_false_s5__m19m (
  out_0r, out_0a0d, out_0a1d,
  inpA_0r, inpA_0a0d, inpA_0a1d,
  inpB_0r, inpB_0a0d, inpB_0a1d
);
  input out_0r;
  output [34:0] out_0a0d;
  output [34:0] out_0a1d;
  output inpA_0r;
  input [34:0] inpA_0a0d;
  input [34:0] inpA_0a1d;
  output inpB_0r;
  input [34:0] inpB_0a0d;
  input [34:0] inpB_0a1d;
  wire [34:0] n1_0n;
  wire [34:0] n0_0n;
  wire [34:0] w1_0n;
  wire [34:0] w0_0n;
  DRAND2 I0 (n0_0n[0], n1_0n[0], w0_0n[0], w1_0n[0], out_0a0d[0], out_0a1d[0]);
  DRAND2 I1 (n0_0n[1], n1_0n[1], w0_0n[1], w1_0n[1], out_0a0d[1], out_0a1d[1]);
  DRAND2 I2 (n0_0n[2], n1_0n[2], w0_0n[2], w1_0n[2], out_0a0d[2], out_0a1d[2]);
  DRAND2 I3 (n0_0n[3], n1_0n[3], w0_0n[3], w1_0n[3], out_0a0d[3], out_0a1d[3]);
  DRAND2 I4 (n0_0n[4], n1_0n[4], w0_0n[4], w1_0n[4], out_0a0d[4], out_0a1d[4]);
  DRAND2 I5 (n0_0n[5], n1_0n[5], w0_0n[5], w1_0n[5], out_0a0d[5], out_0a1d[5]);
  DRAND2 I6 (n0_0n[6], n1_0n[6], w0_0n[6], w1_0n[6], out_0a0d[6], out_0a1d[6]);
  DRAND2 I7 (n0_0n[7], n1_0n[7], w0_0n[7], w1_0n[7], out_0a0d[7], out_0a1d[7]);
  DRAND2 I8 (n0_0n[8], n1_0n[8], w0_0n[8], w1_0n[8], out_0a0d[8], out_0a1d[8]);
  DRAND2 I9 (n0_0n[9], n1_0n[9], w0_0n[9], w1_0n[9], out_0a0d[9], out_0a1d[9]);
  DRAND2 I10 (n0_0n[10], n1_0n[10], w0_0n[10], w1_0n[10], out_0a0d[10], out_0a1d[10]);
  DRAND2 I11 (n0_0n[11], n1_0n[11], w0_0n[11], w1_0n[11], out_0a0d[11], out_0a1d[11]);
  DRAND2 I12 (n0_0n[12], n1_0n[12], w0_0n[12], w1_0n[12], out_0a0d[12], out_0a1d[12]);
  DRAND2 I13 (n0_0n[13], n1_0n[13], w0_0n[13], w1_0n[13], out_0a0d[13], out_0a1d[13]);
  DRAND2 I14 (n0_0n[14], n1_0n[14], w0_0n[14], w1_0n[14], out_0a0d[14], out_0a1d[14]);
  DRAND2 I15 (n0_0n[15], n1_0n[15], w0_0n[15], w1_0n[15], out_0a0d[15], out_0a1d[15]);
  DRAND2 I16 (n0_0n[16], n1_0n[16], w0_0n[16], w1_0n[16], out_0a0d[16], out_0a1d[16]);
  DRAND2 I17 (n0_0n[17], n1_0n[17], w0_0n[17], w1_0n[17], out_0a0d[17], out_0a1d[17]);
  DRAND2 I18 (n0_0n[18], n1_0n[18], w0_0n[18], w1_0n[18], out_0a0d[18], out_0a1d[18]);
  DRAND2 I19 (n0_0n[19], n1_0n[19], w0_0n[19], w1_0n[19], out_0a0d[19], out_0a1d[19]);
  DRAND2 I20 (n0_0n[20], n1_0n[20], w0_0n[20], w1_0n[20], out_0a0d[20], out_0a1d[20]);
  DRAND2 I21 (n0_0n[21], n1_0n[21], w0_0n[21], w1_0n[21], out_0a0d[21], out_0a1d[21]);
  DRAND2 I22 (n0_0n[22], n1_0n[22], w0_0n[22], w1_0n[22], out_0a0d[22], out_0a1d[22]);
  DRAND2 I23 (n0_0n[23], n1_0n[23], w0_0n[23], w1_0n[23], out_0a0d[23], out_0a1d[23]);
  DRAND2 I24 (n0_0n[24], n1_0n[24], w0_0n[24], w1_0n[24], out_0a0d[24], out_0a1d[24]);
  DRAND2 I25 (n0_0n[25], n1_0n[25], w0_0n[25], w1_0n[25], out_0a0d[25], out_0a1d[25]);
  DRAND2 I26 (n0_0n[26], n1_0n[26], w0_0n[26], w1_0n[26], out_0a0d[26], out_0a1d[26]);
  DRAND2 I27 (n0_0n[27], n1_0n[27], w0_0n[27], w1_0n[27], out_0a0d[27], out_0a1d[27]);
  DRAND2 I28 (n0_0n[28], n1_0n[28], w0_0n[28], w1_0n[28], out_0a0d[28], out_0a1d[28]);
  DRAND2 I29 (n0_0n[29], n1_0n[29], w0_0n[29], w1_0n[29], out_0a0d[29], out_0a1d[29]);
  DRAND2 I30 (n0_0n[30], n1_0n[30], w0_0n[30], w1_0n[30], out_0a0d[30], out_0a1d[30]);
  DRAND2 I31 (n0_0n[31], n1_0n[31], w0_0n[31], w1_0n[31], out_0a0d[31], out_0a1d[31]);
  DRAND2 I32 (n0_0n[32], n1_0n[32], w0_0n[32], w1_0n[32], out_0a0d[32], out_0a1d[32]);
  DRAND2 I33 (n0_0n[33], n1_0n[33], w0_0n[33], w1_0n[33], out_0a0d[33], out_0a1d[33]);
  DRAND2 I34 (n0_0n[34], n1_0n[34], w0_0n[34], w1_0n[34], out_0a0d[34], out_0a1d[34]);
  BUFF I35 (n0_0n[0], inpB_0a0d[0]);
  BUFF I36 (n0_0n[1], inpB_0a0d[1]);
  BUFF I37 (n0_0n[2], inpB_0a0d[2]);
  BUFF I38 (n0_0n[3], inpB_0a0d[3]);
  BUFF I39 (n0_0n[4], inpB_0a0d[4]);
  BUFF I40 (n0_0n[5], inpB_0a0d[5]);
  BUFF I41 (n0_0n[6], inpB_0a0d[6]);
  BUFF I42 (n0_0n[7], inpB_0a0d[7]);
  BUFF I43 (n0_0n[8], inpB_0a0d[8]);
  BUFF I44 (n0_0n[9], inpB_0a0d[9]);
  BUFF I45 (n0_0n[10], inpB_0a0d[10]);
  BUFF I46 (n0_0n[11], inpB_0a0d[11]);
  BUFF I47 (n0_0n[12], inpB_0a0d[12]);
  BUFF I48 (n0_0n[13], inpB_0a0d[13]);
  BUFF I49 (n0_0n[14], inpB_0a0d[14]);
  BUFF I50 (n0_0n[15], inpB_0a0d[15]);
  BUFF I51 (n0_0n[16], inpB_0a0d[16]);
  BUFF I52 (n0_0n[17], inpB_0a0d[17]);
  BUFF I53 (n0_0n[18], inpB_0a0d[18]);
  BUFF I54 (n0_0n[19], inpB_0a0d[19]);
  BUFF I55 (n0_0n[20], inpB_0a0d[20]);
  BUFF I56 (n0_0n[21], inpB_0a0d[21]);
  BUFF I57 (n0_0n[22], inpB_0a0d[22]);
  BUFF I58 (n0_0n[23], inpB_0a0d[23]);
  BUFF I59 (n0_0n[24], inpB_0a0d[24]);
  BUFF I60 (n0_0n[25], inpB_0a0d[25]);
  BUFF I61 (n0_0n[26], inpB_0a0d[26]);
  BUFF I62 (n0_0n[27], inpB_0a0d[27]);
  BUFF I63 (n0_0n[28], inpB_0a0d[28]);
  BUFF I64 (n0_0n[29], inpB_0a0d[29]);
  BUFF I65 (n0_0n[30], inpB_0a0d[30]);
  BUFF I66 (n0_0n[31], inpB_0a0d[31]);
  BUFF I67 (n0_0n[32], inpB_0a0d[32]);
  BUFF I68 (n0_0n[33], inpB_0a0d[33]);
  BUFF I69 (n0_0n[34], inpB_0a0d[34]);
  BUFF I70 (n1_0n[0], inpB_0a1d[0]);
  BUFF I71 (n1_0n[1], inpB_0a1d[1]);
  BUFF I72 (n1_0n[2], inpB_0a1d[2]);
  BUFF I73 (n1_0n[3], inpB_0a1d[3]);
  BUFF I74 (n1_0n[4], inpB_0a1d[4]);
  BUFF I75 (n1_0n[5], inpB_0a1d[5]);
  BUFF I76 (n1_0n[6], inpB_0a1d[6]);
  BUFF I77 (n1_0n[7], inpB_0a1d[7]);
  BUFF I78 (n1_0n[8], inpB_0a1d[8]);
  BUFF I79 (n1_0n[9], inpB_0a1d[9]);
  BUFF I80 (n1_0n[10], inpB_0a1d[10]);
  BUFF I81 (n1_0n[11], inpB_0a1d[11]);
  BUFF I82 (n1_0n[12], inpB_0a1d[12]);
  BUFF I83 (n1_0n[13], inpB_0a1d[13]);
  BUFF I84 (n1_0n[14], inpB_0a1d[14]);
  BUFF I85 (n1_0n[15], inpB_0a1d[15]);
  BUFF I86 (n1_0n[16], inpB_0a1d[16]);
  BUFF I87 (n1_0n[17], inpB_0a1d[17]);
  BUFF I88 (n1_0n[18], inpB_0a1d[18]);
  BUFF I89 (n1_0n[19], inpB_0a1d[19]);
  BUFF I90 (n1_0n[20], inpB_0a1d[20]);
  BUFF I91 (n1_0n[21], inpB_0a1d[21]);
  BUFF I92 (n1_0n[22], inpB_0a1d[22]);
  BUFF I93 (n1_0n[23], inpB_0a1d[23]);
  BUFF I94 (n1_0n[24], inpB_0a1d[24]);
  BUFF I95 (n1_0n[25], inpB_0a1d[25]);
  BUFF I96 (n1_0n[26], inpB_0a1d[26]);
  BUFF I97 (n1_0n[27], inpB_0a1d[27]);
  BUFF I98 (n1_0n[28], inpB_0a1d[28]);
  BUFF I99 (n1_0n[29], inpB_0a1d[29]);
  BUFF I100 (n1_0n[30], inpB_0a1d[30]);
  BUFF I101 (n1_0n[31], inpB_0a1d[31]);
  BUFF I102 (n1_0n[32], inpB_0a1d[32]);
  BUFF I103 (n1_0n[33], inpB_0a1d[33]);
  BUFF I104 (n1_0n[34], inpB_0a1d[34]);
  BUFF I105 (w0_0n[0], inpA_0a0d[0]);
  BUFF I106 (w0_0n[1], inpA_0a0d[1]);
  BUFF I107 (w0_0n[2], inpA_0a0d[2]);
  BUFF I108 (w0_0n[3], inpA_0a0d[3]);
  BUFF I109 (w0_0n[4], inpA_0a0d[4]);
  BUFF I110 (w0_0n[5], inpA_0a0d[5]);
  BUFF I111 (w0_0n[6], inpA_0a0d[6]);
  BUFF I112 (w0_0n[7], inpA_0a0d[7]);
  BUFF I113 (w0_0n[8], inpA_0a0d[8]);
  BUFF I114 (w0_0n[9], inpA_0a0d[9]);
  BUFF I115 (w0_0n[10], inpA_0a0d[10]);
  BUFF I116 (w0_0n[11], inpA_0a0d[11]);
  BUFF I117 (w0_0n[12], inpA_0a0d[12]);
  BUFF I118 (w0_0n[13], inpA_0a0d[13]);
  BUFF I119 (w0_0n[14], inpA_0a0d[14]);
  BUFF I120 (w0_0n[15], inpA_0a0d[15]);
  BUFF I121 (w0_0n[16], inpA_0a0d[16]);
  BUFF I122 (w0_0n[17], inpA_0a0d[17]);
  BUFF I123 (w0_0n[18], inpA_0a0d[18]);
  BUFF I124 (w0_0n[19], inpA_0a0d[19]);
  BUFF I125 (w0_0n[20], inpA_0a0d[20]);
  BUFF I126 (w0_0n[21], inpA_0a0d[21]);
  BUFF I127 (w0_0n[22], inpA_0a0d[22]);
  BUFF I128 (w0_0n[23], inpA_0a0d[23]);
  BUFF I129 (w0_0n[24], inpA_0a0d[24]);
  BUFF I130 (w0_0n[25], inpA_0a0d[25]);
  BUFF I131 (w0_0n[26], inpA_0a0d[26]);
  BUFF I132 (w0_0n[27], inpA_0a0d[27]);
  BUFF I133 (w0_0n[28], inpA_0a0d[28]);
  BUFF I134 (w0_0n[29], inpA_0a0d[29]);
  BUFF I135 (w0_0n[30], inpA_0a0d[30]);
  BUFF I136 (w0_0n[31], inpA_0a0d[31]);
  BUFF I137 (w0_0n[32], inpA_0a0d[32]);
  BUFF I138 (w0_0n[33], inpA_0a0d[33]);
  BUFF I139 (w0_0n[34], inpA_0a0d[34]);
  BUFF I140 (w1_0n[0], inpA_0a1d[0]);
  BUFF I141 (w1_0n[1], inpA_0a1d[1]);
  BUFF I142 (w1_0n[2], inpA_0a1d[2]);
  BUFF I143 (w1_0n[3], inpA_0a1d[3]);
  BUFF I144 (w1_0n[4], inpA_0a1d[4]);
  BUFF I145 (w1_0n[5], inpA_0a1d[5]);
  BUFF I146 (w1_0n[6], inpA_0a1d[6]);
  BUFF I147 (w1_0n[7], inpA_0a1d[7]);
  BUFF I148 (w1_0n[8], inpA_0a1d[8]);
  BUFF I149 (w1_0n[9], inpA_0a1d[9]);
  BUFF I150 (w1_0n[10], inpA_0a1d[10]);
  BUFF I151 (w1_0n[11], inpA_0a1d[11]);
  BUFF I152 (w1_0n[12], inpA_0a1d[12]);
  BUFF I153 (w1_0n[13], inpA_0a1d[13]);
  BUFF I154 (w1_0n[14], inpA_0a1d[14]);
  BUFF I155 (w1_0n[15], inpA_0a1d[15]);
  BUFF I156 (w1_0n[16], inpA_0a1d[16]);
  BUFF I157 (w1_0n[17], inpA_0a1d[17]);
  BUFF I158 (w1_0n[18], inpA_0a1d[18]);
  BUFF I159 (w1_0n[19], inpA_0a1d[19]);
  BUFF I160 (w1_0n[20], inpA_0a1d[20]);
  BUFF I161 (w1_0n[21], inpA_0a1d[21]);
  BUFF I162 (w1_0n[22], inpA_0a1d[22]);
  BUFF I163 (w1_0n[23], inpA_0a1d[23]);
  BUFF I164 (w1_0n[24], inpA_0a1d[24]);
  BUFF I165 (w1_0n[25], inpA_0a1d[25]);
  BUFF I166 (w1_0n[26], inpA_0a1d[26]);
  BUFF I167 (w1_0n[27], inpA_0a1d[27]);
  BUFF I168 (w1_0n[28], inpA_0a1d[28]);
  BUFF I169 (w1_0n[29], inpA_0a1d[29]);
  BUFF I170 (w1_0n[30], inpA_0a1d[30]);
  BUFF I171 (w1_0n[31], inpA_0a1d[31]);
  BUFF I172 (w1_0n[32], inpA_0a1d[32]);
  BUFF I173 (w1_0n[33], inpA_0a1d[33]);
  BUFF I174 (w1_0n[34], inpA_0a1d[34]);
  BUFF I175 (inpA_0r, out_0r);
  BUFF I176 (inpB_0r, out_0r);
endmodule

module DROR2 (
  i0_0,
  i0_1,
  i1_0,
  i1_1,
  q_0,
  q_1
);
  input i0_0;
  input i0_1;
  input i1_0;
  input i1_1;
  output q_0;
  output q_1;
  wire n0_0n;
  wire n1_0n;
  wire n2_0n;
  C2 I0 (q_0, i0_0, i1_0);
  OR3 I1 (q_1, n0_0n, n1_0n, n2_0n);
  C2 I2 (n2_0n, i0_1, i1_1);
  C2 I3 (n1_0n, i0_1, i1_0);
  C2 I4 (n0_0n, i0_0, i1_1);
endmodule

module BrzBinaryFunc_35_35_35_s2_Or_s5_false_s5_f_m21m (
  out_0r, out_0a0d, out_0a1d,
  inpA_0r, inpA_0a0d, inpA_0a1d,
  inpB_0r, inpB_0a0d, inpB_0a1d
);
  input out_0r;
  output [34:0] out_0a0d;
  output [34:0] out_0a1d;
  output inpA_0r;
  input [34:0] inpA_0a0d;
  input [34:0] inpA_0a1d;
  output inpB_0r;
  input [34:0] inpB_0a0d;
  input [34:0] inpB_0a1d;
  wire [34:0] n1_0n;
  wire [34:0] n0_0n;
  wire [34:0] w1_0n;
  wire [34:0] w0_0n;
  DROR2 I0 (n0_0n[0], n1_0n[0], w0_0n[0], w1_0n[0], out_0a0d[0], out_0a1d[0]);
  DROR2 I1 (n0_0n[1], n1_0n[1], w0_0n[1], w1_0n[1], out_0a0d[1], out_0a1d[1]);
  DROR2 I2 (n0_0n[2], n1_0n[2], w0_0n[2], w1_0n[2], out_0a0d[2], out_0a1d[2]);
  DROR2 I3 (n0_0n[3], n1_0n[3], w0_0n[3], w1_0n[3], out_0a0d[3], out_0a1d[3]);
  DROR2 I4 (n0_0n[4], n1_0n[4], w0_0n[4], w1_0n[4], out_0a0d[4], out_0a1d[4]);
  DROR2 I5 (n0_0n[5], n1_0n[5], w0_0n[5], w1_0n[5], out_0a0d[5], out_0a1d[5]);
  DROR2 I6 (n0_0n[6], n1_0n[6], w0_0n[6], w1_0n[6], out_0a0d[6], out_0a1d[6]);
  DROR2 I7 (n0_0n[7], n1_0n[7], w0_0n[7], w1_0n[7], out_0a0d[7], out_0a1d[7]);
  DROR2 I8 (n0_0n[8], n1_0n[8], w0_0n[8], w1_0n[8], out_0a0d[8], out_0a1d[8]);
  DROR2 I9 (n0_0n[9], n1_0n[9], w0_0n[9], w1_0n[9], out_0a0d[9], out_0a1d[9]);
  DROR2 I10 (n0_0n[10], n1_0n[10], w0_0n[10], w1_0n[10], out_0a0d[10], out_0a1d[10]);
  DROR2 I11 (n0_0n[11], n1_0n[11], w0_0n[11], w1_0n[11], out_0a0d[11], out_0a1d[11]);
  DROR2 I12 (n0_0n[12], n1_0n[12], w0_0n[12], w1_0n[12], out_0a0d[12], out_0a1d[12]);
  DROR2 I13 (n0_0n[13], n1_0n[13], w0_0n[13], w1_0n[13], out_0a0d[13], out_0a1d[13]);
  DROR2 I14 (n0_0n[14], n1_0n[14], w0_0n[14], w1_0n[14], out_0a0d[14], out_0a1d[14]);
  DROR2 I15 (n0_0n[15], n1_0n[15], w0_0n[15], w1_0n[15], out_0a0d[15], out_0a1d[15]);
  DROR2 I16 (n0_0n[16], n1_0n[16], w0_0n[16], w1_0n[16], out_0a0d[16], out_0a1d[16]);
  DROR2 I17 (n0_0n[17], n1_0n[17], w0_0n[17], w1_0n[17], out_0a0d[17], out_0a1d[17]);
  DROR2 I18 (n0_0n[18], n1_0n[18], w0_0n[18], w1_0n[18], out_0a0d[18], out_0a1d[18]);
  DROR2 I19 (n0_0n[19], n1_0n[19], w0_0n[19], w1_0n[19], out_0a0d[19], out_0a1d[19]);
  DROR2 I20 (n0_0n[20], n1_0n[20], w0_0n[20], w1_0n[20], out_0a0d[20], out_0a1d[20]);
  DROR2 I21 (n0_0n[21], n1_0n[21], w0_0n[21], w1_0n[21], out_0a0d[21], out_0a1d[21]);
  DROR2 I22 (n0_0n[22], n1_0n[22], w0_0n[22], w1_0n[22], out_0a0d[22], out_0a1d[22]);
  DROR2 I23 (n0_0n[23], n1_0n[23], w0_0n[23], w1_0n[23], out_0a0d[23], out_0a1d[23]);
  DROR2 I24 (n0_0n[24], n1_0n[24], w0_0n[24], w1_0n[24], out_0a0d[24], out_0a1d[24]);
  DROR2 I25 (n0_0n[25], n1_0n[25], w0_0n[25], w1_0n[25], out_0a0d[25], out_0a1d[25]);
  DROR2 I26 (n0_0n[26], n1_0n[26], w0_0n[26], w1_0n[26], out_0a0d[26], out_0a1d[26]);
  DROR2 I27 (n0_0n[27], n1_0n[27], w0_0n[27], w1_0n[27], out_0a0d[27], out_0a1d[27]);
  DROR2 I28 (n0_0n[28], n1_0n[28], w0_0n[28], w1_0n[28], out_0a0d[28], out_0a1d[28]);
  DROR2 I29 (n0_0n[29], n1_0n[29], w0_0n[29], w1_0n[29], out_0a0d[29], out_0a1d[29]);
  DROR2 I30 (n0_0n[30], n1_0n[30], w0_0n[30], w1_0n[30], out_0a0d[30], out_0a1d[30]);
  DROR2 I31 (n0_0n[31], n1_0n[31], w0_0n[31], w1_0n[31], out_0a0d[31], out_0a1d[31]);
  DROR2 I32 (n0_0n[32], n1_0n[32], w0_0n[32], w1_0n[32], out_0a0d[32], out_0a1d[32]);
  DROR2 I33 (n0_0n[33], n1_0n[33], w0_0n[33], w1_0n[33], out_0a0d[33], out_0a1d[33]);
  DROR2 I34 (n0_0n[34], n1_0n[34], w0_0n[34], w1_0n[34], out_0a0d[34], out_0a1d[34]);
  BUFF I35 (n0_0n[0], inpB_0a0d[0]);
  BUFF I36 (n0_0n[1], inpB_0a0d[1]);
  BUFF I37 (n0_0n[2], inpB_0a0d[2]);
  BUFF I38 (n0_0n[3], inpB_0a0d[3]);
  BUFF I39 (n0_0n[4], inpB_0a0d[4]);
  BUFF I40 (n0_0n[5], inpB_0a0d[5]);
  BUFF I41 (n0_0n[6], inpB_0a0d[6]);
  BUFF I42 (n0_0n[7], inpB_0a0d[7]);
  BUFF I43 (n0_0n[8], inpB_0a0d[8]);
  BUFF I44 (n0_0n[9], inpB_0a0d[9]);
  BUFF I45 (n0_0n[10], inpB_0a0d[10]);
  BUFF I46 (n0_0n[11], inpB_0a0d[11]);
  BUFF I47 (n0_0n[12], inpB_0a0d[12]);
  BUFF I48 (n0_0n[13], inpB_0a0d[13]);
  BUFF I49 (n0_0n[14], inpB_0a0d[14]);
  BUFF I50 (n0_0n[15], inpB_0a0d[15]);
  BUFF I51 (n0_0n[16], inpB_0a0d[16]);
  BUFF I52 (n0_0n[17], inpB_0a0d[17]);
  BUFF I53 (n0_0n[18], inpB_0a0d[18]);
  BUFF I54 (n0_0n[19], inpB_0a0d[19]);
  BUFF I55 (n0_0n[20], inpB_0a0d[20]);
  BUFF I56 (n0_0n[21], inpB_0a0d[21]);
  BUFF I57 (n0_0n[22], inpB_0a0d[22]);
  BUFF I58 (n0_0n[23], inpB_0a0d[23]);
  BUFF I59 (n0_0n[24], inpB_0a0d[24]);
  BUFF I60 (n0_0n[25], inpB_0a0d[25]);
  BUFF I61 (n0_0n[26], inpB_0a0d[26]);
  BUFF I62 (n0_0n[27], inpB_0a0d[27]);
  BUFF I63 (n0_0n[28], inpB_0a0d[28]);
  BUFF I64 (n0_0n[29], inpB_0a0d[29]);
  BUFF I65 (n0_0n[30], inpB_0a0d[30]);
  BUFF I66 (n0_0n[31], inpB_0a0d[31]);
  BUFF I67 (n0_0n[32], inpB_0a0d[32]);
  BUFF I68 (n0_0n[33], inpB_0a0d[33]);
  BUFF I69 (n0_0n[34], inpB_0a0d[34]);
  BUFF I70 (n1_0n[0], inpB_0a1d[0]);
  BUFF I71 (n1_0n[1], inpB_0a1d[1]);
  BUFF I72 (n1_0n[2], inpB_0a1d[2]);
  BUFF I73 (n1_0n[3], inpB_0a1d[3]);
  BUFF I74 (n1_0n[4], inpB_0a1d[4]);
  BUFF I75 (n1_0n[5], inpB_0a1d[5]);
  BUFF I76 (n1_0n[6], inpB_0a1d[6]);
  BUFF I77 (n1_0n[7], inpB_0a1d[7]);
  BUFF I78 (n1_0n[8], inpB_0a1d[8]);
  BUFF I79 (n1_0n[9], inpB_0a1d[9]);
  BUFF I80 (n1_0n[10], inpB_0a1d[10]);
  BUFF I81 (n1_0n[11], inpB_0a1d[11]);
  BUFF I82 (n1_0n[12], inpB_0a1d[12]);
  BUFF I83 (n1_0n[13], inpB_0a1d[13]);
  BUFF I84 (n1_0n[14], inpB_0a1d[14]);
  BUFF I85 (n1_0n[15], inpB_0a1d[15]);
  BUFF I86 (n1_0n[16], inpB_0a1d[16]);
  BUFF I87 (n1_0n[17], inpB_0a1d[17]);
  BUFF I88 (n1_0n[18], inpB_0a1d[18]);
  BUFF I89 (n1_0n[19], inpB_0a1d[19]);
  BUFF I90 (n1_0n[20], inpB_0a1d[20]);
  BUFF I91 (n1_0n[21], inpB_0a1d[21]);
  BUFF I92 (n1_0n[22], inpB_0a1d[22]);
  BUFF I93 (n1_0n[23], inpB_0a1d[23]);
  BUFF I94 (n1_0n[24], inpB_0a1d[24]);
  BUFF I95 (n1_0n[25], inpB_0a1d[25]);
  BUFF I96 (n1_0n[26], inpB_0a1d[26]);
  BUFF I97 (n1_0n[27], inpB_0a1d[27]);
  BUFF I98 (n1_0n[28], inpB_0a1d[28]);
  BUFF I99 (n1_0n[29], inpB_0a1d[29]);
  BUFF I100 (n1_0n[30], inpB_0a1d[30]);
  BUFF I101 (n1_0n[31], inpB_0a1d[31]);
  BUFF I102 (n1_0n[32], inpB_0a1d[32]);
  BUFF I103 (n1_0n[33], inpB_0a1d[33]);
  BUFF I104 (n1_0n[34], inpB_0a1d[34]);
  BUFF I105 (w0_0n[0], inpA_0a0d[0]);
  BUFF I106 (w0_0n[1], inpA_0a0d[1]);
  BUFF I107 (w0_0n[2], inpA_0a0d[2]);
  BUFF I108 (w0_0n[3], inpA_0a0d[3]);
  BUFF I109 (w0_0n[4], inpA_0a0d[4]);
  BUFF I110 (w0_0n[5], inpA_0a0d[5]);
  BUFF I111 (w0_0n[6], inpA_0a0d[6]);
  BUFF I112 (w0_0n[7], inpA_0a0d[7]);
  BUFF I113 (w0_0n[8], inpA_0a0d[8]);
  BUFF I114 (w0_0n[9], inpA_0a0d[9]);
  BUFF I115 (w0_0n[10], inpA_0a0d[10]);
  BUFF I116 (w0_0n[11], inpA_0a0d[11]);
  BUFF I117 (w0_0n[12], inpA_0a0d[12]);
  BUFF I118 (w0_0n[13], inpA_0a0d[13]);
  BUFF I119 (w0_0n[14], inpA_0a0d[14]);
  BUFF I120 (w0_0n[15], inpA_0a0d[15]);
  BUFF I121 (w0_0n[16], inpA_0a0d[16]);
  BUFF I122 (w0_0n[17], inpA_0a0d[17]);
  BUFF I123 (w0_0n[18], inpA_0a0d[18]);
  BUFF I124 (w0_0n[19], inpA_0a0d[19]);
  BUFF I125 (w0_0n[20], inpA_0a0d[20]);
  BUFF I126 (w0_0n[21], inpA_0a0d[21]);
  BUFF I127 (w0_0n[22], inpA_0a0d[22]);
  BUFF I128 (w0_0n[23], inpA_0a0d[23]);
  BUFF I129 (w0_0n[24], inpA_0a0d[24]);
  BUFF I130 (w0_0n[25], inpA_0a0d[25]);
  BUFF I131 (w0_0n[26], inpA_0a0d[26]);
  BUFF I132 (w0_0n[27], inpA_0a0d[27]);
  BUFF I133 (w0_0n[28], inpA_0a0d[28]);
  BUFF I134 (w0_0n[29], inpA_0a0d[29]);
  BUFF I135 (w0_0n[30], inpA_0a0d[30]);
  BUFF I136 (w0_0n[31], inpA_0a0d[31]);
  BUFF I137 (w0_0n[32], inpA_0a0d[32]);
  BUFF I138 (w0_0n[33], inpA_0a0d[33]);
  BUFF I139 (w0_0n[34], inpA_0a0d[34]);
  BUFF I140 (w1_0n[0], inpA_0a1d[0]);
  BUFF I141 (w1_0n[1], inpA_0a1d[1]);
  BUFF I142 (w1_0n[2], inpA_0a1d[2]);
  BUFF I143 (w1_0n[3], inpA_0a1d[3]);
  BUFF I144 (w1_0n[4], inpA_0a1d[4]);
  BUFF I145 (w1_0n[5], inpA_0a1d[5]);
  BUFF I146 (w1_0n[6], inpA_0a1d[6]);
  BUFF I147 (w1_0n[7], inpA_0a1d[7]);
  BUFF I148 (w1_0n[8], inpA_0a1d[8]);
  BUFF I149 (w1_0n[9], inpA_0a1d[9]);
  BUFF I150 (w1_0n[10], inpA_0a1d[10]);
  BUFF I151 (w1_0n[11], inpA_0a1d[11]);
  BUFF I152 (w1_0n[12], inpA_0a1d[12]);
  BUFF I153 (w1_0n[13], inpA_0a1d[13]);
  BUFF I154 (w1_0n[14], inpA_0a1d[14]);
  BUFF I155 (w1_0n[15], inpA_0a1d[15]);
  BUFF I156 (w1_0n[16], inpA_0a1d[16]);
  BUFF I157 (w1_0n[17], inpA_0a1d[17]);
  BUFF I158 (w1_0n[18], inpA_0a1d[18]);
  BUFF I159 (w1_0n[19], inpA_0a1d[19]);
  BUFF I160 (w1_0n[20], inpA_0a1d[20]);
  BUFF I161 (w1_0n[21], inpA_0a1d[21]);
  BUFF I162 (w1_0n[22], inpA_0a1d[22]);
  BUFF I163 (w1_0n[23], inpA_0a1d[23]);
  BUFF I164 (w1_0n[24], inpA_0a1d[24]);
  BUFF I165 (w1_0n[25], inpA_0a1d[25]);
  BUFF I166 (w1_0n[26], inpA_0a1d[26]);
  BUFF I167 (w1_0n[27], inpA_0a1d[27]);
  BUFF I168 (w1_0n[28], inpA_0a1d[28]);
  BUFF I169 (w1_0n[29], inpA_0a1d[29]);
  BUFF I170 (w1_0n[30], inpA_0a1d[30]);
  BUFF I171 (w1_0n[31], inpA_0a1d[31]);
  BUFF I172 (w1_0n[32], inpA_0a1d[32]);
  BUFF I173 (w1_0n[33], inpA_0a1d[33]);
  BUFF I174 (w1_0n[34], inpA_0a1d[34]);
  BUFF I175 (inpA_0r, out_0r);
  BUFF I176 (inpB_0r, out_0r);
endmodule

module DRXOR2 (
  i0_0,
  i0_1,
  i1_0,
  i1_1,
  q_0,
  q_1
);
  input i0_0;
  input i0_1;
  input i1_0;
  input i1_1;
  output q_0;
  output q_1;
  wire n0_0n;
  wire n1_0n;
  wire n2_0n;
  wire n3_0n;
  OR2 I0 (q_0, n0_0n, n3_0n);
  C2 I1 (n3_0n, i0_1, i1_1);
  C2 I2 (n0_0n, i0_0, i1_0);
  OR2 I3 (q_1, n1_0n, n2_0n);
  C2 I4 (n1_0n, i0_0, i1_1);
  C2 I5 (n2_0n, i0_1, i1_0);
endmodule

module BrzBinaryFunc_35_35_35_s3_Xor_s5_false_s5__m23m (
  out_0r, out_0a0d, out_0a1d,
  inpA_0r, inpA_0a0d, inpA_0a1d,
  inpB_0r, inpB_0a0d, inpB_0a1d
);
  input out_0r;
  output [34:0] out_0a0d;
  output [34:0] out_0a1d;
  output inpA_0r;
  input [34:0] inpA_0a0d;
  input [34:0] inpA_0a1d;
  output inpB_0r;
  input [34:0] inpB_0a0d;
  input [34:0] inpB_0a1d;
  wire [34:0] n1_0n;
  wire [34:0] n0_0n;
  wire [34:0] w1_0n;
  wire [34:0] w0_0n;
  DRXOR2 I0 (n0_0n[0], n1_0n[0], w0_0n[0], w1_0n[0], out_0a0d[0], out_0a1d[0]);
  DRXOR2 I1 (n0_0n[1], n1_0n[1], w0_0n[1], w1_0n[1], out_0a0d[1], out_0a1d[1]);
  DRXOR2 I2 (n0_0n[2], n1_0n[2], w0_0n[2], w1_0n[2], out_0a0d[2], out_0a1d[2]);
  DRXOR2 I3 (n0_0n[3], n1_0n[3], w0_0n[3], w1_0n[3], out_0a0d[3], out_0a1d[3]);
  DRXOR2 I4 (n0_0n[4], n1_0n[4], w0_0n[4], w1_0n[4], out_0a0d[4], out_0a1d[4]);
  DRXOR2 I5 (n0_0n[5], n1_0n[5], w0_0n[5], w1_0n[5], out_0a0d[5], out_0a1d[5]);
  DRXOR2 I6 (n0_0n[6], n1_0n[6], w0_0n[6], w1_0n[6], out_0a0d[6], out_0a1d[6]);
  DRXOR2 I7 (n0_0n[7], n1_0n[7], w0_0n[7], w1_0n[7], out_0a0d[7], out_0a1d[7]);
  DRXOR2 I8 (n0_0n[8], n1_0n[8], w0_0n[8], w1_0n[8], out_0a0d[8], out_0a1d[8]);
  DRXOR2 I9 (n0_0n[9], n1_0n[9], w0_0n[9], w1_0n[9], out_0a0d[9], out_0a1d[9]);
  DRXOR2 I10 (n0_0n[10], n1_0n[10], w0_0n[10], w1_0n[10], out_0a0d[10], out_0a1d[10]);
  DRXOR2 I11 (n0_0n[11], n1_0n[11], w0_0n[11], w1_0n[11], out_0a0d[11], out_0a1d[11]);
  DRXOR2 I12 (n0_0n[12], n1_0n[12], w0_0n[12], w1_0n[12], out_0a0d[12], out_0a1d[12]);
  DRXOR2 I13 (n0_0n[13], n1_0n[13], w0_0n[13], w1_0n[13], out_0a0d[13], out_0a1d[13]);
  DRXOR2 I14 (n0_0n[14], n1_0n[14], w0_0n[14], w1_0n[14], out_0a0d[14], out_0a1d[14]);
  DRXOR2 I15 (n0_0n[15], n1_0n[15], w0_0n[15], w1_0n[15], out_0a0d[15], out_0a1d[15]);
  DRXOR2 I16 (n0_0n[16], n1_0n[16], w0_0n[16], w1_0n[16], out_0a0d[16], out_0a1d[16]);
  DRXOR2 I17 (n0_0n[17], n1_0n[17], w0_0n[17], w1_0n[17], out_0a0d[17], out_0a1d[17]);
  DRXOR2 I18 (n0_0n[18], n1_0n[18], w0_0n[18], w1_0n[18], out_0a0d[18], out_0a1d[18]);
  DRXOR2 I19 (n0_0n[19], n1_0n[19], w0_0n[19], w1_0n[19], out_0a0d[19], out_0a1d[19]);
  DRXOR2 I20 (n0_0n[20], n1_0n[20], w0_0n[20], w1_0n[20], out_0a0d[20], out_0a1d[20]);
  DRXOR2 I21 (n0_0n[21], n1_0n[21], w0_0n[21], w1_0n[21], out_0a0d[21], out_0a1d[21]);
  DRXOR2 I22 (n0_0n[22], n1_0n[22], w0_0n[22], w1_0n[22], out_0a0d[22], out_0a1d[22]);
  DRXOR2 I23 (n0_0n[23], n1_0n[23], w0_0n[23], w1_0n[23], out_0a0d[23], out_0a1d[23]);
  DRXOR2 I24 (n0_0n[24], n1_0n[24], w0_0n[24], w1_0n[24], out_0a0d[24], out_0a1d[24]);
  DRXOR2 I25 (n0_0n[25], n1_0n[25], w0_0n[25], w1_0n[25], out_0a0d[25], out_0a1d[25]);
  DRXOR2 I26 (n0_0n[26], n1_0n[26], w0_0n[26], w1_0n[26], out_0a0d[26], out_0a1d[26]);
  DRXOR2 I27 (n0_0n[27], n1_0n[27], w0_0n[27], w1_0n[27], out_0a0d[27], out_0a1d[27]);
  DRXOR2 I28 (n0_0n[28], n1_0n[28], w0_0n[28], w1_0n[28], out_0a0d[28], out_0a1d[28]);
  DRXOR2 I29 (n0_0n[29], n1_0n[29], w0_0n[29], w1_0n[29], out_0a0d[29], out_0a1d[29]);
  DRXOR2 I30 (n0_0n[30], n1_0n[30], w0_0n[30], w1_0n[30], out_0a0d[30], out_0a1d[30]);
  DRXOR2 I31 (n0_0n[31], n1_0n[31], w0_0n[31], w1_0n[31], out_0a0d[31], out_0a1d[31]);
  DRXOR2 I32 (n0_0n[32], n1_0n[32], w0_0n[32], w1_0n[32], out_0a0d[32], out_0a1d[32]);
  DRXOR2 I33 (n0_0n[33], n1_0n[33], w0_0n[33], w1_0n[33], out_0a0d[33], out_0a1d[33]);
  DRXOR2 I34 (n0_0n[34], n1_0n[34], w0_0n[34], w1_0n[34], out_0a0d[34], out_0a1d[34]);
  BUFF I35 (n0_0n[0], inpB_0a0d[0]);
  BUFF I36 (n0_0n[1], inpB_0a0d[1]);
  BUFF I37 (n0_0n[2], inpB_0a0d[2]);
  BUFF I38 (n0_0n[3], inpB_0a0d[3]);
  BUFF I39 (n0_0n[4], inpB_0a0d[4]);
  BUFF I40 (n0_0n[5], inpB_0a0d[5]);
  BUFF I41 (n0_0n[6], inpB_0a0d[6]);
  BUFF I42 (n0_0n[7], inpB_0a0d[7]);
  BUFF I43 (n0_0n[8], inpB_0a0d[8]);
  BUFF I44 (n0_0n[9], inpB_0a0d[9]);
  BUFF I45 (n0_0n[10], inpB_0a0d[10]);
  BUFF I46 (n0_0n[11], inpB_0a0d[11]);
  BUFF I47 (n0_0n[12], inpB_0a0d[12]);
  BUFF I48 (n0_0n[13], inpB_0a0d[13]);
  BUFF I49 (n0_0n[14], inpB_0a0d[14]);
  BUFF I50 (n0_0n[15], inpB_0a0d[15]);
  BUFF I51 (n0_0n[16], inpB_0a0d[16]);
  BUFF I52 (n0_0n[17], inpB_0a0d[17]);
  BUFF I53 (n0_0n[18], inpB_0a0d[18]);
  BUFF I54 (n0_0n[19], inpB_0a0d[19]);
  BUFF I55 (n0_0n[20], inpB_0a0d[20]);
  BUFF I56 (n0_0n[21], inpB_0a0d[21]);
  BUFF I57 (n0_0n[22], inpB_0a0d[22]);
  BUFF I58 (n0_0n[23], inpB_0a0d[23]);
  BUFF I59 (n0_0n[24], inpB_0a0d[24]);
  BUFF I60 (n0_0n[25], inpB_0a0d[25]);
  BUFF I61 (n0_0n[26], inpB_0a0d[26]);
  BUFF I62 (n0_0n[27], inpB_0a0d[27]);
  BUFF I63 (n0_0n[28], inpB_0a0d[28]);
  BUFF I64 (n0_0n[29], inpB_0a0d[29]);
  BUFF I65 (n0_0n[30], inpB_0a0d[30]);
  BUFF I66 (n0_0n[31], inpB_0a0d[31]);
  BUFF I67 (n0_0n[32], inpB_0a0d[32]);
  BUFF I68 (n0_0n[33], inpB_0a0d[33]);
  BUFF I69 (n0_0n[34], inpB_0a0d[34]);
  BUFF I70 (n1_0n[0], inpB_0a1d[0]);
  BUFF I71 (n1_0n[1], inpB_0a1d[1]);
  BUFF I72 (n1_0n[2], inpB_0a1d[2]);
  BUFF I73 (n1_0n[3], inpB_0a1d[3]);
  BUFF I74 (n1_0n[4], inpB_0a1d[4]);
  BUFF I75 (n1_0n[5], inpB_0a1d[5]);
  BUFF I76 (n1_0n[6], inpB_0a1d[6]);
  BUFF I77 (n1_0n[7], inpB_0a1d[7]);
  BUFF I78 (n1_0n[8], inpB_0a1d[8]);
  BUFF I79 (n1_0n[9], inpB_0a1d[9]);
  BUFF I80 (n1_0n[10], inpB_0a1d[10]);
  BUFF I81 (n1_0n[11], inpB_0a1d[11]);
  BUFF I82 (n1_0n[12], inpB_0a1d[12]);
  BUFF I83 (n1_0n[13], inpB_0a1d[13]);
  BUFF I84 (n1_0n[14], inpB_0a1d[14]);
  BUFF I85 (n1_0n[15], inpB_0a1d[15]);
  BUFF I86 (n1_0n[16], inpB_0a1d[16]);
  BUFF I87 (n1_0n[17], inpB_0a1d[17]);
  BUFF I88 (n1_0n[18], inpB_0a1d[18]);
  BUFF I89 (n1_0n[19], inpB_0a1d[19]);
  BUFF I90 (n1_0n[20], inpB_0a1d[20]);
  BUFF I91 (n1_0n[21], inpB_0a1d[21]);
  BUFF I92 (n1_0n[22], inpB_0a1d[22]);
  BUFF I93 (n1_0n[23], inpB_0a1d[23]);
  BUFF I94 (n1_0n[24], inpB_0a1d[24]);
  BUFF I95 (n1_0n[25], inpB_0a1d[25]);
  BUFF I96 (n1_0n[26], inpB_0a1d[26]);
  BUFF I97 (n1_0n[27], inpB_0a1d[27]);
  BUFF I98 (n1_0n[28], inpB_0a1d[28]);
  BUFF I99 (n1_0n[29], inpB_0a1d[29]);
  BUFF I100 (n1_0n[30], inpB_0a1d[30]);
  BUFF I101 (n1_0n[31], inpB_0a1d[31]);
  BUFF I102 (n1_0n[32], inpB_0a1d[32]);
  BUFF I103 (n1_0n[33], inpB_0a1d[33]);
  BUFF I104 (n1_0n[34], inpB_0a1d[34]);
  BUFF I105 (w0_0n[0], inpA_0a0d[0]);
  BUFF I106 (w0_0n[1], inpA_0a0d[1]);
  BUFF I107 (w0_0n[2], inpA_0a0d[2]);
  BUFF I108 (w0_0n[3], inpA_0a0d[3]);
  BUFF I109 (w0_0n[4], inpA_0a0d[4]);
  BUFF I110 (w0_0n[5], inpA_0a0d[5]);
  BUFF I111 (w0_0n[6], inpA_0a0d[6]);
  BUFF I112 (w0_0n[7], inpA_0a0d[7]);
  BUFF I113 (w0_0n[8], inpA_0a0d[8]);
  BUFF I114 (w0_0n[9], inpA_0a0d[9]);
  BUFF I115 (w0_0n[10], inpA_0a0d[10]);
  BUFF I116 (w0_0n[11], inpA_0a0d[11]);
  BUFF I117 (w0_0n[12], inpA_0a0d[12]);
  BUFF I118 (w0_0n[13], inpA_0a0d[13]);
  BUFF I119 (w0_0n[14], inpA_0a0d[14]);
  BUFF I120 (w0_0n[15], inpA_0a0d[15]);
  BUFF I121 (w0_0n[16], inpA_0a0d[16]);
  BUFF I122 (w0_0n[17], inpA_0a0d[17]);
  BUFF I123 (w0_0n[18], inpA_0a0d[18]);
  BUFF I124 (w0_0n[19], inpA_0a0d[19]);
  BUFF I125 (w0_0n[20], inpA_0a0d[20]);
  BUFF I126 (w0_0n[21], inpA_0a0d[21]);
  BUFF I127 (w0_0n[22], inpA_0a0d[22]);
  BUFF I128 (w0_0n[23], inpA_0a0d[23]);
  BUFF I129 (w0_0n[24], inpA_0a0d[24]);
  BUFF I130 (w0_0n[25], inpA_0a0d[25]);
  BUFF I131 (w0_0n[26], inpA_0a0d[26]);
  BUFF I132 (w0_0n[27], inpA_0a0d[27]);
  BUFF I133 (w0_0n[28], inpA_0a0d[28]);
  BUFF I134 (w0_0n[29], inpA_0a0d[29]);
  BUFF I135 (w0_0n[30], inpA_0a0d[30]);
  BUFF I136 (w0_0n[31], inpA_0a0d[31]);
  BUFF I137 (w0_0n[32], inpA_0a0d[32]);
  BUFF I138 (w0_0n[33], inpA_0a0d[33]);
  BUFF I139 (w0_0n[34], inpA_0a0d[34]);
  BUFF I140 (w1_0n[0], inpA_0a1d[0]);
  BUFF I141 (w1_0n[1], inpA_0a1d[1]);
  BUFF I142 (w1_0n[2], inpA_0a1d[2]);
  BUFF I143 (w1_0n[3], inpA_0a1d[3]);
  BUFF I144 (w1_0n[4], inpA_0a1d[4]);
  BUFF I145 (w1_0n[5], inpA_0a1d[5]);
  BUFF I146 (w1_0n[6], inpA_0a1d[6]);
  BUFF I147 (w1_0n[7], inpA_0a1d[7]);
  BUFF I148 (w1_0n[8], inpA_0a1d[8]);
  BUFF I149 (w1_0n[9], inpA_0a1d[9]);
  BUFF I150 (w1_0n[10], inpA_0a1d[10]);
  BUFF I151 (w1_0n[11], inpA_0a1d[11]);
  BUFF I152 (w1_0n[12], inpA_0a1d[12]);
  BUFF I153 (w1_0n[13], inpA_0a1d[13]);
  BUFF I154 (w1_0n[14], inpA_0a1d[14]);
  BUFF I155 (w1_0n[15], inpA_0a1d[15]);
  BUFF I156 (w1_0n[16], inpA_0a1d[16]);
  BUFF I157 (w1_0n[17], inpA_0a1d[17]);
  BUFF I158 (w1_0n[18], inpA_0a1d[18]);
  BUFF I159 (w1_0n[19], inpA_0a1d[19]);
  BUFF I160 (w1_0n[20], inpA_0a1d[20]);
  BUFF I161 (w1_0n[21], inpA_0a1d[21]);
  BUFF I162 (w1_0n[22], inpA_0a1d[22]);
  BUFF I163 (w1_0n[23], inpA_0a1d[23]);
  BUFF I164 (w1_0n[24], inpA_0a1d[24]);
  BUFF I165 (w1_0n[25], inpA_0a1d[25]);
  BUFF I166 (w1_0n[26], inpA_0a1d[26]);
  BUFF I167 (w1_0n[27], inpA_0a1d[27]);
  BUFF I168 (w1_0n[28], inpA_0a1d[28]);
  BUFF I169 (w1_0n[29], inpA_0a1d[29]);
  BUFF I170 (w1_0n[30], inpA_0a1d[30]);
  BUFF I171 (w1_0n[31], inpA_0a1d[31]);
  BUFF I172 (w1_0n[32], inpA_0a1d[32]);
  BUFF I173 (w1_0n[33], inpA_0a1d[33]);
  BUFF I174 (w1_0n[34], inpA_0a1d[34]);
  BUFF I175 (inpA_0r, out_0r);
  BUFF I176 (inpB_0r, out_0r);
endmodule

module BrzBinaryFuncConstR_1_32_1_s6_Equals_s5_fa_m25m (
  out_0r, out_0a0d, out_0a1d,
  inpA_0r, inpA_0a0d, inpA_0a1d
);
  input out_0r;
  output out_0a0d;
  output out_0a1d;
  output inpA_0r;
  input [31:0] inpA_0a0d;
  input [31:0] inpA_0a1d;
  wire [31:0] compOut1_0n;
  wire [31:0] compOut0_0n;
  wire [30:0] internalA1_0n;
  wire [30:0] internalA0_0n;
  BUFF I0 (out_0a0d, internalA1_0n[0]);
  BUFF I1 (out_0a1d, internalA0_0n[0]);
  DROR2 I2 (compOut0_0n[30], compOut1_0n[30], compOut0_0n[31], compOut1_0n[31], internalA0_0n[30], internalA1_0n[30]);
  DROR2 I3 (compOut0_0n[28], compOut1_0n[28], compOut0_0n[29], compOut1_0n[29], internalA0_0n[29], internalA1_0n[29]);
  DROR2 I4 (internalA0_0n[29], internalA1_0n[29], internalA0_0n[30], internalA1_0n[30], internalA0_0n[28], internalA1_0n[28]);
  DROR2 I5 (compOut0_0n[26], compOut1_0n[26], compOut0_0n[27], compOut1_0n[27], internalA0_0n[27], internalA1_0n[27]);
  DROR2 I6 (compOut0_0n[24], compOut1_0n[24], compOut0_0n[25], compOut1_0n[25], internalA0_0n[26], internalA1_0n[26]);
  DROR2 I7 (internalA0_0n[26], internalA1_0n[26], internalA0_0n[27], internalA1_0n[27], internalA0_0n[25], internalA1_0n[25]);
  DROR2 I8 (internalA0_0n[25], internalA1_0n[25], internalA0_0n[28], internalA1_0n[28], internalA0_0n[24], internalA1_0n[24]);
  DROR2 I9 (compOut0_0n[22], compOut1_0n[22], compOut0_0n[23], compOut1_0n[23], internalA0_0n[23], internalA1_0n[23]);
  DROR2 I10 (compOut0_0n[20], compOut1_0n[20], compOut0_0n[21], compOut1_0n[21], internalA0_0n[22], internalA1_0n[22]);
  DROR2 I11 (internalA0_0n[22], internalA1_0n[22], internalA0_0n[23], internalA1_0n[23], internalA0_0n[21], internalA1_0n[21]);
  DROR2 I12 (compOut0_0n[18], compOut1_0n[18], compOut0_0n[19], compOut1_0n[19], internalA0_0n[20], internalA1_0n[20]);
  DROR2 I13 (compOut0_0n[16], compOut1_0n[16], compOut0_0n[17], compOut1_0n[17], internalA0_0n[19], internalA1_0n[19]);
  DROR2 I14 (internalA0_0n[19], internalA1_0n[19], internalA0_0n[20], internalA1_0n[20], internalA0_0n[18], internalA1_0n[18]);
  DROR2 I15 (internalA0_0n[18], internalA1_0n[18], internalA0_0n[21], internalA1_0n[21], internalA0_0n[17], internalA1_0n[17]);
  DROR2 I16 (internalA0_0n[17], internalA1_0n[17], internalA0_0n[24], internalA1_0n[24], internalA0_0n[16], internalA1_0n[16]);
  DROR2 I17 (compOut0_0n[14], compOut1_0n[14], compOut0_0n[15], compOut1_0n[15], internalA0_0n[15], internalA1_0n[15]);
  DROR2 I18 (compOut0_0n[12], compOut1_0n[12], compOut0_0n[13], compOut1_0n[13], internalA0_0n[14], internalA1_0n[14]);
  DROR2 I19 (internalA0_0n[14], internalA1_0n[14], internalA0_0n[15], internalA1_0n[15], internalA0_0n[13], internalA1_0n[13]);
  DROR2 I20 (compOut0_0n[10], compOut1_0n[10], compOut0_0n[11], compOut1_0n[11], internalA0_0n[12], internalA1_0n[12]);
  DROR2 I21 (compOut0_0n[8], compOut1_0n[8], compOut0_0n[9], compOut1_0n[9], internalA0_0n[11], internalA1_0n[11]);
  DROR2 I22 (internalA0_0n[11], internalA1_0n[11], internalA0_0n[12], internalA1_0n[12], internalA0_0n[10], internalA1_0n[10]);
  DROR2 I23 (internalA0_0n[10], internalA1_0n[10], internalA0_0n[13], internalA1_0n[13], internalA0_0n[9], internalA1_0n[9]);
  DROR2 I24 (compOut0_0n[6], compOut1_0n[6], compOut0_0n[7], compOut1_0n[7], internalA0_0n[8], internalA1_0n[8]);
  DROR2 I25 (compOut0_0n[4], compOut1_0n[4], compOut0_0n[5], compOut1_0n[5], internalA0_0n[7], internalA1_0n[7]);
  DROR2 I26 (internalA0_0n[7], internalA1_0n[7], internalA0_0n[8], internalA1_0n[8], internalA0_0n[6], internalA1_0n[6]);
  DROR2 I27 (compOut0_0n[2], compOut1_0n[2], compOut0_0n[3], compOut1_0n[3], internalA0_0n[5], internalA1_0n[5]);
  DROR2 I28 (compOut0_0n[0], compOut1_0n[0], compOut0_0n[1], compOut1_0n[1], internalA0_0n[4], internalA1_0n[4]);
  DROR2 I29 (internalA0_0n[4], internalA1_0n[4], internalA0_0n[5], internalA1_0n[5], internalA0_0n[3], internalA1_0n[3]);
  DROR2 I30 (internalA0_0n[3], internalA1_0n[3], internalA0_0n[6], internalA1_0n[6], internalA0_0n[2], internalA1_0n[2]);
  DROR2 I31 (internalA0_0n[2], internalA1_0n[2], internalA0_0n[9], internalA1_0n[9], internalA0_0n[1], internalA1_0n[1]);
  DROR2 I32 (internalA0_0n[1], internalA1_0n[1], internalA0_0n[16], internalA1_0n[16], internalA0_0n[0], internalA1_0n[0]);
  BUFF I33 (compOut0_0n[0], inpA_0a0d[0]);
  BUFF I34 (compOut0_0n[1], inpA_0a0d[1]);
  BUFF I35 (compOut0_0n[2], inpA_0a0d[2]);
  BUFF I36 (compOut0_0n[3], inpA_0a0d[3]);
  BUFF I37 (compOut0_0n[4], inpA_0a0d[4]);
  BUFF I38 (compOut0_0n[5], inpA_0a0d[5]);
  BUFF I39 (compOut0_0n[6], inpA_0a0d[6]);
  BUFF I40 (compOut0_0n[7], inpA_0a0d[7]);
  BUFF I41 (compOut0_0n[8], inpA_0a0d[8]);
  BUFF I42 (compOut0_0n[9], inpA_0a0d[9]);
  BUFF I43 (compOut0_0n[10], inpA_0a0d[10]);
  BUFF I44 (compOut0_0n[11], inpA_0a0d[11]);
  BUFF I45 (compOut0_0n[12], inpA_0a0d[12]);
  BUFF I46 (compOut0_0n[13], inpA_0a0d[13]);
  BUFF I47 (compOut0_0n[14], inpA_0a0d[14]);
  BUFF I48 (compOut0_0n[15], inpA_0a0d[15]);
  BUFF I49 (compOut0_0n[16], inpA_0a0d[16]);
  BUFF I50 (compOut0_0n[17], inpA_0a0d[17]);
  BUFF I51 (compOut0_0n[18], inpA_0a0d[18]);
  BUFF I52 (compOut0_0n[19], inpA_0a0d[19]);
  BUFF I53 (compOut0_0n[20], inpA_0a0d[20]);
  BUFF I54 (compOut0_0n[21], inpA_0a0d[21]);
  BUFF I55 (compOut0_0n[22], inpA_0a0d[22]);
  BUFF I56 (compOut0_0n[23], inpA_0a0d[23]);
  BUFF I57 (compOut0_0n[24], inpA_0a0d[24]);
  BUFF I58 (compOut0_0n[25], inpA_0a0d[25]);
  BUFF I59 (compOut0_0n[26], inpA_0a0d[26]);
  BUFF I60 (compOut0_0n[27], inpA_0a0d[27]);
  BUFF I61 (compOut0_0n[28], inpA_0a0d[28]);
  BUFF I62 (compOut0_0n[29], inpA_0a0d[29]);
  BUFF I63 (compOut0_0n[30], inpA_0a0d[30]);
  BUFF I64 (compOut0_0n[31], inpA_0a0d[31]);
  BUFF I65 (compOut1_0n[0], inpA_0a1d[0]);
  BUFF I66 (compOut1_0n[1], inpA_0a1d[1]);
  BUFF I67 (compOut1_0n[2], inpA_0a1d[2]);
  BUFF I68 (compOut1_0n[3], inpA_0a1d[3]);
  BUFF I69 (compOut1_0n[4], inpA_0a1d[4]);
  BUFF I70 (compOut1_0n[5], inpA_0a1d[5]);
  BUFF I71 (compOut1_0n[6], inpA_0a1d[6]);
  BUFF I72 (compOut1_0n[7], inpA_0a1d[7]);
  BUFF I73 (compOut1_0n[8], inpA_0a1d[8]);
  BUFF I74 (compOut1_0n[9], inpA_0a1d[9]);
  BUFF I75 (compOut1_0n[10], inpA_0a1d[10]);
  BUFF I76 (compOut1_0n[11], inpA_0a1d[11]);
  BUFF I77 (compOut1_0n[12], inpA_0a1d[12]);
  BUFF I78 (compOut1_0n[13], inpA_0a1d[13]);
  BUFF I79 (compOut1_0n[14], inpA_0a1d[14]);
  BUFF I80 (compOut1_0n[15], inpA_0a1d[15]);
  BUFF I81 (compOut1_0n[16], inpA_0a1d[16]);
  BUFF I82 (compOut1_0n[17], inpA_0a1d[17]);
  BUFF I83 (compOut1_0n[18], inpA_0a1d[18]);
  BUFF I84 (compOut1_0n[19], inpA_0a1d[19]);
  BUFF I85 (compOut1_0n[20], inpA_0a1d[20]);
  BUFF I86 (compOut1_0n[21], inpA_0a1d[21]);
  BUFF I87 (compOut1_0n[22], inpA_0a1d[22]);
  BUFF I88 (compOut1_0n[23], inpA_0a1d[23]);
  BUFF I89 (compOut1_0n[24], inpA_0a1d[24]);
  BUFF I90 (compOut1_0n[25], inpA_0a1d[25]);
  BUFF I91 (compOut1_0n[26], inpA_0a1d[26]);
  BUFF I92 (compOut1_0n[27], inpA_0a1d[27]);
  BUFF I93 (compOut1_0n[28], inpA_0a1d[28]);
  BUFF I94 (compOut1_0n[29], inpA_0a1d[29]);
  BUFF I95 (compOut1_0n[30], inpA_0a1d[30]);
  BUFF I96 (compOut1_0n[31], inpA_0a1d[31]);
  BUFF I97 (inpA_0r, out_0r);
endmodule

module BrzCall_2 (
  inp_0r, inp_0a,
  inp_1r, inp_1a,
  out_0r, out_0a
);
  input inp_0r;
  output inp_0a;
  input inp_1r;
  output inp_1a;
  output out_0r;
  input out_0a;
  OR2 I0 (out_0r, inp_0r, inp_1r);
  C2 I1 (inp_0a, inp_0r, out_0a);
  C2 I2 (inp_1a, inp_1r, out_0a);
endmodule

module BrzCallDemux_1_3 (
  out_0r, out_0a0d, out_0a1d,
  out_1r, out_1a0d, out_1a1d,
  out_2r, out_2a0d, out_2a1d,
  inp_0r, inp_0a0d, inp_0a1d
);
  input out_0r;
  output out_0a0d;
  output out_0a1d;
  input out_1r;
  output out_1a0d;
  output out_1a1d;
  input out_2r;
  output out_2a0d;
  output out_2a1d;
  output inp_0r;
  input inp_0a0d;
  input inp_0a1d;
  wire [2:0] outReq_0n;
  OR3 I0 (inp_0r, outReq_0n[0], outReq_0n[1], outReq_0n[2]);
  C2 I1 (out_0a1d, outReq_0n[0], inp_0a1d);
  C2 I2 (out_1a1d, outReq_0n[1], inp_0a1d);
  C2 I3 (out_2a1d, outReq_0n[2], inp_0a1d);
  C2 I4 (out_0a0d, outReq_0n[0], inp_0a0d);
  C2 I5 (out_1a0d, outReq_0n[1], inp_0a0d);
  C2 I6 (out_2a0d, outReq_0n[2], inp_0a0d);
  BUFF I7 (outReq_0n[0], out_0r);
  BUFF I8 (outReq_0n[1], out_1r);
  BUFF I9 (outReq_0n[2], out_2r);
endmodule

module BrzCallDemux_32_2 (
  out_0r, out_0a0d, out_0a1d,
  out_1r, out_1a0d, out_1a1d,
  inp_0r, inp_0a0d, inp_0a1d
);
  input out_0r;
  output [31:0] out_0a0d;
  output [31:0] out_0a1d;
  input out_1r;
  output [31:0] out_1a0d;
  output [31:0] out_1a1d;
  output inp_0r;
  input [31:0] inp_0a0d;
  input [31:0] inp_0a1d;
  wire [1:0] outReq_0n;
  OR2 I0 (inp_0r, outReq_0n[0], outReq_0n[1]);
  C2 I1 (out_0a1d[0], outReq_0n[0], inp_0a1d[0]);
  C2 I2 (out_0a1d[1], outReq_0n[0], inp_0a1d[1]);
  C2 I3 (out_0a1d[2], outReq_0n[0], inp_0a1d[2]);
  C2 I4 (out_0a1d[3], outReq_0n[0], inp_0a1d[3]);
  C2 I5 (out_0a1d[4], outReq_0n[0], inp_0a1d[4]);
  C2 I6 (out_0a1d[5], outReq_0n[0], inp_0a1d[5]);
  C2 I7 (out_0a1d[6], outReq_0n[0], inp_0a1d[6]);
  C2 I8 (out_0a1d[7], outReq_0n[0], inp_0a1d[7]);
  C2 I9 (out_0a1d[8], outReq_0n[0], inp_0a1d[8]);
  C2 I10 (out_0a1d[9], outReq_0n[0], inp_0a1d[9]);
  C2 I11 (out_0a1d[10], outReq_0n[0], inp_0a1d[10]);
  C2 I12 (out_0a1d[11], outReq_0n[0], inp_0a1d[11]);
  C2 I13 (out_0a1d[12], outReq_0n[0], inp_0a1d[12]);
  C2 I14 (out_0a1d[13], outReq_0n[0], inp_0a1d[13]);
  C2 I15 (out_0a1d[14], outReq_0n[0], inp_0a1d[14]);
  C2 I16 (out_0a1d[15], outReq_0n[0], inp_0a1d[15]);
  C2 I17 (out_0a1d[16], outReq_0n[0], inp_0a1d[16]);
  C2 I18 (out_0a1d[17], outReq_0n[0], inp_0a1d[17]);
  C2 I19 (out_0a1d[18], outReq_0n[0], inp_0a1d[18]);
  C2 I20 (out_0a1d[19], outReq_0n[0], inp_0a1d[19]);
  C2 I21 (out_0a1d[20], outReq_0n[0], inp_0a1d[20]);
  C2 I22 (out_0a1d[21], outReq_0n[0], inp_0a1d[21]);
  C2 I23 (out_0a1d[22], outReq_0n[0], inp_0a1d[22]);
  C2 I24 (out_0a1d[23], outReq_0n[0], inp_0a1d[23]);
  C2 I25 (out_0a1d[24], outReq_0n[0], inp_0a1d[24]);
  C2 I26 (out_0a1d[25], outReq_0n[0], inp_0a1d[25]);
  C2 I27 (out_0a1d[26], outReq_0n[0], inp_0a1d[26]);
  C2 I28 (out_0a1d[27], outReq_0n[0], inp_0a1d[27]);
  C2 I29 (out_0a1d[28], outReq_0n[0], inp_0a1d[28]);
  C2 I30 (out_0a1d[29], outReq_0n[0], inp_0a1d[29]);
  C2 I31 (out_0a1d[30], outReq_0n[0], inp_0a1d[30]);
  C2 I32 (out_0a1d[31], outReq_0n[0], inp_0a1d[31]);
  C2 I33 (out_1a1d[0], outReq_0n[1], inp_0a1d[0]);
  C2 I34 (out_1a1d[1], outReq_0n[1], inp_0a1d[1]);
  C2 I35 (out_1a1d[2], outReq_0n[1], inp_0a1d[2]);
  C2 I36 (out_1a1d[3], outReq_0n[1], inp_0a1d[3]);
  C2 I37 (out_1a1d[4], outReq_0n[1], inp_0a1d[4]);
  C2 I38 (out_1a1d[5], outReq_0n[1], inp_0a1d[5]);
  C2 I39 (out_1a1d[6], outReq_0n[1], inp_0a1d[6]);
  C2 I40 (out_1a1d[7], outReq_0n[1], inp_0a1d[7]);
  C2 I41 (out_1a1d[8], outReq_0n[1], inp_0a1d[8]);
  C2 I42 (out_1a1d[9], outReq_0n[1], inp_0a1d[9]);
  C2 I43 (out_1a1d[10], outReq_0n[1], inp_0a1d[10]);
  C2 I44 (out_1a1d[11], outReq_0n[1], inp_0a1d[11]);
  C2 I45 (out_1a1d[12], outReq_0n[1], inp_0a1d[12]);
  C2 I46 (out_1a1d[13], outReq_0n[1], inp_0a1d[13]);
  C2 I47 (out_1a1d[14], outReq_0n[1], inp_0a1d[14]);
  C2 I48 (out_1a1d[15], outReq_0n[1], inp_0a1d[15]);
  C2 I49 (out_1a1d[16], outReq_0n[1], inp_0a1d[16]);
  C2 I50 (out_1a1d[17], outReq_0n[1], inp_0a1d[17]);
  C2 I51 (out_1a1d[18], outReq_0n[1], inp_0a1d[18]);
  C2 I52 (out_1a1d[19], outReq_0n[1], inp_0a1d[19]);
  C2 I53 (out_1a1d[20], outReq_0n[1], inp_0a1d[20]);
  C2 I54 (out_1a1d[21], outReq_0n[1], inp_0a1d[21]);
  C2 I55 (out_1a1d[22], outReq_0n[1], inp_0a1d[22]);
  C2 I56 (out_1a1d[23], outReq_0n[1], inp_0a1d[23]);
  C2 I57 (out_1a1d[24], outReq_0n[1], inp_0a1d[24]);
  C2 I58 (out_1a1d[25], outReq_0n[1], inp_0a1d[25]);
  C2 I59 (out_1a1d[26], outReq_0n[1], inp_0a1d[26]);
  C2 I60 (out_1a1d[27], outReq_0n[1], inp_0a1d[27]);
  C2 I61 (out_1a1d[28], outReq_0n[1], inp_0a1d[28]);
  C2 I62 (out_1a1d[29], outReq_0n[1], inp_0a1d[29]);
  C2 I63 (out_1a1d[30], outReq_0n[1], inp_0a1d[30]);
  C2 I64 (out_1a1d[31], outReq_0n[1], inp_0a1d[31]);
  C2 I65 (out_0a0d[0], outReq_0n[0], inp_0a0d[0]);
  C2 I66 (out_0a0d[1], outReq_0n[0], inp_0a0d[1]);
  C2 I67 (out_0a0d[2], outReq_0n[0], inp_0a0d[2]);
  C2 I68 (out_0a0d[3], outReq_0n[0], inp_0a0d[3]);
  C2 I69 (out_0a0d[4], outReq_0n[0], inp_0a0d[4]);
  C2 I70 (out_0a0d[5], outReq_0n[0], inp_0a0d[5]);
  C2 I71 (out_0a0d[6], outReq_0n[0], inp_0a0d[6]);
  C2 I72 (out_0a0d[7], outReq_0n[0], inp_0a0d[7]);
  C2 I73 (out_0a0d[8], outReq_0n[0], inp_0a0d[8]);
  C2 I74 (out_0a0d[9], outReq_0n[0], inp_0a0d[9]);
  C2 I75 (out_0a0d[10], outReq_0n[0], inp_0a0d[10]);
  C2 I76 (out_0a0d[11], outReq_0n[0], inp_0a0d[11]);
  C2 I77 (out_0a0d[12], outReq_0n[0], inp_0a0d[12]);
  C2 I78 (out_0a0d[13], outReq_0n[0], inp_0a0d[13]);
  C2 I79 (out_0a0d[14], outReq_0n[0], inp_0a0d[14]);
  C2 I80 (out_0a0d[15], outReq_0n[0], inp_0a0d[15]);
  C2 I81 (out_0a0d[16], outReq_0n[0], inp_0a0d[16]);
  C2 I82 (out_0a0d[17], outReq_0n[0], inp_0a0d[17]);
  C2 I83 (out_0a0d[18], outReq_0n[0], inp_0a0d[18]);
  C2 I84 (out_0a0d[19], outReq_0n[0], inp_0a0d[19]);
  C2 I85 (out_0a0d[20], outReq_0n[0], inp_0a0d[20]);
  C2 I86 (out_0a0d[21], outReq_0n[0], inp_0a0d[21]);
  C2 I87 (out_0a0d[22], outReq_0n[0], inp_0a0d[22]);
  C2 I88 (out_0a0d[23], outReq_0n[0], inp_0a0d[23]);
  C2 I89 (out_0a0d[24], outReq_0n[0], inp_0a0d[24]);
  C2 I90 (out_0a0d[25], outReq_0n[0], inp_0a0d[25]);
  C2 I91 (out_0a0d[26], outReq_0n[0], inp_0a0d[26]);
  C2 I92 (out_0a0d[27], outReq_0n[0], inp_0a0d[27]);
  C2 I93 (out_0a0d[28], outReq_0n[0], inp_0a0d[28]);
  C2 I94 (out_0a0d[29], outReq_0n[0], inp_0a0d[29]);
  C2 I95 (out_0a0d[30], outReq_0n[0], inp_0a0d[30]);
  C2 I96 (out_0a0d[31], outReq_0n[0], inp_0a0d[31]);
  C2 I97 (out_1a0d[0], outReq_0n[1], inp_0a0d[0]);
  C2 I98 (out_1a0d[1], outReq_0n[1], inp_0a0d[1]);
  C2 I99 (out_1a0d[2], outReq_0n[1], inp_0a0d[2]);
  C2 I100 (out_1a0d[3], outReq_0n[1], inp_0a0d[3]);
  C2 I101 (out_1a0d[4], outReq_0n[1], inp_0a0d[4]);
  C2 I102 (out_1a0d[5], outReq_0n[1], inp_0a0d[5]);
  C2 I103 (out_1a0d[6], outReq_0n[1], inp_0a0d[6]);
  C2 I104 (out_1a0d[7], outReq_0n[1], inp_0a0d[7]);
  C2 I105 (out_1a0d[8], outReq_0n[1], inp_0a0d[8]);
  C2 I106 (out_1a0d[9], outReq_0n[1], inp_0a0d[9]);
  C2 I107 (out_1a0d[10], outReq_0n[1], inp_0a0d[10]);
  C2 I108 (out_1a0d[11], outReq_0n[1], inp_0a0d[11]);
  C2 I109 (out_1a0d[12], outReq_0n[1], inp_0a0d[12]);
  C2 I110 (out_1a0d[13], outReq_0n[1], inp_0a0d[13]);
  C2 I111 (out_1a0d[14], outReq_0n[1], inp_0a0d[14]);
  C2 I112 (out_1a0d[15], outReq_0n[1], inp_0a0d[15]);
  C2 I113 (out_1a0d[16], outReq_0n[1], inp_0a0d[16]);
  C2 I114 (out_1a0d[17], outReq_0n[1], inp_0a0d[17]);
  C2 I115 (out_1a0d[18], outReq_0n[1], inp_0a0d[18]);
  C2 I116 (out_1a0d[19], outReq_0n[1], inp_0a0d[19]);
  C2 I117 (out_1a0d[20], outReq_0n[1], inp_0a0d[20]);
  C2 I118 (out_1a0d[21], outReq_0n[1], inp_0a0d[21]);
  C2 I119 (out_1a0d[22], outReq_0n[1], inp_0a0d[22]);
  C2 I120 (out_1a0d[23], outReq_0n[1], inp_0a0d[23]);
  C2 I121 (out_1a0d[24], outReq_0n[1], inp_0a0d[24]);
  C2 I122 (out_1a0d[25], outReq_0n[1], inp_0a0d[25]);
  C2 I123 (out_1a0d[26], outReq_0n[1], inp_0a0d[26]);
  C2 I124 (out_1a0d[27], outReq_0n[1], inp_0a0d[27]);
  C2 I125 (out_1a0d[28], outReq_0n[1], inp_0a0d[28]);
  C2 I126 (out_1a0d[29], outReq_0n[1], inp_0a0d[29]);
  C2 I127 (out_1a0d[30], outReq_0n[1], inp_0a0d[30]);
  C2 I128 (out_1a0d[31], outReq_0n[1], inp_0a0d[31]);
  BUFF I129 (outReq_0n[0], out_0r);
  BUFF I130 (outReq_0n[1], out_1r);
endmodule

module BrzCallDemux_32_3 (
  out_0r, out_0a0d, out_0a1d,
  out_1r, out_1a0d, out_1a1d,
  out_2r, out_2a0d, out_2a1d,
  inp_0r, inp_0a0d, inp_0a1d
);
  input out_0r;
  output [31:0] out_0a0d;
  output [31:0] out_0a1d;
  input out_1r;
  output [31:0] out_1a0d;
  output [31:0] out_1a1d;
  input out_2r;
  output [31:0] out_2a0d;
  output [31:0] out_2a1d;
  output inp_0r;
  input [31:0] inp_0a0d;
  input [31:0] inp_0a1d;
  wire [2:0] outReq_0n;
  OR3 I0 (inp_0r, outReq_0n[0], outReq_0n[1], outReq_0n[2]);
  C2 I1 (out_0a1d[0], outReq_0n[0], inp_0a1d[0]);
  C2 I2 (out_0a1d[1], outReq_0n[0], inp_0a1d[1]);
  C2 I3 (out_0a1d[2], outReq_0n[0], inp_0a1d[2]);
  C2 I4 (out_0a1d[3], outReq_0n[0], inp_0a1d[3]);
  C2 I5 (out_0a1d[4], outReq_0n[0], inp_0a1d[4]);
  C2 I6 (out_0a1d[5], outReq_0n[0], inp_0a1d[5]);
  C2 I7 (out_0a1d[6], outReq_0n[0], inp_0a1d[6]);
  C2 I8 (out_0a1d[7], outReq_0n[0], inp_0a1d[7]);
  C2 I9 (out_0a1d[8], outReq_0n[0], inp_0a1d[8]);
  C2 I10 (out_0a1d[9], outReq_0n[0], inp_0a1d[9]);
  C2 I11 (out_0a1d[10], outReq_0n[0], inp_0a1d[10]);
  C2 I12 (out_0a1d[11], outReq_0n[0], inp_0a1d[11]);
  C2 I13 (out_0a1d[12], outReq_0n[0], inp_0a1d[12]);
  C2 I14 (out_0a1d[13], outReq_0n[0], inp_0a1d[13]);
  C2 I15 (out_0a1d[14], outReq_0n[0], inp_0a1d[14]);
  C2 I16 (out_0a1d[15], outReq_0n[0], inp_0a1d[15]);
  C2 I17 (out_0a1d[16], outReq_0n[0], inp_0a1d[16]);
  C2 I18 (out_0a1d[17], outReq_0n[0], inp_0a1d[17]);
  C2 I19 (out_0a1d[18], outReq_0n[0], inp_0a1d[18]);
  C2 I20 (out_0a1d[19], outReq_0n[0], inp_0a1d[19]);
  C2 I21 (out_0a1d[20], outReq_0n[0], inp_0a1d[20]);
  C2 I22 (out_0a1d[21], outReq_0n[0], inp_0a1d[21]);
  C2 I23 (out_0a1d[22], outReq_0n[0], inp_0a1d[22]);
  C2 I24 (out_0a1d[23], outReq_0n[0], inp_0a1d[23]);
  C2 I25 (out_0a1d[24], outReq_0n[0], inp_0a1d[24]);
  C2 I26 (out_0a1d[25], outReq_0n[0], inp_0a1d[25]);
  C2 I27 (out_0a1d[26], outReq_0n[0], inp_0a1d[26]);
  C2 I28 (out_0a1d[27], outReq_0n[0], inp_0a1d[27]);
  C2 I29 (out_0a1d[28], outReq_0n[0], inp_0a1d[28]);
  C2 I30 (out_0a1d[29], outReq_0n[0], inp_0a1d[29]);
  C2 I31 (out_0a1d[30], outReq_0n[0], inp_0a1d[30]);
  C2 I32 (out_0a1d[31], outReq_0n[0], inp_0a1d[31]);
  C2 I33 (out_1a1d[0], outReq_0n[1], inp_0a1d[0]);
  C2 I34 (out_1a1d[1], outReq_0n[1], inp_0a1d[1]);
  C2 I35 (out_1a1d[2], outReq_0n[1], inp_0a1d[2]);
  C2 I36 (out_1a1d[3], outReq_0n[1], inp_0a1d[3]);
  C2 I37 (out_1a1d[4], outReq_0n[1], inp_0a1d[4]);
  C2 I38 (out_1a1d[5], outReq_0n[1], inp_0a1d[5]);
  C2 I39 (out_1a1d[6], outReq_0n[1], inp_0a1d[6]);
  C2 I40 (out_1a1d[7], outReq_0n[1], inp_0a1d[7]);
  C2 I41 (out_1a1d[8], outReq_0n[1], inp_0a1d[8]);
  C2 I42 (out_1a1d[9], outReq_0n[1], inp_0a1d[9]);
  C2 I43 (out_1a1d[10], outReq_0n[1], inp_0a1d[10]);
  C2 I44 (out_1a1d[11], outReq_0n[1], inp_0a1d[11]);
  C2 I45 (out_1a1d[12], outReq_0n[1], inp_0a1d[12]);
  C2 I46 (out_1a1d[13], outReq_0n[1], inp_0a1d[13]);
  C2 I47 (out_1a1d[14], outReq_0n[1], inp_0a1d[14]);
  C2 I48 (out_1a1d[15], outReq_0n[1], inp_0a1d[15]);
  C2 I49 (out_1a1d[16], outReq_0n[1], inp_0a1d[16]);
  C2 I50 (out_1a1d[17], outReq_0n[1], inp_0a1d[17]);
  C2 I51 (out_1a1d[18], outReq_0n[1], inp_0a1d[18]);
  C2 I52 (out_1a1d[19], outReq_0n[1], inp_0a1d[19]);
  C2 I53 (out_1a1d[20], outReq_0n[1], inp_0a1d[20]);
  C2 I54 (out_1a1d[21], outReq_0n[1], inp_0a1d[21]);
  C2 I55 (out_1a1d[22], outReq_0n[1], inp_0a1d[22]);
  C2 I56 (out_1a1d[23], outReq_0n[1], inp_0a1d[23]);
  C2 I57 (out_1a1d[24], outReq_0n[1], inp_0a1d[24]);
  C2 I58 (out_1a1d[25], outReq_0n[1], inp_0a1d[25]);
  C2 I59 (out_1a1d[26], outReq_0n[1], inp_0a1d[26]);
  C2 I60 (out_1a1d[27], outReq_0n[1], inp_0a1d[27]);
  C2 I61 (out_1a1d[28], outReq_0n[1], inp_0a1d[28]);
  C2 I62 (out_1a1d[29], outReq_0n[1], inp_0a1d[29]);
  C2 I63 (out_1a1d[30], outReq_0n[1], inp_0a1d[30]);
  C2 I64 (out_1a1d[31], outReq_0n[1], inp_0a1d[31]);
  C2 I65 (out_2a1d[0], outReq_0n[2], inp_0a1d[0]);
  C2 I66 (out_2a1d[1], outReq_0n[2], inp_0a1d[1]);
  C2 I67 (out_2a1d[2], outReq_0n[2], inp_0a1d[2]);
  C2 I68 (out_2a1d[3], outReq_0n[2], inp_0a1d[3]);
  C2 I69 (out_2a1d[4], outReq_0n[2], inp_0a1d[4]);
  C2 I70 (out_2a1d[5], outReq_0n[2], inp_0a1d[5]);
  C2 I71 (out_2a1d[6], outReq_0n[2], inp_0a1d[6]);
  C2 I72 (out_2a1d[7], outReq_0n[2], inp_0a1d[7]);
  C2 I73 (out_2a1d[8], outReq_0n[2], inp_0a1d[8]);
  C2 I74 (out_2a1d[9], outReq_0n[2], inp_0a1d[9]);
  C2 I75 (out_2a1d[10], outReq_0n[2], inp_0a1d[10]);
  C2 I76 (out_2a1d[11], outReq_0n[2], inp_0a1d[11]);
  C2 I77 (out_2a1d[12], outReq_0n[2], inp_0a1d[12]);
  C2 I78 (out_2a1d[13], outReq_0n[2], inp_0a1d[13]);
  C2 I79 (out_2a1d[14], outReq_0n[2], inp_0a1d[14]);
  C2 I80 (out_2a1d[15], outReq_0n[2], inp_0a1d[15]);
  C2 I81 (out_2a1d[16], outReq_0n[2], inp_0a1d[16]);
  C2 I82 (out_2a1d[17], outReq_0n[2], inp_0a1d[17]);
  C2 I83 (out_2a1d[18], outReq_0n[2], inp_0a1d[18]);
  C2 I84 (out_2a1d[19], outReq_0n[2], inp_0a1d[19]);
  C2 I85 (out_2a1d[20], outReq_0n[2], inp_0a1d[20]);
  C2 I86 (out_2a1d[21], outReq_0n[2], inp_0a1d[21]);
  C2 I87 (out_2a1d[22], outReq_0n[2], inp_0a1d[22]);
  C2 I88 (out_2a1d[23], outReq_0n[2], inp_0a1d[23]);
  C2 I89 (out_2a1d[24], outReq_0n[2], inp_0a1d[24]);
  C2 I90 (out_2a1d[25], outReq_0n[2], inp_0a1d[25]);
  C2 I91 (out_2a1d[26], outReq_0n[2], inp_0a1d[26]);
  C2 I92 (out_2a1d[27], outReq_0n[2], inp_0a1d[27]);
  C2 I93 (out_2a1d[28], outReq_0n[2], inp_0a1d[28]);
  C2 I94 (out_2a1d[29], outReq_0n[2], inp_0a1d[29]);
  C2 I95 (out_2a1d[30], outReq_0n[2], inp_0a1d[30]);
  C2 I96 (out_2a1d[31], outReq_0n[2], inp_0a1d[31]);
  C2 I97 (out_0a0d[0], outReq_0n[0], inp_0a0d[0]);
  C2 I98 (out_0a0d[1], outReq_0n[0], inp_0a0d[1]);
  C2 I99 (out_0a0d[2], outReq_0n[0], inp_0a0d[2]);
  C2 I100 (out_0a0d[3], outReq_0n[0], inp_0a0d[3]);
  C2 I101 (out_0a0d[4], outReq_0n[0], inp_0a0d[4]);
  C2 I102 (out_0a0d[5], outReq_0n[0], inp_0a0d[5]);
  C2 I103 (out_0a0d[6], outReq_0n[0], inp_0a0d[6]);
  C2 I104 (out_0a0d[7], outReq_0n[0], inp_0a0d[7]);
  C2 I105 (out_0a0d[8], outReq_0n[0], inp_0a0d[8]);
  C2 I106 (out_0a0d[9], outReq_0n[0], inp_0a0d[9]);
  C2 I107 (out_0a0d[10], outReq_0n[0], inp_0a0d[10]);
  C2 I108 (out_0a0d[11], outReq_0n[0], inp_0a0d[11]);
  C2 I109 (out_0a0d[12], outReq_0n[0], inp_0a0d[12]);
  C2 I110 (out_0a0d[13], outReq_0n[0], inp_0a0d[13]);
  C2 I111 (out_0a0d[14], outReq_0n[0], inp_0a0d[14]);
  C2 I112 (out_0a0d[15], outReq_0n[0], inp_0a0d[15]);
  C2 I113 (out_0a0d[16], outReq_0n[0], inp_0a0d[16]);
  C2 I114 (out_0a0d[17], outReq_0n[0], inp_0a0d[17]);
  C2 I115 (out_0a0d[18], outReq_0n[0], inp_0a0d[18]);
  C2 I116 (out_0a0d[19], outReq_0n[0], inp_0a0d[19]);
  C2 I117 (out_0a0d[20], outReq_0n[0], inp_0a0d[20]);
  C2 I118 (out_0a0d[21], outReq_0n[0], inp_0a0d[21]);
  C2 I119 (out_0a0d[22], outReq_0n[0], inp_0a0d[22]);
  C2 I120 (out_0a0d[23], outReq_0n[0], inp_0a0d[23]);
  C2 I121 (out_0a0d[24], outReq_0n[0], inp_0a0d[24]);
  C2 I122 (out_0a0d[25], outReq_0n[0], inp_0a0d[25]);
  C2 I123 (out_0a0d[26], outReq_0n[0], inp_0a0d[26]);
  C2 I124 (out_0a0d[27], outReq_0n[0], inp_0a0d[27]);
  C2 I125 (out_0a0d[28], outReq_0n[0], inp_0a0d[28]);
  C2 I126 (out_0a0d[29], outReq_0n[0], inp_0a0d[29]);
  C2 I127 (out_0a0d[30], outReq_0n[0], inp_0a0d[30]);
  C2 I128 (out_0a0d[31], outReq_0n[0], inp_0a0d[31]);
  C2 I129 (out_1a0d[0], outReq_0n[1], inp_0a0d[0]);
  C2 I130 (out_1a0d[1], outReq_0n[1], inp_0a0d[1]);
  C2 I131 (out_1a0d[2], outReq_0n[1], inp_0a0d[2]);
  C2 I132 (out_1a0d[3], outReq_0n[1], inp_0a0d[3]);
  C2 I133 (out_1a0d[4], outReq_0n[1], inp_0a0d[4]);
  C2 I134 (out_1a0d[5], outReq_0n[1], inp_0a0d[5]);
  C2 I135 (out_1a0d[6], outReq_0n[1], inp_0a0d[6]);
  C2 I136 (out_1a0d[7], outReq_0n[1], inp_0a0d[7]);
  C2 I137 (out_1a0d[8], outReq_0n[1], inp_0a0d[8]);
  C2 I138 (out_1a0d[9], outReq_0n[1], inp_0a0d[9]);
  C2 I139 (out_1a0d[10], outReq_0n[1], inp_0a0d[10]);
  C2 I140 (out_1a0d[11], outReq_0n[1], inp_0a0d[11]);
  C2 I141 (out_1a0d[12], outReq_0n[1], inp_0a0d[12]);
  C2 I142 (out_1a0d[13], outReq_0n[1], inp_0a0d[13]);
  C2 I143 (out_1a0d[14], outReq_0n[1], inp_0a0d[14]);
  C2 I144 (out_1a0d[15], outReq_0n[1], inp_0a0d[15]);
  C2 I145 (out_1a0d[16], outReq_0n[1], inp_0a0d[16]);
  C2 I146 (out_1a0d[17], outReq_0n[1], inp_0a0d[17]);
  C2 I147 (out_1a0d[18], outReq_0n[1], inp_0a0d[18]);
  C2 I148 (out_1a0d[19], outReq_0n[1], inp_0a0d[19]);
  C2 I149 (out_1a0d[20], outReq_0n[1], inp_0a0d[20]);
  C2 I150 (out_1a0d[21], outReq_0n[1], inp_0a0d[21]);
  C2 I151 (out_1a0d[22], outReq_0n[1], inp_0a0d[22]);
  C2 I152 (out_1a0d[23], outReq_0n[1], inp_0a0d[23]);
  C2 I153 (out_1a0d[24], outReq_0n[1], inp_0a0d[24]);
  C2 I154 (out_1a0d[25], outReq_0n[1], inp_0a0d[25]);
  C2 I155 (out_1a0d[26], outReq_0n[1], inp_0a0d[26]);
  C2 I156 (out_1a0d[27], outReq_0n[1], inp_0a0d[27]);
  C2 I157 (out_1a0d[28], outReq_0n[1], inp_0a0d[28]);
  C2 I158 (out_1a0d[29], outReq_0n[1], inp_0a0d[29]);
  C2 I159 (out_1a0d[30], outReq_0n[1], inp_0a0d[30]);
  C2 I160 (out_1a0d[31], outReq_0n[1], inp_0a0d[31]);
  C2 I161 (out_2a0d[0], outReq_0n[2], inp_0a0d[0]);
  C2 I162 (out_2a0d[1], outReq_0n[2], inp_0a0d[1]);
  C2 I163 (out_2a0d[2], outReq_0n[2], inp_0a0d[2]);
  C2 I164 (out_2a0d[3], outReq_0n[2], inp_0a0d[3]);
  C2 I165 (out_2a0d[4], outReq_0n[2], inp_0a0d[4]);
  C2 I166 (out_2a0d[5], outReq_0n[2], inp_0a0d[5]);
  C2 I167 (out_2a0d[6], outReq_0n[2], inp_0a0d[6]);
  C2 I168 (out_2a0d[7], outReq_0n[2], inp_0a0d[7]);
  C2 I169 (out_2a0d[8], outReq_0n[2], inp_0a0d[8]);
  C2 I170 (out_2a0d[9], outReq_0n[2], inp_0a0d[9]);
  C2 I171 (out_2a0d[10], outReq_0n[2], inp_0a0d[10]);
  C2 I172 (out_2a0d[11], outReq_0n[2], inp_0a0d[11]);
  C2 I173 (out_2a0d[12], outReq_0n[2], inp_0a0d[12]);
  C2 I174 (out_2a0d[13], outReq_0n[2], inp_0a0d[13]);
  C2 I175 (out_2a0d[14], outReq_0n[2], inp_0a0d[14]);
  C2 I176 (out_2a0d[15], outReq_0n[2], inp_0a0d[15]);
  C2 I177 (out_2a0d[16], outReq_0n[2], inp_0a0d[16]);
  C2 I178 (out_2a0d[17], outReq_0n[2], inp_0a0d[17]);
  C2 I179 (out_2a0d[18], outReq_0n[2], inp_0a0d[18]);
  C2 I180 (out_2a0d[19], outReq_0n[2], inp_0a0d[19]);
  C2 I181 (out_2a0d[20], outReq_0n[2], inp_0a0d[20]);
  C2 I182 (out_2a0d[21], outReq_0n[2], inp_0a0d[21]);
  C2 I183 (out_2a0d[22], outReq_0n[2], inp_0a0d[22]);
  C2 I184 (out_2a0d[23], outReq_0n[2], inp_0a0d[23]);
  C2 I185 (out_2a0d[24], outReq_0n[2], inp_0a0d[24]);
  C2 I186 (out_2a0d[25], outReq_0n[2], inp_0a0d[25]);
  C2 I187 (out_2a0d[26], outReq_0n[2], inp_0a0d[26]);
  C2 I188 (out_2a0d[27], outReq_0n[2], inp_0a0d[27]);
  C2 I189 (out_2a0d[28], outReq_0n[2], inp_0a0d[28]);
  C2 I190 (out_2a0d[29], outReq_0n[2], inp_0a0d[29]);
  C2 I191 (out_2a0d[30], outReq_0n[2], inp_0a0d[30]);
  C2 I192 (out_2a0d[31], outReq_0n[2], inp_0a0d[31]);
  BUFF I193 (outReq_0n[0], out_0r);
  BUFF I194 (outReq_0n[1], out_1r);
  BUFF I195 (outReq_0n[2], out_2r);
endmodule

module BrzCallMux_1_2 (
  inp_0r0d, inp_0r1d, inp_0a,
  inp_1r0d, inp_1r1d, inp_1a,
  out_0r0d, out_0r1d, out_0a
);
  input inp_0r0d;
  input inp_0r1d;
  output inp_0a;
  input inp_1r0d;
  input inp_1r1d;
  output inp_1a;
  output out_0r0d;
  output out_0r1d;
  input out_0a;
  wire [1:0] sourceId_0n;
  C2 I0 (inp_0a, sourceId_0n[0], out_0a);
  C2 I1 (inp_1a, sourceId_0n[1], out_0a);
  OR2 I2 (sourceId_0n[0], inp_0r0d, inp_0r1d);
  OR2 I3 (sourceId_0n[1], inp_1r0d, inp_1r1d);
  OR2 I4 (out_0r1d, inp_0r1d, inp_1r1d);
  OR2 I5 (out_0r0d, inp_0r0d, inp_1r0d);
endmodule

module BrzCallMux_1_3 (
  inp_0r0d, inp_0r1d, inp_0a,
  inp_1r0d, inp_1r1d, inp_1a,
  inp_2r0d, inp_2r1d, inp_2a,
  out_0r0d, out_0r1d, out_0a
);
  input inp_0r0d;
  input inp_0r1d;
  output inp_0a;
  input inp_1r0d;
  input inp_1r1d;
  output inp_1a;
  input inp_2r0d;
  input inp_2r1d;
  output inp_2a;
  output out_0r0d;
  output out_0r1d;
  input out_0a;
  wire [2:0] sourceId_0n;
  C2 I0 (inp_0a, sourceId_0n[0], out_0a);
  C2 I1 (inp_1a, sourceId_0n[1], out_0a);
  C2 I2 (inp_2a, sourceId_0n[2], out_0a);
  OR2 I3 (sourceId_0n[0], inp_0r0d, inp_0r1d);
  OR2 I4 (sourceId_0n[1], inp_1r0d, inp_1r1d);
  OR2 I5 (sourceId_0n[2], inp_2r0d, inp_2r1d);
  OR3 I6 (out_0r1d, inp_0r1d, inp_1r1d, inp_2r1d);
  OR3 I7 (out_0r0d, inp_0r0d, inp_1r0d, inp_2r0d);
endmodule

module BrzCallMux_4_2 (
  inp_0r0d, inp_0r1d, inp_0a,
  inp_1r0d, inp_1r1d, inp_1a,
  out_0r0d, out_0r1d, out_0a
);
  input [3:0] inp_0r0d;
  input [3:0] inp_0r1d;
  output inp_0a;
  input [3:0] inp_1r0d;
  input [3:0] inp_1r1d;
  output inp_1a;
  output [3:0] out_0r0d;
  output [3:0] out_0r1d;
  input out_0a;
  wire [1:0] sourceId_0n;
  C2 I0 (inp_0a, sourceId_0n[0], out_0a);
  C2 I1 (inp_1a, sourceId_0n[1], out_0a);
  OR2 I2 (sourceId_0n[0], inp_0r0d[0], inp_0r1d[0]);
  OR2 I3 (sourceId_0n[1], inp_1r0d[0], inp_1r1d[0]);
  OR2 I4 (out_0r1d[0], inp_0r1d[0], inp_1r1d[0]);
  OR2 I5 (out_0r1d[1], inp_0r1d[1], inp_1r1d[1]);
  OR2 I6 (out_0r1d[2], inp_0r1d[2], inp_1r1d[2]);
  OR2 I7 (out_0r1d[3], inp_0r1d[3], inp_1r1d[3]);
  OR2 I8 (out_0r0d[0], inp_0r0d[0], inp_1r0d[0]);
  OR2 I9 (out_0r0d[1], inp_0r0d[1], inp_1r0d[1]);
  OR2 I10 (out_0r0d[2], inp_0r0d[2], inp_1r0d[2]);
  OR2 I11 (out_0r0d[3], inp_0r0d[3], inp_1r0d[3]);
endmodule

module BrzCallMux_10_2 (
  inp_0r0d, inp_0r1d, inp_0a,
  inp_1r0d, inp_1r1d, inp_1a,
  out_0r0d, out_0r1d, out_0a
);
  input [9:0] inp_0r0d;
  input [9:0] inp_0r1d;
  output inp_0a;
  input [9:0] inp_1r0d;
  input [9:0] inp_1r1d;
  output inp_1a;
  output [9:0] out_0r0d;
  output [9:0] out_0r1d;
  input out_0a;
  wire [1:0] sourceId_0n;
  C2 I0 (inp_0a, sourceId_0n[0], out_0a);
  C2 I1 (inp_1a, sourceId_0n[1], out_0a);
  OR2 I2 (sourceId_0n[0], inp_0r0d[0], inp_0r1d[0]);
  OR2 I3 (sourceId_0n[1], inp_1r0d[0], inp_1r1d[0]);
  OR2 I4 (out_0r1d[0], inp_0r1d[0], inp_1r1d[0]);
  OR2 I5 (out_0r1d[1], inp_0r1d[1], inp_1r1d[1]);
  OR2 I6 (out_0r1d[2], inp_0r1d[2], inp_1r1d[2]);
  OR2 I7 (out_0r1d[3], inp_0r1d[3], inp_1r1d[3]);
  OR2 I8 (out_0r1d[4], inp_0r1d[4], inp_1r1d[4]);
  OR2 I9 (out_0r1d[5], inp_0r1d[5], inp_1r1d[5]);
  OR2 I10 (out_0r1d[6], inp_0r1d[6], inp_1r1d[6]);
  OR2 I11 (out_0r1d[7], inp_0r1d[7], inp_1r1d[7]);
  OR2 I12 (out_0r1d[8], inp_0r1d[8], inp_1r1d[8]);
  OR2 I13 (out_0r1d[9], inp_0r1d[9], inp_1r1d[9]);
  OR2 I14 (out_0r0d[0], inp_0r0d[0], inp_1r0d[0]);
  OR2 I15 (out_0r0d[1], inp_0r0d[1], inp_1r0d[1]);
  OR2 I16 (out_0r0d[2], inp_0r0d[2], inp_1r0d[2]);
  OR2 I17 (out_0r0d[3], inp_0r0d[3], inp_1r0d[3]);
  OR2 I18 (out_0r0d[4], inp_0r0d[4], inp_1r0d[4]);
  OR2 I19 (out_0r0d[5], inp_0r0d[5], inp_1r0d[5]);
  OR2 I20 (out_0r0d[6], inp_0r0d[6], inp_1r0d[6]);
  OR2 I21 (out_0r0d[7], inp_0r0d[7], inp_1r0d[7]);
  OR2 I22 (out_0r0d[8], inp_0r0d[8], inp_1r0d[8]);
  OR2 I23 (out_0r0d[9], inp_0r0d[9], inp_1r0d[9]);
endmodule

module BrzCallMux_32_2 (
  inp_0r0d, inp_0r1d, inp_0a,
  inp_1r0d, inp_1r1d, inp_1a,
  out_0r0d, out_0r1d, out_0a
);
  input [31:0] inp_0r0d;
  input [31:0] inp_0r1d;
  output inp_0a;
  input [31:0] inp_1r0d;
  input [31:0] inp_1r1d;
  output inp_1a;
  output [31:0] out_0r0d;
  output [31:0] out_0r1d;
  input out_0a;
  wire [1:0] sourceId_0n;
  C2 I0 (inp_0a, sourceId_0n[0], out_0a);
  C2 I1 (inp_1a, sourceId_0n[1], out_0a);
  OR2 I2 (sourceId_0n[0], inp_0r0d[0], inp_0r1d[0]);
  OR2 I3 (sourceId_0n[1], inp_1r0d[0], inp_1r1d[0]);
  OR2 I4 (out_0r1d[0], inp_0r1d[0], inp_1r1d[0]);
  OR2 I5 (out_0r1d[1], inp_0r1d[1], inp_1r1d[1]);
  OR2 I6 (out_0r1d[2], inp_0r1d[2], inp_1r1d[2]);
  OR2 I7 (out_0r1d[3], inp_0r1d[3], inp_1r1d[3]);
  OR2 I8 (out_0r1d[4], inp_0r1d[4], inp_1r1d[4]);
  OR2 I9 (out_0r1d[5], inp_0r1d[5], inp_1r1d[5]);
  OR2 I10 (out_0r1d[6], inp_0r1d[6], inp_1r1d[6]);
  OR2 I11 (out_0r1d[7], inp_0r1d[7], inp_1r1d[7]);
  OR2 I12 (out_0r1d[8], inp_0r1d[8], inp_1r1d[8]);
  OR2 I13 (out_0r1d[9], inp_0r1d[9], inp_1r1d[9]);
  OR2 I14 (out_0r1d[10], inp_0r1d[10], inp_1r1d[10]);
  OR2 I15 (out_0r1d[11], inp_0r1d[11], inp_1r1d[11]);
  OR2 I16 (out_0r1d[12], inp_0r1d[12], inp_1r1d[12]);
  OR2 I17 (out_0r1d[13], inp_0r1d[13], inp_1r1d[13]);
  OR2 I18 (out_0r1d[14], inp_0r1d[14], inp_1r1d[14]);
  OR2 I19 (out_0r1d[15], inp_0r1d[15], inp_1r1d[15]);
  OR2 I20 (out_0r1d[16], inp_0r1d[16], inp_1r1d[16]);
  OR2 I21 (out_0r1d[17], inp_0r1d[17], inp_1r1d[17]);
  OR2 I22 (out_0r1d[18], inp_0r1d[18], inp_1r1d[18]);
  OR2 I23 (out_0r1d[19], inp_0r1d[19], inp_1r1d[19]);
  OR2 I24 (out_0r1d[20], inp_0r1d[20], inp_1r1d[20]);
  OR2 I25 (out_0r1d[21], inp_0r1d[21], inp_1r1d[21]);
  OR2 I26 (out_0r1d[22], inp_0r1d[22], inp_1r1d[22]);
  OR2 I27 (out_0r1d[23], inp_0r1d[23], inp_1r1d[23]);
  OR2 I28 (out_0r1d[24], inp_0r1d[24], inp_1r1d[24]);
  OR2 I29 (out_0r1d[25], inp_0r1d[25], inp_1r1d[25]);
  OR2 I30 (out_0r1d[26], inp_0r1d[26], inp_1r1d[26]);
  OR2 I31 (out_0r1d[27], inp_0r1d[27], inp_1r1d[27]);
  OR2 I32 (out_0r1d[28], inp_0r1d[28], inp_1r1d[28]);
  OR2 I33 (out_0r1d[29], inp_0r1d[29], inp_1r1d[29]);
  OR2 I34 (out_0r1d[30], inp_0r1d[30], inp_1r1d[30]);
  OR2 I35 (out_0r1d[31], inp_0r1d[31], inp_1r1d[31]);
  OR2 I36 (out_0r0d[0], inp_0r0d[0], inp_1r0d[0]);
  OR2 I37 (out_0r0d[1], inp_0r0d[1], inp_1r0d[1]);
  OR2 I38 (out_0r0d[2], inp_0r0d[2], inp_1r0d[2]);
  OR2 I39 (out_0r0d[3], inp_0r0d[3], inp_1r0d[3]);
  OR2 I40 (out_0r0d[4], inp_0r0d[4], inp_1r0d[4]);
  OR2 I41 (out_0r0d[5], inp_0r0d[5], inp_1r0d[5]);
  OR2 I42 (out_0r0d[6], inp_0r0d[6], inp_1r0d[6]);
  OR2 I43 (out_0r0d[7], inp_0r0d[7], inp_1r0d[7]);
  OR2 I44 (out_0r0d[8], inp_0r0d[8], inp_1r0d[8]);
  OR2 I45 (out_0r0d[9], inp_0r0d[9], inp_1r0d[9]);
  OR2 I46 (out_0r0d[10], inp_0r0d[10], inp_1r0d[10]);
  OR2 I47 (out_0r0d[11], inp_0r0d[11], inp_1r0d[11]);
  OR2 I48 (out_0r0d[12], inp_0r0d[12], inp_1r0d[12]);
  OR2 I49 (out_0r0d[13], inp_0r0d[13], inp_1r0d[13]);
  OR2 I50 (out_0r0d[14], inp_0r0d[14], inp_1r0d[14]);
  OR2 I51 (out_0r0d[15], inp_0r0d[15], inp_1r0d[15]);
  OR2 I52 (out_0r0d[16], inp_0r0d[16], inp_1r0d[16]);
  OR2 I53 (out_0r0d[17], inp_0r0d[17], inp_1r0d[17]);
  OR2 I54 (out_0r0d[18], inp_0r0d[18], inp_1r0d[18]);
  OR2 I55 (out_0r0d[19], inp_0r0d[19], inp_1r0d[19]);
  OR2 I56 (out_0r0d[20], inp_0r0d[20], inp_1r0d[20]);
  OR2 I57 (out_0r0d[21], inp_0r0d[21], inp_1r0d[21]);
  OR2 I58 (out_0r0d[22], inp_0r0d[22], inp_1r0d[22]);
  OR2 I59 (out_0r0d[23], inp_0r0d[23], inp_1r0d[23]);
  OR2 I60 (out_0r0d[24], inp_0r0d[24], inp_1r0d[24]);
  OR2 I61 (out_0r0d[25], inp_0r0d[25], inp_1r0d[25]);
  OR2 I62 (out_0r0d[26], inp_0r0d[26], inp_1r0d[26]);
  OR2 I63 (out_0r0d[27], inp_0r0d[27], inp_1r0d[27]);
  OR2 I64 (out_0r0d[28], inp_0r0d[28], inp_1r0d[28]);
  OR2 I65 (out_0r0d[29], inp_0r0d[29], inp_1r0d[29]);
  OR2 I66 (out_0r0d[30], inp_0r0d[30], inp_1r0d[30]);
  OR2 I67 (out_0r0d[31], inp_0r0d[31], inp_1r0d[31]);
endmodule

module BrzCallMux_32_3 (
  inp_0r0d, inp_0r1d, inp_0a,
  inp_1r0d, inp_1r1d, inp_1a,
  inp_2r0d, inp_2r1d, inp_2a,
  out_0r0d, out_0r1d, out_0a
);
  input [31:0] inp_0r0d;
  input [31:0] inp_0r1d;
  output inp_0a;
  input [31:0] inp_1r0d;
  input [31:0] inp_1r1d;
  output inp_1a;
  input [31:0] inp_2r0d;
  input [31:0] inp_2r1d;
  output inp_2a;
  output [31:0] out_0r0d;
  output [31:0] out_0r1d;
  input out_0a;
  wire [2:0] sourceId_0n;
  C2 I0 (inp_0a, sourceId_0n[0], out_0a);
  C2 I1 (inp_1a, sourceId_0n[1], out_0a);
  C2 I2 (inp_2a, sourceId_0n[2], out_0a);
  OR2 I3 (sourceId_0n[0], inp_0r0d[0], inp_0r1d[0]);
  OR2 I4 (sourceId_0n[1], inp_1r0d[0], inp_1r1d[0]);
  OR2 I5 (sourceId_0n[2], inp_2r0d[0], inp_2r1d[0]);
  OR3 I6 (out_0r1d[0], inp_0r1d[0], inp_1r1d[0], inp_2r1d[0]);
  OR3 I7 (out_0r1d[1], inp_0r1d[1], inp_1r1d[1], inp_2r1d[1]);
  OR3 I8 (out_0r1d[2], inp_0r1d[2], inp_1r1d[2], inp_2r1d[2]);
  OR3 I9 (out_0r1d[3], inp_0r1d[3], inp_1r1d[3], inp_2r1d[3]);
  OR3 I10 (out_0r1d[4], inp_0r1d[4], inp_1r1d[4], inp_2r1d[4]);
  OR3 I11 (out_0r1d[5], inp_0r1d[5], inp_1r1d[5], inp_2r1d[5]);
  OR3 I12 (out_0r1d[6], inp_0r1d[6], inp_1r1d[6], inp_2r1d[6]);
  OR3 I13 (out_0r1d[7], inp_0r1d[7], inp_1r1d[7], inp_2r1d[7]);
  OR3 I14 (out_0r1d[8], inp_0r1d[8], inp_1r1d[8], inp_2r1d[8]);
  OR3 I15 (out_0r1d[9], inp_0r1d[9], inp_1r1d[9], inp_2r1d[9]);
  OR3 I16 (out_0r1d[10], inp_0r1d[10], inp_1r1d[10], inp_2r1d[10]);
  OR3 I17 (out_0r1d[11], inp_0r1d[11], inp_1r1d[11], inp_2r1d[11]);
  OR3 I18 (out_0r1d[12], inp_0r1d[12], inp_1r1d[12], inp_2r1d[12]);
  OR3 I19 (out_0r1d[13], inp_0r1d[13], inp_1r1d[13], inp_2r1d[13]);
  OR3 I20 (out_0r1d[14], inp_0r1d[14], inp_1r1d[14], inp_2r1d[14]);
  OR3 I21 (out_0r1d[15], inp_0r1d[15], inp_1r1d[15], inp_2r1d[15]);
  OR3 I22 (out_0r1d[16], inp_0r1d[16], inp_1r1d[16], inp_2r1d[16]);
  OR3 I23 (out_0r1d[17], inp_0r1d[17], inp_1r1d[17], inp_2r1d[17]);
  OR3 I24 (out_0r1d[18], inp_0r1d[18], inp_1r1d[18], inp_2r1d[18]);
  OR3 I25 (out_0r1d[19], inp_0r1d[19], inp_1r1d[19], inp_2r1d[19]);
  OR3 I26 (out_0r1d[20], inp_0r1d[20], inp_1r1d[20], inp_2r1d[20]);
  OR3 I27 (out_0r1d[21], inp_0r1d[21], inp_1r1d[21], inp_2r1d[21]);
  OR3 I28 (out_0r1d[22], inp_0r1d[22], inp_1r1d[22], inp_2r1d[22]);
  OR3 I29 (out_0r1d[23], inp_0r1d[23], inp_1r1d[23], inp_2r1d[23]);
  OR3 I30 (out_0r1d[24], inp_0r1d[24], inp_1r1d[24], inp_2r1d[24]);
  OR3 I31 (out_0r1d[25], inp_0r1d[25], inp_1r1d[25], inp_2r1d[25]);
  OR3 I32 (out_0r1d[26], inp_0r1d[26], inp_1r1d[26], inp_2r1d[26]);
  OR3 I33 (out_0r1d[27], inp_0r1d[27], inp_1r1d[27], inp_2r1d[27]);
  OR3 I34 (out_0r1d[28], inp_0r1d[28], inp_1r1d[28], inp_2r1d[28]);
  OR3 I35 (out_0r1d[29], inp_0r1d[29], inp_1r1d[29], inp_2r1d[29]);
  OR3 I36 (out_0r1d[30], inp_0r1d[30], inp_1r1d[30], inp_2r1d[30]);
  OR3 I37 (out_0r1d[31], inp_0r1d[31], inp_1r1d[31], inp_2r1d[31]);
  OR3 I38 (out_0r0d[0], inp_0r0d[0], inp_1r0d[0], inp_2r0d[0]);
  OR3 I39 (out_0r0d[1], inp_0r0d[1], inp_1r0d[1], inp_2r0d[1]);
  OR3 I40 (out_0r0d[2], inp_0r0d[2], inp_1r0d[2], inp_2r0d[2]);
  OR3 I41 (out_0r0d[3], inp_0r0d[3], inp_1r0d[3], inp_2r0d[3]);
  OR3 I42 (out_0r0d[4], inp_0r0d[4], inp_1r0d[4], inp_2r0d[4]);
  OR3 I43 (out_0r0d[5], inp_0r0d[5], inp_1r0d[5], inp_2r0d[5]);
  OR3 I44 (out_0r0d[6], inp_0r0d[6], inp_1r0d[6], inp_2r0d[6]);
  OR3 I45 (out_0r0d[7], inp_0r0d[7], inp_1r0d[7], inp_2r0d[7]);
  OR3 I46 (out_0r0d[8], inp_0r0d[8], inp_1r0d[8], inp_2r0d[8]);
  OR3 I47 (out_0r0d[9], inp_0r0d[9], inp_1r0d[9], inp_2r0d[9]);
  OR3 I48 (out_0r0d[10], inp_0r0d[10], inp_1r0d[10], inp_2r0d[10]);
  OR3 I49 (out_0r0d[11], inp_0r0d[11], inp_1r0d[11], inp_2r0d[11]);
  OR3 I50 (out_0r0d[12], inp_0r0d[12], inp_1r0d[12], inp_2r0d[12]);
  OR3 I51 (out_0r0d[13], inp_0r0d[13], inp_1r0d[13], inp_2r0d[13]);
  OR3 I52 (out_0r0d[14], inp_0r0d[14], inp_1r0d[14], inp_2r0d[14]);
  OR3 I53 (out_0r0d[15], inp_0r0d[15], inp_1r0d[15], inp_2r0d[15]);
  OR3 I54 (out_0r0d[16], inp_0r0d[16], inp_1r0d[16], inp_2r0d[16]);
  OR3 I55 (out_0r0d[17], inp_0r0d[17], inp_1r0d[17], inp_2r0d[17]);
  OR3 I56 (out_0r0d[18], inp_0r0d[18], inp_1r0d[18], inp_2r0d[18]);
  OR3 I57 (out_0r0d[19], inp_0r0d[19], inp_1r0d[19], inp_2r0d[19]);
  OR3 I58 (out_0r0d[20], inp_0r0d[20], inp_1r0d[20], inp_2r0d[20]);
  OR3 I59 (out_0r0d[21], inp_0r0d[21], inp_1r0d[21], inp_2r0d[21]);
  OR3 I60 (out_0r0d[22], inp_0r0d[22], inp_1r0d[22], inp_2r0d[22]);
  OR3 I61 (out_0r0d[23], inp_0r0d[23], inp_1r0d[23], inp_2r0d[23]);
  OR3 I62 (out_0r0d[24], inp_0r0d[24], inp_1r0d[24], inp_2r0d[24]);
  OR3 I63 (out_0r0d[25], inp_0r0d[25], inp_1r0d[25], inp_2r0d[25]);
  OR3 I64 (out_0r0d[26], inp_0r0d[26], inp_1r0d[26], inp_2r0d[26]);
  OR3 I65 (out_0r0d[27], inp_0r0d[27], inp_1r0d[27], inp_2r0d[27]);
  OR3 I66 (out_0r0d[28], inp_0r0d[28], inp_1r0d[28], inp_2r0d[28]);
  OR3 I67 (out_0r0d[29], inp_0r0d[29], inp_1r0d[29], inp_2r0d[29]);
  OR3 I68 (out_0r0d[30], inp_0r0d[30], inp_1r0d[30], inp_2r0d[30]);
  OR3 I69 (out_0r0d[31], inp_0r0d[31], inp_1r0d[31], inp_2r0d[31]);
endmodule

module BrzCallMux_35_2 (
  inp_0r0d, inp_0r1d, inp_0a,
  inp_1r0d, inp_1r1d, inp_1a,
  out_0r0d, out_0r1d, out_0a
);
  input [34:0] inp_0r0d;
  input [34:0] inp_0r1d;
  output inp_0a;
  input [34:0] inp_1r0d;
  input [34:0] inp_1r1d;
  output inp_1a;
  output [34:0] out_0r0d;
  output [34:0] out_0r1d;
  input out_0a;
  wire [1:0] sourceId_0n;
  C2 I0 (inp_0a, sourceId_0n[0], out_0a);
  C2 I1 (inp_1a, sourceId_0n[1], out_0a);
  OR2 I2 (sourceId_0n[0], inp_0r0d[0], inp_0r1d[0]);
  OR2 I3 (sourceId_0n[1], inp_1r0d[0], inp_1r1d[0]);
  OR2 I4 (out_0r1d[0], inp_0r1d[0], inp_1r1d[0]);
  OR2 I5 (out_0r1d[1], inp_0r1d[1], inp_1r1d[1]);
  OR2 I6 (out_0r1d[2], inp_0r1d[2], inp_1r1d[2]);
  OR2 I7 (out_0r1d[3], inp_0r1d[3], inp_1r1d[3]);
  OR2 I8 (out_0r1d[4], inp_0r1d[4], inp_1r1d[4]);
  OR2 I9 (out_0r1d[5], inp_0r1d[5], inp_1r1d[5]);
  OR2 I10 (out_0r1d[6], inp_0r1d[6], inp_1r1d[6]);
  OR2 I11 (out_0r1d[7], inp_0r1d[7], inp_1r1d[7]);
  OR2 I12 (out_0r1d[8], inp_0r1d[8], inp_1r1d[8]);
  OR2 I13 (out_0r1d[9], inp_0r1d[9], inp_1r1d[9]);
  OR2 I14 (out_0r1d[10], inp_0r1d[10], inp_1r1d[10]);
  OR2 I15 (out_0r1d[11], inp_0r1d[11], inp_1r1d[11]);
  OR2 I16 (out_0r1d[12], inp_0r1d[12], inp_1r1d[12]);
  OR2 I17 (out_0r1d[13], inp_0r1d[13], inp_1r1d[13]);
  OR2 I18 (out_0r1d[14], inp_0r1d[14], inp_1r1d[14]);
  OR2 I19 (out_0r1d[15], inp_0r1d[15], inp_1r1d[15]);
  OR2 I20 (out_0r1d[16], inp_0r1d[16], inp_1r1d[16]);
  OR2 I21 (out_0r1d[17], inp_0r1d[17], inp_1r1d[17]);
  OR2 I22 (out_0r1d[18], inp_0r1d[18], inp_1r1d[18]);
  OR2 I23 (out_0r1d[19], inp_0r1d[19], inp_1r1d[19]);
  OR2 I24 (out_0r1d[20], inp_0r1d[20], inp_1r1d[20]);
  OR2 I25 (out_0r1d[21], inp_0r1d[21], inp_1r1d[21]);
  OR2 I26 (out_0r1d[22], inp_0r1d[22], inp_1r1d[22]);
  OR2 I27 (out_0r1d[23], inp_0r1d[23], inp_1r1d[23]);
  OR2 I28 (out_0r1d[24], inp_0r1d[24], inp_1r1d[24]);
  OR2 I29 (out_0r1d[25], inp_0r1d[25], inp_1r1d[25]);
  OR2 I30 (out_0r1d[26], inp_0r1d[26], inp_1r1d[26]);
  OR2 I31 (out_0r1d[27], inp_0r1d[27], inp_1r1d[27]);
  OR2 I32 (out_0r1d[28], inp_0r1d[28], inp_1r1d[28]);
  OR2 I33 (out_0r1d[29], inp_0r1d[29], inp_1r1d[29]);
  OR2 I34 (out_0r1d[30], inp_0r1d[30], inp_1r1d[30]);
  OR2 I35 (out_0r1d[31], inp_0r1d[31], inp_1r1d[31]);
  OR2 I36 (out_0r1d[32], inp_0r1d[32], inp_1r1d[32]);
  OR2 I37 (out_0r1d[33], inp_0r1d[33], inp_1r1d[33]);
  OR2 I38 (out_0r1d[34], inp_0r1d[34], inp_1r1d[34]);
  OR2 I39 (out_0r0d[0], inp_0r0d[0], inp_1r0d[0]);
  OR2 I40 (out_0r0d[1], inp_0r0d[1], inp_1r0d[1]);
  OR2 I41 (out_0r0d[2], inp_0r0d[2], inp_1r0d[2]);
  OR2 I42 (out_0r0d[3], inp_0r0d[3], inp_1r0d[3]);
  OR2 I43 (out_0r0d[4], inp_0r0d[4], inp_1r0d[4]);
  OR2 I44 (out_0r0d[5], inp_0r0d[5], inp_1r0d[5]);
  OR2 I45 (out_0r0d[6], inp_0r0d[6], inp_1r0d[6]);
  OR2 I46 (out_0r0d[7], inp_0r0d[7], inp_1r0d[7]);
  OR2 I47 (out_0r0d[8], inp_0r0d[8], inp_1r0d[8]);
  OR2 I48 (out_0r0d[9], inp_0r0d[9], inp_1r0d[9]);
  OR2 I49 (out_0r0d[10], inp_0r0d[10], inp_1r0d[10]);
  OR2 I50 (out_0r0d[11], inp_0r0d[11], inp_1r0d[11]);
  OR2 I51 (out_0r0d[12], inp_0r0d[12], inp_1r0d[12]);
  OR2 I52 (out_0r0d[13], inp_0r0d[13], inp_1r0d[13]);
  OR2 I53 (out_0r0d[14], inp_0r0d[14], inp_1r0d[14]);
  OR2 I54 (out_0r0d[15], inp_0r0d[15], inp_1r0d[15]);
  OR2 I55 (out_0r0d[16], inp_0r0d[16], inp_1r0d[16]);
  OR2 I56 (out_0r0d[17], inp_0r0d[17], inp_1r0d[17]);
  OR2 I57 (out_0r0d[18], inp_0r0d[18], inp_1r0d[18]);
  OR2 I58 (out_0r0d[19], inp_0r0d[19], inp_1r0d[19]);
  OR2 I59 (out_0r0d[20], inp_0r0d[20], inp_1r0d[20]);
  OR2 I60 (out_0r0d[21], inp_0r0d[21], inp_1r0d[21]);
  OR2 I61 (out_0r0d[22], inp_0r0d[22], inp_1r0d[22]);
  OR2 I62 (out_0r0d[23], inp_0r0d[23], inp_1r0d[23]);
  OR2 I63 (out_0r0d[24], inp_0r0d[24], inp_1r0d[24]);
  OR2 I64 (out_0r0d[25], inp_0r0d[25], inp_1r0d[25]);
  OR2 I65 (out_0r0d[26], inp_0r0d[26], inp_1r0d[26]);
  OR2 I66 (out_0r0d[27], inp_0r0d[27], inp_1r0d[27]);
  OR2 I67 (out_0r0d[28], inp_0r0d[28], inp_1r0d[28]);
  OR2 I68 (out_0r0d[29], inp_0r0d[29], inp_1r0d[29]);
  OR2 I69 (out_0r0d[30], inp_0r0d[30], inp_1r0d[30]);
  OR2 I70 (out_0r0d[31], inp_0r0d[31], inp_1r0d[31]);
  OR2 I71 (out_0r0d[32], inp_0r0d[32], inp_1r0d[32]);
  OR2 I72 (out_0r0d[33], inp_0r0d[33], inp_1r0d[33]);
  OR2 I73 (out_0r0d[34], inp_0r0d[34], inp_1r0d[34]);
endmodule

module BrzCallMux_35_9 (
  inp_0r0d, inp_0r1d, inp_0a,
  inp_1r0d, inp_1r1d, inp_1a,
  inp_2r0d, inp_2r1d, inp_2a,
  inp_3r0d, inp_3r1d, inp_3a,
  inp_4r0d, inp_4r1d, inp_4a,
  inp_5r0d, inp_5r1d, inp_5a,
  inp_6r0d, inp_6r1d, inp_6a,
  inp_7r0d, inp_7r1d, inp_7a,
  inp_8r0d, inp_8r1d, inp_8a,
  out_0r0d, out_0r1d, out_0a
);
  input [34:0] inp_0r0d;
  input [34:0] inp_0r1d;
  output inp_0a;
  input [34:0] inp_1r0d;
  input [34:0] inp_1r1d;
  output inp_1a;
  input [34:0] inp_2r0d;
  input [34:0] inp_2r1d;
  output inp_2a;
  input [34:0] inp_3r0d;
  input [34:0] inp_3r1d;
  output inp_3a;
  input [34:0] inp_4r0d;
  input [34:0] inp_4r1d;
  output inp_4a;
  input [34:0] inp_5r0d;
  input [34:0] inp_5r1d;
  output inp_5a;
  input [34:0] inp_6r0d;
  input [34:0] inp_6r1d;
  output inp_6a;
  input [34:0] inp_7r0d;
  input [34:0] inp_7r1d;
  output inp_7a;
  input [34:0] inp_8r0d;
  input [34:0] inp_8r1d;
  output inp_8a;
  output [34:0] out_0r0d;
  output [34:0] out_0r1d;
  input out_0a;
  wire [209:0] internal_0n;
  wire [8:0] sourceId_0n;
  C2 I0 (inp_0a, sourceId_0n[0], out_0a);
  C2 I1 (inp_1a, sourceId_0n[1], out_0a);
  C2 I2 (inp_2a, sourceId_0n[2], out_0a);
  C2 I3 (inp_3a, sourceId_0n[3], out_0a);
  C2 I4 (inp_4a, sourceId_0n[4], out_0a);
  C2 I5 (inp_5a, sourceId_0n[5], out_0a);
  C2 I6 (inp_6a, sourceId_0n[6], out_0a);
  C2 I7 (inp_7a, sourceId_0n[7], out_0a);
  C2 I8 (inp_8a, sourceId_0n[8], out_0a);
  OR2 I9 (sourceId_0n[0], inp_0r0d[0], inp_0r1d[0]);
  OR2 I10 (sourceId_0n[1], inp_1r0d[0], inp_1r1d[0]);
  OR2 I11 (sourceId_0n[2], inp_2r0d[0], inp_2r1d[0]);
  OR2 I12 (sourceId_0n[3], inp_3r0d[0], inp_3r1d[0]);
  OR2 I13 (sourceId_0n[4], inp_4r0d[0], inp_4r1d[0]);
  OR2 I14 (sourceId_0n[5], inp_5r0d[0], inp_5r1d[0]);
  OR2 I15 (sourceId_0n[6], inp_6r0d[0], inp_6r1d[0]);
  OR2 I16 (sourceId_0n[7], inp_7r0d[0], inp_7r1d[0]);
  OR2 I17 (sourceId_0n[8], inp_8r0d[0], inp_8r1d[0]);
  NOR3 I18 (internal_0n[0], inp_0r1d[0], inp_1r1d[0], inp_2r1d[0]);
  NOR3 I19 (internal_0n[1], inp_3r1d[0], inp_4r1d[0], inp_5r1d[0]);
  NOR3 I20 (internal_0n[2], inp_6r1d[0], inp_7r1d[0], inp_8r1d[0]);
  NAND3 I21 (out_0r1d[0], internal_0n[0], internal_0n[1], internal_0n[2]);
  NOR3 I22 (internal_0n[3], inp_0r1d[1], inp_1r1d[1], inp_2r1d[1]);
  NOR3 I23 (internal_0n[4], inp_3r1d[1], inp_4r1d[1], inp_5r1d[1]);
  NOR3 I24 (internal_0n[5], inp_6r1d[1], inp_7r1d[1], inp_8r1d[1]);
  NAND3 I25 (out_0r1d[1], internal_0n[3], internal_0n[4], internal_0n[5]);
  NOR3 I26 (internal_0n[6], inp_0r1d[2], inp_1r1d[2], inp_2r1d[2]);
  NOR3 I27 (internal_0n[7], inp_3r1d[2], inp_4r1d[2], inp_5r1d[2]);
  NOR3 I28 (internal_0n[8], inp_6r1d[2], inp_7r1d[2], inp_8r1d[2]);
  NAND3 I29 (out_0r1d[2], internal_0n[6], internal_0n[7], internal_0n[8]);
  NOR3 I30 (internal_0n[9], inp_0r1d[3], inp_1r1d[3], inp_2r1d[3]);
  NOR3 I31 (internal_0n[10], inp_3r1d[3], inp_4r1d[3], inp_5r1d[3]);
  NOR3 I32 (internal_0n[11], inp_6r1d[3], inp_7r1d[3], inp_8r1d[3]);
  NAND3 I33 (out_0r1d[3], internal_0n[9], internal_0n[10], internal_0n[11]);
  NOR3 I34 (internal_0n[12], inp_0r1d[4], inp_1r1d[4], inp_2r1d[4]);
  NOR3 I35 (internal_0n[13], inp_3r1d[4], inp_4r1d[4], inp_5r1d[4]);
  NOR3 I36 (internal_0n[14], inp_6r1d[4], inp_7r1d[4], inp_8r1d[4]);
  NAND3 I37 (out_0r1d[4], internal_0n[12], internal_0n[13], internal_0n[14]);
  NOR3 I38 (internal_0n[15], inp_0r1d[5], inp_1r1d[5], inp_2r1d[5]);
  NOR3 I39 (internal_0n[16], inp_3r1d[5], inp_4r1d[5], inp_5r1d[5]);
  NOR3 I40 (internal_0n[17], inp_6r1d[5], inp_7r1d[5], inp_8r1d[5]);
  NAND3 I41 (out_0r1d[5], internal_0n[15], internal_0n[16], internal_0n[17]);
  NOR3 I42 (internal_0n[18], inp_0r1d[6], inp_1r1d[6], inp_2r1d[6]);
  NOR3 I43 (internal_0n[19], inp_3r1d[6], inp_4r1d[6], inp_5r1d[6]);
  NOR3 I44 (internal_0n[20], inp_6r1d[6], inp_7r1d[6], inp_8r1d[6]);
  NAND3 I45 (out_0r1d[6], internal_0n[18], internal_0n[19], internal_0n[20]);
  NOR3 I46 (internal_0n[21], inp_0r1d[7], inp_1r1d[7], inp_2r1d[7]);
  NOR3 I47 (internal_0n[22], inp_3r1d[7], inp_4r1d[7], inp_5r1d[7]);
  NOR3 I48 (internal_0n[23], inp_6r1d[7], inp_7r1d[7], inp_8r1d[7]);
  NAND3 I49 (out_0r1d[7], internal_0n[21], internal_0n[22], internal_0n[23]);
  NOR3 I50 (internal_0n[24], inp_0r1d[8], inp_1r1d[8], inp_2r1d[8]);
  NOR3 I51 (internal_0n[25], inp_3r1d[8], inp_4r1d[8], inp_5r1d[8]);
  NOR3 I52 (internal_0n[26], inp_6r1d[8], inp_7r1d[8], inp_8r1d[8]);
  NAND3 I53 (out_0r1d[8], internal_0n[24], internal_0n[25], internal_0n[26]);
  NOR3 I54 (internal_0n[27], inp_0r1d[9], inp_1r1d[9], inp_2r1d[9]);
  NOR3 I55 (internal_0n[28], inp_3r1d[9], inp_4r1d[9], inp_5r1d[9]);
  NOR3 I56 (internal_0n[29], inp_6r1d[9], inp_7r1d[9], inp_8r1d[9]);
  NAND3 I57 (out_0r1d[9], internal_0n[27], internal_0n[28], internal_0n[29]);
  NOR3 I58 (internal_0n[30], inp_0r1d[10], inp_1r1d[10], inp_2r1d[10]);
  NOR3 I59 (internal_0n[31], inp_3r1d[10], inp_4r1d[10], inp_5r1d[10]);
  NOR3 I60 (internal_0n[32], inp_6r1d[10], inp_7r1d[10], inp_8r1d[10]);
  NAND3 I61 (out_0r1d[10], internal_0n[30], internal_0n[31], internal_0n[32]);
  NOR3 I62 (internal_0n[33], inp_0r1d[11], inp_1r1d[11], inp_2r1d[11]);
  NOR3 I63 (internal_0n[34], inp_3r1d[11], inp_4r1d[11], inp_5r1d[11]);
  NOR3 I64 (internal_0n[35], inp_6r1d[11], inp_7r1d[11], inp_8r1d[11]);
  NAND3 I65 (out_0r1d[11], internal_0n[33], internal_0n[34], internal_0n[35]);
  NOR3 I66 (internal_0n[36], inp_0r1d[12], inp_1r1d[12], inp_2r1d[12]);
  NOR3 I67 (internal_0n[37], inp_3r1d[12], inp_4r1d[12], inp_5r1d[12]);
  NOR3 I68 (internal_0n[38], inp_6r1d[12], inp_7r1d[12], inp_8r1d[12]);
  NAND3 I69 (out_0r1d[12], internal_0n[36], internal_0n[37], internal_0n[38]);
  NOR3 I70 (internal_0n[39], inp_0r1d[13], inp_1r1d[13], inp_2r1d[13]);
  NOR3 I71 (internal_0n[40], inp_3r1d[13], inp_4r1d[13], inp_5r1d[13]);
  NOR3 I72 (internal_0n[41], inp_6r1d[13], inp_7r1d[13], inp_8r1d[13]);
  NAND3 I73 (out_0r1d[13], internal_0n[39], internal_0n[40], internal_0n[41]);
  NOR3 I74 (internal_0n[42], inp_0r1d[14], inp_1r1d[14], inp_2r1d[14]);
  NOR3 I75 (internal_0n[43], inp_3r1d[14], inp_4r1d[14], inp_5r1d[14]);
  NOR3 I76 (internal_0n[44], inp_6r1d[14], inp_7r1d[14], inp_8r1d[14]);
  NAND3 I77 (out_0r1d[14], internal_0n[42], internal_0n[43], internal_0n[44]);
  NOR3 I78 (internal_0n[45], inp_0r1d[15], inp_1r1d[15], inp_2r1d[15]);
  NOR3 I79 (internal_0n[46], inp_3r1d[15], inp_4r1d[15], inp_5r1d[15]);
  NOR3 I80 (internal_0n[47], inp_6r1d[15], inp_7r1d[15], inp_8r1d[15]);
  NAND3 I81 (out_0r1d[15], internal_0n[45], internal_0n[46], internal_0n[47]);
  NOR3 I82 (internal_0n[48], inp_0r1d[16], inp_1r1d[16], inp_2r1d[16]);
  NOR3 I83 (internal_0n[49], inp_3r1d[16], inp_4r1d[16], inp_5r1d[16]);
  NOR3 I84 (internal_0n[50], inp_6r1d[16], inp_7r1d[16], inp_8r1d[16]);
  NAND3 I85 (out_0r1d[16], internal_0n[48], internal_0n[49], internal_0n[50]);
  NOR3 I86 (internal_0n[51], inp_0r1d[17], inp_1r1d[17], inp_2r1d[17]);
  NOR3 I87 (internal_0n[52], inp_3r1d[17], inp_4r1d[17], inp_5r1d[17]);
  NOR3 I88 (internal_0n[53], inp_6r1d[17], inp_7r1d[17], inp_8r1d[17]);
  NAND3 I89 (out_0r1d[17], internal_0n[51], internal_0n[52], internal_0n[53]);
  NOR3 I90 (internal_0n[54], inp_0r1d[18], inp_1r1d[18], inp_2r1d[18]);
  NOR3 I91 (internal_0n[55], inp_3r1d[18], inp_4r1d[18], inp_5r1d[18]);
  NOR3 I92 (internal_0n[56], inp_6r1d[18], inp_7r1d[18], inp_8r1d[18]);
  NAND3 I93 (out_0r1d[18], internal_0n[54], internal_0n[55], internal_0n[56]);
  NOR3 I94 (internal_0n[57], inp_0r1d[19], inp_1r1d[19], inp_2r1d[19]);
  NOR3 I95 (internal_0n[58], inp_3r1d[19], inp_4r1d[19], inp_5r1d[19]);
  NOR3 I96 (internal_0n[59], inp_6r1d[19], inp_7r1d[19], inp_8r1d[19]);
  NAND3 I97 (out_0r1d[19], internal_0n[57], internal_0n[58], internal_0n[59]);
  NOR3 I98 (internal_0n[60], inp_0r1d[20], inp_1r1d[20], inp_2r1d[20]);
  NOR3 I99 (internal_0n[61], inp_3r1d[20], inp_4r1d[20], inp_5r1d[20]);
  NOR3 I100 (internal_0n[62], inp_6r1d[20], inp_7r1d[20], inp_8r1d[20]);
  NAND3 I101 (out_0r1d[20], internal_0n[60], internal_0n[61], internal_0n[62]);
  NOR3 I102 (internal_0n[63], inp_0r1d[21], inp_1r1d[21], inp_2r1d[21]);
  NOR3 I103 (internal_0n[64], inp_3r1d[21], inp_4r1d[21], inp_5r1d[21]);
  NOR3 I104 (internal_0n[65], inp_6r1d[21], inp_7r1d[21], inp_8r1d[21]);
  NAND3 I105 (out_0r1d[21], internal_0n[63], internal_0n[64], internal_0n[65]);
  NOR3 I106 (internal_0n[66], inp_0r1d[22], inp_1r1d[22], inp_2r1d[22]);
  NOR3 I107 (internal_0n[67], inp_3r1d[22], inp_4r1d[22], inp_5r1d[22]);
  NOR3 I108 (internal_0n[68], inp_6r1d[22], inp_7r1d[22], inp_8r1d[22]);
  NAND3 I109 (out_0r1d[22], internal_0n[66], internal_0n[67], internal_0n[68]);
  NOR3 I110 (internal_0n[69], inp_0r1d[23], inp_1r1d[23], inp_2r1d[23]);
  NOR3 I111 (internal_0n[70], inp_3r1d[23], inp_4r1d[23], inp_5r1d[23]);
  NOR3 I112 (internal_0n[71], inp_6r1d[23], inp_7r1d[23], inp_8r1d[23]);
  NAND3 I113 (out_0r1d[23], internal_0n[69], internal_0n[70], internal_0n[71]);
  NOR3 I114 (internal_0n[72], inp_0r1d[24], inp_1r1d[24], inp_2r1d[24]);
  NOR3 I115 (internal_0n[73], inp_3r1d[24], inp_4r1d[24], inp_5r1d[24]);
  NOR3 I116 (internal_0n[74], inp_6r1d[24], inp_7r1d[24], inp_8r1d[24]);
  NAND3 I117 (out_0r1d[24], internal_0n[72], internal_0n[73], internal_0n[74]);
  NOR3 I118 (internal_0n[75], inp_0r1d[25], inp_1r1d[25], inp_2r1d[25]);
  NOR3 I119 (internal_0n[76], inp_3r1d[25], inp_4r1d[25], inp_5r1d[25]);
  NOR3 I120 (internal_0n[77], inp_6r1d[25], inp_7r1d[25], inp_8r1d[25]);
  NAND3 I121 (out_0r1d[25], internal_0n[75], internal_0n[76], internal_0n[77]);
  NOR3 I122 (internal_0n[78], inp_0r1d[26], inp_1r1d[26], inp_2r1d[26]);
  NOR3 I123 (internal_0n[79], inp_3r1d[26], inp_4r1d[26], inp_5r1d[26]);
  NOR3 I124 (internal_0n[80], inp_6r1d[26], inp_7r1d[26], inp_8r1d[26]);
  NAND3 I125 (out_0r1d[26], internal_0n[78], internal_0n[79], internal_0n[80]);
  NOR3 I126 (internal_0n[81], inp_0r1d[27], inp_1r1d[27], inp_2r1d[27]);
  NOR3 I127 (internal_0n[82], inp_3r1d[27], inp_4r1d[27], inp_5r1d[27]);
  NOR3 I128 (internal_0n[83], inp_6r1d[27], inp_7r1d[27], inp_8r1d[27]);
  NAND3 I129 (out_0r1d[27], internal_0n[81], internal_0n[82], internal_0n[83]);
  NOR3 I130 (internal_0n[84], inp_0r1d[28], inp_1r1d[28], inp_2r1d[28]);
  NOR3 I131 (internal_0n[85], inp_3r1d[28], inp_4r1d[28], inp_5r1d[28]);
  NOR3 I132 (internal_0n[86], inp_6r1d[28], inp_7r1d[28], inp_8r1d[28]);
  NAND3 I133 (out_0r1d[28], internal_0n[84], internal_0n[85], internal_0n[86]);
  NOR3 I134 (internal_0n[87], inp_0r1d[29], inp_1r1d[29], inp_2r1d[29]);
  NOR3 I135 (internal_0n[88], inp_3r1d[29], inp_4r1d[29], inp_5r1d[29]);
  NOR3 I136 (internal_0n[89], inp_6r1d[29], inp_7r1d[29], inp_8r1d[29]);
  NAND3 I137 (out_0r1d[29], internal_0n[87], internal_0n[88], internal_0n[89]);
  NOR3 I138 (internal_0n[90], inp_0r1d[30], inp_1r1d[30], inp_2r1d[30]);
  NOR3 I139 (internal_0n[91], inp_3r1d[30], inp_4r1d[30], inp_5r1d[30]);
  NOR3 I140 (internal_0n[92], inp_6r1d[30], inp_7r1d[30], inp_8r1d[30]);
  NAND3 I141 (out_0r1d[30], internal_0n[90], internal_0n[91], internal_0n[92]);
  NOR3 I142 (internal_0n[93], inp_0r1d[31], inp_1r1d[31], inp_2r1d[31]);
  NOR3 I143 (internal_0n[94], inp_3r1d[31], inp_4r1d[31], inp_5r1d[31]);
  NOR3 I144 (internal_0n[95], inp_6r1d[31], inp_7r1d[31], inp_8r1d[31]);
  NAND3 I145 (out_0r1d[31], internal_0n[93], internal_0n[94], internal_0n[95]);
  NOR3 I146 (internal_0n[96], inp_0r1d[32], inp_1r1d[32], inp_2r1d[32]);
  NOR3 I147 (internal_0n[97], inp_3r1d[32], inp_4r1d[32], inp_5r1d[32]);
  NOR3 I148 (internal_0n[98], inp_6r1d[32], inp_7r1d[32], inp_8r1d[32]);
  NAND3 I149 (out_0r1d[32], internal_0n[96], internal_0n[97], internal_0n[98]);
  NOR3 I150 (internal_0n[99], inp_0r1d[33], inp_1r1d[33], inp_2r1d[33]);
  NOR3 I151 (internal_0n[100], inp_3r1d[33], inp_4r1d[33], inp_5r1d[33]);
  NOR3 I152 (internal_0n[101], inp_6r1d[33], inp_7r1d[33], inp_8r1d[33]);
  NAND3 I153 (out_0r1d[33], internal_0n[99], internal_0n[100], internal_0n[101]);
  NOR3 I154 (internal_0n[102], inp_0r1d[34], inp_1r1d[34], inp_2r1d[34]);
  NOR3 I155 (internal_0n[103], inp_3r1d[34], inp_4r1d[34], inp_5r1d[34]);
  NOR3 I156 (internal_0n[104], inp_6r1d[34], inp_7r1d[34], inp_8r1d[34]);
  NAND3 I157 (out_0r1d[34], internal_0n[102], internal_0n[103], internal_0n[104]);
  NOR3 I158 (internal_0n[105], inp_0r0d[0], inp_1r0d[0], inp_2r0d[0]);
  NOR3 I159 (internal_0n[106], inp_3r0d[0], inp_4r0d[0], inp_5r0d[0]);
  NOR3 I160 (internal_0n[107], inp_6r0d[0], inp_7r0d[0], inp_8r0d[0]);
  NAND3 I161 (out_0r0d[0], internal_0n[105], internal_0n[106], internal_0n[107]);
  NOR3 I162 (internal_0n[108], inp_0r0d[1], inp_1r0d[1], inp_2r0d[1]);
  NOR3 I163 (internal_0n[109], inp_3r0d[1], inp_4r0d[1], inp_5r0d[1]);
  NOR3 I164 (internal_0n[110], inp_6r0d[1], inp_7r0d[1], inp_8r0d[1]);
  NAND3 I165 (out_0r0d[1], internal_0n[108], internal_0n[109], internal_0n[110]);
  NOR3 I166 (internal_0n[111], inp_0r0d[2], inp_1r0d[2], inp_2r0d[2]);
  NOR3 I167 (internal_0n[112], inp_3r0d[2], inp_4r0d[2], inp_5r0d[2]);
  NOR3 I168 (internal_0n[113], inp_6r0d[2], inp_7r0d[2], inp_8r0d[2]);
  NAND3 I169 (out_0r0d[2], internal_0n[111], internal_0n[112], internal_0n[113]);
  NOR3 I170 (internal_0n[114], inp_0r0d[3], inp_1r0d[3], inp_2r0d[3]);
  NOR3 I171 (internal_0n[115], inp_3r0d[3], inp_4r0d[3], inp_5r0d[3]);
  NOR3 I172 (internal_0n[116], inp_6r0d[3], inp_7r0d[3], inp_8r0d[3]);
  NAND3 I173 (out_0r0d[3], internal_0n[114], internal_0n[115], internal_0n[116]);
  NOR3 I174 (internal_0n[117], inp_0r0d[4], inp_1r0d[4], inp_2r0d[4]);
  NOR3 I175 (internal_0n[118], inp_3r0d[4], inp_4r0d[4], inp_5r0d[4]);
  NOR3 I176 (internal_0n[119], inp_6r0d[4], inp_7r0d[4], inp_8r0d[4]);
  NAND3 I177 (out_0r0d[4], internal_0n[117], internal_0n[118], internal_0n[119]);
  NOR3 I178 (internal_0n[120], inp_0r0d[5], inp_1r0d[5], inp_2r0d[5]);
  NOR3 I179 (internal_0n[121], inp_3r0d[5], inp_4r0d[5], inp_5r0d[5]);
  NOR3 I180 (internal_0n[122], inp_6r0d[5], inp_7r0d[5], inp_8r0d[5]);
  NAND3 I181 (out_0r0d[5], internal_0n[120], internal_0n[121], internal_0n[122]);
  NOR3 I182 (internal_0n[123], inp_0r0d[6], inp_1r0d[6], inp_2r0d[6]);
  NOR3 I183 (internal_0n[124], inp_3r0d[6], inp_4r0d[6], inp_5r0d[6]);
  NOR3 I184 (internal_0n[125], inp_6r0d[6], inp_7r0d[6], inp_8r0d[6]);
  NAND3 I185 (out_0r0d[6], internal_0n[123], internal_0n[124], internal_0n[125]);
  NOR3 I186 (internal_0n[126], inp_0r0d[7], inp_1r0d[7], inp_2r0d[7]);
  NOR3 I187 (internal_0n[127], inp_3r0d[7], inp_4r0d[7], inp_5r0d[7]);
  NOR3 I188 (internal_0n[128], inp_6r0d[7], inp_7r0d[7], inp_8r0d[7]);
  NAND3 I189 (out_0r0d[7], internal_0n[126], internal_0n[127], internal_0n[128]);
  NOR3 I190 (internal_0n[129], inp_0r0d[8], inp_1r0d[8], inp_2r0d[8]);
  NOR3 I191 (internal_0n[130], inp_3r0d[8], inp_4r0d[8], inp_5r0d[8]);
  NOR3 I192 (internal_0n[131], inp_6r0d[8], inp_7r0d[8], inp_8r0d[8]);
  NAND3 I193 (out_0r0d[8], internal_0n[129], internal_0n[130], internal_0n[131]);
  NOR3 I194 (internal_0n[132], inp_0r0d[9], inp_1r0d[9], inp_2r0d[9]);
  NOR3 I195 (internal_0n[133], inp_3r0d[9], inp_4r0d[9], inp_5r0d[9]);
  NOR3 I196 (internal_0n[134], inp_6r0d[9], inp_7r0d[9], inp_8r0d[9]);
  NAND3 I197 (out_0r0d[9], internal_0n[132], internal_0n[133], internal_0n[134]);
  NOR3 I198 (internal_0n[135], inp_0r0d[10], inp_1r0d[10], inp_2r0d[10]);
  NOR3 I199 (internal_0n[136], inp_3r0d[10], inp_4r0d[10], inp_5r0d[10]);
  NOR3 I200 (internal_0n[137], inp_6r0d[10], inp_7r0d[10], inp_8r0d[10]);
  NAND3 I201 (out_0r0d[10], internal_0n[135], internal_0n[136], internal_0n[137]);
  NOR3 I202 (internal_0n[138], inp_0r0d[11], inp_1r0d[11], inp_2r0d[11]);
  NOR3 I203 (internal_0n[139], inp_3r0d[11], inp_4r0d[11], inp_5r0d[11]);
  NOR3 I204 (internal_0n[140], inp_6r0d[11], inp_7r0d[11], inp_8r0d[11]);
  NAND3 I205 (out_0r0d[11], internal_0n[138], internal_0n[139], internal_0n[140]);
  NOR3 I206 (internal_0n[141], inp_0r0d[12], inp_1r0d[12], inp_2r0d[12]);
  NOR3 I207 (internal_0n[142], inp_3r0d[12], inp_4r0d[12], inp_5r0d[12]);
  NOR3 I208 (internal_0n[143], inp_6r0d[12], inp_7r0d[12], inp_8r0d[12]);
  NAND3 I209 (out_0r0d[12], internal_0n[141], internal_0n[142], internal_0n[143]);
  NOR3 I210 (internal_0n[144], inp_0r0d[13], inp_1r0d[13], inp_2r0d[13]);
  NOR3 I211 (internal_0n[145], inp_3r0d[13], inp_4r0d[13], inp_5r0d[13]);
  NOR3 I212 (internal_0n[146], inp_6r0d[13], inp_7r0d[13], inp_8r0d[13]);
  NAND3 I213 (out_0r0d[13], internal_0n[144], internal_0n[145], internal_0n[146]);
  NOR3 I214 (internal_0n[147], inp_0r0d[14], inp_1r0d[14], inp_2r0d[14]);
  NOR3 I215 (internal_0n[148], inp_3r0d[14], inp_4r0d[14], inp_5r0d[14]);
  NOR3 I216 (internal_0n[149], inp_6r0d[14], inp_7r0d[14], inp_8r0d[14]);
  NAND3 I217 (out_0r0d[14], internal_0n[147], internal_0n[148], internal_0n[149]);
  NOR3 I218 (internal_0n[150], inp_0r0d[15], inp_1r0d[15], inp_2r0d[15]);
  NOR3 I219 (internal_0n[151], inp_3r0d[15], inp_4r0d[15], inp_5r0d[15]);
  NOR3 I220 (internal_0n[152], inp_6r0d[15], inp_7r0d[15], inp_8r0d[15]);
  NAND3 I221 (out_0r0d[15], internal_0n[150], internal_0n[151], internal_0n[152]);
  NOR3 I222 (internal_0n[153], inp_0r0d[16], inp_1r0d[16], inp_2r0d[16]);
  NOR3 I223 (internal_0n[154], inp_3r0d[16], inp_4r0d[16], inp_5r0d[16]);
  NOR3 I224 (internal_0n[155], inp_6r0d[16], inp_7r0d[16], inp_8r0d[16]);
  NAND3 I225 (out_0r0d[16], internal_0n[153], internal_0n[154], internal_0n[155]);
  NOR3 I226 (internal_0n[156], inp_0r0d[17], inp_1r0d[17], inp_2r0d[17]);
  NOR3 I227 (internal_0n[157], inp_3r0d[17], inp_4r0d[17], inp_5r0d[17]);
  NOR3 I228 (internal_0n[158], inp_6r0d[17], inp_7r0d[17], inp_8r0d[17]);
  NAND3 I229 (out_0r0d[17], internal_0n[156], internal_0n[157], internal_0n[158]);
  NOR3 I230 (internal_0n[159], inp_0r0d[18], inp_1r0d[18], inp_2r0d[18]);
  NOR3 I231 (internal_0n[160], inp_3r0d[18], inp_4r0d[18], inp_5r0d[18]);
  NOR3 I232 (internal_0n[161], inp_6r0d[18], inp_7r0d[18], inp_8r0d[18]);
  NAND3 I233 (out_0r0d[18], internal_0n[159], internal_0n[160], internal_0n[161]);
  NOR3 I234 (internal_0n[162], inp_0r0d[19], inp_1r0d[19], inp_2r0d[19]);
  NOR3 I235 (internal_0n[163], inp_3r0d[19], inp_4r0d[19], inp_5r0d[19]);
  NOR3 I236 (internal_0n[164], inp_6r0d[19], inp_7r0d[19], inp_8r0d[19]);
  NAND3 I237 (out_0r0d[19], internal_0n[162], internal_0n[163], internal_0n[164]);
  NOR3 I238 (internal_0n[165], inp_0r0d[20], inp_1r0d[20], inp_2r0d[20]);
  NOR3 I239 (internal_0n[166], inp_3r0d[20], inp_4r0d[20], inp_5r0d[20]);
  NOR3 I240 (internal_0n[167], inp_6r0d[20], inp_7r0d[20], inp_8r0d[20]);
  NAND3 I241 (out_0r0d[20], internal_0n[165], internal_0n[166], internal_0n[167]);
  NOR3 I242 (internal_0n[168], inp_0r0d[21], inp_1r0d[21], inp_2r0d[21]);
  NOR3 I243 (internal_0n[169], inp_3r0d[21], inp_4r0d[21], inp_5r0d[21]);
  NOR3 I244 (internal_0n[170], inp_6r0d[21], inp_7r0d[21], inp_8r0d[21]);
  NAND3 I245 (out_0r0d[21], internal_0n[168], internal_0n[169], internal_0n[170]);
  NOR3 I246 (internal_0n[171], inp_0r0d[22], inp_1r0d[22], inp_2r0d[22]);
  NOR3 I247 (internal_0n[172], inp_3r0d[22], inp_4r0d[22], inp_5r0d[22]);
  NOR3 I248 (internal_0n[173], inp_6r0d[22], inp_7r0d[22], inp_8r0d[22]);
  NAND3 I249 (out_0r0d[22], internal_0n[171], internal_0n[172], internal_0n[173]);
  NOR3 I250 (internal_0n[174], inp_0r0d[23], inp_1r0d[23], inp_2r0d[23]);
  NOR3 I251 (internal_0n[175], inp_3r0d[23], inp_4r0d[23], inp_5r0d[23]);
  NOR3 I252 (internal_0n[176], inp_6r0d[23], inp_7r0d[23], inp_8r0d[23]);
  NAND3 I253 (out_0r0d[23], internal_0n[174], internal_0n[175], internal_0n[176]);
  NOR3 I254 (internal_0n[177], inp_0r0d[24], inp_1r0d[24], inp_2r0d[24]);
  NOR3 I255 (internal_0n[178], inp_3r0d[24], inp_4r0d[24], inp_5r0d[24]);
  NOR3 I256 (internal_0n[179], inp_6r0d[24], inp_7r0d[24], inp_8r0d[24]);
  NAND3 I257 (out_0r0d[24], internal_0n[177], internal_0n[178], internal_0n[179]);
  NOR3 I258 (internal_0n[180], inp_0r0d[25], inp_1r0d[25], inp_2r0d[25]);
  NOR3 I259 (internal_0n[181], inp_3r0d[25], inp_4r0d[25], inp_5r0d[25]);
  NOR3 I260 (internal_0n[182], inp_6r0d[25], inp_7r0d[25], inp_8r0d[25]);
  NAND3 I261 (out_0r0d[25], internal_0n[180], internal_0n[181], internal_0n[182]);
  NOR3 I262 (internal_0n[183], inp_0r0d[26], inp_1r0d[26], inp_2r0d[26]);
  NOR3 I263 (internal_0n[184], inp_3r0d[26], inp_4r0d[26], inp_5r0d[26]);
  NOR3 I264 (internal_0n[185], inp_6r0d[26], inp_7r0d[26], inp_8r0d[26]);
  NAND3 I265 (out_0r0d[26], internal_0n[183], internal_0n[184], internal_0n[185]);
  NOR3 I266 (internal_0n[186], inp_0r0d[27], inp_1r0d[27], inp_2r0d[27]);
  NOR3 I267 (internal_0n[187], inp_3r0d[27], inp_4r0d[27], inp_5r0d[27]);
  NOR3 I268 (internal_0n[188], inp_6r0d[27], inp_7r0d[27], inp_8r0d[27]);
  NAND3 I269 (out_0r0d[27], internal_0n[186], internal_0n[187], internal_0n[188]);
  NOR3 I270 (internal_0n[189], inp_0r0d[28], inp_1r0d[28], inp_2r0d[28]);
  NOR3 I271 (internal_0n[190], inp_3r0d[28], inp_4r0d[28], inp_5r0d[28]);
  NOR3 I272 (internal_0n[191], inp_6r0d[28], inp_7r0d[28], inp_8r0d[28]);
  NAND3 I273 (out_0r0d[28], internal_0n[189], internal_0n[190], internal_0n[191]);
  NOR3 I274 (internal_0n[192], inp_0r0d[29], inp_1r0d[29], inp_2r0d[29]);
  NOR3 I275 (internal_0n[193], inp_3r0d[29], inp_4r0d[29], inp_5r0d[29]);
  NOR3 I276 (internal_0n[194], inp_6r0d[29], inp_7r0d[29], inp_8r0d[29]);
  NAND3 I277 (out_0r0d[29], internal_0n[192], internal_0n[193], internal_0n[194]);
  NOR3 I278 (internal_0n[195], inp_0r0d[30], inp_1r0d[30], inp_2r0d[30]);
  NOR3 I279 (internal_0n[196], inp_3r0d[30], inp_4r0d[30], inp_5r0d[30]);
  NOR3 I280 (internal_0n[197], inp_6r0d[30], inp_7r0d[30], inp_8r0d[30]);
  NAND3 I281 (out_0r0d[30], internal_0n[195], internal_0n[196], internal_0n[197]);
  NOR3 I282 (internal_0n[198], inp_0r0d[31], inp_1r0d[31], inp_2r0d[31]);
  NOR3 I283 (internal_0n[199], inp_3r0d[31], inp_4r0d[31], inp_5r0d[31]);
  NOR3 I284 (internal_0n[200], inp_6r0d[31], inp_7r0d[31], inp_8r0d[31]);
  NAND3 I285 (out_0r0d[31], internal_0n[198], internal_0n[199], internal_0n[200]);
  NOR3 I286 (internal_0n[201], inp_0r0d[32], inp_1r0d[32], inp_2r0d[32]);
  NOR3 I287 (internal_0n[202], inp_3r0d[32], inp_4r0d[32], inp_5r0d[32]);
  NOR3 I288 (internal_0n[203], inp_6r0d[32], inp_7r0d[32], inp_8r0d[32]);
  NAND3 I289 (out_0r0d[32], internal_0n[201], internal_0n[202], internal_0n[203]);
  NOR3 I290 (internal_0n[204], inp_0r0d[33], inp_1r0d[33], inp_2r0d[33]);
  NOR3 I291 (internal_0n[205], inp_3r0d[33], inp_4r0d[33], inp_5r0d[33]);
  NOR3 I292 (internal_0n[206], inp_6r0d[33], inp_7r0d[33], inp_8r0d[33]);
  NAND3 I293 (out_0r0d[33], internal_0n[204], internal_0n[205], internal_0n[206]);
  NOR3 I294 (internal_0n[207], inp_0r0d[34], inp_1r0d[34], inp_2r0d[34]);
  NOR3 I295 (internal_0n[208], inp_3r0d[34], inp_4r0d[34], inp_5r0d[34]);
  NOR3 I296 (internal_0n[209], inp_6r0d[34], inp_7r0d[34], inp_8r0d[34]);
  NAND3 I297 (out_0r0d[34], internal_0n[207], internal_0n[208], internal_0n[209]);
endmodule

module BrzCallMux_36_2 (
  inp_0r0d, inp_0r1d, inp_0a,
  inp_1r0d, inp_1r1d, inp_1a,
  out_0r0d, out_0r1d, out_0a
);
  input [35:0] inp_0r0d;
  input [35:0] inp_0r1d;
  output inp_0a;
  input [35:0] inp_1r0d;
  input [35:0] inp_1r1d;
  output inp_1a;
  output [35:0] out_0r0d;
  output [35:0] out_0r1d;
  input out_0a;
  wire [1:0] sourceId_0n;
  C2 I0 (inp_0a, sourceId_0n[0], out_0a);
  C2 I1 (inp_1a, sourceId_0n[1], out_0a);
  OR2 I2 (sourceId_0n[0], inp_0r0d[0], inp_0r1d[0]);
  OR2 I3 (sourceId_0n[1], inp_1r0d[0], inp_1r1d[0]);
  OR2 I4 (out_0r1d[0], inp_0r1d[0], inp_1r1d[0]);
  OR2 I5 (out_0r1d[1], inp_0r1d[1], inp_1r1d[1]);
  OR2 I6 (out_0r1d[2], inp_0r1d[2], inp_1r1d[2]);
  OR2 I7 (out_0r1d[3], inp_0r1d[3], inp_1r1d[3]);
  OR2 I8 (out_0r1d[4], inp_0r1d[4], inp_1r1d[4]);
  OR2 I9 (out_0r1d[5], inp_0r1d[5], inp_1r1d[5]);
  OR2 I10 (out_0r1d[6], inp_0r1d[6], inp_1r1d[6]);
  OR2 I11 (out_0r1d[7], inp_0r1d[7], inp_1r1d[7]);
  OR2 I12 (out_0r1d[8], inp_0r1d[8], inp_1r1d[8]);
  OR2 I13 (out_0r1d[9], inp_0r1d[9], inp_1r1d[9]);
  OR2 I14 (out_0r1d[10], inp_0r1d[10], inp_1r1d[10]);
  OR2 I15 (out_0r1d[11], inp_0r1d[11], inp_1r1d[11]);
  OR2 I16 (out_0r1d[12], inp_0r1d[12], inp_1r1d[12]);
  OR2 I17 (out_0r1d[13], inp_0r1d[13], inp_1r1d[13]);
  OR2 I18 (out_0r1d[14], inp_0r1d[14], inp_1r1d[14]);
  OR2 I19 (out_0r1d[15], inp_0r1d[15], inp_1r1d[15]);
  OR2 I20 (out_0r1d[16], inp_0r1d[16], inp_1r1d[16]);
  OR2 I21 (out_0r1d[17], inp_0r1d[17], inp_1r1d[17]);
  OR2 I22 (out_0r1d[18], inp_0r1d[18], inp_1r1d[18]);
  OR2 I23 (out_0r1d[19], inp_0r1d[19], inp_1r1d[19]);
  OR2 I24 (out_0r1d[20], inp_0r1d[20], inp_1r1d[20]);
  OR2 I25 (out_0r1d[21], inp_0r1d[21], inp_1r1d[21]);
  OR2 I26 (out_0r1d[22], inp_0r1d[22], inp_1r1d[22]);
  OR2 I27 (out_0r1d[23], inp_0r1d[23], inp_1r1d[23]);
  OR2 I28 (out_0r1d[24], inp_0r1d[24], inp_1r1d[24]);
  OR2 I29 (out_0r1d[25], inp_0r1d[25], inp_1r1d[25]);
  OR2 I30 (out_0r1d[26], inp_0r1d[26], inp_1r1d[26]);
  OR2 I31 (out_0r1d[27], inp_0r1d[27], inp_1r1d[27]);
  OR2 I32 (out_0r1d[28], inp_0r1d[28], inp_1r1d[28]);
  OR2 I33 (out_0r1d[29], inp_0r1d[29], inp_1r1d[29]);
  OR2 I34 (out_0r1d[30], inp_0r1d[30], inp_1r1d[30]);
  OR2 I35 (out_0r1d[31], inp_0r1d[31], inp_1r1d[31]);
  OR2 I36 (out_0r1d[32], inp_0r1d[32], inp_1r1d[32]);
  OR2 I37 (out_0r1d[33], inp_0r1d[33], inp_1r1d[33]);
  OR2 I38 (out_0r1d[34], inp_0r1d[34], inp_1r1d[34]);
  OR2 I39 (out_0r1d[35], inp_0r1d[35], inp_1r1d[35]);
  OR2 I40 (out_0r0d[0], inp_0r0d[0], inp_1r0d[0]);
  OR2 I41 (out_0r0d[1], inp_0r0d[1], inp_1r0d[1]);
  OR2 I42 (out_0r0d[2], inp_0r0d[2], inp_1r0d[2]);
  OR2 I43 (out_0r0d[3], inp_0r0d[3], inp_1r0d[3]);
  OR2 I44 (out_0r0d[4], inp_0r0d[4], inp_1r0d[4]);
  OR2 I45 (out_0r0d[5], inp_0r0d[5], inp_1r0d[5]);
  OR2 I46 (out_0r0d[6], inp_0r0d[6], inp_1r0d[6]);
  OR2 I47 (out_0r0d[7], inp_0r0d[7], inp_1r0d[7]);
  OR2 I48 (out_0r0d[8], inp_0r0d[8], inp_1r0d[8]);
  OR2 I49 (out_0r0d[9], inp_0r0d[9], inp_1r0d[9]);
  OR2 I50 (out_0r0d[10], inp_0r0d[10], inp_1r0d[10]);
  OR2 I51 (out_0r0d[11], inp_0r0d[11], inp_1r0d[11]);
  OR2 I52 (out_0r0d[12], inp_0r0d[12], inp_1r0d[12]);
  OR2 I53 (out_0r0d[13], inp_0r0d[13], inp_1r0d[13]);
  OR2 I54 (out_0r0d[14], inp_0r0d[14], inp_1r0d[14]);
  OR2 I55 (out_0r0d[15], inp_0r0d[15], inp_1r0d[15]);
  OR2 I56 (out_0r0d[16], inp_0r0d[16], inp_1r0d[16]);
  OR2 I57 (out_0r0d[17], inp_0r0d[17], inp_1r0d[17]);
  OR2 I58 (out_0r0d[18], inp_0r0d[18], inp_1r0d[18]);
  OR2 I59 (out_0r0d[19], inp_0r0d[19], inp_1r0d[19]);
  OR2 I60 (out_0r0d[20], inp_0r0d[20], inp_1r0d[20]);
  OR2 I61 (out_0r0d[21], inp_0r0d[21], inp_1r0d[21]);
  OR2 I62 (out_0r0d[22], inp_0r0d[22], inp_1r0d[22]);
  OR2 I63 (out_0r0d[23], inp_0r0d[23], inp_1r0d[23]);
  OR2 I64 (out_0r0d[24], inp_0r0d[24], inp_1r0d[24]);
  OR2 I65 (out_0r0d[25], inp_0r0d[25], inp_1r0d[25]);
  OR2 I66 (out_0r0d[26], inp_0r0d[26], inp_1r0d[26]);
  OR2 I67 (out_0r0d[27], inp_0r0d[27], inp_1r0d[27]);
  OR2 I68 (out_0r0d[28], inp_0r0d[28], inp_1r0d[28]);
  OR2 I69 (out_0r0d[29], inp_0r0d[29], inp_1r0d[29]);
  OR2 I70 (out_0r0d[30], inp_0r0d[30], inp_1r0d[30]);
  OR2 I71 (out_0r0d[31], inp_0r0d[31], inp_1r0d[31]);
  OR2 I72 (out_0r0d[32], inp_0r0d[32], inp_1r0d[32]);
  OR2 I73 (out_0r0d[33], inp_0r0d[33], inp_1r0d[33]);
  OR2 I74 (out_0r0d[34], inp_0r0d[34], inp_1r0d[34]);
  OR2 I75 (out_0r0d[35], inp_0r0d[35], inp_1r0d[35]);
endmodule

module BrzCase_1_1_s1_1 (
  inp_0r0d, inp_0r1d, inp_0a,
  activateOut_0r, activateOut_0a
);
  input inp_0r0d;
  input inp_0r1d;
  output inp_0a;
  output activateOut_0r;
  input activateOut_0a;
  wire elseAck_0n;
  wire inpComplete_0n;
  wire inpDone_0n;
  wire outDone_0n;
  wire [1:0] int0_0n;
  C2 I0 (inp_0a, outDone_0n, inpDone_0n);
  OR2 I1 (outDone_0n, activateOut_0a, elseAck_0n);
  BUFF I2 (int0_0n[0], inp_0r0d);
  BUFF I3 (int0_0n[1], inp_0r1d);
  BUFF I4 (elseAck_0n, int0_0n[0]);
  BUFF I5 (activateOut_0r, int0_0n[1]);
  BUFF I6 (inpDone_0n, inpComplete_0n);
  OR2 I7 (inpComplete_0n, inp_0r0d, inp_0r1d);
endmodule

module BrzCase_1_2_s5_0_3b1 (
  inp_0r0d, inp_0r1d, inp_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a
);
  input inp_0r0d;
  input inp_0r1d;
  output inp_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  wire elseAck_0n;
  wire inpComplete_0n;
  wire inpDone_0n;
  wire outDone_0n;
  wire [1:0] int0_0n;
  C2 I0 (inp_0a, outDone_0n, inpDone_0n);
  OR2 I1 (outDone_0n, activateOut_0a, activateOut_1a);
  BUFF I2 (int0_0n[0], inp_0r1d);
  BUFF I3 (int0_0n[1], inp_0r0d);
  BUFF I4 (activateOut_1r, int0_0n[0]);
  BUFF I5 (activateOut_0r, int0_0n[1]);
  BUFF I6 (inpDone_0n, inpComplete_0n);
  OR2 I7 (inpComplete_0n, inp_0r0d, inp_0r1d);
endmodule

module BrzCase_3_2_s25_1_2c3m4_2c2m4_3b5_2c4_2c0 (
  inp_0r0d, inp_0r1d, inp_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a
);
  input [2:0] inp_0r0d;
  input [2:0] inp_0r1d;
  output inp_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  wire elseAck_0n;
  wire [2:0] inpComplete_0n;
  wire inpDone_0n;
  wire outDone_0n;
  wire [3:0] int0_0n;
  C2 I0 (inp_0a, outDone_0n, inpDone_0n);
  OR2 I1 (outDone_0n, activateOut_0a, activateOut_1a);
  C2 I2 (int0_0n[0], inp_0r0d[1], inp_0r0d[0]);
  C2 I3 (int0_0n[1], inp_0r1d[2], inp_0r0d[1]);
  C2 I4 (int0_0n[2], inp_0r0d[2], inp_0r1d[0]);
  BUFF I5 (int0_0n[3], inp_0r1d[1]);
  OR2 I6 (activateOut_1r, int0_0n[0], int0_0n[1]);
  OR2 I7 (activateOut_0r, int0_0n[2], int0_0n[3]);
  C3 I8 (inpDone_0n, inpComplete_0n[0], inpComplete_0n[1], inpComplete_0n[2]);
  OR2 I9 (inpComplete_0n[0], inp_0r0d[0], inp_0r1d[0]);
  OR2 I10 (inpComplete_0n[1], inp_0r0d[1], inp_0r1d[1]);
  OR2 I11 (inpComplete_0n[2], inp_0r0d[2], inp_0r1d[2]);
endmodule

module BrzCase_3_2_s19_3_2c0m6_3b7_2c5_2c1 (
  inp_0r0d, inp_0r1d, inp_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a
);
  input [2:0] inp_0r0d;
  input [2:0] inp_0r1d;
  output inp_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  wire elseAck_0n;
  wire [2:0] inpComplete_0n;
  wire inpDone_0n;
  wire outDone_0n;
  wire [3:0] int0_0n;
  C2 I0 (inp_0a, outDone_0n, inpDone_0n);
  OR2 I1 (outDone_0n, activateOut_0a, activateOut_1a);
  C2 I2 (int0_0n[0], inp_0r0d[2], inp_0r1d[1]);
  C2 I3 (int0_0n[1], inp_0r0d[1], inp_0r1d[0]);
  C2 I4 (int0_0n[2], inp_0r1d[2], inp_0r1d[0]);
  BUFF I5 (int0_0n[3], inp_0r0d[0]);
  OR2 I6 (activateOut_1r, int0_0n[1], int0_0n[2]);
  OR2 I7 (activateOut_0r, int0_0n[0], int0_0n[3]);
  C3 I8 (inpDone_0n, inpComplete_0n[0], inpComplete_0n[1], inpComplete_0n[2]);
  OR2 I9 (inpComplete_0n[0], inp_0r0d[0], inp_0r1d[0]);
  OR2 I10 (inpComplete_0n[1], inp_0r0d[1], inp_0r1d[1]);
  OR2 I11 (inpComplete_0n[2], inp_0r0d[2], inp_0r1d[2]);
endmodule

module BrzCase_4_9_s67_15_2c0_3b2_2c1_3b4_2c3_3b6_m27m (
  inp_0r0d, inp_0r1d, inp_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a,
  activateOut_2r, activateOut_2a,
  activateOut_3r, activateOut_3a,
  activateOut_4r, activateOut_4a,
  activateOut_5r, activateOut_5a,
  activateOut_6r, activateOut_6a,
  activateOut_7r, activateOut_7a,
  activateOut_8r, activateOut_8a
);
  input [3:0] inp_0r0d;
  input [3:0] inp_0r1d;
  output inp_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  output activateOut_2r;
  input activateOut_2a;
  output activateOut_3r;
  input activateOut_3a;
  output activateOut_4r;
  input activateOut_4a;
  output activateOut_5r;
  input activateOut_5a;
  output activateOut_6r;
  input activateOut_6a;
  output activateOut_7r;
  input activateOut_7a;
  output activateOut_8r;
  input activateOut_8a;
  wire [36:0] internal_0n;
  wire elseAck_0n;
  wire [3:0] inpComplete_0n;
  wire inpDone_0n;
  wire outDone_0n;
  wire [15:0] int0_0n;
  C2 I0 (inp_0a, outDone_0n, inpDone_0n);
  NOR3 I1 (internal_0n[0], activateOut_0a, activateOut_1a, activateOut_2a);
  NOR3 I2 (internal_0n[1], activateOut_3a, activateOut_4a, activateOut_5a);
  NOR3 I3 (internal_0n[2], activateOut_6a, activateOut_7a, activateOut_8a);
  NAND3 I4 (outDone_0n, internal_0n[0], internal_0n[1], internal_0n[2]);
  C2 I5 (internal_0n[3], inp_0r1d[3], inp_0r0d[2]);
  C2 I6 (internal_0n[4], inp_0r0d[1], inp_0r0d[0]);
  C2 I7 (int0_0n[0], internal_0n[3], internal_0n[4]);
  C2 I8 (internal_0n[5], inp_0r0d[3], inp_0r1d[2]);
  C2 I9 (internal_0n[6], inp_0r1d[1], inp_0r1d[0]);
  C2 I10 (int0_0n[1], internal_0n[5], internal_0n[6]);
  C2 I11 (internal_0n[7], inp_0r1d[3], inp_0r1d[2]);
  C2 I12 (internal_0n[8], inp_0r1d[1], inp_0r0d[0]);
  C2 I13 (int0_0n[2], internal_0n[7], internal_0n[8]);
  C2 I14 (internal_0n[9], inp_0r1d[3], inp_0r1d[2]);
  C2 I15 (internal_0n[10], inp_0r0d[1], inp_0r1d[0]);
  C2 I16 (int0_0n[3], internal_0n[9], internal_0n[10]);
  C2 I17 (internal_0n[11], inp_0r1d[3], inp_0r1d[2]);
  C2 I18 (internal_0n[12], inp_0r0d[1], inp_0r0d[0]);
  C2 I19 (int0_0n[4], internal_0n[11], internal_0n[12]);
  C2 I20 (internal_0n[13], inp_0r1d[3], inp_0r0d[2]);
  C2 I21 (internal_0n[14], inp_0r1d[1], inp_0r1d[0]);
  C2 I22 (int0_0n[5], internal_0n[13], internal_0n[14]);
  C2 I23 (internal_0n[15], inp_0r1d[3], inp_0r0d[2]);
  C2 I24 (internal_0n[16], inp_0r1d[1], inp_0r0d[0]);
  C2 I25 (int0_0n[6], internal_0n[15], internal_0n[16]);
  C2 I26 (internal_0n[17], inp_0r1d[3], inp_0r0d[2]);
  C2 I27 (internal_0n[18], inp_0r0d[1], inp_0r1d[0]);
  C2 I28 (int0_0n[7], internal_0n[17], internal_0n[18]);
  C2 I29 (internal_0n[19], inp_0r0d[3], inp_0r1d[2]);
  C2 I30 (internal_0n[20], inp_0r1d[1], inp_0r0d[0]);
  C2 I31 (int0_0n[8], internal_0n[19], internal_0n[20]);
  C2 I32 (internal_0n[21], inp_0r0d[3], inp_0r1d[2]);
  C2 I33 (internal_0n[22], inp_0r0d[1], inp_0r1d[0]);
  C2 I34 (int0_0n[9], internal_0n[21], internal_0n[22]);
  C2 I35 (internal_0n[23], inp_0r0d[3], inp_0r1d[2]);
  C2 I36 (internal_0n[24], inp_0r0d[1], inp_0r0d[0]);
  C2 I37 (int0_0n[10], internal_0n[23], internal_0n[24]);
  C2 I38 (internal_0n[25], inp_0r0d[3], inp_0r0d[2]);
  C2 I39 (internal_0n[26], inp_0r1d[1], inp_0r1d[0]);
  C2 I40 (int0_0n[11], internal_0n[25], internal_0n[26]);
  C2 I41 (internal_0n[27], inp_0r0d[3], inp_0r0d[2]);
  C2 I42 (internal_0n[28], inp_0r1d[1], inp_0r0d[0]);
  C2 I43 (int0_0n[12], internal_0n[27], internal_0n[28]);
  C2 I44 (internal_0n[29], inp_0r0d[3], inp_0r0d[2]);
  C2 I45 (internal_0n[30], inp_0r0d[1], inp_0r1d[0]);
  C2 I46 (int0_0n[13], internal_0n[29], internal_0n[30]);
  C2 I47 (internal_0n[31], inp_0r0d[3], inp_0r0d[2]);
  C2 I48 (internal_0n[32], inp_0r0d[1], inp_0r0d[0]);
  C2 I49 (int0_0n[14], internal_0n[31], internal_0n[32]);
  C2 I50 (internal_0n[33], inp_0r1d[3], inp_0r1d[2]);
  C2 I51 (internal_0n[34], inp_0r1d[1], inp_0r1d[0]);
  C2 I52 (int0_0n[15], internal_0n[33], internal_0n[34]);
  OR2 I53 (activateOut_8r, int0_0n[2], int0_0n[3]);
  OR2 I54 (activateOut_7r, int0_0n[4], int0_0n[5]);
  OR2 I55 (activateOut_6r, int0_0n[6], int0_0n[7]);
  BUFF I56 (activateOut_5r, int0_0n[0]);
  BUFF I57 (activateOut_4r, int0_0n[1]);
  OR2 I58 (activateOut_3r, int0_0n[8], int0_0n[9]);
  OR2 I59 (activateOut_2r, int0_0n[10], int0_0n[11]);
  OR2 I60 (activateOut_1r, int0_0n[12], int0_0n[13]);
  OR2 I61 (activateOut_0r, int0_0n[14], int0_0n[15]);
  C2 I62 (internal_0n[35], inpComplete_0n[0], inpComplete_0n[1]);
  C2 I63 (internal_0n[36], inpComplete_0n[2], inpComplete_0n[3]);
  C2 I64 (inpDone_0n, internal_0n[35], internal_0n[36]);
  OR2 I65 (inpComplete_0n[0], inp_0r0d[0], inp_0r1d[0]);
  OR2 I66 (inpComplete_0n[1], inp_0r0d[1], inp_0r1d[1]);
  OR2 I67 (inpComplete_0n[2], inp_0r0d[2], inp_0r1d[2]);
  OR2 I68 (inpComplete_0n[3], inp_0r0d[3], inp_0r1d[3]);
endmodule

module BrzCombine_32_1_31 (
  out_0r, out_0a0d, out_0a1d,
  LSInp_0r, LSInp_0a0d, LSInp_0a1d,
  MSInp_0r, MSInp_0a0d, MSInp_0a1d
);
  input out_0r;
  output [31:0] out_0a0d;
  output [31:0] out_0a1d;
  output LSInp_0r;
  input LSInp_0a0d;
  input LSInp_0a1d;
  output MSInp_0r;
  input [30:0] MSInp_0a0d;
  input [30:0] MSInp_0a1d;
  BUFF I0 (LSInp_0r, out_0r);
  BUFF I1 (MSInp_0r, out_0r);
  BUFF I2 (out_0a0d[0], LSInp_0a0d);
  BUFF I3 (out_0a0d[1], MSInp_0a0d[0]);
  BUFF I4 (out_0a0d[2], MSInp_0a0d[1]);
  BUFF I5 (out_0a0d[3], MSInp_0a0d[2]);
  BUFF I6 (out_0a0d[4], MSInp_0a0d[3]);
  BUFF I7 (out_0a0d[5], MSInp_0a0d[4]);
  BUFF I8 (out_0a0d[6], MSInp_0a0d[5]);
  BUFF I9 (out_0a0d[7], MSInp_0a0d[6]);
  BUFF I10 (out_0a0d[8], MSInp_0a0d[7]);
  BUFF I11 (out_0a0d[9], MSInp_0a0d[8]);
  BUFF I12 (out_0a0d[10], MSInp_0a0d[9]);
  BUFF I13 (out_0a0d[11], MSInp_0a0d[10]);
  BUFF I14 (out_0a0d[12], MSInp_0a0d[11]);
  BUFF I15 (out_0a0d[13], MSInp_0a0d[12]);
  BUFF I16 (out_0a0d[14], MSInp_0a0d[13]);
  BUFF I17 (out_0a0d[15], MSInp_0a0d[14]);
  BUFF I18 (out_0a0d[16], MSInp_0a0d[15]);
  BUFF I19 (out_0a0d[17], MSInp_0a0d[16]);
  BUFF I20 (out_0a0d[18], MSInp_0a0d[17]);
  BUFF I21 (out_0a0d[19], MSInp_0a0d[18]);
  BUFF I22 (out_0a0d[20], MSInp_0a0d[19]);
  BUFF I23 (out_0a0d[21], MSInp_0a0d[20]);
  BUFF I24 (out_0a0d[22], MSInp_0a0d[21]);
  BUFF I25 (out_0a0d[23], MSInp_0a0d[22]);
  BUFF I26 (out_0a0d[24], MSInp_0a0d[23]);
  BUFF I27 (out_0a0d[25], MSInp_0a0d[24]);
  BUFF I28 (out_0a0d[26], MSInp_0a0d[25]);
  BUFF I29 (out_0a0d[27], MSInp_0a0d[26]);
  BUFF I30 (out_0a0d[28], MSInp_0a0d[27]);
  BUFF I31 (out_0a0d[29], MSInp_0a0d[28]);
  BUFF I32 (out_0a0d[30], MSInp_0a0d[29]);
  BUFF I33 (out_0a0d[31], MSInp_0a0d[30]);
  BUFF I34 (out_0a1d[0], LSInp_0a1d);
  BUFF I35 (out_0a1d[1], MSInp_0a1d[0]);
  BUFF I36 (out_0a1d[2], MSInp_0a1d[1]);
  BUFF I37 (out_0a1d[3], MSInp_0a1d[2]);
  BUFF I38 (out_0a1d[4], MSInp_0a1d[3]);
  BUFF I39 (out_0a1d[5], MSInp_0a1d[4]);
  BUFF I40 (out_0a1d[6], MSInp_0a1d[5]);
  BUFF I41 (out_0a1d[7], MSInp_0a1d[6]);
  BUFF I42 (out_0a1d[8], MSInp_0a1d[7]);
  BUFF I43 (out_0a1d[9], MSInp_0a1d[8]);
  BUFF I44 (out_0a1d[10], MSInp_0a1d[9]);
  BUFF I45 (out_0a1d[11], MSInp_0a1d[10]);
  BUFF I46 (out_0a1d[12], MSInp_0a1d[11]);
  BUFF I47 (out_0a1d[13], MSInp_0a1d[12]);
  BUFF I48 (out_0a1d[14], MSInp_0a1d[13]);
  BUFF I49 (out_0a1d[15], MSInp_0a1d[14]);
  BUFF I50 (out_0a1d[16], MSInp_0a1d[15]);
  BUFF I51 (out_0a1d[17], MSInp_0a1d[16]);
  BUFF I52 (out_0a1d[18], MSInp_0a1d[17]);
  BUFF I53 (out_0a1d[19], MSInp_0a1d[18]);
  BUFF I54 (out_0a1d[20], MSInp_0a1d[19]);
  BUFF I55 (out_0a1d[21], MSInp_0a1d[20]);
  BUFF I56 (out_0a1d[22], MSInp_0a1d[21]);
  BUFF I57 (out_0a1d[23], MSInp_0a1d[22]);
  BUFF I58 (out_0a1d[24], MSInp_0a1d[23]);
  BUFF I59 (out_0a1d[25], MSInp_0a1d[24]);
  BUFF I60 (out_0a1d[26], MSInp_0a1d[25]);
  BUFF I61 (out_0a1d[27], MSInp_0a1d[26]);
  BUFF I62 (out_0a1d[28], MSInp_0a1d[27]);
  BUFF I63 (out_0a1d[29], MSInp_0a1d[28]);
  BUFF I64 (out_0a1d[30], MSInp_0a1d[29]);
  BUFF I65 (out_0a1d[31], MSInp_0a1d[30]);
endmodule

module BrzCombine_33_1_32 (
  out_0r, out_0a0d, out_0a1d,
  LSInp_0r, LSInp_0a0d, LSInp_0a1d,
  MSInp_0r, MSInp_0a0d, MSInp_0a1d
);
  input out_0r;
  output [32:0] out_0a0d;
  output [32:0] out_0a1d;
  output LSInp_0r;
  input LSInp_0a0d;
  input LSInp_0a1d;
  output MSInp_0r;
  input [31:0] MSInp_0a0d;
  input [31:0] MSInp_0a1d;
  BUFF I0 (LSInp_0r, out_0r);
  BUFF I1 (MSInp_0r, out_0r);
  BUFF I2 (out_0a0d[0], LSInp_0a0d);
  BUFF I3 (out_0a0d[1], MSInp_0a0d[0]);
  BUFF I4 (out_0a0d[2], MSInp_0a0d[1]);
  BUFF I5 (out_0a0d[3], MSInp_0a0d[2]);
  BUFF I6 (out_0a0d[4], MSInp_0a0d[3]);
  BUFF I7 (out_0a0d[5], MSInp_0a0d[4]);
  BUFF I8 (out_0a0d[6], MSInp_0a0d[5]);
  BUFF I9 (out_0a0d[7], MSInp_0a0d[6]);
  BUFF I10 (out_0a0d[8], MSInp_0a0d[7]);
  BUFF I11 (out_0a0d[9], MSInp_0a0d[8]);
  BUFF I12 (out_0a0d[10], MSInp_0a0d[9]);
  BUFF I13 (out_0a0d[11], MSInp_0a0d[10]);
  BUFF I14 (out_0a0d[12], MSInp_0a0d[11]);
  BUFF I15 (out_0a0d[13], MSInp_0a0d[12]);
  BUFF I16 (out_0a0d[14], MSInp_0a0d[13]);
  BUFF I17 (out_0a0d[15], MSInp_0a0d[14]);
  BUFF I18 (out_0a0d[16], MSInp_0a0d[15]);
  BUFF I19 (out_0a0d[17], MSInp_0a0d[16]);
  BUFF I20 (out_0a0d[18], MSInp_0a0d[17]);
  BUFF I21 (out_0a0d[19], MSInp_0a0d[18]);
  BUFF I22 (out_0a0d[20], MSInp_0a0d[19]);
  BUFF I23 (out_0a0d[21], MSInp_0a0d[20]);
  BUFF I24 (out_0a0d[22], MSInp_0a0d[21]);
  BUFF I25 (out_0a0d[23], MSInp_0a0d[22]);
  BUFF I26 (out_0a0d[24], MSInp_0a0d[23]);
  BUFF I27 (out_0a0d[25], MSInp_0a0d[24]);
  BUFF I28 (out_0a0d[26], MSInp_0a0d[25]);
  BUFF I29 (out_0a0d[27], MSInp_0a0d[26]);
  BUFF I30 (out_0a0d[28], MSInp_0a0d[27]);
  BUFF I31 (out_0a0d[29], MSInp_0a0d[28]);
  BUFF I32 (out_0a0d[30], MSInp_0a0d[29]);
  BUFF I33 (out_0a0d[31], MSInp_0a0d[30]);
  BUFF I34 (out_0a0d[32], MSInp_0a0d[31]);
  BUFF I35 (out_0a1d[0], LSInp_0a1d);
  BUFF I36 (out_0a1d[1], MSInp_0a1d[0]);
  BUFF I37 (out_0a1d[2], MSInp_0a1d[1]);
  BUFF I38 (out_0a1d[3], MSInp_0a1d[2]);
  BUFF I39 (out_0a1d[4], MSInp_0a1d[3]);
  BUFF I40 (out_0a1d[5], MSInp_0a1d[4]);
  BUFF I41 (out_0a1d[6], MSInp_0a1d[5]);
  BUFF I42 (out_0a1d[7], MSInp_0a1d[6]);
  BUFF I43 (out_0a1d[8], MSInp_0a1d[7]);
  BUFF I44 (out_0a1d[9], MSInp_0a1d[8]);
  BUFF I45 (out_0a1d[10], MSInp_0a1d[9]);
  BUFF I46 (out_0a1d[11], MSInp_0a1d[10]);
  BUFF I47 (out_0a1d[12], MSInp_0a1d[11]);
  BUFF I48 (out_0a1d[13], MSInp_0a1d[12]);
  BUFF I49 (out_0a1d[14], MSInp_0a1d[13]);
  BUFF I50 (out_0a1d[15], MSInp_0a1d[14]);
  BUFF I51 (out_0a1d[16], MSInp_0a1d[15]);
  BUFF I52 (out_0a1d[17], MSInp_0a1d[16]);
  BUFF I53 (out_0a1d[18], MSInp_0a1d[17]);
  BUFF I54 (out_0a1d[19], MSInp_0a1d[18]);
  BUFF I55 (out_0a1d[20], MSInp_0a1d[19]);
  BUFF I56 (out_0a1d[21], MSInp_0a1d[20]);
  BUFF I57 (out_0a1d[22], MSInp_0a1d[21]);
  BUFF I58 (out_0a1d[23], MSInp_0a1d[22]);
  BUFF I59 (out_0a1d[24], MSInp_0a1d[23]);
  BUFF I60 (out_0a1d[25], MSInp_0a1d[24]);
  BUFF I61 (out_0a1d[26], MSInp_0a1d[25]);
  BUFF I62 (out_0a1d[27], MSInp_0a1d[26]);
  BUFF I63 (out_0a1d[28], MSInp_0a1d[27]);
  BUFF I64 (out_0a1d[29], MSInp_0a1d[28]);
  BUFF I65 (out_0a1d[30], MSInp_0a1d[29]);
  BUFF I66 (out_0a1d[31], MSInp_0a1d[30]);
  BUFF I67 (out_0a1d[32], MSInp_0a1d[31]);
endmodule

module BrzCombine_33_32_1 (
  out_0r, out_0a0d, out_0a1d,
  LSInp_0r, LSInp_0a0d, LSInp_0a1d,
  MSInp_0r, MSInp_0a0d, MSInp_0a1d
);
  input out_0r;
  output [32:0] out_0a0d;
  output [32:0] out_0a1d;
  output LSInp_0r;
  input [31:0] LSInp_0a0d;
  input [31:0] LSInp_0a1d;
  output MSInp_0r;
  input MSInp_0a0d;
  input MSInp_0a1d;
  BUFF I0 (LSInp_0r, out_0r);
  BUFF I1 (MSInp_0r, out_0r);
  BUFF I2 (out_0a0d[0], LSInp_0a0d[0]);
  BUFF I3 (out_0a0d[1], LSInp_0a0d[1]);
  BUFF I4 (out_0a0d[2], LSInp_0a0d[2]);
  BUFF I5 (out_0a0d[3], LSInp_0a0d[3]);
  BUFF I6 (out_0a0d[4], LSInp_0a0d[4]);
  BUFF I7 (out_0a0d[5], LSInp_0a0d[5]);
  BUFF I8 (out_0a0d[6], LSInp_0a0d[6]);
  BUFF I9 (out_0a0d[7], LSInp_0a0d[7]);
  BUFF I10 (out_0a0d[8], LSInp_0a0d[8]);
  BUFF I11 (out_0a0d[9], LSInp_0a0d[9]);
  BUFF I12 (out_0a0d[10], LSInp_0a0d[10]);
  BUFF I13 (out_0a0d[11], LSInp_0a0d[11]);
  BUFF I14 (out_0a0d[12], LSInp_0a0d[12]);
  BUFF I15 (out_0a0d[13], LSInp_0a0d[13]);
  BUFF I16 (out_0a0d[14], LSInp_0a0d[14]);
  BUFF I17 (out_0a0d[15], LSInp_0a0d[15]);
  BUFF I18 (out_0a0d[16], LSInp_0a0d[16]);
  BUFF I19 (out_0a0d[17], LSInp_0a0d[17]);
  BUFF I20 (out_0a0d[18], LSInp_0a0d[18]);
  BUFF I21 (out_0a0d[19], LSInp_0a0d[19]);
  BUFF I22 (out_0a0d[20], LSInp_0a0d[20]);
  BUFF I23 (out_0a0d[21], LSInp_0a0d[21]);
  BUFF I24 (out_0a0d[22], LSInp_0a0d[22]);
  BUFF I25 (out_0a0d[23], LSInp_0a0d[23]);
  BUFF I26 (out_0a0d[24], LSInp_0a0d[24]);
  BUFF I27 (out_0a0d[25], LSInp_0a0d[25]);
  BUFF I28 (out_0a0d[26], LSInp_0a0d[26]);
  BUFF I29 (out_0a0d[27], LSInp_0a0d[27]);
  BUFF I30 (out_0a0d[28], LSInp_0a0d[28]);
  BUFF I31 (out_0a0d[29], LSInp_0a0d[29]);
  BUFF I32 (out_0a0d[30], LSInp_0a0d[30]);
  BUFF I33 (out_0a0d[31], LSInp_0a0d[31]);
  BUFF I34 (out_0a0d[32], MSInp_0a0d);
  BUFF I35 (out_0a1d[0], LSInp_0a1d[0]);
  BUFF I36 (out_0a1d[1], LSInp_0a1d[1]);
  BUFF I37 (out_0a1d[2], LSInp_0a1d[2]);
  BUFF I38 (out_0a1d[3], LSInp_0a1d[3]);
  BUFF I39 (out_0a1d[4], LSInp_0a1d[4]);
  BUFF I40 (out_0a1d[5], LSInp_0a1d[5]);
  BUFF I41 (out_0a1d[6], LSInp_0a1d[6]);
  BUFF I42 (out_0a1d[7], LSInp_0a1d[7]);
  BUFF I43 (out_0a1d[8], LSInp_0a1d[8]);
  BUFF I44 (out_0a1d[9], LSInp_0a1d[9]);
  BUFF I45 (out_0a1d[10], LSInp_0a1d[10]);
  BUFF I46 (out_0a1d[11], LSInp_0a1d[11]);
  BUFF I47 (out_0a1d[12], LSInp_0a1d[12]);
  BUFF I48 (out_0a1d[13], LSInp_0a1d[13]);
  BUFF I49 (out_0a1d[14], LSInp_0a1d[14]);
  BUFF I50 (out_0a1d[15], LSInp_0a1d[15]);
  BUFF I51 (out_0a1d[16], LSInp_0a1d[16]);
  BUFF I52 (out_0a1d[17], LSInp_0a1d[17]);
  BUFF I53 (out_0a1d[18], LSInp_0a1d[18]);
  BUFF I54 (out_0a1d[19], LSInp_0a1d[19]);
  BUFF I55 (out_0a1d[20], LSInp_0a1d[20]);
  BUFF I56 (out_0a1d[21], LSInp_0a1d[21]);
  BUFF I57 (out_0a1d[22], LSInp_0a1d[22]);
  BUFF I58 (out_0a1d[23], LSInp_0a1d[23]);
  BUFF I59 (out_0a1d[24], LSInp_0a1d[24]);
  BUFF I60 (out_0a1d[25], LSInp_0a1d[25]);
  BUFF I61 (out_0a1d[26], LSInp_0a1d[26]);
  BUFF I62 (out_0a1d[27], LSInp_0a1d[27]);
  BUFF I63 (out_0a1d[28], LSInp_0a1d[28]);
  BUFF I64 (out_0a1d[29], LSInp_0a1d[29]);
  BUFF I65 (out_0a1d[30], LSInp_0a1d[30]);
  BUFF I66 (out_0a1d[31], LSInp_0a1d[31]);
  BUFF I67 (out_0a1d[32], MSInp_0a1d);
endmodule

module BrzCombine_35_1_34 (
  out_0r, out_0a0d, out_0a1d,
  LSInp_0r, LSInp_0a0d, LSInp_0a1d,
  MSInp_0r, MSInp_0a0d, MSInp_0a1d
);
  input out_0r;
  output [34:0] out_0a0d;
  output [34:0] out_0a1d;
  output LSInp_0r;
  input LSInp_0a0d;
  input LSInp_0a1d;
  output MSInp_0r;
  input [33:0] MSInp_0a0d;
  input [33:0] MSInp_0a1d;
  BUFF I0 (LSInp_0r, out_0r);
  BUFF I1 (MSInp_0r, out_0r);
  BUFF I2 (out_0a0d[0], LSInp_0a0d);
  BUFF I3 (out_0a0d[1], MSInp_0a0d[0]);
  BUFF I4 (out_0a0d[2], MSInp_0a0d[1]);
  BUFF I5 (out_0a0d[3], MSInp_0a0d[2]);
  BUFF I6 (out_0a0d[4], MSInp_0a0d[3]);
  BUFF I7 (out_0a0d[5], MSInp_0a0d[4]);
  BUFF I8 (out_0a0d[6], MSInp_0a0d[5]);
  BUFF I9 (out_0a0d[7], MSInp_0a0d[6]);
  BUFF I10 (out_0a0d[8], MSInp_0a0d[7]);
  BUFF I11 (out_0a0d[9], MSInp_0a0d[8]);
  BUFF I12 (out_0a0d[10], MSInp_0a0d[9]);
  BUFF I13 (out_0a0d[11], MSInp_0a0d[10]);
  BUFF I14 (out_0a0d[12], MSInp_0a0d[11]);
  BUFF I15 (out_0a0d[13], MSInp_0a0d[12]);
  BUFF I16 (out_0a0d[14], MSInp_0a0d[13]);
  BUFF I17 (out_0a0d[15], MSInp_0a0d[14]);
  BUFF I18 (out_0a0d[16], MSInp_0a0d[15]);
  BUFF I19 (out_0a0d[17], MSInp_0a0d[16]);
  BUFF I20 (out_0a0d[18], MSInp_0a0d[17]);
  BUFF I21 (out_0a0d[19], MSInp_0a0d[18]);
  BUFF I22 (out_0a0d[20], MSInp_0a0d[19]);
  BUFF I23 (out_0a0d[21], MSInp_0a0d[20]);
  BUFF I24 (out_0a0d[22], MSInp_0a0d[21]);
  BUFF I25 (out_0a0d[23], MSInp_0a0d[22]);
  BUFF I26 (out_0a0d[24], MSInp_0a0d[23]);
  BUFF I27 (out_0a0d[25], MSInp_0a0d[24]);
  BUFF I28 (out_0a0d[26], MSInp_0a0d[25]);
  BUFF I29 (out_0a0d[27], MSInp_0a0d[26]);
  BUFF I30 (out_0a0d[28], MSInp_0a0d[27]);
  BUFF I31 (out_0a0d[29], MSInp_0a0d[28]);
  BUFF I32 (out_0a0d[30], MSInp_0a0d[29]);
  BUFF I33 (out_0a0d[31], MSInp_0a0d[30]);
  BUFF I34 (out_0a0d[32], MSInp_0a0d[31]);
  BUFF I35 (out_0a0d[33], MSInp_0a0d[32]);
  BUFF I36 (out_0a0d[34], MSInp_0a0d[33]);
  BUFF I37 (out_0a1d[0], LSInp_0a1d);
  BUFF I38 (out_0a1d[1], MSInp_0a1d[0]);
  BUFF I39 (out_0a1d[2], MSInp_0a1d[1]);
  BUFF I40 (out_0a1d[3], MSInp_0a1d[2]);
  BUFF I41 (out_0a1d[4], MSInp_0a1d[3]);
  BUFF I42 (out_0a1d[5], MSInp_0a1d[4]);
  BUFF I43 (out_0a1d[6], MSInp_0a1d[5]);
  BUFF I44 (out_0a1d[7], MSInp_0a1d[6]);
  BUFF I45 (out_0a1d[8], MSInp_0a1d[7]);
  BUFF I46 (out_0a1d[9], MSInp_0a1d[8]);
  BUFF I47 (out_0a1d[10], MSInp_0a1d[9]);
  BUFF I48 (out_0a1d[11], MSInp_0a1d[10]);
  BUFF I49 (out_0a1d[12], MSInp_0a1d[11]);
  BUFF I50 (out_0a1d[13], MSInp_0a1d[12]);
  BUFF I51 (out_0a1d[14], MSInp_0a1d[13]);
  BUFF I52 (out_0a1d[15], MSInp_0a1d[14]);
  BUFF I53 (out_0a1d[16], MSInp_0a1d[15]);
  BUFF I54 (out_0a1d[17], MSInp_0a1d[16]);
  BUFF I55 (out_0a1d[18], MSInp_0a1d[17]);
  BUFF I56 (out_0a1d[19], MSInp_0a1d[18]);
  BUFF I57 (out_0a1d[20], MSInp_0a1d[19]);
  BUFF I58 (out_0a1d[21], MSInp_0a1d[20]);
  BUFF I59 (out_0a1d[22], MSInp_0a1d[21]);
  BUFF I60 (out_0a1d[23], MSInp_0a1d[22]);
  BUFF I61 (out_0a1d[24], MSInp_0a1d[23]);
  BUFF I62 (out_0a1d[25], MSInp_0a1d[24]);
  BUFF I63 (out_0a1d[26], MSInp_0a1d[25]);
  BUFF I64 (out_0a1d[27], MSInp_0a1d[26]);
  BUFF I65 (out_0a1d[28], MSInp_0a1d[27]);
  BUFF I66 (out_0a1d[29], MSInp_0a1d[28]);
  BUFF I67 (out_0a1d[30], MSInp_0a1d[29]);
  BUFF I68 (out_0a1d[31], MSInp_0a1d[30]);
  BUFF I69 (out_0a1d[32], MSInp_0a1d[31]);
  BUFF I70 (out_0a1d[33], MSInp_0a1d[32]);
  BUFF I71 (out_0a1d[34], MSInp_0a1d[33]);
endmodule

module BrzCombine_35_2_33 (
  out_0r, out_0a0d, out_0a1d,
  LSInp_0r, LSInp_0a0d, LSInp_0a1d,
  MSInp_0r, MSInp_0a0d, MSInp_0a1d
);
  input out_0r;
  output [34:0] out_0a0d;
  output [34:0] out_0a1d;
  output LSInp_0r;
  input [1:0] LSInp_0a0d;
  input [1:0] LSInp_0a1d;
  output MSInp_0r;
  input [32:0] MSInp_0a0d;
  input [32:0] MSInp_0a1d;
  BUFF I0 (LSInp_0r, out_0r);
  BUFF I1 (MSInp_0r, out_0r);
  BUFF I2 (out_0a0d[0], LSInp_0a0d[0]);
  BUFF I3 (out_0a0d[1], LSInp_0a0d[1]);
  BUFF I4 (out_0a0d[2], MSInp_0a0d[0]);
  BUFF I5 (out_0a0d[3], MSInp_0a0d[1]);
  BUFF I6 (out_0a0d[4], MSInp_0a0d[2]);
  BUFF I7 (out_0a0d[5], MSInp_0a0d[3]);
  BUFF I8 (out_0a0d[6], MSInp_0a0d[4]);
  BUFF I9 (out_0a0d[7], MSInp_0a0d[5]);
  BUFF I10 (out_0a0d[8], MSInp_0a0d[6]);
  BUFF I11 (out_0a0d[9], MSInp_0a0d[7]);
  BUFF I12 (out_0a0d[10], MSInp_0a0d[8]);
  BUFF I13 (out_0a0d[11], MSInp_0a0d[9]);
  BUFF I14 (out_0a0d[12], MSInp_0a0d[10]);
  BUFF I15 (out_0a0d[13], MSInp_0a0d[11]);
  BUFF I16 (out_0a0d[14], MSInp_0a0d[12]);
  BUFF I17 (out_0a0d[15], MSInp_0a0d[13]);
  BUFF I18 (out_0a0d[16], MSInp_0a0d[14]);
  BUFF I19 (out_0a0d[17], MSInp_0a0d[15]);
  BUFF I20 (out_0a0d[18], MSInp_0a0d[16]);
  BUFF I21 (out_0a0d[19], MSInp_0a0d[17]);
  BUFF I22 (out_0a0d[20], MSInp_0a0d[18]);
  BUFF I23 (out_0a0d[21], MSInp_0a0d[19]);
  BUFF I24 (out_0a0d[22], MSInp_0a0d[20]);
  BUFF I25 (out_0a0d[23], MSInp_0a0d[21]);
  BUFF I26 (out_0a0d[24], MSInp_0a0d[22]);
  BUFF I27 (out_0a0d[25], MSInp_0a0d[23]);
  BUFF I28 (out_0a0d[26], MSInp_0a0d[24]);
  BUFF I29 (out_0a0d[27], MSInp_0a0d[25]);
  BUFF I30 (out_0a0d[28], MSInp_0a0d[26]);
  BUFF I31 (out_0a0d[29], MSInp_0a0d[27]);
  BUFF I32 (out_0a0d[30], MSInp_0a0d[28]);
  BUFF I33 (out_0a0d[31], MSInp_0a0d[29]);
  BUFF I34 (out_0a0d[32], MSInp_0a0d[30]);
  BUFF I35 (out_0a0d[33], MSInp_0a0d[31]);
  BUFF I36 (out_0a0d[34], MSInp_0a0d[32]);
  BUFF I37 (out_0a1d[0], LSInp_0a1d[0]);
  BUFF I38 (out_0a1d[1], LSInp_0a1d[1]);
  BUFF I39 (out_0a1d[2], MSInp_0a1d[0]);
  BUFF I40 (out_0a1d[3], MSInp_0a1d[1]);
  BUFF I41 (out_0a1d[4], MSInp_0a1d[2]);
  BUFF I42 (out_0a1d[5], MSInp_0a1d[3]);
  BUFF I43 (out_0a1d[6], MSInp_0a1d[4]);
  BUFF I44 (out_0a1d[7], MSInp_0a1d[5]);
  BUFF I45 (out_0a1d[8], MSInp_0a1d[6]);
  BUFF I46 (out_0a1d[9], MSInp_0a1d[7]);
  BUFF I47 (out_0a1d[10], MSInp_0a1d[8]);
  BUFF I48 (out_0a1d[11], MSInp_0a1d[9]);
  BUFF I49 (out_0a1d[12], MSInp_0a1d[10]);
  BUFF I50 (out_0a1d[13], MSInp_0a1d[11]);
  BUFF I51 (out_0a1d[14], MSInp_0a1d[12]);
  BUFF I52 (out_0a1d[15], MSInp_0a1d[13]);
  BUFF I53 (out_0a1d[16], MSInp_0a1d[14]);
  BUFF I54 (out_0a1d[17], MSInp_0a1d[15]);
  BUFF I55 (out_0a1d[18], MSInp_0a1d[16]);
  BUFF I56 (out_0a1d[19], MSInp_0a1d[17]);
  BUFF I57 (out_0a1d[20], MSInp_0a1d[18]);
  BUFF I58 (out_0a1d[21], MSInp_0a1d[19]);
  BUFF I59 (out_0a1d[22], MSInp_0a1d[20]);
  BUFF I60 (out_0a1d[23], MSInp_0a1d[21]);
  BUFF I61 (out_0a1d[24], MSInp_0a1d[22]);
  BUFF I62 (out_0a1d[25], MSInp_0a1d[23]);
  BUFF I63 (out_0a1d[26], MSInp_0a1d[24]);
  BUFF I64 (out_0a1d[27], MSInp_0a1d[25]);
  BUFF I65 (out_0a1d[28], MSInp_0a1d[26]);
  BUFF I66 (out_0a1d[29], MSInp_0a1d[27]);
  BUFF I67 (out_0a1d[30], MSInp_0a1d[28]);
  BUFF I68 (out_0a1d[31], MSInp_0a1d[29]);
  BUFF I69 (out_0a1d[32], MSInp_0a1d[30]);
  BUFF I70 (out_0a1d[33], MSInp_0a1d[31]);
  BUFF I71 (out_0a1d[34], MSInp_0a1d[32]);
endmodule

module BrzCombine_35_32_3 (
  out_0r, out_0a0d, out_0a1d,
  LSInp_0r, LSInp_0a0d, LSInp_0a1d,
  MSInp_0r, MSInp_0a0d, MSInp_0a1d
);
  input out_0r;
  output [34:0] out_0a0d;
  output [34:0] out_0a1d;
  output LSInp_0r;
  input [31:0] LSInp_0a0d;
  input [31:0] LSInp_0a1d;
  output MSInp_0r;
  input [2:0] MSInp_0a0d;
  input [2:0] MSInp_0a1d;
  BUFF I0 (LSInp_0r, out_0r);
  BUFF I1 (MSInp_0r, out_0r);
  BUFF I2 (out_0a0d[0], LSInp_0a0d[0]);
  BUFF I3 (out_0a0d[1], LSInp_0a0d[1]);
  BUFF I4 (out_0a0d[2], LSInp_0a0d[2]);
  BUFF I5 (out_0a0d[3], LSInp_0a0d[3]);
  BUFF I6 (out_0a0d[4], LSInp_0a0d[4]);
  BUFF I7 (out_0a0d[5], LSInp_0a0d[5]);
  BUFF I8 (out_0a0d[6], LSInp_0a0d[6]);
  BUFF I9 (out_0a0d[7], LSInp_0a0d[7]);
  BUFF I10 (out_0a0d[8], LSInp_0a0d[8]);
  BUFF I11 (out_0a0d[9], LSInp_0a0d[9]);
  BUFF I12 (out_0a0d[10], LSInp_0a0d[10]);
  BUFF I13 (out_0a0d[11], LSInp_0a0d[11]);
  BUFF I14 (out_0a0d[12], LSInp_0a0d[12]);
  BUFF I15 (out_0a0d[13], LSInp_0a0d[13]);
  BUFF I16 (out_0a0d[14], LSInp_0a0d[14]);
  BUFF I17 (out_0a0d[15], LSInp_0a0d[15]);
  BUFF I18 (out_0a0d[16], LSInp_0a0d[16]);
  BUFF I19 (out_0a0d[17], LSInp_0a0d[17]);
  BUFF I20 (out_0a0d[18], LSInp_0a0d[18]);
  BUFF I21 (out_0a0d[19], LSInp_0a0d[19]);
  BUFF I22 (out_0a0d[20], LSInp_0a0d[20]);
  BUFF I23 (out_0a0d[21], LSInp_0a0d[21]);
  BUFF I24 (out_0a0d[22], LSInp_0a0d[22]);
  BUFF I25 (out_0a0d[23], LSInp_0a0d[23]);
  BUFF I26 (out_0a0d[24], LSInp_0a0d[24]);
  BUFF I27 (out_0a0d[25], LSInp_0a0d[25]);
  BUFF I28 (out_0a0d[26], LSInp_0a0d[26]);
  BUFF I29 (out_0a0d[27], LSInp_0a0d[27]);
  BUFF I30 (out_0a0d[28], LSInp_0a0d[28]);
  BUFF I31 (out_0a0d[29], LSInp_0a0d[29]);
  BUFF I32 (out_0a0d[30], LSInp_0a0d[30]);
  BUFF I33 (out_0a0d[31], LSInp_0a0d[31]);
  BUFF I34 (out_0a0d[32], MSInp_0a0d[0]);
  BUFF I35 (out_0a0d[33], MSInp_0a0d[1]);
  BUFF I36 (out_0a0d[34], MSInp_0a0d[2]);
  BUFF I37 (out_0a1d[0], LSInp_0a1d[0]);
  BUFF I38 (out_0a1d[1], LSInp_0a1d[1]);
  BUFF I39 (out_0a1d[2], LSInp_0a1d[2]);
  BUFF I40 (out_0a1d[3], LSInp_0a1d[3]);
  BUFF I41 (out_0a1d[4], LSInp_0a1d[4]);
  BUFF I42 (out_0a1d[5], LSInp_0a1d[5]);
  BUFF I43 (out_0a1d[6], LSInp_0a1d[6]);
  BUFF I44 (out_0a1d[7], LSInp_0a1d[7]);
  BUFF I45 (out_0a1d[8], LSInp_0a1d[8]);
  BUFF I46 (out_0a1d[9], LSInp_0a1d[9]);
  BUFF I47 (out_0a1d[10], LSInp_0a1d[10]);
  BUFF I48 (out_0a1d[11], LSInp_0a1d[11]);
  BUFF I49 (out_0a1d[12], LSInp_0a1d[12]);
  BUFF I50 (out_0a1d[13], LSInp_0a1d[13]);
  BUFF I51 (out_0a1d[14], LSInp_0a1d[14]);
  BUFF I52 (out_0a1d[15], LSInp_0a1d[15]);
  BUFF I53 (out_0a1d[16], LSInp_0a1d[16]);
  BUFF I54 (out_0a1d[17], LSInp_0a1d[17]);
  BUFF I55 (out_0a1d[18], LSInp_0a1d[18]);
  BUFF I56 (out_0a1d[19], LSInp_0a1d[19]);
  BUFF I57 (out_0a1d[20], LSInp_0a1d[20]);
  BUFF I58 (out_0a1d[21], LSInp_0a1d[21]);
  BUFF I59 (out_0a1d[22], LSInp_0a1d[22]);
  BUFF I60 (out_0a1d[23], LSInp_0a1d[23]);
  BUFF I61 (out_0a1d[24], LSInp_0a1d[24]);
  BUFF I62 (out_0a1d[25], LSInp_0a1d[25]);
  BUFF I63 (out_0a1d[26], LSInp_0a1d[26]);
  BUFF I64 (out_0a1d[27], LSInp_0a1d[27]);
  BUFF I65 (out_0a1d[28], LSInp_0a1d[28]);
  BUFF I66 (out_0a1d[29], LSInp_0a1d[29]);
  BUFF I67 (out_0a1d[30], LSInp_0a1d[30]);
  BUFF I68 (out_0a1d[31], LSInp_0a1d[31]);
  BUFF I69 (out_0a1d[32], MSInp_0a1d[0]);
  BUFF I70 (out_0a1d[33], MSInp_0a1d[1]);
  BUFF I71 (out_0a1d[34], MSInp_0a1d[2]);
endmodule

module BrzCombine_35_33_2 (
  out_0r, out_0a0d, out_0a1d,
  LSInp_0r, LSInp_0a0d, LSInp_0a1d,
  MSInp_0r, MSInp_0a0d, MSInp_0a1d
);
  input out_0r;
  output [34:0] out_0a0d;
  output [34:0] out_0a1d;
  output LSInp_0r;
  input [32:0] LSInp_0a0d;
  input [32:0] LSInp_0a1d;
  output MSInp_0r;
  input [1:0] MSInp_0a0d;
  input [1:0] MSInp_0a1d;
  BUFF I0 (LSInp_0r, out_0r);
  BUFF I1 (MSInp_0r, out_0r);
  BUFF I2 (out_0a0d[0], LSInp_0a0d[0]);
  BUFF I3 (out_0a0d[1], LSInp_0a0d[1]);
  BUFF I4 (out_0a0d[2], LSInp_0a0d[2]);
  BUFF I5 (out_0a0d[3], LSInp_0a0d[3]);
  BUFF I6 (out_0a0d[4], LSInp_0a0d[4]);
  BUFF I7 (out_0a0d[5], LSInp_0a0d[5]);
  BUFF I8 (out_0a0d[6], LSInp_0a0d[6]);
  BUFF I9 (out_0a0d[7], LSInp_0a0d[7]);
  BUFF I10 (out_0a0d[8], LSInp_0a0d[8]);
  BUFF I11 (out_0a0d[9], LSInp_0a0d[9]);
  BUFF I12 (out_0a0d[10], LSInp_0a0d[10]);
  BUFF I13 (out_0a0d[11], LSInp_0a0d[11]);
  BUFF I14 (out_0a0d[12], LSInp_0a0d[12]);
  BUFF I15 (out_0a0d[13], LSInp_0a0d[13]);
  BUFF I16 (out_0a0d[14], LSInp_0a0d[14]);
  BUFF I17 (out_0a0d[15], LSInp_0a0d[15]);
  BUFF I18 (out_0a0d[16], LSInp_0a0d[16]);
  BUFF I19 (out_0a0d[17], LSInp_0a0d[17]);
  BUFF I20 (out_0a0d[18], LSInp_0a0d[18]);
  BUFF I21 (out_0a0d[19], LSInp_0a0d[19]);
  BUFF I22 (out_0a0d[20], LSInp_0a0d[20]);
  BUFF I23 (out_0a0d[21], LSInp_0a0d[21]);
  BUFF I24 (out_0a0d[22], LSInp_0a0d[22]);
  BUFF I25 (out_0a0d[23], LSInp_0a0d[23]);
  BUFF I26 (out_0a0d[24], LSInp_0a0d[24]);
  BUFF I27 (out_0a0d[25], LSInp_0a0d[25]);
  BUFF I28 (out_0a0d[26], LSInp_0a0d[26]);
  BUFF I29 (out_0a0d[27], LSInp_0a0d[27]);
  BUFF I30 (out_0a0d[28], LSInp_0a0d[28]);
  BUFF I31 (out_0a0d[29], LSInp_0a0d[29]);
  BUFF I32 (out_0a0d[30], LSInp_0a0d[30]);
  BUFF I33 (out_0a0d[31], LSInp_0a0d[31]);
  BUFF I34 (out_0a0d[32], LSInp_0a0d[32]);
  BUFF I35 (out_0a0d[33], MSInp_0a0d[0]);
  BUFF I36 (out_0a0d[34], MSInp_0a0d[1]);
  BUFF I37 (out_0a1d[0], LSInp_0a1d[0]);
  BUFF I38 (out_0a1d[1], LSInp_0a1d[1]);
  BUFF I39 (out_0a1d[2], LSInp_0a1d[2]);
  BUFF I40 (out_0a1d[3], LSInp_0a1d[3]);
  BUFF I41 (out_0a1d[4], LSInp_0a1d[4]);
  BUFF I42 (out_0a1d[5], LSInp_0a1d[5]);
  BUFF I43 (out_0a1d[6], LSInp_0a1d[6]);
  BUFF I44 (out_0a1d[7], LSInp_0a1d[7]);
  BUFF I45 (out_0a1d[8], LSInp_0a1d[8]);
  BUFF I46 (out_0a1d[9], LSInp_0a1d[9]);
  BUFF I47 (out_0a1d[10], LSInp_0a1d[10]);
  BUFF I48 (out_0a1d[11], LSInp_0a1d[11]);
  BUFF I49 (out_0a1d[12], LSInp_0a1d[12]);
  BUFF I50 (out_0a1d[13], LSInp_0a1d[13]);
  BUFF I51 (out_0a1d[14], LSInp_0a1d[14]);
  BUFF I52 (out_0a1d[15], LSInp_0a1d[15]);
  BUFF I53 (out_0a1d[16], LSInp_0a1d[16]);
  BUFF I54 (out_0a1d[17], LSInp_0a1d[17]);
  BUFF I55 (out_0a1d[18], LSInp_0a1d[18]);
  BUFF I56 (out_0a1d[19], LSInp_0a1d[19]);
  BUFF I57 (out_0a1d[20], LSInp_0a1d[20]);
  BUFF I58 (out_0a1d[21], LSInp_0a1d[21]);
  BUFF I59 (out_0a1d[22], LSInp_0a1d[22]);
  BUFF I60 (out_0a1d[23], LSInp_0a1d[23]);
  BUFF I61 (out_0a1d[24], LSInp_0a1d[24]);
  BUFF I62 (out_0a1d[25], LSInp_0a1d[25]);
  BUFF I63 (out_0a1d[26], LSInp_0a1d[26]);
  BUFF I64 (out_0a1d[27], LSInp_0a1d[27]);
  BUFF I65 (out_0a1d[28], LSInp_0a1d[28]);
  BUFF I66 (out_0a1d[29], LSInp_0a1d[29]);
  BUFF I67 (out_0a1d[30], LSInp_0a1d[30]);
  BUFF I68 (out_0a1d[31], LSInp_0a1d[31]);
  BUFF I69 (out_0a1d[32], LSInp_0a1d[32]);
  BUFF I70 (out_0a1d[33], MSInp_0a1d[0]);
  BUFF I71 (out_0a1d[34], MSInp_0a1d[1]);
endmodule

module BrzCombineEqual_2_1_2 (
  out_0r, out_0a0d, out_0a1d,
  inp_0r, inp_0a0d, inp_0a1d,
  inp_1r, inp_1a0d, inp_1a1d
);
  input out_0r;
  output [1:0] out_0a0d;
  output [1:0] out_0a1d;
  output inp_0r;
  input inp_0a0d;
  input inp_0a1d;
  output inp_1r;
  input inp_1a0d;
  input inp_1a1d;
  wire outReq_0n;
  BUFF I0 (inp_0r, outReq_0n);
  BUFF I1 (inp_1r, outReq_0n);
  BUFF I2 (outReq_0n, out_0r);
  BUFF I3 (out_0a0d[0], inp_0a0d);
  BUFF I4 (out_0a0d[1], inp_1a0d);
  BUFF I5 (out_0a1d[0], inp_0a1d);
  BUFF I6 (out_0a1d[1], inp_1a1d);
endmodule

module BrzConcur_2 (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  wire [1:0] acks_0n;
  wire actReq_0n;
  C2 I0 (activate_0a, acks_0n[0], acks_0n[1]);
  BALSA_TELEM I1 (actReq_0n, acks_0n[0], activateOut_0r, activateOut_0a);
  BALSA_TELEM I2 (actReq_0n, acks_0n[1], activateOut_1r, activateOut_1a);
  BUFF I3 (actReq_0n, activate_0r);
endmodule

module BrzConcur_3 (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a,
  activateOut_2r, activateOut_2a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  output activateOut_2r;
  input activateOut_2a;
  wire [2:0] acks_0n;
  wire actReq_0n;
  C3 I0 (activate_0a, acks_0n[0], acks_0n[1], acks_0n[2]);
  BALSA_TELEM I1 (actReq_0n, acks_0n[0], activateOut_0r, activateOut_0a);
  BALSA_TELEM I2 (actReq_0n, acks_0n[1], activateOut_1r, activateOut_1a);
  BALSA_TELEM I3 (actReq_0n, acks_0n[2], activateOut_2r, activateOut_2a);
  BUFF I4 (actReq_0n, activate_0r);
endmodule

module BrzConcur_4 (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a,
  activateOut_2r, activateOut_2a,
  activateOut_3r, activateOut_3a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  output activateOut_2r;
  input activateOut_2a;
  output activateOut_3r;
  input activateOut_3a;
  wire [1:0] internal_0n;
  wire [3:0] acks_0n;
  wire actReq_0n;
  C2 I0 (internal_0n[0], acks_0n[0], acks_0n[1]);
  C2 I1 (internal_0n[1], acks_0n[2], acks_0n[3]);
  C2 I2 (activate_0a, internal_0n[0], internal_0n[1]);
  BALSA_TELEM I3 (actReq_0n, acks_0n[0], activateOut_0r, activateOut_0a);
  BALSA_TELEM I4 (actReq_0n, acks_0n[1], activateOut_1r, activateOut_1a);
  BALSA_TELEM I5 (actReq_0n, acks_0n[2], activateOut_2r, activateOut_2a);
  BALSA_TELEM I6 (actReq_0n, acks_0n[3], activateOut_3r, activateOut_3a);
  BUFF I7 (actReq_0n, activate_0r);
endmodule

module BrzConcur_5 (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a,
  activateOut_2r, activateOut_2a,
  activateOut_3r, activateOut_3a,
  activateOut_4r, activateOut_4a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  output activateOut_2r;
  input activateOut_2a;
  output activateOut_3r;
  input activateOut_3a;
  output activateOut_4r;
  input activateOut_4a;
  wire [1:0] internal_0n;
  wire [4:0] acks_0n;
  wire actReq_0n;
  C3 I0 (internal_0n[0], acks_0n[0], acks_0n[1], acks_0n[2]);
  C2 I1 (internal_0n[1], acks_0n[3], acks_0n[4]);
  C2 I2 (activate_0a, internal_0n[0], internal_0n[1]);
  BALSA_TELEM I3 (actReq_0n, acks_0n[0], activateOut_0r, activateOut_0a);
  BALSA_TELEM I4 (actReq_0n, acks_0n[1], activateOut_1r, activateOut_1a);
  BALSA_TELEM I5 (actReq_0n, acks_0n[2], activateOut_2r, activateOut_2a);
  BALSA_TELEM I6 (actReq_0n, acks_0n[3], activateOut_3r, activateOut_3a);
  BALSA_TELEM I7 (actReq_0n, acks_0n[4], activateOut_4r, activateOut_4a);
  BUFF I8 (actReq_0n, activate_0r);
endmodule

module BrzConcur_6 (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a,
  activateOut_2r, activateOut_2a,
  activateOut_3r, activateOut_3a,
  activateOut_4r, activateOut_4a,
  activateOut_5r, activateOut_5a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  output activateOut_2r;
  input activateOut_2a;
  output activateOut_3r;
  input activateOut_3a;
  output activateOut_4r;
  input activateOut_4a;
  output activateOut_5r;
  input activateOut_5a;
  wire [1:0] internal_0n;
  wire [5:0] acks_0n;
  wire actReq_0n;
  C3 I0 (internal_0n[0], acks_0n[0], acks_0n[1], acks_0n[2]);
  C3 I1 (internal_0n[1], acks_0n[3], acks_0n[4], acks_0n[5]);
  C2 I2 (activate_0a, internal_0n[0], internal_0n[1]);
  BALSA_TELEM I3 (actReq_0n, acks_0n[0], activateOut_0r, activateOut_0a);
  BALSA_TELEM I4 (actReq_0n, acks_0n[1], activateOut_1r, activateOut_1a);
  BALSA_TELEM I5 (actReq_0n, acks_0n[2], activateOut_2r, activateOut_2a);
  BALSA_TELEM I6 (actReq_0n, acks_0n[3], activateOut_3r, activateOut_3a);
  BALSA_TELEM I7 (actReq_0n, acks_0n[4], activateOut_4r, activateOut_4a);
  BALSA_TELEM I8 (actReq_0n, acks_0n[5], activateOut_5r, activateOut_5a);
  BUFF I9 (actReq_0n, activate_0r);
endmodule

module BrzConcur_8 (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a,
  activateOut_2r, activateOut_2a,
  activateOut_3r, activateOut_3a,
  activateOut_4r, activateOut_4a,
  activateOut_5r, activateOut_5a,
  activateOut_6r, activateOut_6a,
  activateOut_7r, activateOut_7a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  output activateOut_2r;
  input activateOut_2a;
  output activateOut_3r;
  input activateOut_3a;
  output activateOut_4r;
  input activateOut_4a;
  output activateOut_5r;
  input activateOut_5a;
  output activateOut_6r;
  input activateOut_6a;
  output activateOut_7r;
  input activateOut_7a;
  wire [2:0] internal_0n;
  wire [7:0] acks_0n;
  wire actReq_0n;
  C3 I0 (internal_0n[0], acks_0n[0], acks_0n[1], acks_0n[2]);
  C3 I1 (internal_0n[1], acks_0n[3], acks_0n[4], acks_0n[5]);
  C2 I2 (internal_0n[2], acks_0n[6], acks_0n[7]);
  C3 I3 (activate_0a, internal_0n[0], internal_0n[1], internal_0n[2]);
  BALSA_TELEM I4 (actReq_0n, acks_0n[0], activateOut_0r, activateOut_0a);
  BALSA_TELEM I5 (actReq_0n, acks_0n[1], activateOut_1r, activateOut_1a);
  BALSA_TELEM I6 (actReq_0n, acks_0n[2], activateOut_2r, activateOut_2a);
  BALSA_TELEM I7 (actReq_0n, acks_0n[3], activateOut_3r, activateOut_3a);
  BALSA_TELEM I8 (actReq_0n, acks_0n[4], activateOut_4r, activateOut_4a);
  BALSA_TELEM I9 (actReq_0n, acks_0n[5], activateOut_5r, activateOut_5a);
  BALSA_TELEM I10 (actReq_0n, acks_0n[6], activateOut_6r, activateOut_6a);
  BALSA_TELEM I11 (actReq_0n, acks_0n[7], activateOut_7r, activateOut_7a);
  BUFF I12 (actReq_0n, activate_0r);
endmodule

module BrzConcur_14 (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a,
  activateOut_2r, activateOut_2a,
  activateOut_3r, activateOut_3a,
  activateOut_4r, activateOut_4a,
  activateOut_5r, activateOut_5a,
  activateOut_6r, activateOut_6a,
  activateOut_7r, activateOut_7a,
  activateOut_8r, activateOut_8a,
  activateOut_9r, activateOut_9a,
  activateOut_10r, activateOut_10a,
  activateOut_11r, activateOut_11a,
  activateOut_12r, activateOut_12a,
  activateOut_13r, activateOut_13a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  output activateOut_2r;
  input activateOut_2a;
  output activateOut_3r;
  input activateOut_3a;
  output activateOut_4r;
  input activateOut_4a;
  output activateOut_5r;
  input activateOut_5a;
  output activateOut_6r;
  input activateOut_6a;
  output activateOut_7r;
  input activateOut_7a;
  output activateOut_8r;
  input activateOut_8a;
  output activateOut_9r;
  input activateOut_9a;
  output activateOut_10r;
  input activateOut_10a;
  output activateOut_11r;
  input activateOut_11a;
  output activateOut_12r;
  input activateOut_12a;
  output activateOut_13r;
  input activateOut_13a;
  wire [6:0] internal_0n;
  wire [13:0] acks_0n;
  wire actReq_0n;
  C3 I0 (internal_0n[0], acks_0n[0], acks_0n[1], acks_0n[2]);
  C3 I1 (internal_0n[1], acks_0n[3], acks_0n[4], acks_0n[5]);
  C3 I2 (internal_0n[2], acks_0n[6], acks_0n[7], acks_0n[8]);
  C3 I3 (internal_0n[3], acks_0n[9], acks_0n[10], acks_0n[11]);
  C2 I4 (internal_0n[4], acks_0n[12], acks_0n[13]);
  C3 I5 (internal_0n[5], internal_0n[0], internal_0n[1], internal_0n[2]);
  C2 I6 (internal_0n[6], internal_0n[3], internal_0n[4]);
  C2 I7 (activate_0a, internal_0n[5], internal_0n[6]);
  BALSA_TELEM I8 (actReq_0n, acks_0n[0], activateOut_0r, activateOut_0a);
  BALSA_TELEM I9 (actReq_0n, acks_0n[1], activateOut_1r, activateOut_1a);
  BALSA_TELEM I10 (actReq_0n, acks_0n[2], activateOut_2r, activateOut_2a);
  BALSA_TELEM I11 (actReq_0n, acks_0n[3], activateOut_3r, activateOut_3a);
  BALSA_TELEM I12 (actReq_0n, acks_0n[4], activateOut_4r, activateOut_4a);
  BALSA_TELEM I13 (actReq_0n, acks_0n[5], activateOut_5r, activateOut_5a);
  BALSA_TELEM I14 (actReq_0n, acks_0n[6], activateOut_6r, activateOut_6a);
  BALSA_TELEM I15 (actReq_0n, acks_0n[7], activateOut_7r, activateOut_7a);
  BALSA_TELEM I16 (actReq_0n, acks_0n[8], activateOut_8r, activateOut_8a);
  BALSA_TELEM I17 (actReq_0n, acks_0n[9], activateOut_9r, activateOut_9a);
  BALSA_TELEM I18 (actReq_0n, acks_0n[10], activateOut_10r, activateOut_10a);
  BALSA_TELEM I19 (actReq_0n, acks_0n[11], activateOut_11r, activateOut_11a);
  BALSA_TELEM I20 (actReq_0n, acks_0n[12], activateOut_12r, activateOut_12a);
  BALSA_TELEM I21 (actReq_0n, acks_0n[13], activateOut_13r, activateOut_13a);
  BUFF I22 (actReq_0n, activate_0r);
endmodule

module BrzConstant_1_0 (
  out_0r, out_0a0d, out_0a1d
);
  input out_0r;
  output out_0a0d;
  output out_0a1d;
  wire reqOut_0n;
  supply0 gnd;
  BUFF I0 (out_0a1d, gnd);
  BUFF I1 (out_0a0d, reqOut_0n);
  BUFF I2 (reqOut_0n, out_0r);
endmodule

module BrzConstant_1_1 (
  out_0r, out_0a0d, out_0a1d
);
  input out_0r;
  output out_0a0d;
  output out_0a1d;
  wire reqOut_0n;
  supply0 gnd;
  BUFF I0 (out_0a0d, gnd);
  BUFF I1 (out_0a1d, reqOut_0n);
  BUFF I2 (reqOut_0n, out_0r);
endmodule

module BrzConstant_2_0 (
  out_0r, out_0a0d, out_0a1d
);
  input out_0r;
  output [1:0] out_0a0d;
  output [1:0] out_0a1d;
  wire reqOut_0n;
  supply0 gnd;
  BUFF I0 (out_0a1d[0], gnd);
  BUFF I1 (out_0a1d[1], gnd);
  BUFF I2 (out_0a0d[0], reqOut_0n);
  BUFF I3 (out_0a0d[1], reqOut_0n);
  BUFF I4 (reqOut_0n, out_0r);
endmodule

module BrzConstant_10_511 (
  out_0r, out_0a0d, out_0a1d
);
  input out_0r;
  output [9:0] out_0a0d;
  output [9:0] out_0a1d;
  wire reqOut_0n;
  supply0 gnd;
  BUFF I0 (out_0a1d[9], gnd);
  BUFF I1 (out_0a0d[9], reqOut_0n);
  BUFF I2 (out_0a0d[0], gnd);
  BUFF I3 (out_0a0d[1], gnd);
  BUFF I4 (out_0a0d[2], gnd);
  BUFF I5 (out_0a0d[3], gnd);
  BUFF I6 (out_0a0d[4], gnd);
  BUFF I7 (out_0a0d[5], gnd);
  BUFF I8 (out_0a0d[6], gnd);
  BUFF I9 (out_0a0d[7], gnd);
  BUFF I10 (out_0a0d[8], gnd);
  BUFF I11 (out_0a1d[0], reqOut_0n);
  BUFF I12 (out_0a1d[1], reqOut_0n);
  BUFF I13 (out_0a1d[2], reqOut_0n);
  BUFF I14 (out_0a1d[3], reqOut_0n);
  BUFF I15 (out_0a1d[4], reqOut_0n);
  BUFF I16 (out_0a1d[5], reqOut_0n);
  BUFF I17 (out_0a1d[6], reqOut_0n);
  BUFF I18 (out_0a1d[7], reqOut_0n);
  BUFF I19 (out_0a1d[8], reqOut_0n);
  BUFF I20 (reqOut_0n, out_0r);
endmodule

module BrzConstant_32_0 (
  out_0r, out_0a0d, out_0a1d
);
  input out_0r;
  output [31:0] out_0a0d;
  output [31:0] out_0a1d;
  wire reqOut_0n;
  supply0 gnd;
  BUFF I0 (out_0a1d[0], gnd);
  BUFF I1 (out_0a1d[1], gnd);
  BUFF I2 (out_0a1d[2], gnd);
  BUFF I3 (out_0a1d[3], gnd);
  BUFF I4 (out_0a1d[4], gnd);
  BUFF I5 (out_0a1d[5], gnd);
  BUFF I6 (out_0a1d[6], gnd);
  BUFF I7 (out_0a1d[7], gnd);
  BUFF I8 (out_0a1d[8], gnd);
  BUFF I9 (out_0a1d[9], gnd);
  BUFF I10 (out_0a1d[10], gnd);
  BUFF I11 (out_0a1d[11], gnd);
  BUFF I12 (out_0a1d[12], gnd);
  BUFF I13 (out_0a1d[13], gnd);
  BUFF I14 (out_0a1d[14], gnd);
  BUFF I15 (out_0a1d[15], gnd);
  BUFF I16 (out_0a1d[16], gnd);
  BUFF I17 (out_0a1d[17], gnd);
  BUFF I18 (out_0a1d[18], gnd);
  BUFF I19 (out_0a1d[19], gnd);
  BUFF I20 (out_0a1d[20], gnd);
  BUFF I21 (out_0a1d[21], gnd);
  BUFF I22 (out_0a1d[22], gnd);
  BUFF I23 (out_0a1d[23], gnd);
  BUFF I24 (out_0a1d[24], gnd);
  BUFF I25 (out_0a1d[25], gnd);
  BUFF I26 (out_0a1d[26], gnd);
  BUFF I27 (out_0a1d[27], gnd);
  BUFF I28 (out_0a1d[28], gnd);
  BUFF I29 (out_0a1d[29], gnd);
  BUFF I30 (out_0a1d[30], gnd);
  BUFF I31 (out_0a1d[31], gnd);
  BUFF I32 (out_0a0d[0], reqOut_0n);
  BUFF I33 (out_0a0d[1], reqOut_0n);
  BUFF I34 (out_0a0d[2], reqOut_0n);
  BUFF I35 (out_0a0d[3], reqOut_0n);
  BUFF I36 (out_0a0d[4], reqOut_0n);
  BUFF I37 (out_0a0d[5], reqOut_0n);
  BUFF I38 (out_0a0d[6], reqOut_0n);
  BUFF I39 (out_0a0d[7], reqOut_0n);
  BUFF I40 (out_0a0d[8], reqOut_0n);
  BUFF I41 (out_0a0d[9], reqOut_0n);
  BUFF I42 (out_0a0d[10], reqOut_0n);
  BUFF I43 (out_0a0d[11], reqOut_0n);
  BUFF I44 (out_0a0d[12], reqOut_0n);
  BUFF I45 (out_0a0d[13], reqOut_0n);
  BUFF I46 (out_0a0d[14], reqOut_0n);
  BUFF I47 (out_0a0d[15], reqOut_0n);
  BUFF I48 (out_0a0d[16], reqOut_0n);
  BUFF I49 (out_0a0d[17], reqOut_0n);
  BUFF I50 (out_0a0d[18], reqOut_0n);
  BUFF I51 (out_0a0d[19], reqOut_0n);
  BUFF I52 (out_0a0d[20], reqOut_0n);
  BUFF I53 (out_0a0d[21], reqOut_0n);
  BUFF I54 (out_0a0d[22], reqOut_0n);
  BUFF I55 (out_0a0d[23], reqOut_0n);
  BUFF I56 (out_0a0d[24], reqOut_0n);
  BUFF I57 (out_0a0d[25], reqOut_0n);
  BUFF I58 (out_0a0d[26], reqOut_0n);
  BUFF I59 (out_0a0d[27], reqOut_0n);
  BUFF I60 (out_0a0d[28], reqOut_0n);
  BUFF I61 (out_0a0d[29], reqOut_0n);
  BUFF I62 (out_0a0d[30], reqOut_0n);
  BUFF I63 (out_0a0d[31], reqOut_0n);
  BUFF I64 (reqOut_0n, out_0r);
endmodule

module BrzConstant_35_0 (
  out_0r, out_0a0d, out_0a1d
);
  input out_0r;
  output [34:0] out_0a0d;
  output [34:0] out_0a1d;
  wire reqOut_0n;
  supply0 gnd;
  BUFF I0 (out_0a1d[0], gnd);
  BUFF I1 (out_0a1d[1], gnd);
  BUFF I2 (out_0a1d[2], gnd);
  BUFF I3 (out_0a1d[3], gnd);
  BUFF I4 (out_0a1d[4], gnd);
  BUFF I5 (out_0a1d[5], gnd);
  BUFF I6 (out_0a1d[6], gnd);
  BUFF I7 (out_0a1d[7], gnd);
  BUFF I8 (out_0a1d[8], gnd);
  BUFF I9 (out_0a1d[9], gnd);
  BUFF I10 (out_0a1d[10], gnd);
  BUFF I11 (out_0a1d[11], gnd);
  BUFF I12 (out_0a1d[12], gnd);
  BUFF I13 (out_0a1d[13], gnd);
  BUFF I14 (out_0a1d[14], gnd);
  BUFF I15 (out_0a1d[15], gnd);
  BUFF I16 (out_0a1d[16], gnd);
  BUFF I17 (out_0a1d[17], gnd);
  BUFF I18 (out_0a1d[18], gnd);
  BUFF I19 (out_0a1d[19], gnd);
  BUFF I20 (out_0a1d[20], gnd);
  BUFF I21 (out_0a1d[21], gnd);
  BUFF I22 (out_0a1d[22], gnd);
  BUFF I23 (out_0a1d[23], gnd);
  BUFF I24 (out_0a1d[24], gnd);
  BUFF I25 (out_0a1d[25], gnd);
  BUFF I26 (out_0a1d[26], gnd);
  BUFF I27 (out_0a1d[27], gnd);
  BUFF I28 (out_0a1d[28], gnd);
  BUFF I29 (out_0a1d[29], gnd);
  BUFF I30 (out_0a1d[30], gnd);
  BUFF I31 (out_0a1d[31], gnd);
  BUFF I32 (out_0a1d[32], gnd);
  BUFF I33 (out_0a1d[33], gnd);
  BUFF I34 (out_0a1d[34], gnd);
  BUFF I35 (out_0a0d[0], reqOut_0n);
  BUFF I36 (out_0a0d[1], reqOut_0n);
  BUFF I37 (out_0a0d[2], reqOut_0n);
  BUFF I38 (out_0a0d[3], reqOut_0n);
  BUFF I39 (out_0a0d[4], reqOut_0n);
  BUFF I40 (out_0a0d[5], reqOut_0n);
  BUFF I41 (out_0a0d[6], reqOut_0n);
  BUFF I42 (out_0a0d[7], reqOut_0n);
  BUFF I43 (out_0a0d[8], reqOut_0n);
  BUFF I44 (out_0a0d[9], reqOut_0n);
  BUFF I45 (out_0a0d[10], reqOut_0n);
  BUFF I46 (out_0a0d[11], reqOut_0n);
  BUFF I47 (out_0a0d[12], reqOut_0n);
  BUFF I48 (out_0a0d[13], reqOut_0n);
  BUFF I49 (out_0a0d[14], reqOut_0n);
  BUFF I50 (out_0a0d[15], reqOut_0n);
  BUFF I51 (out_0a0d[16], reqOut_0n);
  BUFF I52 (out_0a0d[17], reqOut_0n);
  BUFF I53 (out_0a0d[18], reqOut_0n);
  BUFF I54 (out_0a0d[19], reqOut_0n);
  BUFF I55 (out_0a0d[20], reqOut_0n);
  BUFF I56 (out_0a0d[21], reqOut_0n);
  BUFF I57 (out_0a0d[22], reqOut_0n);
  BUFF I58 (out_0a0d[23], reqOut_0n);
  BUFF I59 (out_0a0d[24], reqOut_0n);
  BUFF I60 (out_0a0d[25], reqOut_0n);
  BUFF I61 (out_0a0d[26], reqOut_0n);
  BUFF I62 (out_0a0d[27], reqOut_0n);
  BUFF I63 (out_0a0d[28], reqOut_0n);
  BUFF I64 (out_0a0d[29], reqOut_0n);
  BUFF I65 (out_0a0d[30], reqOut_0n);
  BUFF I66 (out_0a0d[31], reqOut_0n);
  BUFF I67 (out_0a0d[32], reqOut_0n);
  BUFF I68 (out_0a0d[33], reqOut_0n);
  BUFF I69 (out_0a0d[34], reqOut_0n);
  BUFF I70 (reqOut_0n, out_0r);
endmodule

module BrzConstant_36_0 (
  out_0r, out_0a0d, out_0a1d
);
  input out_0r;
  output [35:0] out_0a0d;
  output [35:0] out_0a1d;
  wire reqOut_0n;
  supply0 gnd;
  BUFF I0 (out_0a1d[0], gnd);
  BUFF I1 (out_0a1d[1], gnd);
  BUFF I2 (out_0a1d[2], gnd);
  BUFF I3 (out_0a1d[3], gnd);
  BUFF I4 (out_0a1d[4], gnd);
  BUFF I5 (out_0a1d[5], gnd);
  BUFF I6 (out_0a1d[6], gnd);
  BUFF I7 (out_0a1d[7], gnd);
  BUFF I8 (out_0a1d[8], gnd);
  BUFF I9 (out_0a1d[9], gnd);
  BUFF I10 (out_0a1d[10], gnd);
  BUFF I11 (out_0a1d[11], gnd);
  BUFF I12 (out_0a1d[12], gnd);
  BUFF I13 (out_0a1d[13], gnd);
  BUFF I14 (out_0a1d[14], gnd);
  BUFF I15 (out_0a1d[15], gnd);
  BUFF I16 (out_0a1d[16], gnd);
  BUFF I17 (out_0a1d[17], gnd);
  BUFF I18 (out_0a1d[18], gnd);
  BUFF I19 (out_0a1d[19], gnd);
  BUFF I20 (out_0a1d[20], gnd);
  BUFF I21 (out_0a1d[21], gnd);
  BUFF I22 (out_0a1d[22], gnd);
  BUFF I23 (out_0a1d[23], gnd);
  BUFF I24 (out_0a1d[24], gnd);
  BUFF I25 (out_0a1d[25], gnd);
  BUFF I26 (out_0a1d[26], gnd);
  BUFF I27 (out_0a1d[27], gnd);
  BUFF I28 (out_0a1d[28], gnd);
  BUFF I29 (out_0a1d[29], gnd);
  BUFF I30 (out_0a1d[30], gnd);
  BUFF I31 (out_0a1d[31], gnd);
  BUFF I32 (out_0a1d[32], gnd);
  BUFF I33 (out_0a1d[33], gnd);
  BUFF I34 (out_0a1d[34], gnd);
  BUFF I35 (out_0a1d[35], gnd);
  BUFF I36 (out_0a0d[0], reqOut_0n);
  BUFF I37 (out_0a0d[1], reqOut_0n);
  BUFF I38 (out_0a0d[2], reqOut_0n);
  BUFF I39 (out_0a0d[3], reqOut_0n);
  BUFF I40 (out_0a0d[4], reqOut_0n);
  BUFF I41 (out_0a0d[5], reqOut_0n);
  BUFF I42 (out_0a0d[6], reqOut_0n);
  BUFF I43 (out_0a0d[7], reqOut_0n);
  BUFF I44 (out_0a0d[8], reqOut_0n);
  BUFF I45 (out_0a0d[9], reqOut_0n);
  BUFF I46 (out_0a0d[10], reqOut_0n);
  BUFF I47 (out_0a0d[11], reqOut_0n);
  BUFF I48 (out_0a0d[12], reqOut_0n);
  BUFF I49 (out_0a0d[13], reqOut_0n);
  BUFF I50 (out_0a0d[14], reqOut_0n);
  BUFF I51 (out_0a0d[15], reqOut_0n);
  BUFF I52 (out_0a0d[16], reqOut_0n);
  BUFF I53 (out_0a0d[17], reqOut_0n);
  BUFF I54 (out_0a0d[18], reqOut_0n);
  BUFF I55 (out_0a0d[19], reqOut_0n);
  BUFF I56 (out_0a0d[20], reqOut_0n);
  BUFF I57 (out_0a0d[21], reqOut_0n);
  BUFF I58 (out_0a0d[22], reqOut_0n);
  BUFF I59 (out_0a0d[23], reqOut_0n);
  BUFF I60 (out_0a0d[24], reqOut_0n);
  BUFF I61 (out_0a0d[25], reqOut_0n);
  BUFF I62 (out_0a0d[26], reqOut_0n);
  BUFF I63 (out_0a0d[27], reqOut_0n);
  BUFF I64 (out_0a0d[28], reqOut_0n);
  BUFF I65 (out_0a0d[29], reqOut_0n);
  BUFF I66 (out_0a0d[30], reqOut_0n);
  BUFF I67 (out_0a0d[31], reqOut_0n);
  BUFF I68 (out_0a0d[32], reqOut_0n);
  BUFF I69 (out_0a0d[33], reqOut_0n);
  BUFF I70 (out_0a0d[34], reqOut_0n);
  BUFF I71 (out_0a0d[35], reqOut_0n);
  BUFF I72 (reqOut_0n, out_0r);
endmodule

module BrzContinue (
  inp_0r, inp_0a
);
  input inp_0r;
  output inp_0a;
  BUFF I0 (inp_0a, inp_0r);
endmodule

module BrzDecisionWait_1 (
  activate_0r, activate_0a,
  inp_0r, inp_0a,
  out_0r, out_0a
);
  input activate_0r;
  output activate_0a;
  input inp_0r;
  output inp_0a;
  output out_0r;
  input out_0a;
  BUFF I0 (activate_0a, out_0a);
  C2 I1 (out_0r, inp_0r, activate_0r);
  BUFF I2 (inp_0a, out_0a);
endmodule

module BrzEncode_1_2_s5_0_3b0 (
  inp_0r, inp_0a,
  inp_1r, inp_1a,
  out_0r0d, out_0r1d, out_0a
);
  input inp_0r;
  output inp_0a;
  input inp_1r;
  output inp_1a;
  output out_0r0d;
  output out_0r1d;
  input out_0a;
  wire [1:0] data_0n;
  wire [1:0] int1_0n;
  supply0 gnd;
  C2 I0 (inp_0a, data_0n[0], out_0a);
  C2 I1 (inp_1a, data_0n[1], out_0a);
  BUFF I2 (int1_0n[0], data_0n[0]);
  BUFF I3 (int1_0n[1], data_0n[1]);
  OR2 I4 (out_0r0d, int1_0n[0], int1_0n[1]);
  BUFF I5 (out_0r1d, gnd);
  BUFF I6 (data_0n[0], inp_0r);
  BUFF I7 (data_0n[1], inp_1r);
endmodule

module BrzEncode_1_2_s5_1_3b0 (
  inp_0r, inp_0a,
  inp_1r, inp_1a,
  out_0r0d, out_0r1d, out_0a
);
  input inp_0r;
  output inp_0a;
  input inp_1r;
  output inp_1a;
  output out_0r0d;
  output out_0r1d;
  input out_0a;
  wire [1:0] data_0n;
  wire int1_0n;
  wire int0_0n;
  C2 I0 (inp_0a, data_0n[0], out_0a);
  C2 I1 (inp_1a, data_0n[1], out_0a);
  BUFF I2 (int1_0n, data_0n[1]);
  BUFF I3 (out_0r0d, int1_0n);
  BUFF I4 (int0_0n, data_0n[0]);
  BUFF I5 (out_0r1d, int0_0n);
  BUFF I6 (data_0n[0], inp_0r);
  BUFF I7 (data_0n[1], inp_1r);
endmodule

module BrzFalseVariable_1_1_s0_ (
  write_0r0d, write_0r1d, write_0a,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d
);
  input write_0r0d;
  input write_0r1d;
  output write_0a;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output read_0a0d;
  output read_0a1d;
  wire cd_0n;
  wire partCD_0n;
  wire store_0n;
  wire store_1n;
  wire readReq_0n;
  wire sigAck_0n;
  wire writeAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_0a1d, store_1n, readReq_0n);
  AND2 I1 (read_0a0d, store_0n, readReq_0n);
  BUFF I2 (readReq_0n, read_0r);
  BUFF I3 (store_1n, write_0r1d);
  BUFF I4 (store_0n, write_0r0d);
  AND2 I5 (writeAck_0n, sigAck_0n, rReqOr_0n);
  INV I6 (rReqOr_0n, readReq_0n);
  BALSA_TELEM I7 (partCD_0n, sigAck_0n, signal_0r, signal_0a);
  BUFF I8 (write_0a, writeAck_0n);
  OR2 I9 (partCD_0n, store_0n, store_1n);
endmodule

module BrzFalseVariable_3_1_s0_ (
  write_0r0d, write_0r1d, write_0a,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d
);
  input [2:0] write_0r0d;
  input [2:0] write_0r1d;
  output write_0a;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output [2:0] read_0a0d;
  output [2:0] read_0a1d;
  wire cd_0n;
  wire [2:0] partCD_0n;
  wire [2:0] store_0n;
  wire [2:0] store_1n;
  wire readReq_0n;
  wire sigAck_0n;
  wire writeAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I1 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I2 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I3 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I4 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I5 (read_0a0d[2], store_0n[2], readReq_0n);
  BUFF I6 (readReq_0n, read_0r);
  BUFF I7 (store_1n[0], write_0r1d[0]);
  BUFF I8 (store_1n[1], write_0r1d[1]);
  BUFF I9 (store_1n[2], write_0r1d[2]);
  BUFF I10 (store_0n[0], write_0r0d[0]);
  BUFF I11 (store_0n[1], write_0r0d[1]);
  BUFF I12 (store_0n[2], write_0r0d[2]);
  AND2 I13 (writeAck_0n, sigAck_0n, rReqOr_0n);
  INV I14 (rReqOr_0n, readReq_0n);
  BALSA_TELEM I15 (partCD_0n[0], sigAck_0n, signal_0r, signal_0a);
  C2 I16 (write_0a, writeAck_0n, cd_0n);
  C2 I17 (cd_0n, partCD_0n[1], partCD_0n[2]);
  OR2 I18 (partCD_0n[0], store_0n[0], store_1n[0]);
  OR2 I19 (partCD_0n[1], store_0n[1], store_1n[1]);
  OR2 I20 (partCD_0n[2], store_0n[2], store_1n[2]);
endmodule

module BrzFalseVariable_32_1_s0_ (
  write_0r0d, write_0r1d, write_0a,
  signal_0r, signal_0a,
  read_0r, read_0a0d, read_0a1d
);
  input [31:0] write_0r0d;
  input [31:0] write_0r1d;
  output write_0a;
  output signal_0r;
  input signal_0a;
  input read_0r;
  output [31:0] read_0a0d;
  output [31:0] read_0a1d;
  wire [16:0] internal_0n;
  wire cd_0n;
  wire [31:0] partCD_0n;
  wire [31:0] store_0n;
  wire [31:0] store_1n;
  wire readReq_0n;
  wire sigAck_0n;
  wire writeAck_0n;
  wire rReqOr_0n;
  AND2 I0 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I1 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I2 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I3 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I4 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I5 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I6 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I7 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I8 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I9 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I10 (read_0a1d[10], store_1n[10], readReq_0n);
  AND2 I11 (read_0a1d[11], store_1n[11], readReq_0n);
  AND2 I12 (read_0a1d[12], store_1n[12], readReq_0n);
  AND2 I13 (read_0a1d[13], store_1n[13], readReq_0n);
  AND2 I14 (read_0a1d[14], store_1n[14], readReq_0n);
  AND2 I15 (read_0a1d[15], store_1n[15], readReq_0n);
  AND2 I16 (read_0a1d[16], store_1n[16], readReq_0n);
  AND2 I17 (read_0a1d[17], store_1n[17], readReq_0n);
  AND2 I18 (read_0a1d[18], store_1n[18], readReq_0n);
  AND2 I19 (read_0a1d[19], store_1n[19], readReq_0n);
  AND2 I20 (read_0a1d[20], store_1n[20], readReq_0n);
  AND2 I21 (read_0a1d[21], store_1n[21], readReq_0n);
  AND2 I22 (read_0a1d[22], store_1n[22], readReq_0n);
  AND2 I23 (read_0a1d[23], store_1n[23], readReq_0n);
  AND2 I24 (read_0a1d[24], store_1n[24], readReq_0n);
  AND2 I25 (read_0a1d[25], store_1n[25], readReq_0n);
  AND2 I26 (read_0a1d[26], store_1n[26], readReq_0n);
  AND2 I27 (read_0a1d[27], store_1n[27], readReq_0n);
  AND2 I28 (read_0a1d[28], store_1n[28], readReq_0n);
  AND2 I29 (read_0a1d[29], store_1n[29], readReq_0n);
  AND2 I30 (read_0a1d[30], store_1n[30], readReq_0n);
  AND2 I31 (read_0a1d[31], store_1n[31], readReq_0n);
  AND2 I32 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I33 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I34 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I35 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I36 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I37 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I38 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I39 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I40 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I41 (read_0a0d[9], store_0n[9], readReq_0n);
  AND2 I42 (read_0a0d[10], store_0n[10], readReq_0n);
  AND2 I43 (read_0a0d[11], store_0n[11], readReq_0n);
  AND2 I44 (read_0a0d[12], store_0n[12], readReq_0n);
  AND2 I45 (read_0a0d[13], store_0n[13], readReq_0n);
  AND2 I46 (read_0a0d[14], store_0n[14], readReq_0n);
  AND2 I47 (read_0a0d[15], store_0n[15], readReq_0n);
  AND2 I48 (read_0a0d[16], store_0n[16], readReq_0n);
  AND2 I49 (read_0a0d[17], store_0n[17], readReq_0n);
  AND2 I50 (read_0a0d[18], store_0n[18], readReq_0n);
  AND2 I51 (read_0a0d[19], store_0n[19], readReq_0n);
  AND2 I52 (read_0a0d[20], store_0n[20], readReq_0n);
  AND2 I53 (read_0a0d[21], store_0n[21], readReq_0n);
  AND2 I54 (read_0a0d[22], store_0n[22], readReq_0n);
  AND2 I55 (read_0a0d[23], store_0n[23], readReq_0n);
  AND2 I56 (read_0a0d[24], store_0n[24], readReq_0n);
  AND2 I57 (read_0a0d[25], store_0n[25], readReq_0n);
  AND2 I58 (read_0a0d[26], store_0n[26], readReq_0n);
  AND2 I59 (read_0a0d[27], store_0n[27], readReq_0n);
  AND2 I60 (read_0a0d[28], store_0n[28], readReq_0n);
  AND2 I61 (read_0a0d[29], store_0n[29], readReq_0n);
  AND2 I62 (read_0a0d[30], store_0n[30], readReq_0n);
  AND2 I63 (read_0a0d[31], store_0n[31], readReq_0n);
  BUFF I64 (readReq_0n, read_0r);
  BUFF I65 (store_1n[0], write_0r1d[0]);
  BUFF I66 (store_1n[1], write_0r1d[1]);
  BUFF I67 (store_1n[2], write_0r1d[2]);
  BUFF I68 (store_1n[3], write_0r1d[3]);
  BUFF I69 (store_1n[4], write_0r1d[4]);
  BUFF I70 (store_1n[5], write_0r1d[5]);
  BUFF I71 (store_1n[6], write_0r1d[6]);
  BUFF I72 (store_1n[7], write_0r1d[7]);
  BUFF I73 (store_1n[8], write_0r1d[8]);
  BUFF I74 (store_1n[9], write_0r1d[9]);
  BUFF I75 (store_1n[10], write_0r1d[10]);
  BUFF I76 (store_1n[11], write_0r1d[11]);
  BUFF I77 (store_1n[12], write_0r1d[12]);
  BUFF I78 (store_1n[13], write_0r1d[13]);
  BUFF I79 (store_1n[14], write_0r1d[14]);
  BUFF I80 (store_1n[15], write_0r1d[15]);
  BUFF I81 (store_1n[16], write_0r1d[16]);
  BUFF I82 (store_1n[17], write_0r1d[17]);
  BUFF I83 (store_1n[18], write_0r1d[18]);
  BUFF I84 (store_1n[19], write_0r1d[19]);
  BUFF I85 (store_1n[20], write_0r1d[20]);
  BUFF I86 (store_1n[21], write_0r1d[21]);
  BUFF I87 (store_1n[22], write_0r1d[22]);
  BUFF I88 (store_1n[23], write_0r1d[23]);
  BUFF I89 (store_1n[24], write_0r1d[24]);
  BUFF I90 (store_1n[25], write_0r1d[25]);
  BUFF I91 (store_1n[26], write_0r1d[26]);
  BUFF I92 (store_1n[27], write_0r1d[27]);
  BUFF I93 (store_1n[28], write_0r1d[28]);
  BUFF I94 (store_1n[29], write_0r1d[29]);
  BUFF I95 (store_1n[30], write_0r1d[30]);
  BUFF I96 (store_1n[31], write_0r1d[31]);
  BUFF I97 (store_0n[0], write_0r0d[0]);
  BUFF I98 (store_0n[1], write_0r0d[1]);
  BUFF I99 (store_0n[2], write_0r0d[2]);
  BUFF I100 (store_0n[3], write_0r0d[3]);
  BUFF I101 (store_0n[4], write_0r0d[4]);
  BUFF I102 (store_0n[5], write_0r0d[5]);
  BUFF I103 (store_0n[6], write_0r0d[6]);
  BUFF I104 (store_0n[7], write_0r0d[7]);
  BUFF I105 (store_0n[8], write_0r0d[8]);
  BUFF I106 (store_0n[9], write_0r0d[9]);
  BUFF I107 (store_0n[10], write_0r0d[10]);
  BUFF I108 (store_0n[11], write_0r0d[11]);
  BUFF I109 (store_0n[12], write_0r0d[12]);
  BUFF I110 (store_0n[13], write_0r0d[13]);
  BUFF I111 (store_0n[14], write_0r0d[14]);
  BUFF I112 (store_0n[15], write_0r0d[15]);
  BUFF I113 (store_0n[16], write_0r0d[16]);
  BUFF I114 (store_0n[17], write_0r0d[17]);
  BUFF I115 (store_0n[18], write_0r0d[18]);
  BUFF I116 (store_0n[19], write_0r0d[19]);
  BUFF I117 (store_0n[20], write_0r0d[20]);
  BUFF I118 (store_0n[21], write_0r0d[21]);
  BUFF I119 (store_0n[22], write_0r0d[22]);
  BUFF I120 (store_0n[23], write_0r0d[23]);
  BUFF I121 (store_0n[24], write_0r0d[24]);
  BUFF I122 (store_0n[25], write_0r0d[25]);
  BUFF I123 (store_0n[26], write_0r0d[26]);
  BUFF I124 (store_0n[27], write_0r0d[27]);
  BUFF I125 (store_0n[28], write_0r0d[28]);
  BUFF I126 (store_0n[29], write_0r0d[29]);
  BUFF I127 (store_0n[30], write_0r0d[30]);
  BUFF I128 (store_0n[31], write_0r0d[31]);
  AND2 I129 (writeAck_0n, sigAck_0n, rReqOr_0n);
  INV I130 (rReqOr_0n, readReq_0n);
  BALSA_TELEM I131 (partCD_0n[0], sigAck_0n, signal_0r, signal_0a);
  C2 I132 (write_0a, writeAck_0n, cd_0n);
  C3 I133 (internal_0n[0], partCD_0n[1], partCD_0n[2], partCD_0n[3]);
  C3 I134 (internal_0n[1], partCD_0n[4], partCD_0n[5], partCD_0n[6]);
  C3 I135 (internal_0n[2], partCD_0n[7], partCD_0n[8], partCD_0n[9]);
  C3 I136 (internal_0n[3], partCD_0n[10], partCD_0n[11], partCD_0n[12]);
  C3 I137 (internal_0n[4], partCD_0n[13], partCD_0n[14], partCD_0n[15]);
  C3 I138 (internal_0n[5], partCD_0n[16], partCD_0n[17], partCD_0n[18]);
  C3 I139 (internal_0n[6], partCD_0n[19], partCD_0n[20], partCD_0n[21]);
  C3 I140 (internal_0n[7], partCD_0n[22], partCD_0n[23], partCD_0n[24]);
  C3 I141 (internal_0n[8], partCD_0n[25], partCD_0n[26], partCD_0n[27]);
  C2 I142 (internal_0n[9], partCD_0n[28], partCD_0n[29]);
  C2 I143 (internal_0n[10], partCD_0n[30], partCD_0n[31]);
  C3 I144 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I145 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I146 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I147 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I148 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I149 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I150 (cd_0n, internal_0n[15], internal_0n[16]);
  OR2 I151 (partCD_0n[0], store_0n[0], store_1n[0]);
  OR2 I152 (partCD_0n[1], store_0n[1], store_1n[1]);
  OR2 I153 (partCD_0n[2], store_0n[2], store_1n[2]);
  OR2 I154 (partCD_0n[3], store_0n[3], store_1n[3]);
  OR2 I155 (partCD_0n[4], store_0n[4], store_1n[4]);
  OR2 I156 (partCD_0n[5], store_0n[5], store_1n[5]);
  OR2 I157 (partCD_0n[6], store_0n[6], store_1n[6]);
  OR2 I158 (partCD_0n[7], store_0n[7], store_1n[7]);
  OR2 I159 (partCD_0n[8], store_0n[8], store_1n[8]);
  OR2 I160 (partCD_0n[9], store_0n[9], store_1n[9]);
  OR2 I161 (partCD_0n[10], store_0n[10], store_1n[10]);
  OR2 I162 (partCD_0n[11], store_0n[11], store_1n[11]);
  OR2 I163 (partCD_0n[12], store_0n[12], store_1n[12]);
  OR2 I164 (partCD_0n[13], store_0n[13], store_1n[13]);
  OR2 I165 (partCD_0n[14], store_0n[14], store_1n[14]);
  OR2 I166 (partCD_0n[15], store_0n[15], store_1n[15]);
  OR2 I167 (partCD_0n[16], store_0n[16], store_1n[16]);
  OR2 I168 (partCD_0n[17], store_0n[17], store_1n[17]);
  OR2 I169 (partCD_0n[18], store_0n[18], store_1n[18]);
  OR2 I170 (partCD_0n[19], store_0n[19], store_1n[19]);
  OR2 I171 (partCD_0n[20], store_0n[20], store_1n[20]);
  OR2 I172 (partCD_0n[21], store_0n[21], store_1n[21]);
  OR2 I173 (partCD_0n[22], store_0n[22], store_1n[22]);
  OR2 I174 (partCD_0n[23], store_0n[23], store_1n[23]);
  OR2 I175 (partCD_0n[24], store_0n[24], store_1n[24]);
  OR2 I176 (partCD_0n[25], store_0n[25], store_1n[25]);
  OR2 I177 (partCD_0n[26], store_0n[26], store_1n[26]);
  OR2 I178 (partCD_0n[27], store_0n[27], store_1n[27]);
  OR2 I179 (partCD_0n[28], store_0n[28], store_1n[28]);
  OR2 I180 (partCD_0n[29], store_0n[29], store_1n[29]);
  OR2 I181 (partCD_0n[30], store_0n[30], store_1n[30]);
  OR2 I182 (partCD_0n[31], store_0n[31], store_1n[31]);
endmodule

module BrzFetch_1_s5_false (
  activate_0r, activate_0a,
  inp_0r, inp_0a0d, inp_0a1d,
  out_0r0d, out_0r1d, out_0a
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input inp_0a0d;
  input inp_0a1d;
  output out_0r0d;
  output out_0r1d;
  input out_0a;
  BUFF I0 (inp_0r, activate_0r);
  BUFF I1 (out_0r0d, inp_0a0d);
  BUFF I2 (out_0r1d, inp_0a1d);
  BUFF I3 (activate_0a, out_0a);
endmodule

module BrzFetch_1_s4_true (
  activate_0r, activate_0a,
  inp_0r, inp_0a0d, inp_0a1d,
  out_0r0d, out_0r1d, out_0a
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input inp_0a0d;
  input inp_0a1d;
  output out_0r0d;
  output out_0r1d;
  input out_0a;
  BUFF I0 (inp_0r, activate_0r);
  BUFF I1 (out_0r0d, inp_0a0d);
  BUFF I2 (out_0r1d, inp_0a1d);
  BUFF I3 (activate_0a, out_0a);
endmodule

module BrzFetch_3_s5_false (
  activate_0r, activate_0a,
  inp_0r, inp_0a0d, inp_0a1d,
  out_0r0d, out_0r1d, out_0a
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input [2:0] inp_0a0d;
  input [2:0] inp_0a1d;
  output [2:0] out_0r0d;
  output [2:0] out_0r1d;
  input out_0a;
  BUFF I0 (inp_0r, activate_0r);
  BUFF I1 (out_0r0d[0], inp_0a0d[0]);
  BUFF I2 (out_0r0d[1], inp_0a0d[1]);
  BUFF I3 (out_0r0d[2], inp_0a0d[2]);
  BUFF I4 (out_0r1d[0], inp_0a1d[0]);
  BUFF I5 (out_0r1d[1], inp_0a1d[1]);
  BUFF I6 (out_0r1d[2], inp_0a1d[2]);
  BUFF I7 (activate_0a, out_0a);
endmodule

module BrzFetch_4_s5_false (
  activate_0r, activate_0a,
  inp_0r, inp_0a0d, inp_0a1d,
  out_0r0d, out_0r1d, out_0a
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input [3:0] inp_0a0d;
  input [3:0] inp_0a1d;
  output [3:0] out_0r0d;
  output [3:0] out_0r1d;
  input out_0a;
  BUFF I0 (inp_0r, activate_0r);
  BUFF I1 (out_0r0d[0], inp_0a0d[0]);
  BUFF I2 (out_0r0d[1], inp_0a0d[1]);
  BUFF I3 (out_0r0d[2], inp_0a0d[2]);
  BUFF I4 (out_0r0d[3], inp_0a0d[3]);
  BUFF I5 (out_0r1d[0], inp_0a1d[0]);
  BUFF I6 (out_0r1d[1], inp_0a1d[1]);
  BUFF I7 (out_0r1d[2], inp_0a1d[2]);
  BUFF I8 (out_0r1d[3], inp_0a1d[3]);
  BUFF I9 (activate_0a, out_0a);
endmodule

module BrzFetch_10_s5_false (
  activate_0r, activate_0a,
  inp_0r, inp_0a0d, inp_0a1d,
  out_0r0d, out_0r1d, out_0a
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input [9:0] inp_0a0d;
  input [9:0] inp_0a1d;
  output [9:0] out_0r0d;
  output [9:0] out_0r1d;
  input out_0a;
  BUFF I0 (inp_0r, activate_0r);
  BUFF I1 (out_0r0d[0], inp_0a0d[0]);
  BUFF I2 (out_0r0d[1], inp_0a0d[1]);
  BUFF I3 (out_0r0d[2], inp_0a0d[2]);
  BUFF I4 (out_0r0d[3], inp_0a0d[3]);
  BUFF I5 (out_0r0d[4], inp_0a0d[4]);
  BUFF I6 (out_0r0d[5], inp_0a0d[5]);
  BUFF I7 (out_0r0d[6], inp_0a0d[6]);
  BUFF I8 (out_0r0d[7], inp_0a0d[7]);
  BUFF I9 (out_0r0d[8], inp_0a0d[8]);
  BUFF I10 (out_0r0d[9], inp_0a0d[9]);
  BUFF I11 (out_0r1d[0], inp_0a1d[0]);
  BUFF I12 (out_0r1d[1], inp_0a1d[1]);
  BUFF I13 (out_0r1d[2], inp_0a1d[2]);
  BUFF I14 (out_0r1d[3], inp_0a1d[3]);
  BUFF I15 (out_0r1d[4], inp_0a1d[4]);
  BUFF I16 (out_0r1d[5], inp_0a1d[5]);
  BUFF I17 (out_0r1d[6], inp_0a1d[6]);
  BUFF I18 (out_0r1d[7], inp_0a1d[7]);
  BUFF I19 (out_0r1d[8], inp_0a1d[8]);
  BUFF I20 (out_0r1d[9], inp_0a1d[9]);
  BUFF I21 (activate_0a, out_0a);
endmodule

module BrzFetch_32_s5_false (
  activate_0r, activate_0a,
  inp_0r, inp_0a0d, inp_0a1d,
  out_0r0d, out_0r1d, out_0a
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input [31:0] inp_0a0d;
  input [31:0] inp_0a1d;
  output [31:0] out_0r0d;
  output [31:0] out_0r1d;
  input out_0a;
  BUFF I0 (inp_0r, activate_0r);
  BUFF I1 (out_0r0d[0], inp_0a0d[0]);
  BUFF I2 (out_0r0d[1], inp_0a0d[1]);
  BUFF I3 (out_0r0d[2], inp_0a0d[2]);
  BUFF I4 (out_0r0d[3], inp_0a0d[3]);
  BUFF I5 (out_0r0d[4], inp_0a0d[4]);
  BUFF I6 (out_0r0d[5], inp_0a0d[5]);
  BUFF I7 (out_0r0d[6], inp_0a0d[6]);
  BUFF I8 (out_0r0d[7], inp_0a0d[7]);
  BUFF I9 (out_0r0d[8], inp_0a0d[8]);
  BUFF I10 (out_0r0d[9], inp_0a0d[9]);
  BUFF I11 (out_0r0d[10], inp_0a0d[10]);
  BUFF I12 (out_0r0d[11], inp_0a0d[11]);
  BUFF I13 (out_0r0d[12], inp_0a0d[12]);
  BUFF I14 (out_0r0d[13], inp_0a0d[13]);
  BUFF I15 (out_0r0d[14], inp_0a0d[14]);
  BUFF I16 (out_0r0d[15], inp_0a0d[15]);
  BUFF I17 (out_0r0d[16], inp_0a0d[16]);
  BUFF I18 (out_0r0d[17], inp_0a0d[17]);
  BUFF I19 (out_0r0d[18], inp_0a0d[18]);
  BUFF I20 (out_0r0d[19], inp_0a0d[19]);
  BUFF I21 (out_0r0d[20], inp_0a0d[20]);
  BUFF I22 (out_0r0d[21], inp_0a0d[21]);
  BUFF I23 (out_0r0d[22], inp_0a0d[22]);
  BUFF I24 (out_0r0d[23], inp_0a0d[23]);
  BUFF I25 (out_0r0d[24], inp_0a0d[24]);
  BUFF I26 (out_0r0d[25], inp_0a0d[25]);
  BUFF I27 (out_0r0d[26], inp_0a0d[26]);
  BUFF I28 (out_0r0d[27], inp_0a0d[27]);
  BUFF I29 (out_0r0d[28], inp_0a0d[28]);
  BUFF I30 (out_0r0d[29], inp_0a0d[29]);
  BUFF I31 (out_0r0d[30], inp_0a0d[30]);
  BUFF I32 (out_0r0d[31], inp_0a0d[31]);
  BUFF I33 (out_0r1d[0], inp_0a1d[0]);
  BUFF I34 (out_0r1d[1], inp_0a1d[1]);
  BUFF I35 (out_0r1d[2], inp_0a1d[2]);
  BUFF I36 (out_0r1d[3], inp_0a1d[3]);
  BUFF I37 (out_0r1d[4], inp_0a1d[4]);
  BUFF I38 (out_0r1d[5], inp_0a1d[5]);
  BUFF I39 (out_0r1d[6], inp_0a1d[6]);
  BUFF I40 (out_0r1d[7], inp_0a1d[7]);
  BUFF I41 (out_0r1d[8], inp_0a1d[8]);
  BUFF I42 (out_0r1d[9], inp_0a1d[9]);
  BUFF I43 (out_0r1d[10], inp_0a1d[10]);
  BUFF I44 (out_0r1d[11], inp_0a1d[11]);
  BUFF I45 (out_0r1d[12], inp_0a1d[12]);
  BUFF I46 (out_0r1d[13], inp_0a1d[13]);
  BUFF I47 (out_0r1d[14], inp_0a1d[14]);
  BUFF I48 (out_0r1d[15], inp_0a1d[15]);
  BUFF I49 (out_0r1d[16], inp_0a1d[16]);
  BUFF I50 (out_0r1d[17], inp_0a1d[17]);
  BUFF I51 (out_0r1d[18], inp_0a1d[18]);
  BUFF I52 (out_0r1d[19], inp_0a1d[19]);
  BUFF I53 (out_0r1d[20], inp_0a1d[20]);
  BUFF I54 (out_0r1d[21], inp_0a1d[21]);
  BUFF I55 (out_0r1d[22], inp_0a1d[22]);
  BUFF I56 (out_0r1d[23], inp_0a1d[23]);
  BUFF I57 (out_0r1d[24], inp_0a1d[24]);
  BUFF I58 (out_0r1d[25], inp_0a1d[25]);
  BUFF I59 (out_0r1d[26], inp_0a1d[26]);
  BUFF I60 (out_0r1d[27], inp_0a1d[27]);
  BUFF I61 (out_0r1d[28], inp_0a1d[28]);
  BUFF I62 (out_0r1d[29], inp_0a1d[29]);
  BUFF I63 (out_0r1d[30], inp_0a1d[30]);
  BUFF I64 (out_0r1d[31], inp_0a1d[31]);
  BUFF I65 (activate_0a, out_0a);
endmodule

module BrzFetch_32_s4_true (
  activate_0r, activate_0a,
  inp_0r, inp_0a0d, inp_0a1d,
  out_0r0d, out_0r1d, out_0a
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input [31:0] inp_0a0d;
  input [31:0] inp_0a1d;
  output [31:0] out_0r0d;
  output [31:0] out_0r1d;
  input out_0a;
  BUFF I0 (inp_0r, activate_0r);
  BUFF I1 (out_0r0d[0], inp_0a0d[0]);
  BUFF I2 (out_0r0d[1], inp_0a0d[1]);
  BUFF I3 (out_0r0d[2], inp_0a0d[2]);
  BUFF I4 (out_0r0d[3], inp_0a0d[3]);
  BUFF I5 (out_0r0d[4], inp_0a0d[4]);
  BUFF I6 (out_0r0d[5], inp_0a0d[5]);
  BUFF I7 (out_0r0d[6], inp_0a0d[6]);
  BUFF I8 (out_0r0d[7], inp_0a0d[7]);
  BUFF I9 (out_0r0d[8], inp_0a0d[8]);
  BUFF I10 (out_0r0d[9], inp_0a0d[9]);
  BUFF I11 (out_0r0d[10], inp_0a0d[10]);
  BUFF I12 (out_0r0d[11], inp_0a0d[11]);
  BUFF I13 (out_0r0d[12], inp_0a0d[12]);
  BUFF I14 (out_0r0d[13], inp_0a0d[13]);
  BUFF I15 (out_0r0d[14], inp_0a0d[14]);
  BUFF I16 (out_0r0d[15], inp_0a0d[15]);
  BUFF I17 (out_0r0d[16], inp_0a0d[16]);
  BUFF I18 (out_0r0d[17], inp_0a0d[17]);
  BUFF I19 (out_0r0d[18], inp_0a0d[18]);
  BUFF I20 (out_0r0d[19], inp_0a0d[19]);
  BUFF I21 (out_0r0d[20], inp_0a0d[20]);
  BUFF I22 (out_0r0d[21], inp_0a0d[21]);
  BUFF I23 (out_0r0d[22], inp_0a0d[22]);
  BUFF I24 (out_0r0d[23], inp_0a0d[23]);
  BUFF I25 (out_0r0d[24], inp_0a0d[24]);
  BUFF I26 (out_0r0d[25], inp_0a0d[25]);
  BUFF I27 (out_0r0d[26], inp_0a0d[26]);
  BUFF I28 (out_0r0d[27], inp_0a0d[27]);
  BUFF I29 (out_0r0d[28], inp_0a0d[28]);
  BUFF I30 (out_0r0d[29], inp_0a0d[29]);
  BUFF I31 (out_0r0d[30], inp_0a0d[30]);
  BUFF I32 (out_0r0d[31], inp_0a0d[31]);
  BUFF I33 (out_0r1d[0], inp_0a1d[0]);
  BUFF I34 (out_0r1d[1], inp_0a1d[1]);
  BUFF I35 (out_0r1d[2], inp_0a1d[2]);
  BUFF I36 (out_0r1d[3], inp_0a1d[3]);
  BUFF I37 (out_0r1d[4], inp_0a1d[4]);
  BUFF I38 (out_0r1d[5], inp_0a1d[5]);
  BUFF I39 (out_0r1d[6], inp_0a1d[6]);
  BUFF I40 (out_0r1d[7], inp_0a1d[7]);
  BUFF I41 (out_0r1d[8], inp_0a1d[8]);
  BUFF I42 (out_0r1d[9], inp_0a1d[9]);
  BUFF I43 (out_0r1d[10], inp_0a1d[10]);
  BUFF I44 (out_0r1d[11], inp_0a1d[11]);
  BUFF I45 (out_0r1d[12], inp_0a1d[12]);
  BUFF I46 (out_0r1d[13], inp_0a1d[13]);
  BUFF I47 (out_0r1d[14], inp_0a1d[14]);
  BUFF I48 (out_0r1d[15], inp_0a1d[15]);
  BUFF I49 (out_0r1d[16], inp_0a1d[16]);
  BUFF I50 (out_0r1d[17], inp_0a1d[17]);
  BUFF I51 (out_0r1d[18], inp_0a1d[18]);
  BUFF I52 (out_0r1d[19], inp_0a1d[19]);
  BUFF I53 (out_0r1d[20], inp_0a1d[20]);
  BUFF I54 (out_0r1d[21], inp_0a1d[21]);
  BUFF I55 (out_0r1d[22], inp_0a1d[22]);
  BUFF I56 (out_0r1d[23], inp_0a1d[23]);
  BUFF I57 (out_0r1d[24], inp_0a1d[24]);
  BUFF I58 (out_0r1d[25], inp_0a1d[25]);
  BUFF I59 (out_0r1d[26], inp_0a1d[26]);
  BUFF I60 (out_0r1d[27], inp_0a1d[27]);
  BUFF I61 (out_0r1d[28], inp_0a1d[28]);
  BUFF I62 (out_0r1d[29], inp_0a1d[29]);
  BUFF I63 (out_0r1d[30], inp_0a1d[30]);
  BUFF I64 (out_0r1d[31], inp_0a1d[31]);
  BUFF I65 (activate_0a, out_0a);
endmodule

module BrzFetch_33_s5_false (
  activate_0r, activate_0a,
  inp_0r, inp_0a0d, inp_0a1d,
  out_0r0d, out_0r1d, out_0a
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input [32:0] inp_0a0d;
  input [32:0] inp_0a1d;
  output [32:0] out_0r0d;
  output [32:0] out_0r1d;
  input out_0a;
  BUFF I0 (inp_0r, activate_0r);
  BUFF I1 (out_0r0d[0], inp_0a0d[0]);
  BUFF I2 (out_0r0d[1], inp_0a0d[1]);
  BUFF I3 (out_0r0d[2], inp_0a0d[2]);
  BUFF I4 (out_0r0d[3], inp_0a0d[3]);
  BUFF I5 (out_0r0d[4], inp_0a0d[4]);
  BUFF I6 (out_0r0d[5], inp_0a0d[5]);
  BUFF I7 (out_0r0d[6], inp_0a0d[6]);
  BUFF I8 (out_0r0d[7], inp_0a0d[7]);
  BUFF I9 (out_0r0d[8], inp_0a0d[8]);
  BUFF I10 (out_0r0d[9], inp_0a0d[9]);
  BUFF I11 (out_0r0d[10], inp_0a0d[10]);
  BUFF I12 (out_0r0d[11], inp_0a0d[11]);
  BUFF I13 (out_0r0d[12], inp_0a0d[12]);
  BUFF I14 (out_0r0d[13], inp_0a0d[13]);
  BUFF I15 (out_0r0d[14], inp_0a0d[14]);
  BUFF I16 (out_0r0d[15], inp_0a0d[15]);
  BUFF I17 (out_0r0d[16], inp_0a0d[16]);
  BUFF I18 (out_0r0d[17], inp_0a0d[17]);
  BUFF I19 (out_0r0d[18], inp_0a0d[18]);
  BUFF I20 (out_0r0d[19], inp_0a0d[19]);
  BUFF I21 (out_0r0d[20], inp_0a0d[20]);
  BUFF I22 (out_0r0d[21], inp_0a0d[21]);
  BUFF I23 (out_0r0d[22], inp_0a0d[22]);
  BUFF I24 (out_0r0d[23], inp_0a0d[23]);
  BUFF I25 (out_0r0d[24], inp_0a0d[24]);
  BUFF I26 (out_0r0d[25], inp_0a0d[25]);
  BUFF I27 (out_0r0d[26], inp_0a0d[26]);
  BUFF I28 (out_0r0d[27], inp_0a0d[27]);
  BUFF I29 (out_0r0d[28], inp_0a0d[28]);
  BUFF I30 (out_0r0d[29], inp_0a0d[29]);
  BUFF I31 (out_0r0d[30], inp_0a0d[30]);
  BUFF I32 (out_0r0d[31], inp_0a0d[31]);
  BUFF I33 (out_0r0d[32], inp_0a0d[32]);
  BUFF I34 (out_0r1d[0], inp_0a1d[0]);
  BUFF I35 (out_0r1d[1], inp_0a1d[1]);
  BUFF I36 (out_0r1d[2], inp_0a1d[2]);
  BUFF I37 (out_0r1d[3], inp_0a1d[3]);
  BUFF I38 (out_0r1d[4], inp_0a1d[4]);
  BUFF I39 (out_0r1d[5], inp_0a1d[5]);
  BUFF I40 (out_0r1d[6], inp_0a1d[6]);
  BUFF I41 (out_0r1d[7], inp_0a1d[7]);
  BUFF I42 (out_0r1d[8], inp_0a1d[8]);
  BUFF I43 (out_0r1d[9], inp_0a1d[9]);
  BUFF I44 (out_0r1d[10], inp_0a1d[10]);
  BUFF I45 (out_0r1d[11], inp_0a1d[11]);
  BUFF I46 (out_0r1d[12], inp_0a1d[12]);
  BUFF I47 (out_0r1d[13], inp_0a1d[13]);
  BUFF I48 (out_0r1d[14], inp_0a1d[14]);
  BUFF I49 (out_0r1d[15], inp_0a1d[15]);
  BUFF I50 (out_0r1d[16], inp_0a1d[16]);
  BUFF I51 (out_0r1d[17], inp_0a1d[17]);
  BUFF I52 (out_0r1d[18], inp_0a1d[18]);
  BUFF I53 (out_0r1d[19], inp_0a1d[19]);
  BUFF I54 (out_0r1d[20], inp_0a1d[20]);
  BUFF I55 (out_0r1d[21], inp_0a1d[21]);
  BUFF I56 (out_0r1d[22], inp_0a1d[22]);
  BUFF I57 (out_0r1d[23], inp_0a1d[23]);
  BUFF I58 (out_0r1d[24], inp_0a1d[24]);
  BUFF I59 (out_0r1d[25], inp_0a1d[25]);
  BUFF I60 (out_0r1d[26], inp_0a1d[26]);
  BUFF I61 (out_0r1d[27], inp_0a1d[27]);
  BUFF I62 (out_0r1d[28], inp_0a1d[28]);
  BUFF I63 (out_0r1d[29], inp_0a1d[29]);
  BUFF I64 (out_0r1d[30], inp_0a1d[30]);
  BUFF I65 (out_0r1d[31], inp_0a1d[31]);
  BUFF I66 (out_0r1d[32], inp_0a1d[32]);
  BUFF I67 (activate_0a, out_0a);
endmodule

module BrzFetch_34_s5_false (
  activate_0r, activate_0a,
  inp_0r, inp_0a0d, inp_0a1d,
  out_0r0d, out_0r1d, out_0a
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input [33:0] inp_0a0d;
  input [33:0] inp_0a1d;
  output [33:0] out_0r0d;
  output [33:0] out_0r1d;
  input out_0a;
  BUFF I0 (inp_0r, activate_0r);
  BUFF I1 (out_0r0d[0], inp_0a0d[0]);
  BUFF I2 (out_0r0d[1], inp_0a0d[1]);
  BUFF I3 (out_0r0d[2], inp_0a0d[2]);
  BUFF I4 (out_0r0d[3], inp_0a0d[3]);
  BUFF I5 (out_0r0d[4], inp_0a0d[4]);
  BUFF I6 (out_0r0d[5], inp_0a0d[5]);
  BUFF I7 (out_0r0d[6], inp_0a0d[6]);
  BUFF I8 (out_0r0d[7], inp_0a0d[7]);
  BUFF I9 (out_0r0d[8], inp_0a0d[8]);
  BUFF I10 (out_0r0d[9], inp_0a0d[9]);
  BUFF I11 (out_0r0d[10], inp_0a0d[10]);
  BUFF I12 (out_0r0d[11], inp_0a0d[11]);
  BUFF I13 (out_0r0d[12], inp_0a0d[12]);
  BUFF I14 (out_0r0d[13], inp_0a0d[13]);
  BUFF I15 (out_0r0d[14], inp_0a0d[14]);
  BUFF I16 (out_0r0d[15], inp_0a0d[15]);
  BUFF I17 (out_0r0d[16], inp_0a0d[16]);
  BUFF I18 (out_0r0d[17], inp_0a0d[17]);
  BUFF I19 (out_0r0d[18], inp_0a0d[18]);
  BUFF I20 (out_0r0d[19], inp_0a0d[19]);
  BUFF I21 (out_0r0d[20], inp_0a0d[20]);
  BUFF I22 (out_0r0d[21], inp_0a0d[21]);
  BUFF I23 (out_0r0d[22], inp_0a0d[22]);
  BUFF I24 (out_0r0d[23], inp_0a0d[23]);
  BUFF I25 (out_0r0d[24], inp_0a0d[24]);
  BUFF I26 (out_0r0d[25], inp_0a0d[25]);
  BUFF I27 (out_0r0d[26], inp_0a0d[26]);
  BUFF I28 (out_0r0d[27], inp_0a0d[27]);
  BUFF I29 (out_0r0d[28], inp_0a0d[28]);
  BUFF I30 (out_0r0d[29], inp_0a0d[29]);
  BUFF I31 (out_0r0d[30], inp_0a0d[30]);
  BUFF I32 (out_0r0d[31], inp_0a0d[31]);
  BUFF I33 (out_0r0d[32], inp_0a0d[32]);
  BUFF I34 (out_0r0d[33], inp_0a0d[33]);
  BUFF I35 (out_0r1d[0], inp_0a1d[0]);
  BUFF I36 (out_0r1d[1], inp_0a1d[1]);
  BUFF I37 (out_0r1d[2], inp_0a1d[2]);
  BUFF I38 (out_0r1d[3], inp_0a1d[3]);
  BUFF I39 (out_0r1d[4], inp_0a1d[4]);
  BUFF I40 (out_0r1d[5], inp_0a1d[5]);
  BUFF I41 (out_0r1d[6], inp_0a1d[6]);
  BUFF I42 (out_0r1d[7], inp_0a1d[7]);
  BUFF I43 (out_0r1d[8], inp_0a1d[8]);
  BUFF I44 (out_0r1d[9], inp_0a1d[9]);
  BUFF I45 (out_0r1d[10], inp_0a1d[10]);
  BUFF I46 (out_0r1d[11], inp_0a1d[11]);
  BUFF I47 (out_0r1d[12], inp_0a1d[12]);
  BUFF I48 (out_0r1d[13], inp_0a1d[13]);
  BUFF I49 (out_0r1d[14], inp_0a1d[14]);
  BUFF I50 (out_0r1d[15], inp_0a1d[15]);
  BUFF I51 (out_0r1d[16], inp_0a1d[16]);
  BUFF I52 (out_0r1d[17], inp_0a1d[17]);
  BUFF I53 (out_0r1d[18], inp_0a1d[18]);
  BUFF I54 (out_0r1d[19], inp_0a1d[19]);
  BUFF I55 (out_0r1d[20], inp_0a1d[20]);
  BUFF I56 (out_0r1d[21], inp_0a1d[21]);
  BUFF I57 (out_0r1d[22], inp_0a1d[22]);
  BUFF I58 (out_0r1d[23], inp_0a1d[23]);
  BUFF I59 (out_0r1d[24], inp_0a1d[24]);
  BUFF I60 (out_0r1d[25], inp_0a1d[25]);
  BUFF I61 (out_0r1d[26], inp_0a1d[26]);
  BUFF I62 (out_0r1d[27], inp_0a1d[27]);
  BUFF I63 (out_0r1d[28], inp_0a1d[28]);
  BUFF I64 (out_0r1d[29], inp_0a1d[29]);
  BUFF I65 (out_0r1d[30], inp_0a1d[30]);
  BUFF I66 (out_0r1d[31], inp_0a1d[31]);
  BUFF I67 (out_0r1d[32], inp_0a1d[32]);
  BUFF I68 (out_0r1d[33], inp_0a1d[33]);
  BUFF I69 (activate_0a, out_0a);
endmodule

module BrzFetch_35_s5_false (
  activate_0r, activate_0a,
  inp_0r, inp_0a0d, inp_0a1d,
  out_0r0d, out_0r1d, out_0a
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input [34:0] inp_0a0d;
  input [34:0] inp_0a1d;
  output [34:0] out_0r0d;
  output [34:0] out_0r1d;
  input out_0a;
  BUFF I0 (inp_0r, activate_0r);
  BUFF I1 (out_0r0d[0], inp_0a0d[0]);
  BUFF I2 (out_0r0d[1], inp_0a0d[1]);
  BUFF I3 (out_0r0d[2], inp_0a0d[2]);
  BUFF I4 (out_0r0d[3], inp_0a0d[3]);
  BUFF I5 (out_0r0d[4], inp_0a0d[4]);
  BUFF I6 (out_0r0d[5], inp_0a0d[5]);
  BUFF I7 (out_0r0d[6], inp_0a0d[6]);
  BUFF I8 (out_0r0d[7], inp_0a0d[7]);
  BUFF I9 (out_0r0d[8], inp_0a0d[8]);
  BUFF I10 (out_0r0d[9], inp_0a0d[9]);
  BUFF I11 (out_0r0d[10], inp_0a0d[10]);
  BUFF I12 (out_0r0d[11], inp_0a0d[11]);
  BUFF I13 (out_0r0d[12], inp_0a0d[12]);
  BUFF I14 (out_0r0d[13], inp_0a0d[13]);
  BUFF I15 (out_0r0d[14], inp_0a0d[14]);
  BUFF I16 (out_0r0d[15], inp_0a0d[15]);
  BUFF I17 (out_0r0d[16], inp_0a0d[16]);
  BUFF I18 (out_0r0d[17], inp_0a0d[17]);
  BUFF I19 (out_0r0d[18], inp_0a0d[18]);
  BUFF I20 (out_0r0d[19], inp_0a0d[19]);
  BUFF I21 (out_0r0d[20], inp_0a0d[20]);
  BUFF I22 (out_0r0d[21], inp_0a0d[21]);
  BUFF I23 (out_0r0d[22], inp_0a0d[22]);
  BUFF I24 (out_0r0d[23], inp_0a0d[23]);
  BUFF I25 (out_0r0d[24], inp_0a0d[24]);
  BUFF I26 (out_0r0d[25], inp_0a0d[25]);
  BUFF I27 (out_0r0d[26], inp_0a0d[26]);
  BUFF I28 (out_0r0d[27], inp_0a0d[27]);
  BUFF I29 (out_0r0d[28], inp_0a0d[28]);
  BUFF I30 (out_0r0d[29], inp_0a0d[29]);
  BUFF I31 (out_0r0d[30], inp_0a0d[30]);
  BUFF I32 (out_0r0d[31], inp_0a0d[31]);
  BUFF I33 (out_0r0d[32], inp_0a0d[32]);
  BUFF I34 (out_0r0d[33], inp_0a0d[33]);
  BUFF I35 (out_0r0d[34], inp_0a0d[34]);
  BUFF I36 (out_0r1d[0], inp_0a1d[0]);
  BUFF I37 (out_0r1d[1], inp_0a1d[1]);
  BUFF I38 (out_0r1d[2], inp_0a1d[2]);
  BUFF I39 (out_0r1d[3], inp_0a1d[3]);
  BUFF I40 (out_0r1d[4], inp_0a1d[4]);
  BUFF I41 (out_0r1d[5], inp_0a1d[5]);
  BUFF I42 (out_0r1d[6], inp_0a1d[6]);
  BUFF I43 (out_0r1d[7], inp_0a1d[7]);
  BUFF I44 (out_0r1d[8], inp_0a1d[8]);
  BUFF I45 (out_0r1d[9], inp_0a1d[9]);
  BUFF I46 (out_0r1d[10], inp_0a1d[10]);
  BUFF I47 (out_0r1d[11], inp_0a1d[11]);
  BUFF I48 (out_0r1d[12], inp_0a1d[12]);
  BUFF I49 (out_0r1d[13], inp_0a1d[13]);
  BUFF I50 (out_0r1d[14], inp_0a1d[14]);
  BUFF I51 (out_0r1d[15], inp_0a1d[15]);
  BUFF I52 (out_0r1d[16], inp_0a1d[16]);
  BUFF I53 (out_0r1d[17], inp_0a1d[17]);
  BUFF I54 (out_0r1d[18], inp_0a1d[18]);
  BUFF I55 (out_0r1d[19], inp_0a1d[19]);
  BUFF I56 (out_0r1d[20], inp_0a1d[20]);
  BUFF I57 (out_0r1d[21], inp_0a1d[21]);
  BUFF I58 (out_0r1d[22], inp_0a1d[22]);
  BUFF I59 (out_0r1d[23], inp_0a1d[23]);
  BUFF I60 (out_0r1d[24], inp_0a1d[24]);
  BUFF I61 (out_0r1d[25], inp_0a1d[25]);
  BUFF I62 (out_0r1d[26], inp_0a1d[26]);
  BUFF I63 (out_0r1d[27], inp_0a1d[27]);
  BUFF I64 (out_0r1d[28], inp_0a1d[28]);
  BUFF I65 (out_0r1d[29], inp_0a1d[29]);
  BUFF I66 (out_0r1d[30], inp_0a1d[30]);
  BUFF I67 (out_0r1d[31], inp_0a1d[31]);
  BUFF I68 (out_0r1d[32], inp_0a1d[32]);
  BUFF I69 (out_0r1d[33], inp_0a1d[33]);
  BUFF I70 (out_0r1d[34], inp_0a1d[34]);
  BUFF I71 (activate_0a, out_0a);
endmodule

module BrzFetch_35_s4_true (
  activate_0r, activate_0a,
  inp_0r, inp_0a0d, inp_0a1d,
  out_0r0d, out_0r1d, out_0a
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input [34:0] inp_0a0d;
  input [34:0] inp_0a1d;
  output [34:0] out_0r0d;
  output [34:0] out_0r1d;
  input out_0a;
  BUFF I0 (inp_0r, activate_0r);
  BUFF I1 (out_0r0d[0], inp_0a0d[0]);
  BUFF I2 (out_0r0d[1], inp_0a0d[1]);
  BUFF I3 (out_0r0d[2], inp_0a0d[2]);
  BUFF I4 (out_0r0d[3], inp_0a0d[3]);
  BUFF I5 (out_0r0d[4], inp_0a0d[4]);
  BUFF I6 (out_0r0d[5], inp_0a0d[5]);
  BUFF I7 (out_0r0d[6], inp_0a0d[6]);
  BUFF I8 (out_0r0d[7], inp_0a0d[7]);
  BUFF I9 (out_0r0d[8], inp_0a0d[8]);
  BUFF I10 (out_0r0d[9], inp_0a0d[9]);
  BUFF I11 (out_0r0d[10], inp_0a0d[10]);
  BUFF I12 (out_0r0d[11], inp_0a0d[11]);
  BUFF I13 (out_0r0d[12], inp_0a0d[12]);
  BUFF I14 (out_0r0d[13], inp_0a0d[13]);
  BUFF I15 (out_0r0d[14], inp_0a0d[14]);
  BUFF I16 (out_0r0d[15], inp_0a0d[15]);
  BUFF I17 (out_0r0d[16], inp_0a0d[16]);
  BUFF I18 (out_0r0d[17], inp_0a0d[17]);
  BUFF I19 (out_0r0d[18], inp_0a0d[18]);
  BUFF I20 (out_0r0d[19], inp_0a0d[19]);
  BUFF I21 (out_0r0d[20], inp_0a0d[20]);
  BUFF I22 (out_0r0d[21], inp_0a0d[21]);
  BUFF I23 (out_0r0d[22], inp_0a0d[22]);
  BUFF I24 (out_0r0d[23], inp_0a0d[23]);
  BUFF I25 (out_0r0d[24], inp_0a0d[24]);
  BUFF I26 (out_0r0d[25], inp_0a0d[25]);
  BUFF I27 (out_0r0d[26], inp_0a0d[26]);
  BUFF I28 (out_0r0d[27], inp_0a0d[27]);
  BUFF I29 (out_0r0d[28], inp_0a0d[28]);
  BUFF I30 (out_0r0d[29], inp_0a0d[29]);
  BUFF I31 (out_0r0d[30], inp_0a0d[30]);
  BUFF I32 (out_0r0d[31], inp_0a0d[31]);
  BUFF I33 (out_0r0d[32], inp_0a0d[32]);
  BUFF I34 (out_0r0d[33], inp_0a0d[33]);
  BUFF I35 (out_0r0d[34], inp_0a0d[34]);
  BUFF I36 (out_0r1d[0], inp_0a1d[0]);
  BUFF I37 (out_0r1d[1], inp_0a1d[1]);
  BUFF I38 (out_0r1d[2], inp_0a1d[2]);
  BUFF I39 (out_0r1d[3], inp_0a1d[3]);
  BUFF I40 (out_0r1d[4], inp_0a1d[4]);
  BUFF I41 (out_0r1d[5], inp_0a1d[5]);
  BUFF I42 (out_0r1d[6], inp_0a1d[6]);
  BUFF I43 (out_0r1d[7], inp_0a1d[7]);
  BUFF I44 (out_0r1d[8], inp_0a1d[8]);
  BUFF I45 (out_0r1d[9], inp_0a1d[9]);
  BUFF I46 (out_0r1d[10], inp_0a1d[10]);
  BUFF I47 (out_0r1d[11], inp_0a1d[11]);
  BUFF I48 (out_0r1d[12], inp_0a1d[12]);
  BUFF I49 (out_0r1d[13], inp_0a1d[13]);
  BUFF I50 (out_0r1d[14], inp_0a1d[14]);
  BUFF I51 (out_0r1d[15], inp_0a1d[15]);
  BUFF I52 (out_0r1d[16], inp_0a1d[16]);
  BUFF I53 (out_0r1d[17], inp_0a1d[17]);
  BUFF I54 (out_0r1d[18], inp_0a1d[18]);
  BUFF I55 (out_0r1d[19], inp_0a1d[19]);
  BUFF I56 (out_0r1d[20], inp_0a1d[20]);
  BUFF I57 (out_0r1d[21], inp_0a1d[21]);
  BUFF I58 (out_0r1d[22], inp_0a1d[22]);
  BUFF I59 (out_0r1d[23], inp_0a1d[23]);
  BUFF I60 (out_0r1d[24], inp_0a1d[24]);
  BUFF I61 (out_0r1d[25], inp_0a1d[25]);
  BUFF I62 (out_0r1d[26], inp_0a1d[26]);
  BUFF I63 (out_0r1d[27], inp_0a1d[27]);
  BUFF I64 (out_0r1d[28], inp_0a1d[28]);
  BUFF I65 (out_0r1d[29], inp_0a1d[29]);
  BUFF I66 (out_0r1d[30], inp_0a1d[30]);
  BUFF I67 (out_0r1d[31], inp_0a1d[31]);
  BUFF I68 (out_0r1d[32], inp_0a1d[32]);
  BUFF I69 (out_0r1d[33], inp_0a1d[33]);
  BUFF I70 (out_0r1d[34], inp_0a1d[34]);
  BUFF I71 (activate_0a, out_0a);
endmodule

module BrzFetch_36_s5_false (
  activate_0r, activate_0a,
  inp_0r, inp_0a0d, inp_0a1d,
  out_0r0d, out_0r1d, out_0a
);
  input activate_0r;
  output activate_0a;
  output inp_0r;
  input [35:0] inp_0a0d;
  input [35:0] inp_0a1d;
  output [35:0] out_0r0d;
  output [35:0] out_0r1d;
  input out_0a;
  BUFF I0 (inp_0r, activate_0r);
  BUFF I1 (out_0r0d[0], inp_0a0d[0]);
  BUFF I2 (out_0r0d[1], inp_0a0d[1]);
  BUFF I3 (out_0r0d[2], inp_0a0d[2]);
  BUFF I4 (out_0r0d[3], inp_0a0d[3]);
  BUFF I5 (out_0r0d[4], inp_0a0d[4]);
  BUFF I6 (out_0r0d[5], inp_0a0d[5]);
  BUFF I7 (out_0r0d[6], inp_0a0d[6]);
  BUFF I8 (out_0r0d[7], inp_0a0d[7]);
  BUFF I9 (out_0r0d[8], inp_0a0d[8]);
  BUFF I10 (out_0r0d[9], inp_0a0d[9]);
  BUFF I11 (out_0r0d[10], inp_0a0d[10]);
  BUFF I12 (out_0r0d[11], inp_0a0d[11]);
  BUFF I13 (out_0r0d[12], inp_0a0d[12]);
  BUFF I14 (out_0r0d[13], inp_0a0d[13]);
  BUFF I15 (out_0r0d[14], inp_0a0d[14]);
  BUFF I16 (out_0r0d[15], inp_0a0d[15]);
  BUFF I17 (out_0r0d[16], inp_0a0d[16]);
  BUFF I18 (out_0r0d[17], inp_0a0d[17]);
  BUFF I19 (out_0r0d[18], inp_0a0d[18]);
  BUFF I20 (out_0r0d[19], inp_0a0d[19]);
  BUFF I21 (out_0r0d[20], inp_0a0d[20]);
  BUFF I22 (out_0r0d[21], inp_0a0d[21]);
  BUFF I23 (out_0r0d[22], inp_0a0d[22]);
  BUFF I24 (out_0r0d[23], inp_0a0d[23]);
  BUFF I25 (out_0r0d[24], inp_0a0d[24]);
  BUFF I26 (out_0r0d[25], inp_0a0d[25]);
  BUFF I27 (out_0r0d[26], inp_0a0d[26]);
  BUFF I28 (out_0r0d[27], inp_0a0d[27]);
  BUFF I29 (out_0r0d[28], inp_0a0d[28]);
  BUFF I30 (out_0r0d[29], inp_0a0d[29]);
  BUFF I31 (out_0r0d[30], inp_0a0d[30]);
  BUFF I32 (out_0r0d[31], inp_0a0d[31]);
  BUFF I33 (out_0r0d[32], inp_0a0d[32]);
  BUFF I34 (out_0r0d[33], inp_0a0d[33]);
  BUFF I35 (out_0r0d[34], inp_0a0d[34]);
  BUFF I36 (out_0r0d[35], inp_0a0d[35]);
  BUFF I37 (out_0r1d[0], inp_0a1d[0]);
  BUFF I38 (out_0r1d[1], inp_0a1d[1]);
  BUFF I39 (out_0r1d[2], inp_0a1d[2]);
  BUFF I40 (out_0r1d[3], inp_0a1d[3]);
  BUFF I41 (out_0r1d[4], inp_0a1d[4]);
  BUFF I42 (out_0r1d[5], inp_0a1d[5]);
  BUFF I43 (out_0r1d[6], inp_0a1d[6]);
  BUFF I44 (out_0r1d[7], inp_0a1d[7]);
  BUFF I45 (out_0r1d[8], inp_0a1d[8]);
  BUFF I46 (out_0r1d[9], inp_0a1d[9]);
  BUFF I47 (out_0r1d[10], inp_0a1d[10]);
  BUFF I48 (out_0r1d[11], inp_0a1d[11]);
  BUFF I49 (out_0r1d[12], inp_0a1d[12]);
  BUFF I50 (out_0r1d[13], inp_0a1d[13]);
  BUFF I51 (out_0r1d[14], inp_0a1d[14]);
  BUFF I52 (out_0r1d[15], inp_0a1d[15]);
  BUFF I53 (out_0r1d[16], inp_0a1d[16]);
  BUFF I54 (out_0r1d[17], inp_0a1d[17]);
  BUFF I55 (out_0r1d[18], inp_0a1d[18]);
  BUFF I56 (out_0r1d[19], inp_0a1d[19]);
  BUFF I57 (out_0r1d[20], inp_0a1d[20]);
  BUFF I58 (out_0r1d[21], inp_0a1d[21]);
  BUFF I59 (out_0r1d[22], inp_0a1d[22]);
  BUFF I60 (out_0r1d[23], inp_0a1d[23]);
  BUFF I61 (out_0r1d[24], inp_0a1d[24]);
  BUFF I62 (out_0r1d[25], inp_0a1d[25]);
  BUFF I63 (out_0r1d[26], inp_0a1d[26]);
  BUFF I64 (out_0r1d[27], inp_0a1d[27]);
  BUFF I65 (out_0r1d[28], inp_0a1d[28]);
  BUFF I66 (out_0r1d[29], inp_0a1d[29]);
  BUFF I67 (out_0r1d[30], inp_0a1d[30]);
  BUFF I68 (out_0r1d[31], inp_0a1d[31]);
  BUFF I69 (out_0r1d[32], inp_0a1d[32]);
  BUFF I70 (out_0r1d[33], inp_0a1d[33]);
  BUFF I71 (out_0r1d[34], inp_0a1d[34]);
  BUFF I72 (out_0r1d[35], inp_0a1d[35]);
  BUFF I73 (activate_0a, out_0a);
endmodule

module BrzFork_2 (
  inp_0r, inp_0a,
  out_0r, out_0a,
  out_1r, out_1a
);
  input inp_0r;
  output inp_0a;
  output out_0r;
  input out_0a;
  output out_1r;
  input out_1a;
  C2 I0 (inp_0a, out_0a, out_1a);
  BUFF I1 (out_0r, inp_0r);
  BUFF I2 (out_1r, inp_0r);
endmodule

module BrzFork_3 (
  inp_0r, inp_0a,
  out_0r, out_0a,
  out_1r, out_1a,
  out_2r, out_2a
);
  input inp_0r;
  output inp_0a;
  output out_0r;
  input out_0a;
  output out_1r;
  input out_1a;
  output out_2r;
  input out_2a;
  C3 I0 (inp_0a, out_0a, out_1a, out_2a);
  BUFF I1 (out_0r, inp_0r);
  BUFF I2 (out_1r, inp_0r);
  BUFF I3 (out_2r, inp_0r);
endmodule

module BrzFork_4 (
  inp_0r, inp_0a,
  out_0r, out_0a,
  out_1r, out_1a,
  out_2r, out_2a,
  out_3r, out_3a
);
  input inp_0r;
  output inp_0a;
  output out_0r;
  input out_0a;
  output out_1r;
  input out_1a;
  output out_2r;
  input out_2a;
  output out_3r;
  input out_3a;
  wire [1:0] internal_0n;
  C2 I0 (internal_0n[0], out_0a, out_1a);
  C2 I1 (internal_0n[1], out_2a, out_3a);
  C2 I2 (inp_0a, internal_0n[0], internal_0n[1]);
  BUFF I3 (out_0r, inp_0r);
  BUFF I4 (out_1r, inp_0r);
  BUFF I5 (out_2r, inp_0r);
  BUFF I6 (out_3r, inp_0r);
endmodule

module BrzFork_5 (
  inp_0r, inp_0a,
  out_0r, out_0a,
  out_1r, out_1a,
  out_2r, out_2a,
  out_3r, out_3a,
  out_4r, out_4a
);
  input inp_0r;
  output inp_0a;
  output out_0r;
  input out_0a;
  output out_1r;
  input out_1a;
  output out_2r;
  input out_2a;
  output out_3r;
  input out_3a;
  output out_4r;
  input out_4a;
  wire [1:0] internal_0n;
  C3 I0 (internal_0n[0], out_0a, out_1a, out_2a);
  C2 I1 (internal_0n[1], out_3a, out_4a);
  C2 I2 (inp_0a, internal_0n[0], internal_0n[1]);
  BUFF I3 (out_0r, inp_0r);
  BUFF I4 (out_1r, inp_0r);
  BUFF I5 (out_2r, inp_0r);
  BUFF I6 (out_3r, inp_0r);
  BUFF I7 (out_4r, inp_0r);
endmodule

module BrzLoop (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  wire nReq_0n;
  supply0 gnd;
  INV I0 (nReq_0n, activate_0r);
  NOR2 I1 (activateOut_0r, nReq_0n, activateOut_0a);
  BUFF I2 (activate_0a, gnd);
endmodule

module BrzPassivatorPush_1_1 (
  out_0r, out_0a0d, out_0a1d,
  inp_0r0d, inp_0r1d, inp_0a
);
  input out_0r;
  output out_0a0d;
  output out_0a1d;
  input inp_0r0d;
  input inp_0r1d;
  output inp_0a;
  wire poutReq_0n;
  wire poutReqB_0n;
  wire outComplete_0n;
  wire outData_0n;
  wire outData_1n;
  BUFF I0 (inp_0a, outComplete_0n);
  OR2 I1 (outComplete_0n, outData_0n, outData_1n);
  C2 I2 (outData_1n, inp_0r1d, poutReqB_0n);
  C2 I3 (outData_0n, inp_0r0d, poutReqB_0n);
  BUFF I4 (poutReq_0n, out_0r);
  BUFF I5 (poutReqB_0n, poutReq_0n);
  BUFF I6 (out_0a1d, outData_1n);
  BUFF I7 (out_0a0d, outData_0n);
endmodule

module BrzPassivatorPush_3_1 (
  out_0r, out_0a0d, out_0a1d,
  inp_0r0d, inp_0r1d, inp_0a
);
  input out_0r;
  output [2:0] out_0a0d;
  output [2:0] out_0a1d;
  input [2:0] inp_0r0d;
  input [2:0] inp_0r1d;
  output inp_0a;
  wire poutReq_0n;
  wire poutReqB_0n;
  wire [2:0] outComplete_0n;
  wire [2:0] outData_0n;
  wire [2:0] outData_1n;
  C3 I0 (inp_0a, outComplete_0n[0], outComplete_0n[1], outComplete_0n[2]);
  OR2 I1 (outComplete_0n[0], outData_0n[0], outData_1n[0]);
  OR2 I2 (outComplete_0n[1], outData_0n[1], outData_1n[1]);
  OR2 I3 (outComplete_0n[2], outData_0n[2], outData_1n[2]);
  C2 I4 (outData_1n[0], inp_0r1d[0], poutReqB_0n);
  C2 I5 (outData_1n[1], inp_0r1d[1], poutReqB_0n);
  C2 I6 (outData_1n[2], inp_0r1d[2], poutReqB_0n);
  C2 I7 (outData_0n[0], inp_0r0d[0], poutReqB_0n);
  C2 I8 (outData_0n[1], inp_0r0d[1], poutReqB_0n);
  C2 I9 (outData_0n[2], inp_0r0d[2], poutReqB_0n);
  BUFF I10 (poutReq_0n, out_0r);
  BUFF I11 (poutReqB_0n, poutReq_0n);
  BUFF I12 (out_0a1d[0], outData_1n[0]);
  BUFF I13 (out_0a1d[1], outData_1n[1]);
  BUFF I14 (out_0a1d[2], outData_1n[2]);
  BUFF I15 (out_0a0d[0], outData_0n[0]);
  BUFF I16 (out_0a0d[1], outData_0n[1]);
  BUFF I17 (out_0a0d[2], outData_0n[2]);
endmodule

module BrzPassivatorPush_32_1 (
  out_0r, out_0a0d, out_0a1d,
  inp_0r0d, inp_0r1d, inp_0a
);
  input out_0r;
  output [31:0] out_0a0d;
  output [31:0] out_0a1d;
  input [31:0] inp_0r0d;
  input [31:0] inp_0r1d;
  output inp_0a;
  wire [16:0] internal_0n;
  wire poutReq_0n;
  wire poutReqB_0n;
  wire [31:0] outComplete_0n;
  wire [31:0] outData_0n;
  wire [31:0] outData_1n;
  C3 I0 (internal_0n[0], outComplete_0n[0], outComplete_0n[1], outComplete_0n[2]);
  C3 I1 (internal_0n[1], outComplete_0n[3], outComplete_0n[4], outComplete_0n[5]);
  C3 I2 (internal_0n[2], outComplete_0n[6], outComplete_0n[7], outComplete_0n[8]);
  C3 I3 (internal_0n[3], outComplete_0n[9], outComplete_0n[10], outComplete_0n[11]);
  C3 I4 (internal_0n[4], outComplete_0n[12], outComplete_0n[13], outComplete_0n[14]);
  C3 I5 (internal_0n[5], outComplete_0n[15], outComplete_0n[16], outComplete_0n[17]);
  C3 I6 (internal_0n[6], outComplete_0n[18], outComplete_0n[19], outComplete_0n[20]);
  C3 I7 (internal_0n[7], outComplete_0n[21], outComplete_0n[22], outComplete_0n[23]);
  C3 I8 (internal_0n[8], outComplete_0n[24], outComplete_0n[25], outComplete_0n[26]);
  C3 I9 (internal_0n[9], outComplete_0n[27], outComplete_0n[28], outComplete_0n[29]);
  C2 I10 (internal_0n[10], outComplete_0n[30], outComplete_0n[31]);
  C3 I11 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I12 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I13 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I14 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I15 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I16 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I17 (inp_0a, internal_0n[15], internal_0n[16]);
  OR2 I18 (outComplete_0n[0], outData_0n[0], outData_1n[0]);
  OR2 I19 (outComplete_0n[1], outData_0n[1], outData_1n[1]);
  OR2 I20 (outComplete_0n[2], outData_0n[2], outData_1n[2]);
  OR2 I21 (outComplete_0n[3], outData_0n[3], outData_1n[3]);
  OR2 I22 (outComplete_0n[4], outData_0n[4], outData_1n[4]);
  OR2 I23 (outComplete_0n[5], outData_0n[5], outData_1n[5]);
  OR2 I24 (outComplete_0n[6], outData_0n[6], outData_1n[6]);
  OR2 I25 (outComplete_0n[7], outData_0n[7], outData_1n[7]);
  OR2 I26 (outComplete_0n[8], outData_0n[8], outData_1n[8]);
  OR2 I27 (outComplete_0n[9], outData_0n[9], outData_1n[9]);
  OR2 I28 (outComplete_0n[10], outData_0n[10], outData_1n[10]);
  OR2 I29 (outComplete_0n[11], outData_0n[11], outData_1n[11]);
  OR2 I30 (outComplete_0n[12], outData_0n[12], outData_1n[12]);
  OR2 I31 (outComplete_0n[13], outData_0n[13], outData_1n[13]);
  OR2 I32 (outComplete_0n[14], outData_0n[14], outData_1n[14]);
  OR2 I33 (outComplete_0n[15], outData_0n[15], outData_1n[15]);
  OR2 I34 (outComplete_0n[16], outData_0n[16], outData_1n[16]);
  OR2 I35 (outComplete_0n[17], outData_0n[17], outData_1n[17]);
  OR2 I36 (outComplete_0n[18], outData_0n[18], outData_1n[18]);
  OR2 I37 (outComplete_0n[19], outData_0n[19], outData_1n[19]);
  OR2 I38 (outComplete_0n[20], outData_0n[20], outData_1n[20]);
  OR2 I39 (outComplete_0n[21], outData_0n[21], outData_1n[21]);
  OR2 I40 (outComplete_0n[22], outData_0n[22], outData_1n[22]);
  OR2 I41 (outComplete_0n[23], outData_0n[23], outData_1n[23]);
  OR2 I42 (outComplete_0n[24], outData_0n[24], outData_1n[24]);
  OR2 I43 (outComplete_0n[25], outData_0n[25], outData_1n[25]);
  OR2 I44 (outComplete_0n[26], outData_0n[26], outData_1n[26]);
  OR2 I45 (outComplete_0n[27], outData_0n[27], outData_1n[27]);
  OR2 I46 (outComplete_0n[28], outData_0n[28], outData_1n[28]);
  OR2 I47 (outComplete_0n[29], outData_0n[29], outData_1n[29]);
  OR2 I48 (outComplete_0n[30], outData_0n[30], outData_1n[30]);
  OR2 I49 (outComplete_0n[31], outData_0n[31], outData_1n[31]);
  C2 I50 (outData_1n[0], inp_0r1d[0], poutReqB_0n);
  C2 I51 (outData_1n[1], inp_0r1d[1], poutReqB_0n);
  C2 I52 (outData_1n[2], inp_0r1d[2], poutReqB_0n);
  C2 I53 (outData_1n[3], inp_0r1d[3], poutReqB_0n);
  C2 I54 (outData_1n[4], inp_0r1d[4], poutReqB_0n);
  C2 I55 (outData_1n[5], inp_0r1d[5], poutReqB_0n);
  C2 I56 (outData_1n[6], inp_0r1d[6], poutReqB_0n);
  C2 I57 (outData_1n[7], inp_0r1d[7], poutReqB_0n);
  C2 I58 (outData_1n[8], inp_0r1d[8], poutReqB_0n);
  C2 I59 (outData_1n[9], inp_0r1d[9], poutReqB_0n);
  C2 I60 (outData_1n[10], inp_0r1d[10], poutReqB_0n);
  C2 I61 (outData_1n[11], inp_0r1d[11], poutReqB_0n);
  C2 I62 (outData_1n[12], inp_0r1d[12], poutReqB_0n);
  C2 I63 (outData_1n[13], inp_0r1d[13], poutReqB_0n);
  C2 I64 (outData_1n[14], inp_0r1d[14], poutReqB_0n);
  C2 I65 (outData_1n[15], inp_0r1d[15], poutReqB_0n);
  C2 I66 (outData_1n[16], inp_0r1d[16], poutReqB_0n);
  C2 I67 (outData_1n[17], inp_0r1d[17], poutReqB_0n);
  C2 I68 (outData_1n[18], inp_0r1d[18], poutReqB_0n);
  C2 I69 (outData_1n[19], inp_0r1d[19], poutReqB_0n);
  C2 I70 (outData_1n[20], inp_0r1d[20], poutReqB_0n);
  C2 I71 (outData_1n[21], inp_0r1d[21], poutReqB_0n);
  C2 I72 (outData_1n[22], inp_0r1d[22], poutReqB_0n);
  C2 I73 (outData_1n[23], inp_0r1d[23], poutReqB_0n);
  C2 I74 (outData_1n[24], inp_0r1d[24], poutReqB_0n);
  C2 I75 (outData_1n[25], inp_0r1d[25], poutReqB_0n);
  C2 I76 (outData_1n[26], inp_0r1d[26], poutReqB_0n);
  C2 I77 (outData_1n[27], inp_0r1d[27], poutReqB_0n);
  C2 I78 (outData_1n[28], inp_0r1d[28], poutReqB_0n);
  C2 I79 (outData_1n[29], inp_0r1d[29], poutReqB_0n);
  C2 I80 (outData_1n[30], inp_0r1d[30], poutReqB_0n);
  C2 I81 (outData_1n[31], inp_0r1d[31], poutReqB_0n);
  C2 I82 (outData_0n[0], inp_0r0d[0], poutReqB_0n);
  C2 I83 (outData_0n[1], inp_0r0d[1], poutReqB_0n);
  C2 I84 (outData_0n[2], inp_0r0d[2], poutReqB_0n);
  C2 I85 (outData_0n[3], inp_0r0d[3], poutReqB_0n);
  C2 I86 (outData_0n[4], inp_0r0d[4], poutReqB_0n);
  C2 I87 (outData_0n[5], inp_0r0d[5], poutReqB_0n);
  C2 I88 (outData_0n[6], inp_0r0d[6], poutReqB_0n);
  C2 I89 (outData_0n[7], inp_0r0d[7], poutReqB_0n);
  C2 I90 (outData_0n[8], inp_0r0d[8], poutReqB_0n);
  C2 I91 (outData_0n[9], inp_0r0d[9], poutReqB_0n);
  C2 I92 (outData_0n[10], inp_0r0d[10], poutReqB_0n);
  C2 I93 (outData_0n[11], inp_0r0d[11], poutReqB_0n);
  C2 I94 (outData_0n[12], inp_0r0d[12], poutReqB_0n);
  C2 I95 (outData_0n[13], inp_0r0d[13], poutReqB_0n);
  C2 I96 (outData_0n[14], inp_0r0d[14], poutReqB_0n);
  C2 I97 (outData_0n[15], inp_0r0d[15], poutReqB_0n);
  C2 I98 (outData_0n[16], inp_0r0d[16], poutReqB_0n);
  C2 I99 (outData_0n[17], inp_0r0d[17], poutReqB_0n);
  C2 I100 (outData_0n[18], inp_0r0d[18], poutReqB_0n);
  C2 I101 (outData_0n[19], inp_0r0d[19], poutReqB_0n);
  C2 I102 (outData_0n[20], inp_0r0d[20], poutReqB_0n);
  C2 I103 (outData_0n[21], inp_0r0d[21], poutReqB_0n);
  C2 I104 (outData_0n[22], inp_0r0d[22], poutReqB_0n);
  C2 I105 (outData_0n[23], inp_0r0d[23], poutReqB_0n);
  C2 I106 (outData_0n[24], inp_0r0d[24], poutReqB_0n);
  C2 I107 (outData_0n[25], inp_0r0d[25], poutReqB_0n);
  C2 I108 (outData_0n[26], inp_0r0d[26], poutReqB_0n);
  C2 I109 (outData_0n[27], inp_0r0d[27], poutReqB_0n);
  C2 I110 (outData_0n[28], inp_0r0d[28], poutReqB_0n);
  C2 I111 (outData_0n[29], inp_0r0d[29], poutReqB_0n);
  C2 I112 (outData_0n[30], inp_0r0d[30], poutReqB_0n);
  C2 I113 (outData_0n[31], inp_0r0d[31], poutReqB_0n);
  BUFF I114 (poutReq_0n, out_0r);
  BUFF I115 (poutReqB_0n, poutReq_0n);
  BUFF I116 (out_0a1d[0], outData_1n[0]);
  BUFF I117 (out_0a1d[1], outData_1n[1]);
  BUFF I118 (out_0a1d[2], outData_1n[2]);
  BUFF I119 (out_0a1d[3], outData_1n[3]);
  BUFF I120 (out_0a1d[4], outData_1n[4]);
  BUFF I121 (out_0a1d[5], outData_1n[5]);
  BUFF I122 (out_0a1d[6], outData_1n[6]);
  BUFF I123 (out_0a1d[7], outData_1n[7]);
  BUFF I124 (out_0a1d[8], outData_1n[8]);
  BUFF I125 (out_0a1d[9], outData_1n[9]);
  BUFF I126 (out_0a1d[10], outData_1n[10]);
  BUFF I127 (out_0a1d[11], outData_1n[11]);
  BUFF I128 (out_0a1d[12], outData_1n[12]);
  BUFF I129 (out_0a1d[13], outData_1n[13]);
  BUFF I130 (out_0a1d[14], outData_1n[14]);
  BUFF I131 (out_0a1d[15], outData_1n[15]);
  BUFF I132 (out_0a1d[16], outData_1n[16]);
  BUFF I133 (out_0a1d[17], outData_1n[17]);
  BUFF I134 (out_0a1d[18], outData_1n[18]);
  BUFF I135 (out_0a1d[19], outData_1n[19]);
  BUFF I136 (out_0a1d[20], outData_1n[20]);
  BUFF I137 (out_0a1d[21], outData_1n[21]);
  BUFF I138 (out_0a1d[22], outData_1n[22]);
  BUFF I139 (out_0a1d[23], outData_1n[23]);
  BUFF I140 (out_0a1d[24], outData_1n[24]);
  BUFF I141 (out_0a1d[25], outData_1n[25]);
  BUFF I142 (out_0a1d[26], outData_1n[26]);
  BUFF I143 (out_0a1d[27], outData_1n[27]);
  BUFF I144 (out_0a1d[28], outData_1n[28]);
  BUFF I145 (out_0a1d[29], outData_1n[29]);
  BUFF I146 (out_0a1d[30], outData_1n[30]);
  BUFF I147 (out_0a1d[31], outData_1n[31]);
  BUFF I148 (out_0a0d[0], outData_0n[0]);
  BUFF I149 (out_0a0d[1], outData_0n[1]);
  BUFF I150 (out_0a0d[2], outData_0n[2]);
  BUFF I151 (out_0a0d[3], outData_0n[3]);
  BUFF I152 (out_0a0d[4], outData_0n[4]);
  BUFF I153 (out_0a0d[5], outData_0n[5]);
  BUFF I154 (out_0a0d[6], outData_0n[6]);
  BUFF I155 (out_0a0d[7], outData_0n[7]);
  BUFF I156 (out_0a0d[8], outData_0n[8]);
  BUFF I157 (out_0a0d[9], outData_0n[9]);
  BUFF I158 (out_0a0d[10], outData_0n[10]);
  BUFF I159 (out_0a0d[11], outData_0n[11]);
  BUFF I160 (out_0a0d[12], outData_0n[12]);
  BUFF I161 (out_0a0d[13], outData_0n[13]);
  BUFF I162 (out_0a0d[14], outData_0n[14]);
  BUFF I163 (out_0a0d[15], outData_0n[15]);
  BUFF I164 (out_0a0d[16], outData_0n[16]);
  BUFF I165 (out_0a0d[17], outData_0n[17]);
  BUFF I166 (out_0a0d[18], outData_0n[18]);
  BUFF I167 (out_0a0d[19], outData_0n[19]);
  BUFF I168 (out_0a0d[20], outData_0n[20]);
  BUFF I169 (out_0a0d[21], outData_0n[21]);
  BUFF I170 (out_0a0d[22], outData_0n[22]);
  BUFF I171 (out_0a0d[23], outData_0n[23]);
  BUFF I172 (out_0a0d[24], outData_0n[24]);
  BUFF I173 (out_0a0d[25], outData_0n[25]);
  BUFF I174 (out_0a0d[26], outData_0n[26]);
  BUFF I175 (out_0a0d[27], outData_0n[27]);
  BUFF I176 (out_0a0d[28], outData_0n[28]);
  BUFF I177 (out_0a0d[29], outData_0n[29]);
  BUFF I178 (out_0a0d[30], outData_0n[30]);
  BUFF I179 (out_0a0d[31], outData_0n[31]);
endmodule

module BrzPassivatorPush_33_1 (
  out_0r, out_0a0d, out_0a1d,
  inp_0r0d, inp_0r1d, inp_0a
);
  input out_0r;
  output [32:0] out_0a0d;
  output [32:0] out_0a1d;
  input [32:0] inp_0r0d;
  input [32:0] inp_0r1d;
  output inp_0a;
  wire [16:0] internal_0n;
  wire poutReq_0n;
  wire poutReqB_0n;
  wire [32:0] outComplete_0n;
  wire [32:0] outData_0n;
  wire [32:0] outData_1n;
  C3 I0 (internal_0n[0], outComplete_0n[0], outComplete_0n[1], outComplete_0n[2]);
  C3 I1 (internal_0n[1], outComplete_0n[3], outComplete_0n[4], outComplete_0n[5]);
  C3 I2 (internal_0n[2], outComplete_0n[6], outComplete_0n[7], outComplete_0n[8]);
  C3 I3 (internal_0n[3], outComplete_0n[9], outComplete_0n[10], outComplete_0n[11]);
  C3 I4 (internal_0n[4], outComplete_0n[12], outComplete_0n[13], outComplete_0n[14]);
  C3 I5 (internal_0n[5], outComplete_0n[15], outComplete_0n[16], outComplete_0n[17]);
  C3 I6 (internal_0n[6], outComplete_0n[18], outComplete_0n[19], outComplete_0n[20]);
  C3 I7 (internal_0n[7], outComplete_0n[21], outComplete_0n[22], outComplete_0n[23]);
  C3 I8 (internal_0n[8], outComplete_0n[24], outComplete_0n[25], outComplete_0n[26]);
  C3 I9 (internal_0n[9], outComplete_0n[27], outComplete_0n[28], outComplete_0n[29]);
  C3 I10 (internal_0n[10], outComplete_0n[30], outComplete_0n[31], outComplete_0n[32]);
  C3 I11 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I12 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I13 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I14 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I15 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I16 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I17 (inp_0a, internal_0n[15], internal_0n[16]);
  OR2 I18 (outComplete_0n[0], outData_0n[0], outData_1n[0]);
  OR2 I19 (outComplete_0n[1], outData_0n[1], outData_1n[1]);
  OR2 I20 (outComplete_0n[2], outData_0n[2], outData_1n[2]);
  OR2 I21 (outComplete_0n[3], outData_0n[3], outData_1n[3]);
  OR2 I22 (outComplete_0n[4], outData_0n[4], outData_1n[4]);
  OR2 I23 (outComplete_0n[5], outData_0n[5], outData_1n[5]);
  OR2 I24 (outComplete_0n[6], outData_0n[6], outData_1n[6]);
  OR2 I25 (outComplete_0n[7], outData_0n[7], outData_1n[7]);
  OR2 I26 (outComplete_0n[8], outData_0n[8], outData_1n[8]);
  OR2 I27 (outComplete_0n[9], outData_0n[9], outData_1n[9]);
  OR2 I28 (outComplete_0n[10], outData_0n[10], outData_1n[10]);
  OR2 I29 (outComplete_0n[11], outData_0n[11], outData_1n[11]);
  OR2 I30 (outComplete_0n[12], outData_0n[12], outData_1n[12]);
  OR2 I31 (outComplete_0n[13], outData_0n[13], outData_1n[13]);
  OR2 I32 (outComplete_0n[14], outData_0n[14], outData_1n[14]);
  OR2 I33 (outComplete_0n[15], outData_0n[15], outData_1n[15]);
  OR2 I34 (outComplete_0n[16], outData_0n[16], outData_1n[16]);
  OR2 I35 (outComplete_0n[17], outData_0n[17], outData_1n[17]);
  OR2 I36 (outComplete_0n[18], outData_0n[18], outData_1n[18]);
  OR2 I37 (outComplete_0n[19], outData_0n[19], outData_1n[19]);
  OR2 I38 (outComplete_0n[20], outData_0n[20], outData_1n[20]);
  OR2 I39 (outComplete_0n[21], outData_0n[21], outData_1n[21]);
  OR2 I40 (outComplete_0n[22], outData_0n[22], outData_1n[22]);
  OR2 I41 (outComplete_0n[23], outData_0n[23], outData_1n[23]);
  OR2 I42 (outComplete_0n[24], outData_0n[24], outData_1n[24]);
  OR2 I43 (outComplete_0n[25], outData_0n[25], outData_1n[25]);
  OR2 I44 (outComplete_0n[26], outData_0n[26], outData_1n[26]);
  OR2 I45 (outComplete_0n[27], outData_0n[27], outData_1n[27]);
  OR2 I46 (outComplete_0n[28], outData_0n[28], outData_1n[28]);
  OR2 I47 (outComplete_0n[29], outData_0n[29], outData_1n[29]);
  OR2 I48 (outComplete_0n[30], outData_0n[30], outData_1n[30]);
  OR2 I49 (outComplete_0n[31], outData_0n[31], outData_1n[31]);
  OR2 I50 (outComplete_0n[32], outData_0n[32], outData_1n[32]);
  C2 I51 (outData_1n[0], inp_0r1d[0], poutReqB_0n);
  C2 I52 (outData_1n[1], inp_0r1d[1], poutReqB_0n);
  C2 I53 (outData_1n[2], inp_0r1d[2], poutReqB_0n);
  C2 I54 (outData_1n[3], inp_0r1d[3], poutReqB_0n);
  C2 I55 (outData_1n[4], inp_0r1d[4], poutReqB_0n);
  C2 I56 (outData_1n[5], inp_0r1d[5], poutReqB_0n);
  C2 I57 (outData_1n[6], inp_0r1d[6], poutReqB_0n);
  C2 I58 (outData_1n[7], inp_0r1d[7], poutReqB_0n);
  C2 I59 (outData_1n[8], inp_0r1d[8], poutReqB_0n);
  C2 I60 (outData_1n[9], inp_0r1d[9], poutReqB_0n);
  C2 I61 (outData_1n[10], inp_0r1d[10], poutReqB_0n);
  C2 I62 (outData_1n[11], inp_0r1d[11], poutReqB_0n);
  C2 I63 (outData_1n[12], inp_0r1d[12], poutReqB_0n);
  C2 I64 (outData_1n[13], inp_0r1d[13], poutReqB_0n);
  C2 I65 (outData_1n[14], inp_0r1d[14], poutReqB_0n);
  C2 I66 (outData_1n[15], inp_0r1d[15], poutReqB_0n);
  C2 I67 (outData_1n[16], inp_0r1d[16], poutReqB_0n);
  C2 I68 (outData_1n[17], inp_0r1d[17], poutReqB_0n);
  C2 I69 (outData_1n[18], inp_0r1d[18], poutReqB_0n);
  C2 I70 (outData_1n[19], inp_0r1d[19], poutReqB_0n);
  C2 I71 (outData_1n[20], inp_0r1d[20], poutReqB_0n);
  C2 I72 (outData_1n[21], inp_0r1d[21], poutReqB_0n);
  C2 I73 (outData_1n[22], inp_0r1d[22], poutReqB_0n);
  C2 I74 (outData_1n[23], inp_0r1d[23], poutReqB_0n);
  C2 I75 (outData_1n[24], inp_0r1d[24], poutReqB_0n);
  C2 I76 (outData_1n[25], inp_0r1d[25], poutReqB_0n);
  C2 I77 (outData_1n[26], inp_0r1d[26], poutReqB_0n);
  C2 I78 (outData_1n[27], inp_0r1d[27], poutReqB_0n);
  C2 I79 (outData_1n[28], inp_0r1d[28], poutReqB_0n);
  C2 I80 (outData_1n[29], inp_0r1d[29], poutReqB_0n);
  C2 I81 (outData_1n[30], inp_0r1d[30], poutReqB_0n);
  C2 I82 (outData_1n[31], inp_0r1d[31], poutReqB_0n);
  C2 I83 (outData_1n[32], inp_0r1d[32], poutReqB_0n);
  C2 I84 (outData_0n[0], inp_0r0d[0], poutReqB_0n);
  C2 I85 (outData_0n[1], inp_0r0d[1], poutReqB_0n);
  C2 I86 (outData_0n[2], inp_0r0d[2], poutReqB_0n);
  C2 I87 (outData_0n[3], inp_0r0d[3], poutReqB_0n);
  C2 I88 (outData_0n[4], inp_0r0d[4], poutReqB_0n);
  C2 I89 (outData_0n[5], inp_0r0d[5], poutReqB_0n);
  C2 I90 (outData_0n[6], inp_0r0d[6], poutReqB_0n);
  C2 I91 (outData_0n[7], inp_0r0d[7], poutReqB_0n);
  C2 I92 (outData_0n[8], inp_0r0d[8], poutReqB_0n);
  C2 I93 (outData_0n[9], inp_0r0d[9], poutReqB_0n);
  C2 I94 (outData_0n[10], inp_0r0d[10], poutReqB_0n);
  C2 I95 (outData_0n[11], inp_0r0d[11], poutReqB_0n);
  C2 I96 (outData_0n[12], inp_0r0d[12], poutReqB_0n);
  C2 I97 (outData_0n[13], inp_0r0d[13], poutReqB_0n);
  C2 I98 (outData_0n[14], inp_0r0d[14], poutReqB_0n);
  C2 I99 (outData_0n[15], inp_0r0d[15], poutReqB_0n);
  C2 I100 (outData_0n[16], inp_0r0d[16], poutReqB_0n);
  C2 I101 (outData_0n[17], inp_0r0d[17], poutReqB_0n);
  C2 I102 (outData_0n[18], inp_0r0d[18], poutReqB_0n);
  C2 I103 (outData_0n[19], inp_0r0d[19], poutReqB_0n);
  C2 I104 (outData_0n[20], inp_0r0d[20], poutReqB_0n);
  C2 I105 (outData_0n[21], inp_0r0d[21], poutReqB_0n);
  C2 I106 (outData_0n[22], inp_0r0d[22], poutReqB_0n);
  C2 I107 (outData_0n[23], inp_0r0d[23], poutReqB_0n);
  C2 I108 (outData_0n[24], inp_0r0d[24], poutReqB_0n);
  C2 I109 (outData_0n[25], inp_0r0d[25], poutReqB_0n);
  C2 I110 (outData_0n[26], inp_0r0d[26], poutReqB_0n);
  C2 I111 (outData_0n[27], inp_0r0d[27], poutReqB_0n);
  C2 I112 (outData_0n[28], inp_0r0d[28], poutReqB_0n);
  C2 I113 (outData_0n[29], inp_0r0d[29], poutReqB_0n);
  C2 I114 (outData_0n[30], inp_0r0d[30], poutReqB_0n);
  C2 I115 (outData_0n[31], inp_0r0d[31], poutReqB_0n);
  C2 I116 (outData_0n[32], inp_0r0d[32], poutReqB_0n);
  BUFF I117 (poutReq_0n, out_0r);
  BUFF I118 (poutReqB_0n, poutReq_0n);
  BUFF I119 (out_0a1d[0], outData_1n[0]);
  BUFF I120 (out_0a1d[1], outData_1n[1]);
  BUFF I121 (out_0a1d[2], outData_1n[2]);
  BUFF I122 (out_0a1d[3], outData_1n[3]);
  BUFF I123 (out_0a1d[4], outData_1n[4]);
  BUFF I124 (out_0a1d[5], outData_1n[5]);
  BUFF I125 (out_0a1d[6], outData_1n[6]);
  BUFF I126 (out_0a1d[7], outData_1n[7]);
  BUFF I127 (out_0a1d[8], outData_1n[8]);
  BUFF I128 (out_0a1d[9], outData_1n[9]);
  BUFF I129 (out_0a1d[10], outData_1n[10]);
  BUFF I130 (out_0a1d[11], outData_1n[11]);
  BUFF I131 (out_0a1d[12], outData_1n[12]);
  BUFF I132 (out_0a1d[13], outData_1n[13]);
  BUFF I133 (out_0a1d[14], outData_1n[14]);
  BUFF I134 (out_0a1d[15], outData_1n[15]);
  BUFF I135 (out_0a1d[16], outData_1n[16]);
  BUFF I136 (out_0a1d[17], outData_1n[17]);
  BUFF I137 (out_0a1d[18], outData_1n[18]);
  BUFF I138 (out_0a1d[19], outData_1n[19]);
  BUFF I139 (out_0a1d[20], outData_1n[20]);
  BUFF I140 (out_0a1d[21], outData_1n[21]);
  BUFF I141 (out_0a1d[22], outData_1n[22]);
  BUFF I142 (out_0a1d[23], outData_1n[23]);
  BUFF I143 (out_0a1d[24], outData_1n[24]);
  BUFF I144 (out_0a1d[25], outData_1n[25]);
  BUFF I145 (out_0a1d[26], outData_1n[26]);
  BUFF I146 (out_0a1d[27], outData_1n[27]);
  BUFF I147 (out_0a1d[28], outData_1n[28]);
  BUFF I148 (out_0a1d[29], outData_1n[29]);
  BUFF I149 (out_0a1d[30], outData_1n[30]);
  BUFF I150 (out_0a1d[31], outData_1n[31]);
  BUFF I151 (out_0a1d[32], outData_1n[32]);
  BUFF I152 (out_0a0d[0], outData_0n[0]);
  BUFF I153 (out_0a0d[1], outData_0n[1]);
  BUFF I154 (out_0a0d[2], outData_0n[2]);
  BUFF I155 (out_0a0d[3], outData_0n[3]);
  BUFF I156 (out_0a0d[4], outData_0n[4]);
  BUFF I157 (out_0a0d[5], outData_0n[5]);
  BUFF I158 (out_0a0d[6], outData_0n[6]);
  BUFF I159 (out_0a0d[7], outData_0n[7]);
  BUFF I160 (out_0a0d[8], outData_0n[8]);
  BUFF I161 (out_0a0d[9], outData_0n[9]);
  BUFF I162 (out_0a0d[10], outData_0n[10]);
  BUFF I163 (out_0a0d[11], outData_0n[11]);
  BUFF I164 (out_0a0d[12], outData_0n[12]);
  BUFF I165 (out_0a0d[13], outData_0n[13]);
  BUFF I166 (out_0a0d[14], outData_0n[14]);
  BUFF I167 (out_0a0d[15], outData_0n[15]);
  BUFF I168 (out_0a0d[16], outData_0n[16]);
  BUFF I169 (out_0a0d[17], outData_0n[17]);
  BUFF I170 (out_0a0d[18], outData_0n[18]);
  BUFF I171 (out_0a0d[19], outData_0n[19]);
  BUFF I172 (out_0a0d[20], outData_0n[20]);
  BUFF I173 (out_0a0d[21], outData_0n[21]);
  BUFF I174 (out_0a0d[22], outData_0n[22]);
  BUFF I175 (out_0a0d[23], outData_0n[23]);
  BUFF I176 (out_0a0d[24], outData_0n[24]);
  BUFF I177 (out_0a0d[25], outData_0n[25]);
  BUFF I178 (out_0a0d[26], outData_0n[26]);
  BUFF I179 (out_0a0d[27], outData_0n[27]);
  BUFF I180 (out_0a0d[28], outData_0n[28]);
  BUFF I181 (out_0a0d[29], outData_0n[29]);
  BUFF I182 (out_0a0d[30], outData_0n[30]);
  BUFF I183 (out_0a0d[31], outData_0n[31]);
  BUFF I184 (out_0a0d[32], outData_0n[32]);
endmodule

module BrzPassivatorPush_34_1 (
  out_0r, out_0a0d, out_0a1d,
  inp_0r0d, inp_0r1d, inp_0a
);
  input out_0r;
  output [33:0] out_0a0d;
  output [33:0] out_0a1d;
  input [33:0] inp_0r0d;
  input [33:0] inp_0r1d;
  output inp_0a;
  wire [17:0] internal_0n;
  wire poutReq_0n;
  wire poutReqB_0n;
  wire [33:0] outComplete_0n;
  wire [33:0] outData_0n;
  wire [33:0] outData_1n;
  C3 I0 (internal_0n[0], outComplete_0n[0], outComplete_0n[1], outComplete_0n[2]);
  C3 I1 (internal_0n[1], outComplete_0n[3], outComplete_0n[4], outComplete_0n[5]);
  C3 I2 (internal_0n[2], outComplete_0n[6], outComplete_0n[7], outComplete_0n[8]);
  C3 I3 (internal_0n[3], outComplete_0n[9], outComplete_0n[10], outComplete_0n[11]);
  C3 I4 (internal_0n[4], outComplete_0n[12], outComplete_0n[13], outComplete_0n[14]);
  C3 I5 (internal_0n[5], outComplete_0n[15], outComplete_0n[16], outComplete_0n[17]);
  C3 I6 (internal_0n[6], outComplete_0n[18], outComplete_0n[19], outComplete_0n[20]);
  C3 I7 (internal_0n[7], outComplete_0n[21], outComplete_0n[22], outComplete_0n[23]);
  C3 I8 (internal_0n[8], outComplete_0n[24], outComplete_0n[25], outComplete_0n[26]);
  C3 I9 (internal_0n[9], outComplete_0n[27], outComplete_0n[28], outComplete_0n[29]);
  C2 I10 (internal_0n[10], outComplete_0n[30], outComplete_0n[31]);
  C2 I11 (internal_0n[11], outComplete_0n[32], outComplete_0n[33]);
  C3 I12 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I13 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I14 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I15 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I16 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I17 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I18 (inp_0a, internal_0n[16], internal_0n[17]);
  OR2 I19 (outComplete_0n[0], outData_0n[0], outData_1n[0]);
  OR2 I20 (outComplete_0n[1], outData_0n[1], outData_1n[1]);
  OR2 I21 (outComplete_0n[2], outData_0n[2], outData_1n[2]);
  OR2 I22 (outComplete_0n[3], outData_0n[3], outData_1n[3]);
  OR2 I23 (outComplete_0n[4], outData_0n[4], outData_1n[4]);
  OR2 I24 (outComplete_0n[5], outData_0n[5], outData_1n[5]);
  OR2 I25 (outComplete_0n[6], outData_0n[6], outData_1n[6]);
  OR2 I26 (outComplete_0n[7], outData_0n[7], outData_1n[7]);
  OR2 I27 (outComplete_0n[8], outData_0n[8], outData_1n[8]);
  OR2 I28 (outComplete_0n[9], outData_0n[9], outData_1n[9]);
  OR2 I29 (outComplete_0n[10], outData_0n[10], outData_1n[10]);
  OR2 I30 (outComplete_0n[11], outData_0n[11], outData_1n[11]);
  OR2 I31 (outComplete_0n[12], outData_0n[12], outData_1n[12]);
  OR2 I32 (outComplete_0n[13], outData_0n[13], outData_1n[13]);
  OR2 I33 (outComplete_0n[14], outData_0n[14], outData_1n[14]);
  OR2 I34 (outComplete_0n[15], outData_0n[15], outData_1n[15]);
  OR2 I35 (outComplete_0n[16], outData_0n[16], outData_1n[16]);
  OR2 I36 (outComplete_0n[17], outData_0n[17], outData_1n[17]);
  OR2 I37 (outComplete_0n[18], outData_0n[18], outData_1n[18]);
  OR2 I38 (outComplete_0n[19], outData_0n[19], outData_1n[19]);
  OR2 I39 (outComplete_0n[20], outData_0n[20], outData_1n[20]);
  OR2 I40 (outComplete_0n[21], outData_0n[21], outData_1n[21]);
  OR2 I41 (outComplete_0n[22], outData_0n[22], outData_1n[22]);
  OR2 I42 (outComplete_0n[23], outData_0n[23], outData_1n[23]);
  OR2 I43 (outComplete_0n[24], outData_0n[24], outData_1n[24]);
  OR2 I44 (outComplete_0n[25], outData_0n[25], outData_1n[25]);
  OR2 I45 (outComplete_0n[26], outData_0n[26], outData_1n[26]);
  OR2 I46 (outComplete_0n[27], outData_0n[27], outData_1n[27]);
  OR2 I47 (outComplete_0n[28], outData_0n[28], outData_1n[28]);
  OR2 I48 (outComplete_0n[29], outData_0n[29], outData_1n[29]);
  OR2 I49 (outComplete_0n[30], outData_0n[30], outData_1n[30]);
  OR2 I50 (outComplete_0n[31], outData_0n[31], outData_1n[31]);
  OR2 I51 (outComplete_0n[32], outData_0n[32], outData_1n[32]);
  OR2 I52 (outComplete_0n[33], outData_0n[33], outData_1n[33]);
  C2 I53 (outData_1n[0], inp_0r1d[0], poutReqB_0n);
  C2 I54 (outData_1n[1], inp_0r1d[1], poutReqB_0n);
  C2 I55 (outData_1n[2], inp_0r1d[2], poutReqB_0n);
  C2 I56 (outData_1n[3], inp_0r1d[3], poutReqB_0n);
  C2 I57 (outData_1n[4], inp_0r1d[4], poutReqB_0n);
  C2 I58 (outData_1n[5], inp_0r1d[5], poutReqB_0n);
  C2 I59 (outData_1n[6], inp_0r1d[6], poutReqB_0n);
  C2 I60 (outData_1n[7], inp_0r1d[7], poutReqB_0n);
  C2 I61 (outData_1n[8], inp_0r1d[8], poutReqB_0n);
  C2 I62 (outData_1n[9], inp_0r1d[9], poutReqB_0n);
  C2 I63 (outData_1n[10], inp_0r1d[10], poutReqB_0n);
  C2 I64 (outData_1n[11], inp_0r1d[11], poutReqB_0n);
  C2 I65 (outData_1n[12], inp_0r1d[12], poutReqB_0n);
  C2 I66 (outData_1n[13], inp_0r1d[13], poutReqB_0n);
  C2 I67 (outData_1n[14], inp_0r1d[14], poutReqB_0n);
  C2 I68 (outData_1n[15], inp_0r1d[15], poutReqB_0n);
  C2 I69 (outData_1n[16], inp_0r1d[16], poutReqB_0n);
  C2 I70 (outData_1n[17], inp_0r1d[17], poutReqB_0n);
  C2 I71 (outData_1n[18], inp_0r1d[18], poutReqB_0n);
  C2 I72 (outData_1n[19], inp_0r1d[19], poutReqB_0n);
  C2 I73 (outData_1n[20], inp_0r1d[20], poutReqB_0n);
  C2 I74 (outData_1n[21], inp_0r1d[21], poutReqB_0n);
  C2 I75 (outData_1n[22], inp_0r1d[22], poutReqB_0n);
  C2 I76 (outData_1n[23], inp_0r1d[23], poutReqB_0n);
  C2 I77 (outData_1n[24], inp_0r1d[24], poutReqB_0n);
  C2 I78 (outData_1n[25], inp_0r1d[25], poutReqB_0n);
  C2 I79 (outData_1n[26], inp_0r1d[26], poutReqB_0n);
  C2 I80 (outData_1n[27], inp_0r1d[27], poutReqB_0n);
  C2 I81 (outData_1n[28], inp_0r1d[28], poutReqB_0n);
  C2 I82 (outData_1n[29], inp_0r1d[29], poutReqB_0n);
  C2 I83 (outData_1n[30], inp_0r1d[30], poutReqB_0n);
  C2 I84 (outData_1n[31], inp_0r1d[31], poutReqB_0n);
  C2 I85 (outData_1n[32], inp_0r1d[32], poutReqB_0n);
  C2 I86 (outData_1n[33], inp_0r1d[33], poutReqB_0n);
  C2 I87 (outData_0n[0], inp_0r0d[0], poutReqB_0n);
  C2 I88 (outData_0n[1], inp_0r0d[1], poutReqB_0n);
  C2 I89 (outData_0n[2], inp_0r0d[2], poutReqB_0n);
  C2 I90 (outData_0n[3], inp_0r0d[3], poutReqB_0n);
  C2 I91 (outData_0n[4], inp_0r0d[4], poutReqB_0n);
  C2 I92 (outData_0n[5], inp_0r0d[5], poutReqB_0n);
  C2 I93 (outData_0n[6], inp_0r0d[6], poutReqB_0n);
  C2 I94 (outData_0n[7], inp_0r0d[7], poutReqB_0n);
  C2 I95 (outData_0n[8], inp_0r0d[8], poutReqB_0n);
  C2 I96 (outData_0n[9], inp_0r0d[9], poutReqB_0n);
  C2 I97 (outData_0n[10], inp_0r0d[10], poutReqB_0n);
  C2 I98 (outData_0n[11], inp_0r0d[11], poutReqB_0n);
  C2 I99 (outData_0n[12], inp_0r0d[12], poutReqB_0n);
  C2 I100 (outData_0n[13], inp_0r0d[13], poutReqB_0n);
  C2 I101 (outData_0n[14], inp_0r0d[14], poutReqB_0n);
  C2 I102 (outData_0n[15], inp_0r0d[15], poutReqB_0n);
  C2 I103 (outData_0n[16], inp_0r0d[16], poutReqB_0n);
  C2 I104 (outData_0n[17], inp_0r0d[17], poutReqB_0n);
  C2 I105 (outData_0n[18], inp_0r0d[18], poutReqB_0n);
  C2 I106 (outData_0n[19], inp_0r0d[19], poutReqB_0n);
  C2 I107 (outData_0n[20], inp_0r0d[20], poutReqB_0n);
  C2 I108 (outData_0n[21], inp_0r0d[21], poutReqB_0n);
  C2 I109 (outData_0n[22], inp_0r0d[22], poutReqB_0n);
  C2 I110 (outData_0n[23], inp_0r0d[23], poutReqB_0n);
  C2 I111 (outData_0n[24], inp_0r0d[24], poutReqB_0n);
  C2 I112 (outData_0n[25], inp_0r0d[25], poutReqB_0n);
  C2 I113 (outData_0n[26], inp_0r0d[26], poutReqB_0n);
  C2 I114 (outData_0n[27], inp_0r0d[27], poutReqB_0n);
  C2 I115 (outData_0n[28], inp_0r0d[28], poutReqB_0n);
  C2 I116 (outData_0n[29], inp_0r0d[29], poutReqB_0n);
  C2 I117 (outData_0n[30], inp_0r0d[30], poutReqB_0n);
  C2 I118 (outData_0n[31], inp_0r0d[31], poutReqB_0n);
  C2 I119 (outData_0n[32], inp_0r0d[32], poutReqB_0n);
  C2 I120 (outData_0n[33], inp_0r0d[33], poutReqB_0n);
  BUFF I121 (poutReq_0n, out_0r);
  BUFF I122 (poutReqB_0n, poutReq_0n);
  BUFF I123 (out_0a1d[0], outData_1n[0]);
  BUFF I124 (out_0a1d[1], outData_1n[1]);
  BUFF I125 (out_0a1d[2], outData_1n[2]);
  BUFF I126 (out_0a1d[3], outData_1n[3]);
  BUFF I127 (out_0a1d[4], outData_1n[4]);
  BUFF I128 (out_0a1d[5], outData_1n[5]);
  BUFF I129 (out_0a1d[6], outData_1n[6]);
  BUFF I130 (out_0a1d[7], outData_1n[7]);
  BUFF I131 (out_0a1d[8], outData_1n[8]);
  BUFF I132 (out_0a1d[9], outData_1n[9]);
  BUFF I133 (out_0a1d[10], outData_1n[10]);
  BUFF I134 (out_0a1d[11], outData_1n[11]);
  BUFF I135 (out_0a1d[12], outData_1n[12]);
  BUFF I136 (out_0a1d[13], outData_1n[13]);
  BUFF I137 (out_0a1d[14], outData_1n[14]);
  BUFF I138 (out_0a1d[15], outData_1n[15]);
  BUFF I139 (out_0a1d[16], outData_1n[16]);
  BUFF I140 (out_0a1d[17], outData_1n[17]);
  BUFF I141 (out_0a1d[18], outData_1n[18]);
  BUFF I142 (out_0a1d[19], outData_1n[19]);
  BUFF I143 (out_0a1d[20], outData_1n[20]);
  BUFF I144 (out_0a1d[21], outData_1n[21]);
  BUFF I145 (out_0a1d[22], outData_1n[22]);
  BUFF I146 (out_0a1d[23], outData_1n[23]);
  BUFF I147 (out_0a1d[24], outData_1n[24]);
  BUFF I148 (out_0a1d[25], outData_1n[25]);
  BUFF I149 (out_0a1d[26], outData_1n[26]);
  BUFF I150 (out_0a1d[27], outData_1n[27]);
  BUFF I151 (out_0a1d[28], outData_1n[28]);
  BUFF I152 (out_0a1d[29], outData_1n[29]);
  BUFF I153 (out_0a1d[30], outData_1n[30]);
  BUFF I154 (out_0a1d[31], outData_1n[31]);
  BUFF I155 (out_0a1d[32], outData_1n[32]);
  BUFF I156 (out_0a1d[33], outData_1n[33]);
  BUFF I157 (out_0a0d[0], outData_0n[0]);
  BUFF I158 (out_0a0d[1], outData_0n[1]);
  BUFF I159 (out_0a0d[2], outData_0n[2]);
  BUFF I160 (out_0a0d[3], outData_0n[3]);
  BUFF I161 (out_0a0d[4], outData_0n[4]);
  BUFF I162 (out_0a0d[5], outData_0n[5]);
  BUFF I163 (out_0a0d[6], outData_0n[6]);
  BUFF I164 (out_0a0d[7], outData_0n[7]);
  BUFF I165 (out_0a0d[8], outData_0n[8]);
  BUFF I166 (out_0a0d[9], outData_0n[9]);
  BUFF I167 (out_0a0d[10], outData_0n[10]);
  BUFF I168 (out_0a0d[11], outData_0n[11]);
  BUFF I169 (out_0a0d[12], outData_0n[12]);
  BUFF I170 (out_0a0d[13], outData_0n[13]);
  BUFF I171 (out_0a0d[14], outData_0n[14]);
  BUFF I172 (out_0a0d[15], outData_0n[15]);
  BUFF I173 (out_0a0d[16], outData_0n[16]);
  BUFF I174 (out_0a0d[17], outData_0n[17]);
  BUFF I175 (out_0a0d[18], outData_0n[18]);
  BUFF I176 (out_0a0d[19], outData_0n[19]);
  BUFF I177 (out_0a0d[20], outData_0n[20]);
  BUFF I178 (out_0a0d[21], outData_0n[21]);
  BUFF I179 (out_0a0d[22], outData_0n[22]);
  BUFF I180 (out_0a0d[23], outData_0n[23]);
  BUFF I181 (out_0a0d[24], outData_0n[24]);
  BUFF I182 (out_0a0d[25], outData_0n[25]);
  BUFF I183 (out_0a0d[26], outData_0n[26]);
  BUFF I184 (out_0a0d[27], outData_0n[27]);
  BUFF I185 (out_0a0d[28], outData_0n[28]);
  BUFF I186 (out_0a0d[29], outData_0n[29]);
  BUFF I187 (out_0a0d[30], outData_0n[30]);
  BUFF I188 (out_0a0d[31], outData_0n[31]);
  BUFF I189 (out_0a0d[32], outData_0n[32]);
  BUFF I190 (out_0a0d[33], outData_0n[33]);
endmodule

module BrzPassivatorPush_35_1 (
  out_0r, out_0a0d, out_0a1d,
  inp_0r0d, inp_0r1d, inp_0a
);
  input out_0r;
  output [34:0] out_0a0d;
  output [34:0] out_0a1d;
  input [34:0] inp_0r0d;
  input [34:0] inp_0r1d;
  output inp_0a;
  wire [17:0] internal_0n;
  wire poutReq_0n;
  wire poutReqB_0n;
  wire [34:0] outComplete_0n;
  wire [34:0] outData_0n;
  wire [34:0] outData_1n;
  C3 I0 (internal_0n[0], outComplete_0n[0], outComplete_0n[1], outComplete_0n[2]);
  C3 I1 (internal_0n[1], outComplete_0n[3], outComplete_0n[4], outComplete_0n[5]);
  C3 I2 (internal_0n[2], outComplete_0n[6], outComplete_0n[7], outComplete_0n[8]);
  C3 I3 (internal_0n[3], outComplete_0n[9], outComplete_0n[10], outComplete_0n[11]);
  C3 I4 (internal_0n[4], outComplete_0n[12], outComplete_0n[13], outComplete_0n[14]);
  C3 I5 (internal_0n[5], outComplete_0n[15], outComplete_0n[16], outComplete_0n[17]);
  C3 I6 (internal_0n[6], outComplete_0n[18], outComplete_0n[19], outComplete_0n[20]);
  C3 I7 (internal_0n[7], outComplete_0n[21], outComplete_0n[22], outComplete_0n[23]);
  C3 I8 (internal_0n[8], outComplete_0n[24], outComplete_0n[25], outComplete_0n[26]);
  C3 I9 (internal_0n[9], outComplete_0n[27], outComplete_0n[28], outComplete_0n[29]);
  C3 I10 (internal_0n[10], outComplete_0n[30], outComplete_0n[31], outComplete_0n[32]);
  C2 I11 (internal_0n[11], outComplete_0n[33], outComplete_0n[34]);
  C3 I12 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I13 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I14 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I15 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I16 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I17 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I18 (inp_0a, internal_0n[16], internal_0n[17]);
  OR2 I19 (outComplete_0n[0], outData_0n[0], outData_1n[0]);
  OR2 I20 (outComplete_0n[1], outData_0n[1], outData_1n[1]);
  OR2 I21 (outComplete_0n[2], outData_0n[2], outData_1n[2]);
  OR2 I22 (outComplete_0n[3], outData_0n[3], outData_1n[3]);
  OR2 I23 (outComplete_0n[4], outData_0n[4], outData_1n[4]);
  OR2 I24 (outComplete_0n[5], outData_0n[5], outData_1n[5]);
  OR2 I25 (outComplete_0n[6], outData_0n[6], outData_1n[6]);
  OR2 I26 (outComplete_0n[7], outData_0n[7], outData_1n[7]);
  OR2 I27 (outComplete_0n[8], outData_0n[8], outData_1n[8]);
  OR2 I28 (outComplete_0n[9], outData_0n[9], outData_1n[9]);
  OR2 I29 (outComplete_0n[10], outData_0n[10], outData_1n[10]);
  OR2 I30 (outComplete_0n[11], outData_0n[11], outData_1n[11]);
  OR2 I31 (outComplete_0n[12], outData_0n[12], outData_1n[12]);
  OR2 I32 (outComplete_0n[13], outData_0n[13], outData_1n[13]);
  OR2 I33 (outComplete_0n[14], outData_0n[14], outData_1n[14]);
  OR2 I34 (outComplete_0n[15], outData_0n[15], outData_1n[15]);
  OR2 I35 (outComplete_0n[16], outData_0n[16], outData_1n[16]);
  OR2 I36 (outComplete_0n[17], outData_0n[17], outData_1n[17]);
  OR2 I37 (outComplete_0n[18], outData_0n[18], outData_1n[18]);
  OR2 I38 (outComplete_0n[19], outData_0n[19], outData_1n[19]);
  OR2 I39 (outComplete_0n[20], outData_0n[20], outData_1n[20]);
  OR2 I40 (outComplete_0n[21], outData_0n[21], outData_1n[21]);
  OR2 I41 (outComplete_0n[22], outData_0n[22], outData_1n[22]);
  OR2 I42 (outComplete_0n[23], outData_0n[23], outData_1n[23]);
  OR2 I43 (outComplete_0n[24], outData_0n[24], outData_1n[24]);
  OR2 I44 (outComplete_0n[25], outData_0n[25], outData_1n[25]);
  OR2 I45 (outComplete_0n[26], outData_0n[26], outData_1n[26]);
  OR2 I46 (outComplete_0n[27], outData_0n[27], outData_1n[27]);
  OR2 I47 (outComplete_0n[28], outData_0n[28], outData_1n[28]);
  OR2 I48 (outComplete_0n[29], outData_0n[29], outData_1n[29]);
  OR2 I49 (outComplete_0n[30], outData_0n[30], outData_1n[30]);
  OR2 I50 (outComplete_0n[31], outData_0n[31], outData_1n[31]);
  OR2 I51 (outComplete_0n[32], outData_0n[32], outData_1n[32]);
  OR2 I52 (outComplete_0n[33], outData_0n[33], outData_1n[33]);
  OR2 I53 (outComplete_0n[34], outData_0n[34], outData_1n[34]);
  C2 I54 (outData_1n[0], inp_0r1d[0], poutReqB_0n);
  C2 I55 (outData_1n[1], inp_0r1d[1], poutReqB_0n);
  C2 I56 (outData_1n[2], inp_0r1d[2], poutReqB_0n);
  C2 I57 (outData_1n[3], inp_0r1d[3], poutReqB_0n);
  C2 I58 (outData_1n[4], inp_0r1d[4], poutReqB_0n);
  C2 I59 (outData_1n[5], inp_0r1d[5], poutReqB_0n);
  C2 I60 (outData_1n[6], inp_0r1d[6], poutReqB_0n);
  C2 I61 (outData_1n[7], inp_0r1d[7], poutReqB_0n);
  C2 I62 (outData_1n[8], inp_0r1d[8], poutReqB_0n);
  C2 I63 (outData_1n[9], inp_0r1d[9], poutReqB_0n);
  C2 I64 (outData_1n[10], inp_0r1d[10], poutReqB_0n);
  C2 I65 (outData_1n[11], inp_0r1d[11], poutReqB_0n);
  C2 I66 (outData_1n[12], inp_0r1d[12], poutReqB_0n);
  C2 I67 (outData_1n[13], inp_0r1d[13], poutReqB_0n);
  C2 I68 (outData_1n[14], inp_0r1d[14], poutReqB_0n);
  C2 I69 (outData_1n[15], inp_0r1d[15], poutReqB_0n);
  C2 I70 (outData_1n[16], inp_0r1d[16], poutReqB_0n);
  C2 I71 (outData_1n[17], inp_0r1d[17], poutReqB_0n);
  C2 I72 (outData_1n[18], inp_0r1d[18], poutReqB_0n);
  C2 I73 (outData_1n[19], inp_0r1d[19], poutReqB_0n);
  C2 I74 (outData_1n[20], inp_0r1d[20], poutReqB_0n);
  C2 I75 (outData_1n[21], inp_0r1d[21], poutReqB_0n);
  C2 I76 (outData_1n[22], inp_0r1d[22], poutReqB_0n);
  C2 I77 (outData_1n[23], inp_0r1d[23], poutReqB_0n);
  C2 I78 (outData_1n[24], inp_0r1d[24], poutReqB_0n);
  C2 I79 (outData_1n[25], inp_0r1d[25], poutReqB_0n);
  C2 I80 (outData_1n[26], inp_0r1d[26], poutReqB_0n);
  C2 I81 (outData_1n[27], inp_0r1d[27], poutReqB_0n);
  C2 I82 (outData_1n[28], inp_0r1d[28], poutReqB_0n);
  C2 I83 (outData_1n[29], inp_0r1d[29], poutReqB_0n);
  C2 I84 (outData_1n[30], inp_0r1d[30], poutReqB_0n);
  C2 I85 (outData_1n[31], inp_0r1d[31], poutReqB_0n);
  C2 I86 (outData_1n[32], inp_0r1d[32], poutReqB_0n);
  C2 I87 (outData_1n[33], inp_0r1d[33], poutReqB_0n);
  C2 I88 (outData_1n[34], inp_0r1d[34], poutReqB_0n);
  C2 I89 (outData_0n[0], inp_0r0d[0], poutReqB_0n);
  C2 I90 (outData_0n[1], inp_0r0d[1], poutReqB_0n);
  C2 I91 (outData_0n[2], inp_0r0d[2], poutReqB_0n);
  C2 I92 (outData_0n[3], inp_0r0d[3], poutReqB_0n);
  C2 I93 (outData_0n[4], inp_0r0d[4], poutReqB_0n);
  C2 I94 (outData_0n[5], inp_0r0d[5], poutReqB_0n);
  C2 I95 (outData_0n[6], inp_0r0d[6], poutReqB_0n);
  C2 I96 (outData_0n[7], inp_0r0d[7], poutReqB_0n);
  C2 I97 (outData_0n[8], inp_0r0d[8], poutReqB_0n);
  C2 I98 (outData_0n[9], inp_0r0d[9], poutReqB_0n);
  C2 I99 (outData_0n[10], inp_0r0d[10], poutReqB_0n);
  C2 I100 (outData_0n[11], inp_0r0d[11], poutReqB_0n);
  C2 I101 (outData_0n[12], inp_0r0d[12], poutReqB_0n);
  C2 I102 (outData_0n[13], inp_0r0d[13], poutReqB_0n);
  C2 I103 (outData_0n[14], inp_0r0d[14], poutReqB_0n);
  C2 I104 (outData_0n[15], inp_0r0d[15], poutReqB_0n);
  C2 I105 (outData_0n[16], inp_0r0d[16], poutReqB_0n);
  C2 I106 (outData_0n[17], inp_0r0d[17], poutReqB_0n);
  C2 I107 (outData_0n[18], inp_0r0d[18], poutReqB_0n);
  C2 I108 (outData_0n[19], inp_0r0d[19], poutReqB_0n);
  C2 I109 (outData_0n[20], inp_0r0d[20], poutReqB_0n);
  C2 I110 (outData_0n[21], inp_0r0d[21], poutReqB_0n);
  C2 I111 (outData_0n[22], inp_0r0d[22], poutReqB_0n);
  C2 I112 (outData_0n[23], inp_0r0d[23], poutReqB_0n);
  C2 I113 (outData_0n[24], inp_0r0d[24], poutReqB_0n);
  C2 I114 (outData_0n[25], inp_0r0d[25], poutReqB_0n);
  C2 I115 (outData_0n[26], inp_0r0d[26], poutReqB_0n);
  C2 I116 (outData_0n[27], inp_0r0d[27], poutReqB_0n);
  C2 I117 (outData_0n[28], inp_0r0d[28], poutReqB_0n);
  C2 I118 (outData_0n[29], inp_0r0d[29], poutReqB_0n);
  C2 I119 (outData_0n[30], inp_0r0d[30], poutReqB_0n);
  C2 I120 (outData_0n[31], inp_0r0d[31], poutReqB_0n);
  C2 I121 (outData_0n[32], inp_0r0d[32], poutReqB_0n);
  C2 I122 (outData_0n[33], inp_0r0d[33], poutReqB_0n);
  C2 I123 (outData_0n[34], inp_0r0d[34], poutReqB_0n);
  BUFF I124 (poutReq_0n, out_0r);
  BUFF I125 (poutReqB_0n, poutReq_0n);
  BUFF I126 (out_0a1d[0], outData_1n[0]);
  BUFF I127 (out_0a1d[1], outData_1n[1]);
  BUFF I128 (out_0a1d[2], outData_1n[2]);
  BUFF I129 (out_0a1d[3], outData_1n[3]);
  BUFF I130 (out_0a1d[4], outData_1n[4]);
  BUFF I131 (out_0a1d[5], outData_1n[5]);
  BUFF I132 (out_0a1d[6], outData_1n[6]);
  BUFF I133 (out_0a1d[7], outData_1n[7]);
  BUFF I134 (out_0a1d[8], outData_1n[8]);
  BUFF I135 (out_0a1d[9], outData_1n[9]);
  BUFF I136 (out_0a1d[10], outData_1n[10]);
  BUFF I137 (out_0a1d[11], outData_1n[11]);
  BUFF I138 (out_0a1d[12], outData_1n[12]);
  BUFF I139 (out_0a1d[13], outData_1n[13]);
  BUFF I140 (out_0a1d[14], outData_1n[14]);
  BUFF I141 (out_0a1d[15], outData_1n[15]);
  BUFF I142 (out_0a1d[16], outData_1n[16]);
  BUFF I143 (out_0a1d[17], outData_1n[17]);
  BUFF I144 (out_0a1d[18], outData_1n[18]);
  BUFF I145 (out_0a1d[19], outData_1n[19]);
  BUFF I146 (out_0a1d[20], outData_1n[20]);
  BUFF I147 (out_0a1d[21], outData_1n[21]);
  BUFF I148 (out_0a1d[22], outData_1n[22]);
  BUFF I149 (out_0a1d[23], outData_1n[23]);
  BUFF I150 (out_0a1d[24], outData_1n[24]);
  BUFF I151 (out_0a1d[25], outData_1n[25]);
  BUFF I152 (out_0a1d[26], outData_1n[26]);
  BUFF I153 (out_0a1d[27], outData_1n[27]);
  BUFF I154 (out_0a1d[28], outData_1n[28]);
  BUFF I155 (out_0a1d[29], outData_1n[29]);
  BUFF I156 (out_0a1d[30], outData_1n[30]);
  BUFF I157 (out_0a1d[31], outData_1n[31]);
  BUFF I158 (out_0a1d[32], outData_1n[32]);
  BUFF I159 (out_0a1d[33], outData_1n[33]);
  BUFF I160 (out_0a1d[34], outData_1n[34]);
  BUFF I161 (out_0a0d[0], outData_0n[0]);
  BUFF I162 (out_0a0d[1], outData_0n[1]);
  BUFF I163 (out_0a0d[2], outData_0n[2]);
  BUFF I164 (out_0a0d[3], outData_0n[3]);
  BUFF I165 (out_0a0d[4], outData_0n[4]);
  BUFF I166 (out_0a0d[5], outData_0n[5]);
  BUFF I167 (out_0a0d[6], outData_0n[6]);
  BUFF I168 (out_0a0d[7], outData_0n[7]);
  BUFF I169 (out_0a0d[8], outData_0n[8]);
  BUFF I170 (out_0a0d[9], outData_0n[9]);
  BUFF I171 (out_0a0d[10], outData_0n[10]);
  BUFF I172 (out_0a0d[11], outData_0n[11]);
  BUFF I173 (out_0a0d[12], outData_0n[12]);
  BUFF I174 (out_0a0d[13], outData_0n[13]);
  BUFF I175 (out_0a0d[14], outData_0n[14]);
  BUFF I176 (out_0a0d[15], outData_0n[15]);
  BUFF I177 (out_0a0d[16], outData_0n[16]);
  BUFF I178 (out_0a0d[17], outData_0n[17]);
  BUFF I179 (out_0a0d[18], outData_0n[18]);
  BUFF I180 (out_0a0d[19], outData_0n[19]);
  BUFF I181 (out_0a0d[20], outData_0n[20]);
  BUFF I182 (out_0a0d[21], outData_0n[21]);
  BUFF I183 (out_0a0d[22], outData_0n[22]);
  BUFF I184 (out_0a0d[23], outData_0n[23]);
  BUFF I185 (out_0a0d[24], outData_0n[24]);
  BUFF I186 (out_0a0d[25], outData_0n[25]);
  BUFF I187 (out_0a0d[26], outData_0n[26]);
  BUFF I188 (out_0a0d[27], outData_0n[27]);
  BUFF I189 (out_0a0d[28], outData_0n[28]);
  BUFF I190 (out_0a0d[29], outData_0n[29]);
  BUFF I191 (out_0a0d[30], outData_0n[30]);
  BUFF I192 (out_0a0d[31], outData_0n[31]);
  BUFF I193 (out_0a0d[32], outData_0n[32]);
  BUFF I194 (out_0a0d[33], outData_0n[33]);
  BUFF I195 (out_0a0d[34], outData_0n[34]);
endmodule

module BrzPassivatorPush_36_1 (
  out_0r, out_0a0d, out_0a1d,
  inp_0r0d, inp_0r1d, inp_0a
);
  input out_0r;
  output [35:0] out_0a0d;
  output [35:0] out_0a1d;
  input [35:0] inp_0r0d;
  input [35:0] inp_0r1d;
  output inp_0a;
  wire [17:0] internal_0n;
  wire poutReq_0n;
  wire poutReqB_0n;
  wire [35:0] outComplete_0n;
  wire [35:0] outData_0n;
  wire [35:0] outData_1n;
  C3 I0 (internal_0n[0], outComplete_0n[0], outComplete_0n[1], outComplete_0n[2]);
  C3 I1 (internal_0n[1], outComplete_0n[3], outComplete_0n[4], outComplete_0n[5]);
  C3 I2 (internal_0n[2], outComplete_0n[6], outComplete_0n[7], outComplete_0n[8]);
  C3 I3 (internal_0n[3], outComplete_0n[9], outComplete_0n[10], outComplete_0n[11]);
  C3 I4 (internal_0n[4], outComplete_0n[12], outComplete_0n[13], outComplete_0n[14]);
  C3 I5 (internal_0n[5], outComplete_0n[15], outComplete_0n[16], outComplete_0n[17]);
  C3 I6 (internal_0n[6], outComplete_0n[18], outComplete_0n[19], outComplete_0n[20]);
  C3 I7 (internal_0n[7], outComplete_0n[21], outComplete_0n[22], outComplete_0n[23]);
  C3 I8 (internal_0n[8], outComplete_0n[24], outComplete_0n[25], outComplete_0n[26]);
  C3 I9 (internal_0n[9], outComplete_0n[27], outComplete_0n[28], outComplete_0n[29]);
  C3 I10 (internal_0n[10], outComplete_0n[30], outComplete_0n[31], outComplete_0n[32]);
  C3 I11 (internal_0n[11], outComplete_0n[33], outComplete_0n[34], outComplete_0n[35]);
  C3 I12 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I13 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I14 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I15 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I16 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I17 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I18 (inp_0a, internal_0n[16], internal_0n[17]);
  OR2 I19 (outComplete_0n[0], outData_0n[0], outData_1n[0]);
  OR2 I20 (outComplete_0n[1], outData_0n[1], outData_1n[1]);
  OR2 I21 (outComplete_0n[2], outData_0n[2], outData_1n[2]);
  OR2 I22 (outComplete_0n[3], outData_0n[3], outData_1n[3]);
  OR2 I23 (outComplete_0n[4], outData_0n[4], outData_1n[4]);
  OR2 I24 (outComplete_0n[5], outData_0n[5], outData_1n[5]);
  OR2 I25 (outComplete_0n[6], outData_0n[6], outData_1n[6]);
  OR2 I26 (outComplete_0n[7], outData_0n[7], outData_1n[7]);
  OR2 I27 (outComplete_0n[8], outData_0n[8], outData_1n[8]);
  OR2 I28 (outComplete_0n[9], outData_0n[9], outData_1n[9]);
  OR2 I29 (outComplete_0n[10], outData_0n[10], outData_1n[10]);
  OR2 I30 (outComplete_0n[11], outData_0n[11], outData_1n[11]);
  OR2 I31 (outComplete_0n[12], outData_0n[12], outData_1n[12]);
  OR2 I32 (outComplete_0n[13], outData_0n[13], outData_1n[13]);
  OR2 I33 (outComplete_0n[14], outData_0n[14], outData_1n[14]);
  OR2 I34 (outComplete_0n[15], outData_0n[15], outData_1n[15]);
  OR2 I35 (outComplete_0n[16], outData_0n[16], outData_1n[16]);
  OR2 I36 (outComplete_0n[17], outData_0n[17], outData_1n[17]);
  OR2 I37 (outComplete_0n[18], outData_0n[18], outData_1n[18]);
  OR2 I38 (outComplete_0n[19], outData_0n[19], outData_1n[19]);
  OR2 I39 (outComplete_0n[20], outData_0n[20], outData_1n[20]);
  OR2 I40 (outComplete_0n[21], outData_0n[21], outData_1n[21]);
  OR2 I41 (outComplete_0n[22], outData_0n[22], outData_1n[22]);
  OR2 I42 (outComplete_0n[23], outData_0n[23], outData_1n[23]);
  OR2 I43 (outComplete_0n[24], outData_0n[24], outData_1n[24]);
  OR2 I44 (outComplete_0n[25], outData_0n[25], outData_1n[25]);
  OR2 I45 (outComplete_0n[26], outData_0n[26], outData_1n[26]);
  OR2 I46 (outComplete_0n[27], outData_0n[27], outData_1n[27]);
  OR2 I47 (outComplete_0n[28], outData_0n[28], outData_1n[28]);
  OR2 I48 (outComplete_0n[29], outData_0n[29], outData_1n[29]);
  OR2 I49 (outComplete_0n[30], outData_0n[30], outData_1n[30]);
  OR2 I50 (outComplete_0n[31], outData_0n[31], outData_1n[31]);
  OR2 I51 (outComplete_0n[32], outData_0n[32], outData_1n[32]);
  OR2 I52 (outComplete_0n[33], outData_0n[33], outData_1n[33]);
  OR2 I53 (outComplete_0n[34], outData_0n[34], outData_1n[34]);
  OR2 I54 (outComplete_0n[35], outData_0n[35], outData_1n[35]);
  C2 I55 (outData_1n[0], inp_0r1d[0], poutReqB_0n);
  C2 I56 (outData_1n[1], inp_0r1d[1], poutReqB_0n);
  C2 I57 (outData_1n[2], inp_0r1d[2], poutReqB_0n);
  C2 I58 (outData_1n[3], inp_0r1d[3], poutReqB_0n);
  C2 I59 (outData_1n[4], inp_0r1d[4], poutReqB_0n);
  C2 I60 (outData_1n[5], inp_0r1d[5], poutReqB_0n);
  C2 I61 (outData_1n[6], inp_0r1d[6], poutReqB_0n);
  C2 I62 (outData_1n[7], inp_0r1d[7], poutReqB_0n);
  C2 I63 (outData_1n[8], inp_0r1d[8], poutReqB_0n);
  C2 I64 (outData_1n[9], inp_0r1d[9], poutReqB_0n);
  C2 I65 (outData_1n[10], inp_0r1d[10], poutReqB_0n);
  C2 I66 (outData_1n[11], inp_0r1d[11], poutReqB_0n);
  C2 I67 (outData_1n[12], inp_0r1d[12], poutReqB_0n);
  C2 I68 (outData_1n[13], inp_0r1d[13], poutReqB_0n);
  C2 I69 (outData_1n[14], inp_0r1d[14], poutReqB_0n);
  C2 I70 (outData_1n[15], inp_0r1d[15], poutReqB_0n);
  C2 I71 (outData_1n[16], inp_0r1d[16], poutReqB_0n);
  C2 I72 (outData_1n[17], inp_0r1d[17], poutReqB_0n);
  C2 I73 (outData_1n[18], inp_0r1d[18], poutReqB_0n);
  C2 I74 (outData_1n[19], inp_0r1d[19], poutReqB_0n);
  C2 I75 (outData_1n[20], inp_0r1d[20], poutReqB_0n);
  C2 I76 (outData_1n[21], inp_0r1d[21], poutReqB_0n);
  C2 I77 (outData_1n[22], inp_0r1d[22], poutReqB_0n);
  C2 I78 (outData_1n[23], inp_0r1d[23], poutReqB_0n);
  C2 I79 (outData_1n[24], inp_0r1d[24], poutReqB_0n);
  C2 I80 (outData_1n[25], inp_0r1d[25], poutReqB_0n);
  C2 I81 (outData_1n[26], inp_0r1d[26], poutReqB_0n);
  C2 I82 (outData_1n[27], inp_0r1d[27], poutReqB_0n);
  C2 I83 (outData_1n[28], inp_0r1d[28], poutReqB_0n);
  C2 I84 (outData_1n[29], inp_0r1d[29], poutReqB_0n);
  C2 I85 (outData_1n[30], inp_0r1d[30], poutReqB_0n);
  C2 I86 (outData_1n[31], inp_0r1d[31], poutReqB_0n);
  C2 I87 (outData_1n[32], inp_0r1d[32], poutReqB_0n);
  C2 I88 (outData_1n[33], inp_0r1d[33], poutReqB_0n);
  C2 I89 (outData_1n[34], inp_0r1d[34], poutReqB_0n);
  C2 I90 (outData_1n[35], inp_0r1d[35], poutReqB_0n);
  C2 I91 (outData_0n[0], inp_0r0d[0], poutReqB_0n);
  C2 I92 (outData_0n[1], inp_0r0d[1], poutReqB_0n);
  C2 I93 (outData_0n[2], inp_0r0d[2], poutReqB_0n);
  C2 I94 (outData_0n[3], inp_0r0d[3], poutReqB_0n);
  C2 I95 (outData_0n[4], inp_0r0d[4], poutReqB_0n);
  C2 I96 (outData_0n[5], inp_0r0d[5], poutReqB_0n);
  C2 I97 (outData_0n[6], inp_0r0d[6], poutReqB_0n);
  C2 I98 (outData_0n[7], inp_0r0d[7], poutReqB_0n);
  C2 I99 (outData_0n[8], inp_0r0d[8], poutReqB_0n);
  C2 I100 (outData_0n[9], inp_0r0d[9], poutReqB_0n);
  C2 I101 (outData_0n[10], inp_0r0d[10], poutReqB_0n);
  C2 I102 (outData_0n[11], inp_0r0d[11], poutReqB_0n);
  C2 I103 (outData_0n[12], inp_0r0d[12], poutReqB_0n);
  C2 I104 (outData_0n[13], inp_0r0d[13], poutReqB_0n);
  C2 I105 (outData_0n[14], inp_0r0d[14], poutReqB_0n);
  C2 I106 (outData_0n[15], inp_0r0d[15], poutReqB_0n);
  C2 I107 (outData_0n[16], inp_0r0d[16], poutReqB_0n);
  C2 I108 (outData_0n[17], inp_0r0d[17], poutReqB_0n);
  C2 I109 (outData_0n[18], inp_0r0d[18], poutReqB_0n);
  C2 I110 (outData_0n[19], inp_0r0d[19], poutReqB_0n);
  C2 I111 (outData_0n[20], inp_0r0d[20], poutReqB_0n);
  C2 I112 (outData_0n[21], inp_0r0d[21], poutReqB_0n);
  C2 I113 (outData_0n[22], inp_0r0d[22], poutReqB_0n);
  C2 I114 (outData_0n[23], inp_0r0d[23], poutReqB_0n);
  C2 I115 (outData_0n[24], inp_0r0d[24], poutReqB_0n);
  C2 I116 (outData_0n[25], inp_0r0d[25], poutReqB_0n);
  C2 I117 (outData_0n[26], inp_0r0d[26], poutReqB_0n);
  C2 I118 (outData_0n[27], inp_0r0d[27], poutReqB_0n);
  C2 I119 (outData_0n[28], inp_0r0d[28], poutReqB_0n);
  C2 I120 (outData_0n[29], inp_0r0d[29], poutReqB_0n);
  C2 I121 (outData_0n[30], inp_0r0d[30], poutReqB_0n);
  C2 I122 (outData_0n[31], inp_0r0d[31], poutReqB_0n);
  C2 I123 (outData_0n[32], inp_0r0d[32], poutReqB_0n);
  C2 I124 (outData_0n[33], inp_0r0d[33], poutReqB_0n);
  C2 I125 (outData_0n[34], inp_0r0d[34], poutReqB_0n);
  C2 I126 (outData_0n[35], inp_0r0d[35], poutReqB_0n);
  BUFF I127 (poutReq_0n, out_0r);
  BUFF I128 (poutReqB_0n, poutReq_0n);
  BUFF I129 (out_0a1d[0], outData_1n[0]);
  BUFF I130 (out_0a1d[1], outData_1n[1]);
  BUFF I131 (out_0a1d[2], outData_1n[2]);
  BUFF I132 (out_0a1d[3], outData_1n[3]);
  BUFF I133 (out_0a1d[4], outData_1n[4]);
  BUFF I134 (out_0a1d[5], outData_1n[5]);
  BUFF I135 (out_0a1d[6], outData_1n[6]);
  BUFF I136 (out_0a1d[7], outData_1n[7]);
  BUFF I137 (out_0a1d[8], outData_1n[8]);
  BUFF I138 (out_0a1d[9], outData_1n[9]);
  BUFF I139 (out_0a1d[10], outData_1n[10]);
  BUFF I140 (out_0a1d[11], outData_1n[11]);
  BUFF I141 (out_0a1d[12], outData_1n[12]);
  BUFF I142 (out_0a1d[13], outData_1n[13]);
  BUFF I143 (out_0a1d[14], outData_1n[14]);
  BUFF I144 (out_0a1d[15], outData_1n[15]);
  BUFF I145 (out_0a1d[16], outData_1n[16]);
  BUFF I146 (out_0a1d[17], outData_1n[17]);
  BUFF I147 (out_0a1d[18], outData_1n[18]);
  BUFF I148 (out_0a1d[19], outData_1n[19]);
  BUFF I149 (out_0a1d[20], outData_1n[20]);
  BUFF I150 (out_0a1d[21], outData_1n[21]);
  BUFF I151 (out_0a1d[22], outData_1n[22]);
  BUFF I152 (out_0a1d[23], outData_1n[23]);
  BUFF I153 (out_0a1d[24], outData_1n[24]);
  BUFF I154 (out_0a1d[25], outData_1n[25]);
  BUFF I155 (out_0a1d[26], outData_1n[26]);
  BUFF I156 (out_0a1d[27], outData_1n[27]);
  BUFF I157 (out_0a1d[28], outData_1n[28]);
  BUFF I158 (out_0a1d[29], outData_1n[29]);
  BUFF I159 (out_0a1d[30], outData_1n[30]);
  BUFF I160 (out_0a1d[31], outData_1n[31]);
  BUFF I161 (out_0a1d[32], outData_1n[32]);
  BUFF I162 (out_0a1d[33], outData_1n[33]);
  BUFF I163 (out_0a1d[34], outData_1n[34]);
  BUFF I164 (out_0a1d[35], outData_1n[35]);
  BUFF I165 (out_0a0d[0], outData_0n[0]);
  BUFF I166 (out_0a0d[1], outData_0n[1]);
  BUFF I167 (out_0a0d[2], outData_0n[2]);
  BUFF I168 (out_0a0d[3], outData_0n[3]);
  BUFF I169 (out_0a0d[4], outData_0n[4]);
  BUFF I170 (out_0a0d[5], outData_0n[5]);
  BUFF I171 (out_0a0d[6], outData_0n[6]);
  BUFF I172 (out_0a0d[7], outData_0n[7]);
  BUFF I173 (out_0a0d[8], outData_0n[8]);
  BUFF I174 (out_0a0d[9], outData_0n[9]);
  BUFF I175 (out_0a0d[10], outData_0n[10]);
  BUFF I176 (out_0a0d[11], outData_0n[11]);
  BUFF I177 (out_0a0d[12], outData_0n[12]);
  BUFF I178 (out_0a0d[13], outData_0n[13]);
  BUFF I179 (out_0a0d[14], outData_0n[14]);
  BUFF I180 (out_0a0d[15], outData_0n[15]);
  BUFF I181 (out_0a0d[16], outData_0n[16]);
  BUFF I182 (out_0a0d[17], outData_0n[17]);
  BUFF I183 (out_0a0d[18], outData_0n[18]);
  BUFF I184 (out_0a0d[19], outData_0n[19]);
  BUFF I185 (out_0a0d[20], outData_0n[20]);
  BUFF I186 (out_0a0d[21], outData_0n[21]);
  BUFF I187 (out_0a0d[22], outData_0n[22]);
  BUFF I188 (out_0a0d[23], outData_0n[23]);
  BUFF I189 (out_0a0d[24], outData_0n[24]);
  BUFF I190 (out_0a0d[25], outData_0n[25]);
  BUFF I191 (out_0a0d[26], outData_0n[26]);
  BUFF I192 (out_0a0d[27], outData_0n[27]);
  BUFF I193 (out_0a0d[28], outData_0n[28]);
  BUFF I194 (out_0a0d[29], outData_0n[29]);
  BUFF I195 (out_0a0d[30], outData_0n[30]);
  BUFF I196 (out_0a0d[31], outData_0n[31]);
  BUFF I197 (out_0a0d[32], outData_0n[32]);
  BUFF I198 (out_0a0d[33], outData_0n[33]);
  BUFF I199 (out_0a0d[34], outData_0n[34]);
  BUFF I200 (out_0a0d[35], outData_0n[35]);
endmodule

module BALSA_SELEM (
  Ar,
  Aa,
  Br,
  Ba
);
  input Ar;
  output Aa;
  output Br;
  input Ba;
  wire s;
  AND2 I0 (Br, Ar, s);
  NOR2 I1 (Aa, Ba, s);
  NC2P I2 (s, Ar, Ba);
endmodule

module BrzSequenceOptimised_2_s1_S (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  wire [1:0] sreq_0n;
  BUFF I0 (activate_0a, activateOut_1a);
  BUFF I1 (activateOut_1r, sreq_0n[1]);
  BUFF I2 (sreq_0n[0], activate_0r);
  BALSA_SELEM I3 (sreq_0n[0], sreq_0n[1], activateOut_0r, activateOut_0a);
endmodule

module BrzSequenceOptimised_2_s1_T (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  wire [1:0] sreq_0n;
  BUFF I0 (activate_0a, activateOut_1a);
  BUFF I1 (activateOut_1r, sreq_0n[1]);
  BUFF I2 (sreq_0n[0], activate_0r);
  BALSA_TELEM I3 (sreq_0n[0], sreq_0n[1], activateOut_0r, activateOut_0a);
endmodule

module BrzSequenceOptimised_5_s4_SSSS (
  activate_0r, activate_0a,
  activateOut_0r, activateOut_0a,
  activateOut_1r, activateOut_1a,
  activateOut_2r, activateOut_2a,
  activateOut_3r, activateOut_3a,
  activateOut_4r, activateOut_4a
);
  input activate_0r;
  output activate_0a;
  output activateOut_0r;
  input activateOut_0a;
  output activateOut_1r;
  input activateOut_1a;
  output activateOut_2r;
  input activateOut_2a;
  output activateOut_3r;
  input activateOut_3a;
  output activateOut_4r;
  input activateOut_4a;
  wire [4:0] sreq_0n;
  BUFF I0 (activate_0a, activateOut_4a);
  BUFF I1 (activateOut_4r, sreq_0n[4]);
  BUFF I2 (sreq_0n[0], activate_0r);
  BALSA_SELEM I3 (sreq_0n[3], sreq_0n[4], activateOut_3r, activateOut_3a);
  BALSA_SELEM I4 (sreq_0n[2], sreq_0n[3], activateOut_2r, activateOut_2a);
  BALSA_SELEM I5 (sreq_0n[1], sreq_0n[2], activateOut_1r, activateOut_1a);
  BALSA_SELEM I6 (sreq_0n[0], sreq_0n[1], activateOut_0r, activateOut_0a);
endmodule

module BrzSynch_2 (
  inp_0r, inp_0a,
  inp_1r, inp_1a,
  out_0r, out_0a
);
  input inp_0r;
  output inp_0a;
  input inp_1r;
  output inp_1a;
  output out_0r;
  input out_0a;
  wire inpAck_0n;
  C2 I0 (out_0r, inp_0r, inp_1r);
  BUFF I1 (inpAck_0n, out_0a);
  BUFF I2 (inp_0a, inpAck_0n);
  BUFF I3 (inp_1a, inpAck_0n);
endmodule

module BrzSynch_3 (
  inp_0r, inp_0a,
  inp_1r, inp_1a,
  inp_2r, inp_2a,
  out_0r, out_0a
);
  input inp_0r;
  output inp_0a;
  input inp_1r;
  output inp_1a;
  input inp_2r;
  output inp_2a;
  output out_0r;
  input out_0a;
  wire inpAck_0n;
  C3 I0 (out_0r, inp_0r, inp_1r, inp_2r);
  BUFF I1 (inpAck_0n, out_0a);
  BUFF I2 (inp_0a, inpAck_0n);
  BUFF I3 (inp_1a, inpAck_0n);
  BUFF I4 (inp_2a, inpAck_0n);
endmodule

module BrzSynch_4 (
  inp_0r, inp_0a,
  inp_1r, inp_1a,
  inp_2r, inp_2a,
  inp_3r, inp_3a,
  out_0r, out_0a
);
  input inp_0r;
  output inp_0a;
  input inp_1r;
  output inp_1a;
  input inp_2r;
  output inp_2a;
  input inp_3r;
  output inp_3a;
  output out_0r;
  input out_0a;
  wire [1:0] internal_0n;
  wire inpAck_0n;
  C2 I0 (internal_0n[0], inp_0r, inp_1r);
  C2 I1 (internal_0n[1], inp_2r, inp_3r);
  C2 I2 (out_0r, internal_0n[0], internal_0n[1]);
  BUFF I3 (inpAck_0n, out_0a);
  BUFF I4 (inp_0a, inpAck_0n);
  BUFF I5 (inp_1a, inpAck_0n);
  BUFF I6 (inp_2a, inpAck_0n);
  BUFF I7 (inp_3a, inpAck_0n);
endmodule

module BrzSynch_5 (
  inp_0r, inp_0a,
  inp_1r, inp_1a,
  inp_2r, inp_2a,
  inp_3r, inp_3a,
  inp_4r, inp_4a,
  out_0r, out_0a
);
  input inp_0r;
  output inp_0a;
  input inp_1r;
  output inp_1a;
  input inp_2r;
  output inp_2a;
  input inp_3r;
  output inp_3a;
  input inp_4r;
  output inp_4a;
  output out_0r;
  input out_0a;
  wire [1:0] internal_0n;
  wire inpAck_0n;
  C3 I0 (internal_0n[0], inp_0r, inp_1r, inp_2r);
  C2 I1 (internal_0n[1], inp_3r, inp_4r);
  C2 I2 (out_0r, internal_0n[0], internal_0n[1]);
  BUFF I3 (inpAck_0n, out_0a);
  BUFF I4 (inp_0a, inpAck_0n);
  BUFF I5 (inp_1a, inpAck_0n);
  BUFF I6 (inp_2a, inpAck_0n);
  BUFF I7 (inp_3a, inpAck_0n);
  BUFF I8 (inp_4a, inpAck_0n);
endmodule

module BrzUnaryFunc_35_35_s6_Invert_s5_false (
  out_0r, out_0a0d, out_0a1d,
  inp_0r, inp_0a0d, inp_0a1d
);
  input out_0r;
  output [34:0] out_0a0d;
  output [34:0] out_0a1d;
  output inp_0r;
  input [34:0] inp_0a0d;
  input [34:0] inp_0a1d;
  wire [35:0] c1_0n;
  wire [35:0] c0_0n;
  wire s1_0n;
  wire s0_0n;
  BUFF I0 (out_0a0d[0], inp_0a1d[0]);
  BUFF I1 (out_0a0d[1], inp_0a1d[1]);
  BUFF I2 (out_0a0d[2], inp_0a1d[2]);
  BUFF I3 (out_0a0d[3], inp_0a1d[3]);
  BUFF I4 (out_0a0d[4], inp_0a1d[4]);
  BUFF I5 (out_0a0d[5], inp_0a1d[5]);
  BUFF I6 (out_0a0d[6], inp_0a1d[6]);
  BUFF I7 (out_0a0d[7], inp_0a1d[7]);
  BUFF I8 (out_0a0d[8], inp_0a1d[8]);
  BUFF I9 (out_0a0d[9], inp_0a1d[9]);
  BUFF I10 (out_0a0d[10], inp_0a1d[10]);
  BUFF I11 (out_0a0d[11], inp_0a1d[11]);
  BUFF I12 (out_0a0d[12], inp_0a1d[12]);
  BUFF I13 (out_0a0d[13], inp_0a1d[13]);
  BUFF I14 (out_0a0d[14], inp_0a1d[14]);
  BUFF I15 (out_0a0d[15], inp_0a1d[15]);
  BUFF I16 (out_0a0d[16], inp_0a1d[16]);
  BUFF I17 (out_0a0d[17], inp_0a1d[17]);
  BUFF I18 (out_0a0d[18], inp_0a1d[18]);
  BUFF I19 (out_0a0d[19], inp_0a1d[19]);
  BUFF I20 (out_0a0d[20], inp_0a1d[20]);
  BUFF I21 (out_0a0d[21], inp_0a1d[21]);
  BUFF I22 (out_0a0d[22], inp_0a1d[22]);
  BUFF I23 (out_0a0d[23], inp_0a1d[23]);
  BUFF I24 (out_0a0d[24], inp_0a1d[24]);
  BUFF I25 (out_0a0d[25], inp_0a1d[25]);
  BUFF I26 (out_0a0d[26], inp_0a1d[26]);
  BUFF I27 (out_0a0d[27], inp_0a1d[27]);
  BUFF I28 (out_0a0d[28], inp_0a1d[28]);
  BUFF I29 (out_0a0d[29], inp_0a1d[29]);
  BUFF I30 (out_0a0d[30], inp_0a1d[30]);
  BUFF I31 (out_0a0d[31], inp_0a1d[31]);
  BUFF I32 (out_0a0d[32], inp_0a1d[32]);
  BUFF I33 (out_0a0d[33], inp_0a1d[33]);
  BUFF I34 (out_0a0d[34], inp_0a1d[34]);
  BUFF I35 (out_0a1d[0], inp_0a0d[0]);
  BUFF I36 (out_0a1d[1], inp_0a0d[1]);
  BUFF I37 (out_0a1d[2], inp_0a0d[2]);
  BUFF I38 (out_0a1d[3], inp_0a0d[3]);
  BUFF I39 (out_0a1d[4], inp_0a0d[4]);
  BUFF I40 (out_0a1d[5], inp_0a0d[5]);
  BUFF I41 (out_0a1d[6], inp_0a0d[6]);
  BUFF I42 (out_0a1d[7], inp_0a0d[7]);
  BUFF I43 (out_0a1d[8], inp_0a0d[8]);
  BUFF I44 (out_0a1d[9], inp_0a0d[9]);
  BUFF I45 (out_0a1d[10], inp_0a0d[10]);
  BUFF I46 (out_0a1d[11], inp_0a0d[11]);
  BUFF I47 (out_0a1d[12], inp_0a0d[12]);
  BUFF I48 (out_0a1d[13], inp_0a0d[13]);
  BUFF I49 (out_0a1d[14], inp_0a0d[14]);
  BUFF I50 (out_0a1d[15], inp_0a0d[15]);
  BUFF I51 (out_0a1d[16], inp_0a0d[16]);
  BUFF I52 (out_0a1d[17], inp_0a0d[17]);
  BUFF I53 (out_0a1d[18], inp_0a0d[18]);
  BUFF I54 (out_0a1d[19], inp_0a0d[19]);
  BUFF I55 (out_0a1d[20], inp_0a0d[20]);
  BUFF I56 (out_0a1d[21], inp_0a0d[21]);
  BUFF I57 (out_0a1d[22], inp_0a0d[22]);
  BUFF I58 (out_0a1d[23], inp_0a0d[23]);
  BUFF I59 (out_0a1d[24], inp_0a0d[24]);
  BUFF I60 (out_0a1d[25], inp_0a0d[25]);
  BUFF I61 (out_0a1d[26], inp_0a0d[26]);
  BUFF I62 (out_0a1d[27], inp_0a0d[27]);
  BUFF I63 (out_0a1d[28], inp_0a0d[28]);
  BUFF I64 (out_0a1d[29], inp_0a0d[29]);
  BUFF I65 (out_0a1d[30], inp_0a0d[30]);
  BUFF I66 (out_0a1d[31], inp_0a0d[31]);
  BUFF I67 (out_0a1d[32], inp_0a0d[32]);
  BUFF I68 (out_0a1d[33], inp_0a0d[33]);
  BUFF I69 (out_0a1d[34], inp_0a0d[34]);
  BUFF I70 (inp_0r, out_0r);
endmodule

module AO22 (
  q,
  i0,
  i1,
  i2,
  i3
);
  output q;
  input i0;
  input i1;
  input i2;
  input i3;
  wire [1:0] int_0n;
  OR2 I0 (q, int_0n[0], int_0n[1]);
  AND2 I1 (int_0n[1], i2, i3);
  AND2 I2 (int_0n[0], i0, i1);
endmodule

module DRLATCH (
  in_0,
  in_1,
  in_a,
  out_0,
  out_1
);
  input in_0;
  input in_1;
  output in_a;
  output out_0;
  output out_1;

`ifdef balsa_simulate
  initial begin
    force out_0 = 1;
    #`balsa_init_time;
    release out_0;
    if (out_0 !== 1)
        $display ("module %m: signal out_0 not correctly initialised");
  end
`endif

  AO22 I0 (in_a, in_0, out_0, in_1, out_1);
  NOR2 I1 (out_0, in_1, out_1);
  NOR2 I2 (out_1, in_0, out_0);
endmodule

module BrzVariable_1_1_s0_ (
  write_0r0d, write_0r1d, write_0a,
  read_0r, read_0a0d, read_0a1d
);
  input write_0r0d;
  input write_0r1d;
  output write_0a;
  input read_0r;
  output read_0a0d;
  output read_0a1d;
  wire store_0n;
  wire store_1n;
  wire ldata_0n;
  wire ldata_1n;
  wire wack_0n;
  wire readReq_0n;
  AND2 I0 (read_0a1d, store_1n, readReq_0n);
  AND2 I1 (read_0a0d, store_0n, readReq_0n);
  BUFF I2 (readReq_0n, read_0r);
  BUFF I3 (store_0n, ldata_0n);
  BUFF I4 (store_1n, ldata_1n);
  BUFF I5 (write_0a, wack_0n);
  DRLATCH I6 (write_0r0d, write_0r1d, wack_0n, ldata_0n, ldata_1n);
endmodule

module BrzVariable_1_2_s0_ (
  write_0r0d, write_0r1d, write_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d
);
  input write_0r0d;
  input write_0r1d;
  output write_0a;
  input read_0r;
  output read_0a0d;
  output read_0a1d;
  input read_1r;
  output read_1a0d;
  output read_1a1d;
  wire store_0n;
  wire store_1n;
  wire ldata_0n;
  wire ldata_1n;
  wire wack_0n;
  wire readReq_0n;
  wire readReq_1n;
  AND2 I0 (read_1a1d, store_1n, readReq_1n);
  AND2 I1 (read_1a0d, store_0n, readReq_1n);
  AND2 I2 (read_0a1d, store_1n, readReq_0n);
  AND2 I3 (read_0a0d, store_0n, readReq_0n);
  BUFF I4 (readReq_0n, read_0r);
  BUFF I5 (readReq_1n, read_1r);
  BUFF I6 (store_0n, ldata_0n);
  BUFF I7 (store_1n, ldata_1n);
  BUFF I8 (write_0a, wack_0n);
  DRLATCH I9 (write_0r0d, write_0r1d, wack_0n, ldata_0n, ldata_1n);
endmodule

module BrzVariable_1_3_s0_ (
  write_0r0d, write_0r1d, write_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d,
  read_2r, read_2a0d, read_2a1d
);
  input write_0r0d;
  input write_0r1d;
  output write_0a;
  input read_0r;
  output read_0a0d;
  output read_0a1d;
  input read_1r;
  output read_1a0d;
  output read_1a1d;
  input read_2r;
  output read_2a0d;
  output read_2a1d;
  wire store_0n;
  wire store_1n;
  wire ldata_0n;
  wire ldata_1n;
  wire wack_0n;
  wire readReq_0n;
  wire readReq_1n;
  wire readReq_2n;
  AND2 I0 (read_2a1d, store_1n, readReq_2n);
  AND2 I1 (read_2a0d, store_0n, readReq_2n);
  AND2 I2 (read_1a1d, store_1n, readReq_1n);
  AND2 I3 (read_1a0d, store_0n, readReq_1n);
  AND2 I4 (read_0a1d, store_1n, readReq_0n);
  AND2 I5 (read_0a0d, store_0n, readReq_0n);
  BUFF I6 (readReq_0n, read_0r);
  BUFF I7 (readReq_1n, read_1r);
  BUFF I8 (readReq_2n, read_2r);
  BUFF I9 (store_0n, ldata_0n);
  BUFF I10 (store_1n, ldata_1n);
  BUFF I11 (write_0a, wack_0n);
  DRLATCH I12 (write_0r0d, write_0r1d, wack_0n, ldata_0n, ldata_1n);
endmodule

module BrzVariable_4_3_s8_3_2e_2e3 (
  write_0r0d, write_0r1d, write_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d,
  read_2r, read_2a0d, read_2a1d
);
  input [3:0] write_0r0d;
  input [3:0] write_0r1d;
  output write_0a;
  input read_0r;
  output read_0a0d;
  output read_0a1d;
  input read_1r;
  output [3:0] read_1a0d;
  output [3:0] read_1a1d;
  input read_2r;
  output [3:0] read_2a0d;
  output [3:0] read_2a1d;
  wire [1:0] internal_0n;
  wire [3:0] store_0n;
  wire [3:0] store_1n;
  wire [3:0] ldata_0n;
  wire [3:0] ldata_1n;
  wire [3:0] wack_0n;
  wire readReq_0n;
  wire readReq_1n;
  wire readReq_2n;
  AND2 I0 (read_2a1d[0], store_1n[0], readReq_2n);
  AND2 I1 (read_2a1d[1], store_1n[1], readReq_2n);
  AND2 I2 (read_2a1d[2], store_1n[2], readReq_2n);
  AND2 I3 (read_2a1d[3], store_1n[3], readReq_2n);
  AND2 I4 (read_2a0d[0], store_0n[0], readReq_2n);
  AND2 I5 (read_2a0d[1], store_0n[1], readReq_2n);
  AND2 I6 (read_2a0d[2], store_0n[2], readReq_2n);
  AND2 I7 (read_2a0d[3], store_0n[3], readReq_2n);
  AND2 I8 (read_1a1d[0], store_1n[0], readReq_1n);
  AND2 I9 (read_1a1d[1], store_1n[1], readReq_1n);
  AND2 I10 (read_1a1d[2], store_1n[2], readReq_1n);
  AND2 I11 (read_1a1d[3], store_1n[3], readReq_1n);
  AND2 I12 (read_1a0d[0], store_0n[0], readReq_1n);
  AND2 I13 (read_1a0d[1], store_0n[1], readReq_1n);
  AND2 I14 (read_1a0d[2], store_0n[2], readReq_1n);
  AND2 I15 (read_1a0d[3], store_0n[3], readReq_1n);
  AND2 I16 (read_0a1d, store_1n[3], readReq_0n);
  AND2 I17 (read_0a0d, store_0n[3], readReq_0n);
  BUFF I18 (readReq_0n, read_0r);
  BUFF I19 (readReq_1n, read_1r);
  BUFF I20 (readReq_2n, read_2r);
  BUFF I21 (store_0n[0], ldata_0n[0]);
  BUFF I22 (store_0n[1], ldata_0n[1]);
  BUFF I23 (store_0n[2], ldata_0n[2]);
  BUFF I24 (store_0n[3], ldata_0n[3]);
  BUFF I25 (store_1n[0], ldata_1n[0]);
  BUFF I26 (store_1n[1], ldata_1n[1]);
  BUFF I27 (store_1n[2], ldata_1n[2]);
  BUFF I28 (store_1n[3], ldata_1n[3]);
  C2 I29 (internal_0n[0], wack_0n[0], wack_0n[1]);
  C2 I30 (internal_0n[1], wack_0n[2], wack_0n[3]);
  C2 I31 (write_0a, internal_0n[0], internal_0n[1]);
  DRLATCH I32 (write_0r0d[0], write_0r1d[0], wack_0n[0], ldata_0n[0], ldata_1n[0]);
  DRLATCH I33 (write_0r0d[1], write_0r1d[1], wack_0n[1], ldata_0n[1], ldata_1n[1]);
  DRLATCH I34 (write_0r0d[2], write_0r1d[2], wack_0n[2], ldata_0n[2], ldata_1n[2]);
  DRLATCH I35 (write_0r0d[3], write_0r1d[3], wack_0n[3], ldata_0n[3], ldata_1n[3]);
endmodule

module BrzVariable_10_1_s0_ (
  write_0r0d, write_0r1d, write_0a,
  read_0r, read_0a0d, read_0a1d
);
  input [9:0] write_0r0d;
  input [9:0] write_0r1d;
  output write_0a;
  input read_0r;
  output [9:0] read_0a0d;
  output [9:0] read_0a1d;
  wire [5:0] internal_0n;
  wire [9:0] store_0n;
  wire [9:0] store_1n;
  wire [9:0] ldata_0n;
  wire [9:0] ldata_1n;
  wire [9:0] wack_0n;
  wire readReq_0n;
  AND2 I0 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I1 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I2 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I3 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I4 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I5 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I6 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I7 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I8 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I9 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I10 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I11 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I12 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I13 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I14 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I15 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I16 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I17 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I18 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I19 (read_0a0d[9], store_0n[9], readReq_0n);
  BUFF I20 (readReq_0n, read_0r);
  BUFF I21 (store_0n[0], ldata_0n[0]);
  BUFF I22 (store_0n[1], ldata_0n[1]);
  BUFF I23 (store_0n[2], ldata_0n[2]);
  BUFF I24 (store_0n[3], ldata_0n[3]);
  BUFF I25 (store_0n[4], ldata_0n[4]);
  BUFF I26 (store_0n[5], ldata_0n[5]);
  BUFF I27 (store_0n[6], ldata_0n[6]);
  BUFF I28 (store_0n[7], ldata_0n[7]);
  BUFF I29 (store_0n[8], ldata_0n[8]);
  BUFF I30 (store_0n[9], ldata_0n[9]);
  BUFF I31 (store_1n[0], ldata_1n[0]);
  BUFF I32 (store_1n[1], ldata_1n[1]);
  BUFF I33 (store_1n[2], ldata_1n[2]);
  BUFF I34 (store_1n[3], ldata_1n[3]);
  BUFF I35 (store_1n[4], ldata_1n[4]);
  BUFF I36 (store_1n[5], ldata_1n[5]);
  BUFF I37 (store_1n[6], ldata_1n[6]);
  BUFF I38 (store_1n[7], ldata_1n[7]);
  BUFF I39 (store_1n[8], ldata_1n[8]);
  BUFF I40 (store_1n[9], ldata_1n[9]);
  C3 I41 (internal_0n[0], wack_0n[0], wack_0n[1], wack_0n[2]);
  C3 I42 (internal_0n[1], wack_0n[3], wack_0n[4], wack_0n[5]);
  C2 I43 (internal_0n[2], wack_0n[6], wack_0n[7]);
  C2 I44 (internal_0n[3], wack_0n[8], wack_0n[9]);
  C2 I45 (internal_0n[4], internal_0n[0], internal_0n[1]);
  C2 I46 (internal_0n[5], internal_0n[2], internal_0n[3]);
  C2 I47 (write_0a, internal_0n[4], internal_0n[5]);
  DRLATCH I48 (write_0r0d[0], write_0r1d[0], wack_0n[0], ldata_0n[0], ldata_1n[0]);
  DRLATCH I49 (write_0r0d[1], write_0r1d[1], wack_0n[1], ldata_0n[1], ldata_1n[1]);
  DRLATCH I50 (write_0r0d[2], write_0r1d[2], wack_0n[2], ldata_0n[2], ldata_1n[2]);
  DRLATCH I51 (write_0r0d[3], write_0r1d[3], wack_0n[3], ldata_0n[3], ldata_1n[3]);
  DRLATCH I52 (write_0r0d[4], write_0r1d[4], wack_0n[4], ldata_0n[4], ldata_1n[4]);
  DRLATCH I53 (write_0r0d[5], write_0r1d[5], wack_0n[5], ldata_0n[5], ldata_1n[5]);
  DRLATCH I54 (write_0r0d[6], write_0r1d[6], wack_0n[6], ldata_0n[6], ldata_1n[6]);
  DRLATCH I55 (write_0r0d[7], write_0r1d[7], wack_0n[7], ldata_0n[7], ldata_1n[7]);
  DRLATCH I56 (write_0r0d[8], write_0r1d[8], wack_0n[8], ldata_0n[8], ldata_1n[8]);
  DRLATCH I57 (write_0r0d[9], write_0r1d[9], wack_0n[9], ldata_0n[9], ldata_1n[9]);
endmodule

module BrzVariable_10_2_s19_0_2e_2e0_3b1_2e_2e9 (
  write_0r0d, write_0r1d, write_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d
);
  input [9:0] write_0r0d;
  input [9:0] write_0r1d;
  output write_0a;
  input read_0r;
  output read_0a0d;
  output read_0a1d;
  input read_1r;
  output [8:0] read_1a0d;
  output [8:0] read_1a1d;
  wire [5:0] internal_0n;
  wire [9:0] store_0n;
  wire [9:0] store_1n;
  wire [9:0] ldata_0n;
  wire [9:0] ldata_1n;
  wire [9:0] wack_0n;
  wire readReq_0n;
  wire readReq_1n;
  AND2 I0 (read_1a1d[0], store_1n[1], readReq_1n);
  AND2 I1 (read_1a1d[1], store_1n[2], readReq_1n);
  AND2 I2 (read_1a1d[2], store_1n[3], readReq_1n);
  AND2 I3 (read_1a1d[3], store_1n[4], readReq_1n);
  AND2 I4 (read_1a1d[4], store_1n[5], readReq_1n);
  AND2 I5 (read_1a1d[5], store_1n[6], readReq_1n);
  AND2 I6 (read_1a1d[6], store_1n[7], readReq_1n);
  AND2 I7 (read_1a1d[7], store_1n[8], readReq_1n);
  AND2 I8 (read_1a1d[8], store_1n[9], readReq_1n);
  AND2 I9 (read_1a0d[0], store_0n[1], readReq_1n);
  AND2 I10 (read_1a0d[1], store_0n[2], readReq_1n);
  AND2 I11 (read_1a0d[2], store_0n[3], readReq_1n);
  AND2 I12 (read_1a0d[3], store_0n[4], readReq_1n);
  AND2 I13 (read_1a0d[4], store_0n[5], readReq_1n);
  AND2 I14 (read_1a0d[5], store_0n[6], readReq_1n);
  AND2 I15 (read_1a0d[6], store_0n[7], readReq_1n);
  AND2 I16 (read_1a0d[7], store_0n[8], readReq_1n);
  AND2 I17 (read_1a0d[8], store_0n[9], readReq_1n);
  AND2 I18 (read_0a1d, store_1n[0], readReq_0n);
  AND2 I19 (read_0a0d, store_0n[0], readReq_0n);
  BUFF I20 (readReq_0n, read_0r);
  BUFF I21 (readReq_1n, read_1r);
  BUFF I22 (store_0n[0], ldata_0n[0]);
  BUFF I23 (store_0n[1], ldata_0n[1]);
  BUFF I24 (store_0n[2], ldata_0n[2]);
  BUFF I25 (store_0n[3], ldata_0n[3]);
  BUFF I26 (store_0n[4], ldata_0n[4]);
  BUFF I27 (store_0n[5], ldata_0n[5]);
  BUFF I28 (store_0n[6], ldata_0n[6]);
  BUFF I29 (store_0n[7], ldata_0n[7]);
  BUFF I30 (store_0n[8], ldata_0n[8]);
  BUFF I31 (store_0n[9], ldata_0n[9]);
  BUFF I32 (store_1n[0], ldata_1n[0]);
  BUFF I33 (store_1n[1], ldata_1n[1]);
  BUFF I34 (store_1n[2], ldata_1n[2]);
  BUFF I35 (store_1n[3], ldata_1n[3]);
  BUFF I36 (store_1n[4], ldata_1n[4]);
  BUFF I37 (store_1n[5], ldata_1n[5]);
  BUFF I38 (store_1n[6], ldata_1n[6]);
  BUFF I39 (store_1n[7], ldata_1n[7]);
  BUFF I40 (store_1n[8], ldata_1n[8]);
  BUFF I41 (store_1n[9], ldata_1n[9]);
  C3 I42 (internal_0n[0], wack_0n[0], wack_0n[1], wack_0n[2]);
  C3 I43 (internal_0n[1], wack_0n[3], wack_0n[4], wack_0n[5]);
  C2 I44 (internal_0n[2], wack_0n[6], wack_0n[7]);
  C2 I45 (internal_0n[3], wack_0n[8], wack_0n[9]);
  C2 I46 (internal_0n[4], internal_0n[0], internal_0n[1]);
  C2 I47 (internal_0n[5], internal_0n[2], internal_0n[3]);
  C2 I48 (write_0a, internal_0n[4], internal_0n[5]);
  DRLATCH I49 (write_0r0d[0], write_0r1d[0], wack_0n[0], ldata_0n[0], ldata_1n[0]);
  DRLATCH I50 (write_0r0d[1], write_0r1d[1], wack_0n[1], ldata_0n[1], ldata_1n[1]);
  DRLATCH I51 (write_0r0d[2], write_0r1d[2], wack_0n[2], ldata_0n[2], ldata_1n[2]);
  DRLATCH I52 (write_0r0d[3], write_0r1d[3], wack_0n[3], ldata_0n[3], ldata_1n[3]);
  DRLATCH I53 (write_0r0d[4], write_0r1d[4], wack_0n[4], ldata_0n[4], ldata_1n[4]);
  DRLATCH I54 (write_0r0d[5], write_0r1d[5], wack_0n[5], ldata_0n[5], ldata_1n[5]);
  DRLATCH I55 (write_0r0d[6], write_0r1d[6], wack_0n[6], ldata_0n[6], ldata_1n[6]);
  DRLATCH I56 (write_0r0d[7], write_0r1d[7], wack_0n[7], ldata_0n[7], ldata_1n[7]);
  DRLATCH I57 (write_0r0d[8], write_0r1d[8], wack_0n[8], ldata_0n[8], ldata_1n[8]);
  DRLATCH I58 (write_0r0d[9], write_0r1d[9], wack_0n[9], ldata_0n[9], ldata_1n[9]);
endmodule

module BrzVariable_32_2_s0_ (
  write_0r0d, write_0r1d, write_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d
);
  input [31:0] write_0r0d;
  input [31:0] write_0r1d;
  output write_0a;
  input read_0r;
  output [31:0] read_0a0d;
  output [31:0] read_0a1d;
  input read_1r;
  output [31:0] read_1a0d;
  output [31:0] read_1a1d;
  wire [16:0] internal_0n;
  wire [31:0] store_0n;
  wire [31:0] store_1n;
  wire [31:0] ldata_0n;
  wire [31:0] ldata_1n;
  wire [31:0] wack_0n;
  wire readReq_0n;
  wire readReq_1n;
  AND2 I0 (read_1a1d[0], store_1n[0], readReq_1n);
  AND2 I1 (read_1a1d[1], store_1n[1], readReq_1n);
  AND2 I2 (read_1a1d[2], store_1n[2], readReq_1n);
  AND2 I3 (read_1a1d[3], store_1n[3], readReq_1n);
  AND2 I4 (read_1a1d[4], store_1n[4], readReq_1n);
  AND2 I5 (read_1a1d[5], store_1n[5], readReq_1n);
  AND2 I6 (read_1a1d[6], store_1n[6], readReq_1n);
  AND2 I7 (read_1a1d[7], store_1n[7], readReq_1n);
  AND2 I8 (read_1a1d[8], store_1n[8], readReq_1n);
  AND2 I9 (read_1a1d[9], store_1n[9], readReq_1n);
  AND2 I10 (read_1a1d[10], store_1n[10], readReq_1n);
  AND2 I11 (read_1a1d[11], store_1n[11], readReq_1n);
  AND2 I12 (read_1a1d[12], store_1n[12], readReq_1n);
  AND2 I13 (read_1a1d[13], store_1n[13], readReq_1n);
  AND2 I14 (read_1a1d[14], store_1n[14], readReq_1n);
  AND2 I15 (read_1a1d[15], store_1n[15], readReq_1n);
  AND2 I16 (read_1a1d[16], store_1n[16], readReq_1n);
  AND2 I17 (read_1a1d[17], store_1n[17], readReq_1n);
  AND2 I18 (read_1a1d[18], store_1n[18], readReq_1n);
  AND2 I19 (read_1a1d[19], store_1n[19], readReq_1n);
  AND2 I20 (read_1a1d[20], store_1n[20], readReq_1n);
  AND2 I21 (read_1a1d[21], store_1n[21], readReq_1n);
  AND2 I22 (read_1a1d[22], store_1n[22], readReq_1n);
  AND2 I23 (read_1a1d[23], store_1n[23], readReq_1n);
  AND2 I24 (read_1a1d[24], store_1n[24], readReq_1n);
  AND2 I25 (read_1a1d[25], store_1n[25], readReq_1n);
  AND2 I26 (read_1a1d[26], store_1n[26], readReq_1n);
  AND2 I27 (read_1a1d[27], store_1n[27], readReq_1n);
  AND2 I28 (read_1a1d[28], store_1n[28], readReq_1n);
  AND2 I29 (read_1a1d[29], store_1n[29], readReq_1n);
  AND2 I30 (read_1a1d[30], store_1n[30], readReq_1n);
  AND2 I31 (read_1a1d[31], store_1n[31], readReq_1n);
  AND2 I32 (read_1a0d[0], store_0n[0], readReq_1n);
  AND2 I33 (read_1a0d[1], store_0n[1], readReq_1n);
  AND2 I34 (read_1a0d[2], store_0n[2], readReq_1n);
  AND2 I35 (read_1a0d[3], store_0n[3], readReq_1n);
  AND2 I36 (read_1a0d[4], store_0n[4], readReq_1n);
  AND2 I37 (read_1a0d[5], store_0n[5], readReq_1n);
  AND2 I38 (read_1a0d[6], store_0n[6], readReq_1n);
  AND2 I39 (read_1a0d[7], store_0n[7], readReq_1n);
  AND2 I40 (read_1a0d[8], store_0n[8], readReq_1n);
  AND2 I41 (read_1a0d[9], store_0n[9], readReq_1n);
  AND2 I42 (read_1a0d[10], store_0n[10], readReq_1n);
  AND2 I43 (read_1a0d[11], store_0n[11], readReq_1n);
  AND2 I44 (read_1a0d[12], store_0n[12], readReq_1n);
  AND2 I45 (read_1a0d[13], store_0n[13], readReq_1n);
  AND2 I46 (read_1a0d[14], store_0n[14], readReq_1n);
  AND2 I47 (read_1a0d[15], store_0n[15], readReq_1n);
  AND2 I48 (read_1a0d[16], store_0n[16], readReq_1n);
  AND2 I49 (read_1a0d[17], store_0n[17], readReq_1n);
  AND2 I50 (read_1a0d[18], store_0n[18], readReq_1n);
  AND2 I51 (read_1a0d[19], store_0n[19], readReq_1n);
  AND2 I52 (read_1a0d[20], store_0n[20], readReq_1n);
  AND2 I53 (read_1a0d[21], store_0n[21], readReq_1n);
  AND2 I54 (read_1a0d[22], store_0n[22], readReq_1n);
  AND2 I55 (read_1a0d[23], store_0n[23], readReq_1n);
  AND2 I56 (read_1a0d[24], store_0n[24], readReq_1n);
  AND2 I57 (read_1a0d[25], store_0n[25], readReq_1n);
  AND2 I58 (read_1a0d[26], store_0n[26], readReq_1n);
  AND2 I59 (read_1a0d[27], store_0n[27], readReq_1n);
  AND2 I60 (read_1a0d[28], store_0n[28], readReq_1n);
  AND2 I61 (read_1a0d[29], store_0n[29], readReq_1n);
  AND2 I62 (read_1a0d[30], store_0n[30], readReq_1n);
  AND2 I63 (read_1a0d[31], store_0n[31], readReq_1n);
  AND2 I64 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I65 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I66 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I67 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I68 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I69 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I70 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I71 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I72 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I73 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I74 (read_0a1d[10], store_1n[10], readReq_0n);
  AND2 I75 (read_0a1d[11], store_1n[11], readReq_0n);
  AND2 I76 (read_0a1d[12], store_1n[12], readReq_0n);
  AND2 I77 (read_0a1d[13], store_1n[13], readReq_0n);
  AND2 I78 (read_0a1d[14], store_1n[14], readReq_0n);
  AND2 I79 (read_0a1d[15], store_1n[15], readReq_0n);
  AND2 I80 (read_0a1d[16], store_1n[16], readReq_0n);
  AND2 I81 (read_0a1d[17], store_1n[17], readReq_0n);
  AND2 I82 (read_0a1d[18], store_1n[18], readReq_0n);
  AND2 I83 (read_0a1d[19], store_1n[19], readReq_0n);
  AND2 I84 (read_0a1d[20], store_1n[20], readReq_0n);
  AND2 I85 (read_0a1d[21], store_1n[21], readReq_0n);
  AND2 I86 (read_0a1d[22], store_1n[22], readReq_0n);
  AND2 I87 (read_0a1d[23], store_1n[23], readReq_0n);
  AND2 I88 (read_0a1d[24], store_1n[24], readReq_0n);
  AND2 I89 (read_0a1d[25], store_1n[25], readReq_0n);
  AND2 I90 (read_0a1d[26], store_1n[26], readReq_0n);
  AND2 I91 (read_0a1d[27], store_1n[27], readReq_0n);
  AND2 I92 (read_0a1d[28], store_1n[28], readReq_0n);
  AND2 I93 (read_0a1d[29], store_1n[29], readReq_0n);
  AND2 I94 (read_0a1d[30], store_1n[30], readReq_0n);
  AND2 I95 (read_0a1d[31], store_1n[31], readReq_0n);
  AND2 I96 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I97 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I98 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I99 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I100 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I101 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I102 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I103 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I104 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I105 (read_0a0d[9], store_0n[9], readReq_0n);
  AND2 I106 (read_0a0d[10], store_0n[10], readReq_0n);
  AND2 I107 (read_0a0d[11], store_0n[11], readReq_0n);
  AND2 I108 (read_0a0d[12], store_0n[12], readReq_0n);
  AND2 I109 (read_0a0d[13], store_0n[13], readReq_0n);
  AND2 I110 (read_0a0d[14], store_0n[14], readReq_0n);
  AND2 I111 (read_0a0d[15], store_0n[15], readReq_0n);
  AND2 I112 (read_0a0d[16], store_0n[16], readReq_0n);
  AND2 I113 (read_0a0d[17], store_0n[17], readReq_0n);
  AND2 I114 (read_0a0d[18], store_0n[18], readReq_0n);
  AND2 I115 (read_0a0d[19], store_0n[19], readReq_0n);
  AND2 I116 (read_0a0d[20], store_0n[20], readReq_0n);
  AND2 I117 (read_0a0d[21], store_0n[21], readReq_0n);
  AND2 I118 (read_0a0d[22], store_0n[22], readReq_0n);
  AND2 I119 (read_0a0d[23], store_0n[23], readReq_0n);
  AND2 I120 (read_0a0d[24], store_0n[24], readReq_0n);
  AND2 I121 (read_0a0d[25], store_0n[25], readReq_0n);
  AND2 I122 (read_0a0d[26], store_0n[26], readReq_0n);
  AND2 I123 (read_0a0d[27], store_0n[27], readReq_0n);
  AND2 I124 (read_0a0d[28], store_0n[28], readReq_0n);
  AND2 I125 (read_0a0d[29], store_0n[29], readReq_0n);
  AND2 I126 (read_0a0d[30], store_0n[30], readReq_0n);
  AND2 I127 (read_0a0d[31], store_0n[31], readReq_0n);
  BUFF I128 (readReq_0n, read_0r);
  BUFF I129 (readReq_1n, read_1r);
  BUFF I130 (store_0n[0], ldata_0n[0]);
  BUFF I131 (store_0n[1], ldata_0n[1]);
  BUFF I132 (store_0n[2], ldata_0n[2]);
  BUFF I133 (store_0n[3], ldata_0n[3]);
  BUFF I134 (store_0n[4], ldata_0n[4]);
  BUFF I135 (store_0n[5], ldata_0n[5]);
  BUFF I136 (store_0n[6], ldata_0n[6]);
  BUFF I137 (store_0n[7], ldata_0n[7]);
  BUFF I138 (store_0n[8], ldata_0n[8]);
  BUFF I139 (store_0n[9], ldata_0n[9]);
  BUFF I140 (store_0n[10], ldata_0n[10]);
  BUFF I141 (store_0n[11], ldata_0n[11]);
  BUFF I142 (store_0n[12], ldata_0n[12]);
  BUFF I143 (store_0n[13], ldata_0n[13]);
  BUFF I144 (store_0n[14], ldata_0n[14]);
  BUFF I145 (store_0n[15], ldata_0n[15]);
  BUFF I146 (store_0n[16], ldata_0n[16]);
  BUFF I147 (store_0n[17], ldata_0n[17]);
  BUFF I148 (store_0n[18], ldata_0n[18]);
  BUFF I149 (store_0n[19], ldata_0n[19]);
  BUFF I150 (store_0n[20], ldata_0n[20]);
  BUFF I151 (store_0n[21], ldata_0n[21]);
  BUFF I152 (store_0n[22], ldata_0n[22]);
  BUFF I153 (store_0n[23], ldata_0n[23]);
  BUFF I154 (store_0n[24], ldata_0n[24]);
  BUFF I155 (store_0n[25], ldata_0n[25]);
  BUFF I156 (store_0n[26], ldata_0n[26]);
  BUFF I157 (store_0n[27], ldata_0n[27]);
  BUFF I158 (store_0n[28], ldata_0n[28]);
  BUFF I159 (store_0n[29], ldata_0n[29]);
  BUFF I160 (store_0n[30], ldata_0n[30]);
  BUFF I161 (store_0n[31], ldata_0n[31]);
  BUFF I162 (store_1n[0], ldata_1n[0]);
  BUFF I163 (store_1n[1], ldata_1n[1]);
  BUFF I164 (store_1n[2], ldata_1n[2]);
  BUFF I165 (store_1n[3], ldata_1n[3]);
  BUFF I166 (store_1n[4], ldata_1n[4]);
  BUFF I167 (store_1n[5], ldata_1n[5]);
  BUFF I168 (store_1n[6], ldata_1n[6]);
  BUFF I169 (store_1n[7], ldata_1n[7]);
  BUFF I170 (store_1n[8], ldata_1n[8]);
  BUFF I171 (store_1n[9], ldata_1n[9]);
  BUFF I172 (store_1n[10], ldata_1n[10]);
  BUFF I173 (store_1n[11], ldata_1n[11]);
  BUFF I174 (store_1n[12], ldata_1n[12]);
  BUFF I175 (store_1n[13], ldata_1n[13]);
  BUFF I176 (store_1n[14], ldata_1n[14]);
  BUFF I177 (store_1n[15], ldata_1n[15]);
  BUFF I178 (store_1n[16], ldata_1n[16]);
  BUFF I179 (store_1n[17], ldata_1n[17]);
  BUFF I180 (store_1n[18], ldata_1n[18]);
  BUFF I181 (store_1n[19], ldata_1n[19]);
  BUFF I182 (store_1n[20], ldata_1n[20]);
  BUFF I183 (store_1n[21], ldata_1n[21]);
  BUFF I184 (store_1n[22], ldata_1n[22]);
  BUFF I185 (store_1n[23], ldata_1n[23]);
  BUFF I186 (store_1n[24], ldata_1n[24]);
  BUFF I187 (store_1n[25], ldata_1n[25]);
  BUFF I188 (store_1n[26], ldata_1n[26]);
  BUFF I189 (store_1n[27], ldata_1n[27]);
  BUFF I190 (store_1n[28], ldata_1n[28]);
  BUFF I191 (store_1n[29], ldata_1n[29]);
  BUFF I192 (store_1n[30], ldata_1n[30]);
  BUFF I193 (store_1n[31], ldata_1n[31]);
  C3 I194 (internal_0n[0], wack_0n[0], wack_0n[1], wack_0n[2]);
  C3 I195 (internal_0n[1], wack_0n[3], wack_0n[4], wack_0n[5]);
  C3 I196 (internal_0n[2], wack_0n[6], wack_0n[7], wack_0n[8]);
  C3 I197 (internal_0n[3], wack_0n[9], wack_0n[10], wack_0n[11]);
  C3 I198 (internal_0n[4], wack_0n[12], wack_0n[13], wack_0n[14]);
  C3 I199 (internal_0n[5], wack_0n[15], wack_0n[16], wack_0n[17]);
  C3 I200 (internal_0n[6], wack_0n[18], wack_0n[19], wack_0n[20]);
  C3 I201 (internal_0n[7], wack_0n[21], wack_0n[22], wack_0n[23]);
  C3 I202 (internal_0n[8], wack_0n[24], wack_0n[25], wack_0n[26]);
  C3 I203 (internal_0n[9], wack_0n[27], wack_0n[28], wack_0n[29]);
  C2 I204 (internal_0n[10], wack_0n[30], wack_0n[31]);
  C3 I205 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I206 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I207 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I208 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I209 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I210 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I211 (write_0a, internal_0n[15], internal_0n[16]);
  DRLATCH I212 (write_0r0d[0], write_0r1d[0], wack_0n[0], ldata_0n[0], ldata_1n[0]);
  DRLATCH I213 (write_0r0d[1], write_0r1d[1], wack_0n[1], ldata_0n[1], ldata_1n[1]);
  DRLATCH I214 (write_0r0d[2], write_0r1d[2], wack_0n[2], ldata_0n[2], ldata_1n[2]);
  DRLATCH I215 (write_0r0d[3], write_0r1d[3], wack_0n[3], ldata_0n[3], ldata_1n[3]);
  DRLATCH I216 (write_0r0d[4], write_0r1d[4], wack_0n[4], ldata_0n[4], ldata_1n[4]);
  DRLATCH I217 (write_0r0d[5], write_0r1d[5], wack_0n[5], ldata_0n[5], ldata_1n[5]);
  DRLATCH I218 (write_0r0d[6], write_0r1d[6], wack_0n[6], ldata_0n[6], ldata_1n[6]);
  DRLATCH I219 (write_0r0d[7], write_0r1d[7], wack_0n[7], ldata_0n[7], ldata_1n[7]);
  DRLATCH I220 (write_0r0d[8], write_0r1d[8], wack_0n[8], ldata_0n[8], ldata_1n[8]);
  DRLATCH I221 (write_0r0d[9], write_0r1d[9], wack_0n[9], ldata_0n[9], ldata_1n[9]);
  DRLATCH I222 (write_0r0d[10], write_0r1d[10], wack_0n[10], ldata_0n[10], ldata_1n[10]);
  DRLATCH I223 (write_0r0d[11], write_0r1d[11], wack_0n[11], ldata_0n[11], ldata_1n[11]);
  DRLATCH I224 (write_0r0d[12], write_0r1d[12], wack_0n[12], ldata_0n[12], ldata_1n[12]);
  DRLATCH I225 (write_0r0d[13], write_0r1d[13], wack_0n[13], ldata_0n[13], ldata_1n[13]);
  DRLATCH I226 (write_0r0d[14], write_0r1d[14], wack_0n[14], ldata_0n[14], ldata_1n[14]);
  DRLATCH I227 (write_0r0d[15], write_0r1d[15], wack_0n[15], ldata_0n[15], ldata_1n[15]);
  DRLATCH I228 (write_0r0d[16], write_0r1d[16], wack_0n[16], ldata_0n[16], ldata_1n[16]);
  DRLATCH I229 (write_0r0d[17], write_0r1d[17], wack_0n[17], ldata_0n[17], ldata_1n[17]);
  DRLATCH I230 (write_0r0d[18], write_0r1d[18], wack_0n[18], ldata_0n[18], ldata_1n[18]);
  DRLATCH I231 (write_0r0d[19], write_0r1d[19], wack_0n[19], ldata_0n[19], ldata_1n[19]);
  DRLATCH I232 (write_0r0d[20], write_0r1d[20], wack_0n[20], ldata_0n[20], ldata_1n[20]);
  DRLATCH I233 (write_0r0d[21], write_0r1d[21], wack_0n[21], ldata_0n[21], ldata_1n[21]);
  DRLATCH I234 (write_0r0d[22], write_0r1d[22], wack_0n[22], ldata_0n[22], ldata_1n[22]);
  DRLATCH I235 (write_0r0d[23], write_0r1d[23], wack_0n[23], ldata_0n[23], ldata_1n[23]);
  DRLATCH I236 (write_0r0d[24], write_0r1d[24], wack_0n[24], ldata_0n[24], ldata_1n[24]);
  DRLATCH I237 (write_0r0d[25], write_0r1d[25], wack_0n[25], ldata_0n[25], ldata_1n[25]);
  DRLATCH I238 (write_0r0d[26], write_0r1d[26], wack_0n[26], ldata_0n[26], ldata_1n[26]);
  DRLATCH I239 (write_0r0d[27], write_0r1d[27], wack_0n[27], ldata_0n[27], ldata_1n[27]);
  DRLATCH I240 (write_0r0d[28], write_0r1d[28], wack_0n[28], ldata_0n[28], ldata_1n[28]);
  DRLATCH I241 (write_0r0d[29], write_0r1d[29], wack_0n[29], ldata_0n[29], ldata_1n[29]);
  DRLATCH I242 (write_0r0d[30], write_0r1d[30], wack_0n[30], ldata_0n[30], ldata_1n[30]);
  DRLATCH I243 (write_0r0d[31], write_0r1d[31], wack_0n[31], ldata_0n[31], ldata_1n[31]);
endmodule

module BrzVariable_32_3_s16__3b_3b31_2e_2e31 (
  write_0r0d, write_0r1d, write_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d,
  read_2r, read_2a0d, read_2a1d
);
  input [31:0] write_0r0d;
  input [31:0] write_0r1d;
  output write_0a;
  input read_0r;
  output [31:0] read_0a0d;
  output [31:0] read_0a1d;
  input read_1r;
  output [31:0] read_1a0d;
  output [31:0] read_1a1d;
  input read_2r;
  output read_2a0d;
  output read_2a1d;
  wire [16:0] internal_0n;
  wire [31:0] store_0n;
  wire [31:0] store_1n;
  wire [31:0] ldata_0n;
  wire [31:0] ldata_1n;
  wire [31:0] wack_0n;
  wire readReq_0n;
  wire readReq_1n;
  wire readReq_2n;
  AND2 I0 (read_2a1d, store_1n[31], readReq_2n);
  AND2 I1 (read_2a0d, store_0n[31], readReq_2n);
  AND2 I2 (read_1a1d[0], store_1n[0], readReq_1n);
  AND2 I3 (read_1a1d[1], store_1n[1], readReq_1n);
  AND2 I4 (read_1a1d[2], store_1n[2], readReq_1n);
  AND2 I5 (read_1a1d[3], store_1n[3], readReq_1n);
  AND2 I6 (read_1a1d[4], store_1n[4], readReq_1n);
  AND2 I7 (read_1a1d[5], store_1n[5], readReq_1n);
  AND2 I8 (read_1a1d[6], store_1n[6], readReq_1n);
  AND2 I9 (read_1a1d[7], store_1n[7], readReq_1n);
  AND2 I10 (read_1a1d[8], store_1n[8], readReq_1n);
  AND2 I11 (read_1a1d[9], store_1n[9], readReq_1n);
  AND2 I12 (read_1a1d[10], store_1n[10], readReq_1n);
  AND2 I13 (read_1a1d[11], store_1n[11], readReq_1n);
  AND2 I14 (read_1a1d[12], store_1n[12], readReq_1n);
  AND2 I15 (read_1a1d[13], store_1n[13], readReq_1n);
  AND2 I16 (read_1a1d[14], store_1n[14], readReq_1n);
  AND2 I17 (read_1a1d[15], store_1n[15], readReq_1n);
  AND2 I18 (read_1a1d[16], store_1n[16], readReq_1n);
  AND2 I19 (read_1a1d[17], store_1n[17], readReq_1n);
  AND2 I20 (read_1a1d[18], store_1n[18], readReq_1n);
  AND2 I21 (read_1a1d[19], store_1n[19], readReq_1n);
  AND2 I22 (read_1a1d[20], store_1n[20], readReq_1n);
  AND2 I23 (read_1a1d[21], store_1n[21], readReq_1n);
  AND2 I24 (read_1a1d[22], store_1n[22], readReq_1n);
  AND2 I25 (read_1a1d[23], store_1n[23], readReq_1n);
  AND2 I26 (read_1a1d[24], store_1n[24], readReq_1n);
  AND2 I27 (read_1a1d[25], store_1n[25], readReq_1n);
  AND2 I28 (read_1a1d[26], store_1n[26], readReq_1n);
  AND2 I29 (read_1a1d[27], store_1n[27], readReq_1n);
  AND2 I30 (read_1a1d[28], store_1n[28], readReq_1n);
  AND2 I31 (read_1a1d[29], store_1n[29], readReq_1n);
  AND2 I32 (read_1a1d[30], store_1n[30], readReq_1n);
  AND2 I33 (read_1a1d[31], store_1n[31], readReq_1n);
  AND2 I34 (read_1a0d[0], store_0n[0], readReq_1n);
  AND2 I35 (read_1a0d[1], store_0n[1], readReq_1n);
  AND2 I36 (read_1a0d[2], store_0n[2], readReq_1n);
  AND2 I37 (read_1a0d[3], store_0n[3], readReq_1n);
  AND2 I38 (read_1a0d[4], store_0n[4], readReq_1n);
  AND2 I39 (read_1a0d[5], store_0n[5], readReq_1n);
  AND2 I40 (read_1a0d[6], store_0n[6], readReq_1n);
  AND2 I41 (read_1a0d[7], store_0n[7], readReq_1n);
  AND2 I42 (read_1a0d[8], store_0n[8], readReq_1n);
  AND2 I43 (read_1a0d[9], store_0n[9], readReq_1n);
  AND2 I44 (read_1a0d[10], store_0n[10], readReq_1n);
  AND2 I45 (read_1a0d[11], store_0n[11], readReq_1n);
  AND2 I46 (read_1a0d[12], store_0n[12], readReq_1n);
  AND2 I47 (read_1a0d[13], store_0n[13], readReq_1n);
  AND2 I48 (read_1a0d[14], store_0n[14], readReq_1n);
  AND2 I49 (read_1a0d[15], store_0n[15], readReq_1n);
  AND2 I50 (read_1a0d[16], store_0n[16], readReq_1n);
  AND2 I51 (read_1a0d[17], store_0n[17], readReq_1n);
  AND2 I52 (read_1a0d[18], store_0n[18], readReq_1n);
  AND2 I53 (read_1a0d[19], store_0n[19], readReq_1n);
  AND2 I54 (read_1a0d[20], store_0n[20], readReq_1n);
  AND2 I55 (read_1a0d[21], store_0n[21], readReq_1n);
  AND2 I56 (read_1a0d[22], store_0n[22], readReq_1n);
  AND2 I57 (read_1a0d[23], store_0n[23], readReq_1n);
  AND2 I58 (read_1a0d[24], store_0n[24], readReq_1n);
  AND2 I59 (read_1a0d[25], store_0n[25], readReq_1n);
  AND2 I60 (read_1a0d[26], store_0n[26], readReq_1n);
  AND2 I61 (read_1a0d[27], store_0n[27], readReq_1n);
  AND2 I62 (read_1a0d[28], store_0n[28], readReq_1n);
  AND2 I63 (read_1a0d[29], store_0n[29], readReq_1n);
  AND2 I64 (read_1a0d[30], store_0n[30], readReq_1n);
  AND2 I65 (read_1a0d[31], store_0n[31], readReq_1n);
  AND2 I66 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I67 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I68 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I69 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I70 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I71 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I72 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I73 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I74 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I75 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I76 (read_0a1d[10], store_1n[10], readReq_0n);
  AND2 I77 (read_0a1d[11], store_1n[11], readReq_0n);
  AND2 I78 (read_0a1d[12], store_1n[12], readReq_0n);
  AND2 I79 (read_0a1d[13], store_1n[13], readReq_0n);
  AND2 I80 (read_0a1d[14], store_1n[14], readReq_0n);
  AND2 I81 (read_0a1d[15], store_1n[15], readReq_0n);
  AND2 I82 (read_0a1d[16], store_1n[16], readReq_0n);
  AND2 I83 (read_0a1d[17], store_1n[17], readReq_0n);
  AND2 I84 (read_0a1d[18], store_1n[18], readReq_0n);
  AND2 I85 (read_0a1d[19], store_1n[19], readReq_0n);
  AND2 I86 (read_0a1d[20], store_1n[20], readReq_0n);
  AND2 I87 (read_0a1d[21], store_1n[21], readReq_0n);
  AND2 I88 (read_0a1d[22], store_1n[22], readReq_0n);
  AND2 I89 (read_0a1d[23], store_1n[23], readReq_0n);
  AND2 I90 (read_0a1d[24], store_1n[24], readReq_0n);
  AND2 I91 (read_0a1d[25], store_1n[25], readReq_0n);
  AND2 I92 (read_0a1d[26], store_1n[26], readReq_0n);
  AND2 I93 (read_0a1d[27], store_1n[27], readReq_0n);
  AND2 I94 (read_0a1d[28], store_1n[28], readReq_0n);
  AND2 I95 (read_0a1d[29], store_1n[29], readReq_0n);
  AND2 I96 (read_0a1d[30], store_1n[30], readReq_0n);
  AND2 I97 (read_0a1d[31], store_1n[31], readReq_0n);
  AND2 I98 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I99 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I100 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I101 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I102 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I103 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I104 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I105 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I106 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I107 (read_0a0d[9], store_0n[9], readReq_0n);
  AND2 I108 (read_0a0d[10], store_0n[10], readReq_0n);
  AND2 I109 (read_0a0d[11], store_0n[11], readReq_0n);
  AND2 I110 (read_0a0d[12], store_0n[12], readReq_0n);
  AND2 I111 (read_0a0d[13], store_0n[13], readReq_0n);
  AND2 I112 (read_0a0d[14], store_0n[14], readReq_0n);
  AND2 I113 (read_0a0d[15], store_0n[15], readReq_0n);
  AND2 I114 (read_0a0d[16], store_0n[16], readReq_0n);
  AND2 I115 (read_0a0d[17], store_0n[17], readReq_0n);
  AND2 I116 (read_0a0d[18], store_0n[18], readReq_0n);
  AND2 I117 (read_0a0d[19], store_0n[19], readReq_0n);
  AND2 I118 (read_0a0d[20], store_0n[20], readReq_0n);
  AND2 I119 (read_0a0d[21], store_0n[21], readReq_0n);
  AND2 I120 (read_0a0d[22], store_0n[22], readReq_0n);
  AND2 I121 (read_0a0d[23], store_0n[23], readReq_0n);
  AND2 I122 (read_0a0d[24], store_0n[24], readReq_0n);
  AND2 I123 (read_0a0d[25], store_0n[25], readReq_0n);
  AND2 I124 (read_0a0d[26], store_0n[26], readReq_0n);
  AND2 I125 (read_0a0d[27], store_0n[27], readReq_0n);
  AND2 I126 (read_0a0d[28], store_0n[28], readReq_0n);
  AND2 I127 (read_0a0d[29], store_0n[29], readReq_0n);
  AND2 I128 (read_0a0d[30], store_0n[30], readReq_0n);
  AND2 I129 (read_0a0d[31], store_0n[31], readReq_0n);
  BUFF I130 (readReq_0n, read_0r);
  BUFF I131 (readReq_1n, read_1r);
  BUFF I132 (readReq_2n, read_2r);
  BUFF I133 (store_0n[0], ldata_0n[0]);
  BUFF I134 (store_0n[1], ldata_0n[1]);
  BUFF I135 (store_0n[2], ldata_0n[2]);
  BUFF I136 (store_0n[3], ldata_0n[3]);
  BUFF I137 (store_0n[4], ldata_0n[4]);
  BUFF I138 (store_0n[5], ldata_0n[5]);
  BUFF I139 (store_0n[6], ldata_0n[6]);
  BUFF I140 (store_0n[7], ldata_0n[7]);
  BUFF I141 (store_0n[8], ldata_0n[8]);
  BUFF I142 (store_0n[9], ldata_0n[9]);
  BUFF I143 (store_0n[10], ldata_0n[10]);
  BUFF I144 (store_0n[11], ldata_0n[11]);
  BUFF I145 (store_0n[12], ldata_0n[12]);
  BUFF I146 (store_0n[13], ldata_0n[13]);
  BUFF I147 (store_0n[14], ldata_0n[14]);
  BUFF I148 (store_0n[15], ldata_0n[15]);
  BUFF I149 (store_0n[16], ldata_0n[16]);
  BUFF I150 (store_0n[17], ldata_0n[17]);
  BUFF I151 (store_0n[18], ldata_0n[18]);
  BUFF I152 (store_0n[19], ldata_0n[19]);
  BUFF I153 (store_0n[20], ldata_0n[20]);
  BUFF I154 (store_0n[21], ldata_0n[21]);
  BUFF I155 (store_0n[22], ldata_0n[22]);
  BUFF I156 (store_0n[23], ldata_0n[23]);
  BUFF I157 (store_0n[24], ldata_0n[24]);
  BUFF I158 (store_0n[25], ldata_0n[25]);
  BUFF I159 (store_0n[26], ldata_0n[26]);
  BUFF I160 (store_0n[27], ldata_0n[27]);
  BUFF I161 (store_0n[28], ldata_0n[28]);
  BUFF I162 (store_0n[29], ldata_0n[29]);
  BUFF I163 (store_0n[30], ldata_0n[30]);
  BUFF I164 (store_0n[31], ldata_0n[31]);
  BUFF I165 (store_1n[0], ldata_1n[0]);
  BUFF I166 (store_1n[1], ldata_1n[1]);
  BUFF I167 (store_1n[2], ldata_1n[2]);
  BUFF I168 (store_1n[3], ldata_1n[3]);
  BUFF I169 (store_1n[4], ldata_1n[4]);
  BUFF I170 (store_1n[5], ldata_1n[5]);
  BUFF I171 (store_1n[6], ldata_1n[6]);
  BUFF I172 (store_1n[7], ldata_1n[7]);
  BUFF I173 (store_1n[8], ldata_1n[8]);
  BUFF I174 (store_1n[9], ldata_1n[9]);
  BUFF I175 (store_1n[10], ldata_1n[10]);
  BUFF I176 (store_1n[11], ldata_1n[11]);
  BUFF I177 (store_1n[12], ldata_1n[12]);
  BUFF I178 (store_1n[13], ldata_1n[13]);
  BUFF I179 (store_1n[14], ldata_1n[14]);
  BUFF I180 (store_1n[15], ldata_1n[15]);
  BUFF I181 (store_1n[16], ldata_1n[16]);
  BUFF I182 (store_1n[17], ldata_1n[17]);
  BUFF I183 (store_1n[18], ldata_1n[18]);
  BUFF I184 (store_1n[19], ldata_1n[19]);
  BUFF I185 (store_1n[20], ldata_1n[20]);
  BUFF I186 (store_1n[21], ldata_1n[21]);
  BUFF I187 (store_1n[22], ldata_1n[22]);
  BUFF I188 (store_1n[23], ldata_1n[23]);
  BUFF I189 (store_1n[24], ldata_1n[24]);
  BUFF I190 (store_1n[25], ldata_1n[25]);
  BUFF I191 (store_1n[26], ldata_1n[26]);
  BUFF I192 (store_1n[27], ldata_1n[27]);
  BUFF I193 (store_1n[28], ldata_1n[28]);
  BUFF I194 (store_1n[29], ldata_1n[29]);
  BUFF I195 (store_1n[30], ldata_1n[30]);
  BUFF I196 (store_1n[31], ldata_1n[31]);
  C3 I197 (internal_0n[0], wack_0n[0], wack_0n[1], wack_0n[2]);
  C3 I198 (internal_0n[1], wack_0n[3], wack_0n[4], wack_0n[5]);
  C3 I199 (internal_0n[2], wack_0n[6], wack_0n[7], wack_0n[8]);
  C3 I200 (internal_0n[3], wack_0n[9], wack_0n[10], wack_0n[11]);
  C3 I201 (internal_0n[4], wack_0n[12], wack_0n[13], wack_0n[14]);
  C3 I202 (internal_0n[5], wack_0n[15], wack_0n[16], wack_0n[17]);
  C3 I203 (internal_0n[6], wack_0n[18], wack_0n[19], wack_0n[20]);
  C3 I204 (internal_0n[7], wack_0n[21], wack_0n[22], wack_0n[23]);
  C3 I205 (internal_0n[8], wack_0n[24], wack_0n[25], wack_0n[26]);
  C3 I206 (internal_0n[9], wack_0n[27], wack_0n[28], wack_0n[29]);
  C2 I207 (internal_0n[10], wack_0n[30], wack_0n[31]);
  C3 I208 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I209 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I210 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I211 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I212 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I213 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I214 (write_0a, internal_0n[15], internal_0n[16]);
  DRLATCH I215 (write_0r0d[0], write_0r1d[0], wack_0n[0], ldata_0n[0], ldata_1n[0]);
  DRLATCH I216 (write_0r0d[1], write_0r1d[1], wack_0n[1], ldata_0n[1], ldata_1n[1]);
  DRLATCH I217 (write_0r0d[2], write_0r1d[2], wack_0n[2], ldata_0n[2], ldata_1n[2]);
  DRLATCH I218 (write_0r0d[3], write_0r1d[3], wack_0n[3], ldata_0n[3], ldata_1n[3]);
  DRLATCH I219 (write_0r0d[4], write_0r1d[4], wack_0n[4], ldata_0n[4], ldata_1n[4]);
  DRLATCH I220 (write_0r0d[5], write_0r1d[5], wack_0n[5], ldata_0n[5], ldata_1n[5]);
  DRLATCH I221 (write_0r0d[6], write_0r1d[6], wack_0n[6], ldata_0n[6], ldata_1n[6]);
  DRLATCH I222 (write_0r0d[7], write_0r1d[7], wack_0n[7], ldata_0n[7], ldata_1n[7]);
  DRLATCH I223 (write_0r0d[8], write_0r1d[8], wack_0n[8], ldata_0n[8], ldata_1n[8]);
  DRLATCH I224 (write_0r0d[9], write_0r1d[9], wack_0n[9], ldata_0n[9], ldata_1n[9]);
  DRLATCH I225 (write_0r0d[10], write_0r1d[10], wack_0n[10], ldata_0n[10], ldata_1n[10]);
  DRLATCH I226 (write_0r0d[11], write_0r1d[11], wack_0n[11], ldata_0n[11], ldata_1n[11]);
  DRLATCH I227 (write_0r0d[12], write_0r1d[12], wack_0n[12], ldata_0n[12], ldata_1n[12]);
  DRLATCH I228 (write_0r0d[13], write_0r1d[13], wack_0n[13], ldata_0n[13], ldata_1n[13]);
  DRLATCH I229 (write_0r0d[14], write_0r1d[14], wack_0n[14], ldata_0n[14], ldata_1n[14]);
  DRLATCH I230 (write_0r0d[15], write_0r1d[15], wack_0n[15], ldata_0n[15], ldata_1n[15]);
  DRLATCH I231 (write_0r0d[16], write_0r1d[16], wack_0n[16], ldata_0n[16], ldata_1n[16]);
  DRLATCH I232 (write_0r0d[17], write_0r1d[17], wack_0n[17], ldata_0n[17], ldata_1n[17]);
  DRLATCH I233 (write_0r0d[18], write_0r1d[18], wack_0n[18], ldata_0n[18], ldata_1n[18]);
  DRLATCH I234 (write_0r0d[19], write_0r1d[19], wack_0n[19], ldata_0n[19], ldata_1n[19]);
  DRLATCH I235 (write_0r0d[20], write_0r1d[20], wack_0n[20], ldata_0n[20], ldata_1n[20]);
  DRLATCH I236 (write_0r0d[21], write_0r1d[21], wack_0n[21], ldata_0n[21], ldata_1n[21]);
  DRLATCH I237 (write_0r0d[22], write_0r1d[22], wack_0n[22], ldata_0n[22], ldata_1n[22]);
  DRLATCH I238 (write_0r0d[23], write_0r1d[23], wack_0n[23], ldata_0n[23], ldata_1n[23]);
  DRLATCH I239 (write_0r0d[24], write_0r1d[24], wack_0n[24], ldata_0n[24], ldata_1n[24]);
  DRLATCH I240 (write_0r0d[25], write_0r1d[25], wack_0n[25], ldata_0n[25], ldata_1n[25]);
  DRLATCH I241 (write_0r0d[26], write_0r1d[26], wack_0n[26], ldata_0n[26], ldata_1n[26]);
  DRLATCH I242 (write_0r0d[27], write_0r1d[27], wack_0n[27], ldata_0n[27], ldata_1n[27]);
  DRLATCH I243 (write_0r0d[28], write_0r1d[28], wack_0n[28], ldata_0n[28], ldata_1n[28]);
  DRLATCH I244 (write_0r0d[29], write_0r1d[29], wack_0n[29], ldata_0n[29], ldata_1n[29]);
  DRLATCH I245 (write_0r0d[30], write_0r1d[30], wack_0n[30], ldata_0n[30], ldata_1n[30]);
  DRLATCH I246 (write_0r0d[31], write_0r1d[31], wack_0n[31], ldata_0n[31], ldata_1n[31]);
endmodule

module BrzVariable_35_1_s0_ (
  write_0r0d, write_0r1d, write_0a,
  read_0r, read_0a0d, read_0a1d
);
  input [34:0] write_0r0d;
  input [34:0] write_0r1d;
  output write_0a;
  input read_0r;
  output [34:0] read_0a0d;
  output [34:0] read_0a1d;
  wire [17:0] internal_0n;
  wire [34:0] store_0n;
  wire [34:0] store_1n;
  wire [34:0] ldata_0n;
  wire [34:0] ldata_1n;
  wire [34:0] wack_0n;
  wire readReq_0n;
  AND2 I0 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I1 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I2 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I3 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I4 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I5 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I6 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I7 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I8 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I9 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I10 (read_0a1d[10], store_1n[10], readReq_0n);
  AND2 I11 (read_0a1d[11], store_1n[11], readReq_0n);
  AND2 I12 (read_0a1d[12], store_1n[12], readReq_0n);
  AND2 I13 (read_0a1d[13], store_1n[13], readReq_0n);
  AND2 I14 (read_0a1d[14], store_1n[14], readReq_0n);
  AND2 I15 (read_0a1d[15], store_1n[15], readReq_0n);
  AND2 I16 (read_0a1d[16], store_1n[16], readReq_0n);
  AND2 I17 (read_0a1d[17], store_1n[17], readReq_0n);
  AND2 I18 (read_0a1d[18], store_1n[18], readReq_0n);
  AND2 I19 (read_0a1d[19], store_1n[19], readReq_0n);
  AND2 I20 (read_0a1d[20], store_1n[20], readReq_0n);
  AND2 I21 (read_0a1d[21], store_1n[21], readReq_0n);
  AND2 I22 (read_0a1d[22], store_1n[22], readReq_0n);
  AND2 I23 (read_0a1d[23], store_1n[23], readReq_0n);
  AND2 I24 (read_0a1d[24], store_1n[24], readReq_0n);
  AND2 I25 (read_0a1d[25], store_1n[25], readReq_0n);
  AND2 I26 (read_0a1d[26], store_1n[26], readReq_0n);
  AND2 I27 (read_0a1d[27], store_1n[27], readReq_0n);
  AND2 I28 (read_0a1d[28], store_1n[28], readReq_0n);
  AND2 I29 (read_0a1d[29], store_1n[29], readReq_0n);
  AND2 I30 (read_0a1d[30], store_1n[30], readReq_0n);
  AND2 I31 (read_0a1d[31], store_1n[31], readReq_0n);
  AND2 I32 (read_0a1d[32], store_1n[32], readReq_0n);
  AND2 I33 (read_0a1d[33], store_1n[33], readReq_0n);
  AND2 I34 (read_0a1d[34], store_1n[34], readReq_0n);
  AND2 I35 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I36 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I37 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I38 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I39 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I40 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I41 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I42 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I43 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I44 (read_0a0d[9], store_0n[9], readReq_0n);
  AND2 I45 (read_0a0d[10], store_0n[10], readReq_0n);
  AND2 I46 (read_0a0d[11], store_0n[11], readReq_0n);
  AND2 I47 (read_0a0d[12], store_0n[12], readReq_0n);
  AND2 I48 (read_0a0d[13], store_0n[13], readReq_0n);
  AND2 I49 (read_0a0d[14], store_0n[14], readReq_0n);
  AND2 I50 (read_0a0d[15], store_0n[15], readReq_0n);
  AND2 I51 (read_0a0d[16], store_0n[16], readReq_0n);
  AND2 I52 (read_0a0d[17], store_0n[17], readReq_0n);
  AND2 I53 (read_0a0d[18], store_0n[18], readReq_0n);
  AND2 I54 (read_0a0d[19], store_0n[19], readReq_0n);
  AND2 I55 (read_0a0d[20], store_0n[20], readReq_0n);
  AND2 I56 (read_0a0d[21], store_0n[21], readReq_0n);
  AND2 I57 (read_0a0d[22], store_0n[22], readReq_0n);
  AND2 I58 (read_0a0d[23], store_0n[23], readReq_0n);
  AND2 I59 (read_0a0d[24], store_0n[24], readReq_0n);
  AND2 I60 (read_0a0d[25], store_0n[25], readReq_0n);
  AND2 I61 (read_0a0d[26], store_0n[26], readReq_0n);
  AND2 I62 (read_0a0d[27], store_0n[27], readReq_0n);
  AND2 I63 (read_0a0d[28], store_0n[28], readReq_0n);
  AND2 I64 (read_0a0d[29], store_0n[29], readReq_0n);
  AND2 I65 (read_0a0d[30], store_0n[30], readReq_0n);
  AND2 I66 (read_0a0d[31], store_0n[31], readReq_0n);
  AND2 I67 (read_0a0d[32], store_0n[32], readReq_0n);
  AND2 I68 (read_0a0d[33], store_0n[33], readReq_0n);
  AND2 I69 (read_0a0d[34], store_0n[34], readReq_0n);
  BUFF I70 (readReq_0n, read_0r);
  BUFF I71 (store_0n[0], ldata_0n[0]);
  BUFF I72 (store_0n[1], ldata_0n[1]);
  BUFF I73 (store_0n[2], ldata_0n[2]);
  BUFF I74 (store_0n[3], ldata_0n[3]);
  BUFF I75 (store_0n[4], ldata_0n[4]);
  BUFF I76 (store_0n[5], ldata_0n[5]);
  BUFF I77 (store_0n[6], ldata_0n[6]);
  BUFF I78 (store_0n[7], ldata_0n[7]);
  BUFF I79 (store_0n[8], ldata_0n[8]);
  BUFF I80 (store_0n[9], ldata_0n[9]);
  BUFF I81 (store_0n[10], ldata_0n[10]);
  BUFF I82 (store_0n[11], ldata_0n[11]);
  BUFF I83 (store_0n[12], ldata_0n[12]);
  BUFF I84 (store_0n[13], ldata_0n[13]);
  BUFF I85 (store_0n[14], ldata_0n[14]);
  BUFF I86 (store_0n[15], ldata_0n[15]);
  BUFF I87 (store_0n[16], ldata_0n[16]);
  BUFF I88 (store_0n[17], ldata_0n[17]);
  BUFF I89 (store_0n[18], ldata_0n[18]);
  BUFF I90 (store_0n[19], ldata_0n[19]);
  BUFF I91 (store_0n[20], ldata_0n[20]);
  BUFF I92 (store_0n[21], ldata_0n[21]);
  BUFF I93 (store_0n[22], ldata_0n[22]);
  BUFF I94 (store_0n[23], ldata_0n[23]);
  BUFF I95 (store_0n[24], ldata_0n[24]);
  BUFF I96 (store_0n[25], ldata_0n[25]);
  BUFF I97 (store_0n[26], ldata_0n[26]);
  BUFF I98 (store_0n[27], ldata_0n[27]);
  BUFF I99 (store_0n[28], ldata_0n[28]);
  BUFF I100 (store_0n[29], ldata_0n[29]);
  BUFF I101 (store_0n[30], ldata_0n[30]);
  BUFF I102 (store_0n[31], ldata_0n[31]);
  BUFF I103 (store_0n[32], ldata_0n[32]);
  BUFF I104 (store_0n[33], ldata_0n[33]);
  BUFF I105 (store_0n[34], ldata_0n[34]);
  BUFF I106 (store_1n[0], ldata_1n[0]);
  BUFF I107 (store_1n[1], ldata_1n[1]);
  BUFF I108 (store_1n[2], ldata_1n[2]);
  BUFF I109 (store_1n[3], ldata_1n[3]);
  BUFF I110 (store_1n[4], ldata_1n[4]);
  BUFF I111 (store_1n[5], ldata_1n[5]);
  BUFF I112 (store_1n[6], ldata_1n[6]);
  BUFF I113 (store_1n[7], ldata_1n[7]);
  BUFF I114 (store_1n[8], ldata_1n[8]);
  BUFF I115 (store_1n[9], ldata_1n[9]);
  BUFF I116 (store_1n[10], ldata_1n[10]);
  BUFF I117 (store_1n[11], ldata_1n[11]);
  BUFF I118 (store_1n[12], ldata_1n[12]);
  BUFF I119 (store_1n[13], ldata_1n[13]);
  BUFF I120 (store_1n[14], ldata_1n[14]);
  BUFF I121 (store_1n[15], ldata_1n[15]);
  BUFF I122 (store_1n[16], ldata_1n[16]);
  BUFF I123 (store_1n[17], ldata_1n[17]);
  BUFF I124 (store_1n[18], ldata_1n[18]);
  BUFF I125 (store_1n[19], ldata_1n[19]);
  BUFF I126 (store_1n[20], ldata_1n[20]);
  BUFF I127 (store_1n[21], ldata_1n[21]);
  BUFF I128 (store_1n[22], ldata_1n[22]);
  BUFF I129 (store_1n[23], ldata_1n[23]);
  BUFF I130 (store_1n[24], ldata_1n[24]);
  BUFF I131 (store_1n[25], ldata_1n[25]);
  BUFF I132 (store_1n[26], ldata_1n[26]);
  BUFF I133 (store_1n[27], ldata_1n[27]);
  BUFF I134 (store_1n[28], ldata_1n[28]);
  BUFF I135 (store_1n[29], ldata_1n[29]);
  BUFF I136 (store_1n[30], ldata_1n[30]);
  BUFF I137 (store_1n[31], ldata_1n[31]);
  BUFF I138 (store_1n[32], ldata_1n[32]);
  BUFF I139 (store_1n[33], ldata_1n[33]);
  BUFF I140 (store_1n[34], ldata_1n[34]);
  C3 I141 (internal_0n[0], wack_0n[0], wack_0n[1], wack_0n[2]);
  C3 I142 (internal_0n[1], wack_0n[3], wack_0n[4], wack_0n[5]);
  C3 I143 (internal_0n[2], wack_0n[6], wack_0n[7], wack_0n[8]);
  C3 I144 (internal_0n[3], wack_0n[9], wack_0n[10], wack_0n[11]);
  C3 I145 (internal_0n[4], wack_0n[12], wack_0n[13], wack_0n[14]);
  C3 I146 (internal_0n[5], wack_0n[15], wack_0n[16], wack_0n[17]);
  C3 I147 (internal_0n[6], wack_0n[18], wack_0n[19], wack_0n[20]);
  C3 I148 (internal_0n[7], wack_0n[21], wack_0n[22], wack_0n[23]);
  C3 I149 (internal_0n[8], wack_0n[24], wack_0n[25], wack_0n[26]);
  C3 I150 (internal_0n[9], wack_0n[27], wack_0n[28], wack_0n[29]);
  C3 I151 (internal_0n[10], wack_0n[30], wack_0n[31], wack_0n[32]);
  C2 I152 (internal_0n[11], wack_0n[33], wack_0n[34]);
  C3 I153 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I154 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I155 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I156 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I157 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I158 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I159 (write_0a, internal_0n[16], internal_0n[17]);
  DRLATCH I160 (write_0r0d[0], write_0r1d[0], wack_0n[0], ldata_0n[0], ldata_1n[0]);
  DRLATCH I161 (write_0r0d[1], write_0r1d[1], wack_0n[1], ldata_0n[1], ldata_1n[1]);
  DRLATCH I162 (write_0r0d[2], write_0r1d[2], wack_0n[2], ldata_0n[2], ldata_1n[2]);
  DRLATCH I163 (write_0r0d[3], write_0r1d[3], wack_0n[3], ldata_0n[3], ldata_1n[3]);
  DRLATCH I164 (write_0r0d[4], write_0r1d[4], wack_0n[4], ldata_0n[4], ldata_1n[4]);
  DRLATCH I165 (write_0r0d[5], write_0r1d[5], wack_0n[5], ldata_0n[5], ldata_1n[5]);
  DRLATCH I166 (write_0r0d[6], write_0r1d[6], wack_0n[6], ldata_0n[6], ldata_1n[6]);
  DRLATCH I167 (write_0r0d[7], write_0r1d[7], wack_0n[7], ldata_0n[7], ldata_1n[7]);
  DRLATCH I168 (write_0r0d[8], write_0r1d[8], wack_0n[8], ldata_0n[8], ldata_1n[8]);
  DRLATCH I169 (write_0r0d[9], write_0r1d[9], wack_0n[9], ldata_0n[9], ldata_1n[9]);
  DRLATCH I170 (write_0r0d[10], write_0r1d[10], wack_0n[10], ldata_0n[10], ldata_1n[10]);
  DRLATCH I171 (write_0r0d[11], write_0r1d[11], wack_0n[11], ldata_0n[11], ldata_1n[11]);
  DRLATCH I172 (write_0r0d[12], write_0r1d[12], wack_0n[12], ldata_0n[12], ldata_1n[12]);
  DRLATCH I173 (write_0r0d[13], write_0r1d[13], wack_0n[13], ldata_0n[13], ldata_1n[13]);
  DRLATCH I174 (write_0r0d[14], write_0r1d[14], wack_0n[14], ldata_0n[14], ldata_1n[14]);
  DRLATCH I175 (write_0r0d[15], write_0r1d[15], wack_0n[15], ldata_0n[15], ldata_1n[15]);
  DRLATCH I176 (write_0r0d[16], write_0r1d[16], wack_0n[16], ldata_0n[16], ldata_1n[16]);
  DRLATCH I177 (write_0r0d[17], write_0r1d[17], wack_0n[17], ldata_0n[17], ldata_1n[17]);
  DRLATCH I178 (write_0r0d[18], write_0r1d[18], wack_0n[18], ldata_0n[18], ldata_1n[18]);
  DRLATCH I179 (write_0r0d[19], write_0r1d[19], wack_0n[19], ldata_0n[19], ldata_1n[19]);
  DRLATCH I180 (write_0r0d[20], write_0r1d[20], wack_0n[20], ldata_0n[20], ldata_1n[20]);
  DRLATCH I181 (write_0r0d[21], write_0r1d[21], wack_0n[21], ldata_0n[21], ldata_1n[21]);
  DRLATCH I182 (write_0r0d[22], write_0r1d[22], wack_0n[22], ldata_0n[22], ldata_1n[22]);
  DRLATCH I183 (write_0r0d[23], write_0r1d[23], wack_0n[23], ldata_0n[23], ldata_1n[23]);
  DRLATCH I184 (write_0r0d[24], write_0r1d[24], wack_0n[24], ldata_0n[24], ldata_1n[24]);
  DRLATCH I185 (write_0r0d[25], write_0r1d[25], wack_0n[25], ldata_0n[25], ldata_1n[25]);
  DRLATCH I186 (write_0r0d[26], write_0r1d[26], wack_0n[26], ldata_0n[26], ldata_1n[26]);
  DRLATCH I187 (write_0r0d[27], write_0r1d[27], wack_0n[27], ldata_0n[27], ldata_1n[27]);
  DRLATCH I188 (write_0r0d[28], write_0r1d[28], wack_0n[28], ldata_0n[28], ldata_1n[28]);
  DRLATCH I189 (write_0r0d[29], write_0r1d[29], wack_0n[29], ldata_0n[29], ldata_1n[29]);
  DRLATCH I190 (write_0r0d[30], write_0r1d[30], wack_0n[30], ldata_0n[30], ldata_1n[30]);
  DRLATCH I191 (write_0r0d[31], write_0r1d[31], wack_0n[31], ldata_0n[31], ldata_1n[31]);
  DRLATCH I192 (write_0r0d[32], write_0r1d[32], wack_0n[32], ldata_0n[32], ldata_1n[32]);
  DRLATCH I193 (write_0r0d[33], write_0r1d[33], wack_0n[33], ldata_0n[33], ldata_1n[33]);
  DRLATCH I194 (write_0r0d[34], write_0r1d[34], wack_0n[34], ldata_0n[34], ldata_1n[34]);
endmodule

module BrzVariable_35_2_s0_ (
  write_0r0d, write_0r1d, write_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d
);
  input [34:0] write_0r0d;
  input [34:0] write_0r1d;
  output write_0a;
  input read_0r;
  output [34:0] read_0a0d;
  output [34:0] read_0a1d;
  input read_1r;
  output [34:0] read_1a0d;
  output [34:0] read_1a1d;
  wire [17:0] internal_0n;
  wire [34:0] store_0n;
  wire [34:0] store_1n;
  wire [34:0] ldata_0n;
  wire [34:0] ldata_1n;
  wire [34:0] wack_0n;
  wire readReq_0n;
  wire readReq_1n;
  AND2 I0 (read_1a1d[0], store_1n[0], readReq_1n);
  AND2 I1 (read_1a1d[1], store_1n[1], readReq_1n);
  AND2 I2 (read_1a1d[2], store_1n[2], readReq_1n);
  AND2 I3 (read_1a1d[3], store_1n[3], readReq_1n);
  AND2 I4 (read_1a1d[4], store_1n[4], readReq_1n);
  AND2 I5 (read_1a1d[5], store_1n[5], readReq_1n);
  AND2 I6 (read_1a1d[6], store_1n[6], readReq_1n);
  AND2 I7 (read_1a1d[7], store_1n[7], readReq_1n);
  AND2 I8 (read_1a1d[8], store_1n[8], readReq_1n);
  AND2 I9 (read_1a1d[9], store_1n[9], readReq_1n);
  AND2 I10 (read_1a1d[10], store_1n[10], readReq_1n);
  AND2 I11 (read_1a1d[11], store_1n[11], readReq_1n);
  AND2 I12 (read_1a1d[12], store_1n[12], readReq_1n);
  AND2 I13 (read_1a1d[13], store_1n[13], readReq_1n);
  AND2 I14 (read_1a1d[14], store_1n[14], readReq_1n);
  AND2 I15 (read_1a1d[15], store_1n[15], readReq_1n);
  AND2 I16 (read_1a1d[16], store_1n[16], readReq_1n);
  AND2 I17 (read_1a1d[17], store_1n[17], readReq_1n);
  AND2 I18 (read_1a1d[18], store_1n[18], readReq_1n);
  AND2 I19 (read_1a1d[19], store_1n[19], readReq_1n);
  AND2 I20 (read_1a1d[20], store_1n[20], readReq_1n);
  AND2 I21 (read_1a1d[21], store_1n[21], readReq_1n);
  AND2 I22 (read_1a1d[22], store_1n[22], readReq_1n);
  AND2 I23 (read_1a1d[23], store_1n[23], readReq_1n);
  AND2 I24 (read_1a1d[24], store_1n[24], readReq_1n);
  AND2 I25 (read_1a1d[25], store_1n[25], readReq_1n);
  AND2 I26 (read_1a1d[26], store_1n[26], readReq_1n);
  AND2 I27 (read_1a1d[27], store_1n[27], readReq_1n);
  AND2 I28 (read_1a1d[28], store_1n[28], readReq_1n);
  AND2 I29 (read_1a1d[29], store_1n[29], readReq_1n);
  AND2 I30 (read_1a1d[30], store_1n[30], readReq_1n);
  AND2 I31 (read_1a1d[31], store_1n[31], readReq_1n);
  AND2 I32 (read_1a1d[32], store_1n[32], readReq_1n);
  AND2 I33 (read_1a1d[33], store_1n[33], readReq_1n);
  AND2 I34 (read_1a1d[34], store_1n[34], readReq_1n);
  AND2 I35 (read_1a0d[0], store_0n[0], readReq_1n);
  AND2 I36 (read_1a0d[1], store_0n[1], readReq_1n);
  AND2 I37 (read_1a0d[2], store_0n[2], readReq_1n);
  AND2 I38 (read_1a0d[3], store_0n[3], readReq_1n);
  AND2 I39 (read_1a0d[4], store_0n[4], readReq_1n);
  AND2 I40 (read_1a0d[5], store_0n[5], readReq_1n);
  AND2 I41 (read_1a0d[6], store_0n[6], readReq_1n);
  AND2 I42 (read_1a0d[7], store_0n[7], readReq_1n);
  AND2 I43 (read_1a0d[8], store_0n[8], readReq_1n);
  AND2 I44 (read_1a0d[9], store_0n[9], readReq_1n);
  AND2 I45 (read_1a0d[10], store_0n[10], readReq_1n);
  AND2 I46 (read_1a0d[11], store_0n[11], readReq_1n);
  AND2 I47 (read_1a0d[12], store_0n[12], readReq_1n);
  AND2 I48 (read_1a0d[13], store_0n[13], readReq_1n);
  AND2 I49 (read_1a0d[14], store_0n[14], readReq_1n);
  AND2 I50 (read_1a0d[15], store_0n[15], readReq_1n);
  AND2 I51 (read_1a0d[16], store_0n[16], readReq_1n);
  AND2 I52 (read_1a0d[17], store_0n[17], readReq_1n);
  AND2 I53 (read_1a0d[18], store_0n[18], readReq_1n);
  AND2 I54 (read_1a0d[19], store_0n[19], readReq_1n);
  AND2 I55 (read_1a0d[20], store_0n[20], readReq_1n);
  AND2 I56 (read_1a0d[21], store_0n[21], readReq_1n);
  AND2 I57 (read_1a0d[22], store_0n[22], readReq_1n);
  AND2 I58 (read_1a0d[23], store_0n[23], readReq_1n);
  AND2 I59 (read_1a0d[24], store_0n[24], readReq_1n);
  AND2 I60 (read_1a0d[25], store_0n[25], readReq_1n);
  AND2 I61 (read_1a0d[26], store_0n[26], readReq_1n);
  AND2 I62 (read_1a0d[27], store_0n[27], readReq_1n);
  AND2 I63 (read_1a0d[28], store_0n[28], readReq_1n);
  AND2 I64 (read_1a0d[29], store_0n[29], readReq_1n);
  AND2 I65 (read_1a0d[30], store_0n[30], readReq_1n);
  AND2 I66 (read_1a0d[31], store_0n[31], readReq_1n);
  AND2 I67 (read_1a0d[32], store_0n[32], readReq_1n);
  AND2 I68 (read_1a0d[33], store_0n[33], readReq_1n);
  AND2 I69 (read_1a0d[34], store_0n[34], readReq_1n);
  AND2 I70 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I71 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I72 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I73 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I74 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I75 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I76 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I77 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I78 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I79 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I80 (read_0a1d[10], store_1n[10], readReq_0n);
  AND2 I81 (read_0a1d[11], store_1n[11], readReq_0n);
  AND2 I82 (read_0a1d[12], store_1n[12], readReq_0n);
  AND2 I83 (read_0a1d[13], store_1n[13], readReq_0n);
  AND2 I84 (read_0a1d[14], store_1n[14], readReq_0n);
  AND2 I85 (read_0a1d[15], store_1n[15], readReq_0n);
  AND2 I86 (read_0a1d[16], store_1n[16], readReq_0n);
  AND2 I87 (read_0a1d[17], store_1n[17], readReq_0n);
  AND2 I88 (read_0a1d[18], store_1n[18], readReq_0n);
  AND2 I89 (read_0a1d[19], store_1n[19], readReq_0n);
  AND2 I90 (read_0a1d[20], store_1n[20], readReq_0n);
  AND2 I91 (read_0a1d[21], store_1n[21], readReq_0n);
  AND2 I92 (read_0a1d[22], store_1n[22], readReq_0n);
  AND2 I93 (read_0a1d[23], store_1n[23], readReq_0n);
  AND2 I94 (read_0a1d[24], store_1n[24], readReq_0n);
  AND2 I95 (read_0a1d[25], store_1n[25], readReq_0n);
  AND2 I96 (read_0a1d[26], store_1n[26], readReq_0n);
  AND2 I97 (read_0a1d[27], store_1n[27], readReq_0n);
  AND2 I98 (read_0a1d[28], store_1n[28], readReq_0n);
  AND2 I99 (read_0a1d[29], store_1n[29], readReq_0n);
  AND2 I100 (read_0a1d[30], store_1n[30], readReq_0n);
  AND2 I101 (read_0a1d[31], store_1n[31], readReq_0n);
  AND2 I102 (read_0a1d[32], store_1n[32], readReq_0n);
  AND2 I103 (read_0a1d[33], store_1n[33], readReq_0n);
  AND2 I104 (read_0a1d[34], store_1n[34], readReq_0n);
  AND2 I105 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I106 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I107 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I108 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I109 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I110 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I111 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I112 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I113 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I114 (read_0a0d[9], store_0n[9], readReq_0n);
  AND2 I115 (read_0a0d[10], store_0n[10], readReq_0n);
  AND2 I116 (read_0a0d[11], store_0n[11], readReq_0n);
  AND2 I117 (read_0a0d[12], store_0n[12], readReq_0n);
  AND2 I118 (read_0a0d[13], store_0n[13], readReq_0n);
  AND2 I119 (read_0a0d[14], store_0n[14], readReq_0n);
  AND2 I120 (read_0a0d[15], store_0n[15], readReq_0n);
  AND2 I121 (read_0a0d[16], store_0n[16], readReq_0n);
  AND2 I122 (read_0a0d[17], store_0n[17], readReq_0n);
  AND2 I123 (read_0a0d[18], store_0n[18], readReq_0n);
  AND2 I124 (read_0a0d[19], store_0n[19], readReq_0n);
  AND2 I125 (read_0a0d[20], store_0n[20], readReq_0n);
  AND2 I126 (read_0a0d[21], store_0n[21], readReq_0n);
  AND2 I127 (read_0a0d[22], store_0n[22], readReq_0n);
  AND2 I128 (read_0a0d[23], store_0n[23], readReq_0n);
  AND2 I129 (read_0a0d[24], store_0n[24], readReq_0n);
  AND2 I130 (read_0a0d[25], store_0n[25], readReq_0n);
  AND2 I131 (read_0a0d[26], store_0n[26], readReq_0n);
  AND2 I132 (read_0a0d[27], store_0n[27], readReq_0n);
  AND2 I133 (read_0a0d[28], store_0n[28], readReq_0n);
  AND2 I134 (read_0a0d[29], store_0n[29], readReq_0n);
  AND2 I135 (read_0a0d[30], store_0n[30], readReq_0n);
  AND2 I136 (read_0a0d[31], store_0n[31], readReq_0n);
  AND2 I137 (read_0a0d[32], store_0n[32], readReq_0n);
  AND2 I138 (read_0a0d[33], store_0n[33], readReq_0n);
  AND2 I139 (read_0a0d[34], store_0n[34], readReq_0n);
  BUFF I140 (readReq_0n, read_0r);
  BUFF I141 (readReq_1n, read_1r);
  BUFF I142 (store_0n[0], ldata_0n[0]);
  BUFF I143 (store_0n[1], ldata_0n[1]);
  BUFF I144 (store_0n[2], ldata_0n[2]);
  BUFF I145 (store_0n[3], ldata_0n[3]);
  BUFF I146 (store_0n[4], ldata_0n[4]);
  BUFF I147 (store_0n[5], ldata_0n[5]);
  BUFF I148 (store_0n[6], ldata_0n[6]);
  BUFF I149 (store_0n[7], ldata_0n[7]);
  BUFF I150 (store_0n[8], ldata_0n[8]);
  BUFF I151 (store_0n[9], ldata_0n[9]);
  BUFF I152 (store_0n[10], ldata_0n[10]);
  BUFF I153 (store_0n[11], ldata_0n[11]);
  BUFF I154 (store_0n[12], ldata_0n[12]);
  BUFF I155 (store_0n[13], ldata_0n[13]);
  BUFF I156 (store_0n[14], ldata_0n[14]);
  BUFF I157 (store_0n[15], ldata_0n[15]);
  BUFF I158 (store_0n[16], ldata_0n[16]);
  BUFF I159 (store_0n[17], ldata_0n[17]);
  BUFF I160 (store_0n[18], ldata_0n[18]);
  BUFF I161 (store_0n[19], ldata_0n[19]);
  BUFF I162 (store_0n[20], ldata_0n[20]);
  BUFF I163 (store_0n[21], ldata_0n[21]);
  BUFF I164 (store_0n[22], ldata_0n[22]);
  BUFF I165 (store_0n[23], ldata_0n[23]);
  BUFF I166 (store_0n[24], ldata_0n[24]);
  BUFF I167 (store_0n[25], ldata_0n[25]);
  BUFF I168 (store_0n[26], ldata_0n[26]);
  BUFF I169 (store_0n[27], ldata_0n[27]);
  BUFF I170 (store_0n[28], ldata_0n[28]);
  BUFF I171 (store_0n[29], ldata_0n[29]);
  BUFF I172 (store_0n[30], ldata_0n[30]);
  BUFF I173 (store_0n[31], ldata_0n[31]);
  BUFF I174 (store_0n[32], ldata_0n[32]);
  BUFF I175 (store_0n[33], ldata_0n[33]);
  BUFF I176 (store_0n[34], ldata_0n[34]);
  BUFF I177 (store_1n[0], ldata_1n[0]);
  BUFF I178 (store_1n[1], ldata_1n[1]);
  BUFF I179 (store_1n[2], ldata_1n[2]);
  BUFF I180 (store_1n[3], ldata_1n[3]);
  BUFF I181 (store_1n[4], ldata_1n[4]);
  BUFF I182 (store_1n[5], ldata_1n[5]);
  BUFF I183 (store_1n[6], ldata_1n[6]);
  BUFF I184 (store_1n[7], ldata_1n[7]);
  BUFF I185 (store_1n[8], ldata_1n[8]);
  BUFF I186 (store_1n[9], ldata_1n[9]);
  BUFF I187 (store_1n[10], ldata_1n[10]);
  BUFF I188 (store_1n[11], ldata_1n[11]);
  BUFF I189 (store_1n[12], ldata_1n[12]);
  BUFF I190 (store_1n[13], ldata_1n[13]);
  BUFF I191 (store_1n[14], ldata_1n[14]);
  BUFF I192 (store_1n[15], ldata_1n[15]);
  BUFF I193 (store_1n[16], ldata_1n[16]);
  BUFF I194 (store_1n[17], ldata_1n[17]);
  BUFF I195 (store_1n[18], ldata_1n[18]);
  BUFF I196 (store_1n[19], ldata_1n[19]);
  BUFF I197 (store_1n[20], ldata_1n[20]);
  BUFF I198 (store_1n[21], ldata_1n[21]);
  BUFF I199 (store_1n[22], ldata_1n[22]);
  BUFF I200 (store_1n[23], ldata_1n[23]);
  BUFF I201 (store_1n[24], ldata_1n[24]);
  BUFF I202 (store_1n[25], ldata_1n[25]);
  BUFF I203 (store_1n[26], ldata_1n[26]);
  BUFF I204 (store_1n[27], ldata_1n[27]);
  BUFF I205 (store_1n[28], ldata_1n[28]);
  BUFF I206 (store_1n[29], ldata_1n[29]);
  BUFF I207 (store_1n[30], ldata_1n[30]);
  BUFF I208 (store_1n[31], ldata_1n[31]);
  BUFF I209 (store_1n[32], ldata_1n[32]);
  BUFF I210 (store_1n[33], ldata_1n[33]);
  BUFF I211 (store_1n[34], ldata_1n[34]);
  C3 I212 (internal_0n[0], wack_0n[0], wack_0n[1], wack_0n[2]);
  C3 I213 (internal_0n[1], wack_0n[3], wack_0n[4], wack_0n[5]);
  C3 I214 (internal_0n[2], wack_0n[6], wack_0n[7], wack_0n[8]);
  C3 I215 (internal_0n[3], wack_0n[9], wack_0n[10], wack_0n[11]);
  C3 I216 (internal_0n[4], wack_0n[12], wack_0n[13], wack_0n[14]);
  C3 I217 (internal_0n[5], wack_0n[15], wack_0n[16], wack_0n[17]);
  C3 I218 (internal_0n[6], wack_0n[18], wack_0n[19], wack_0n[20]);
  C3 I219 (internal_0n[7], wack_0n[21], wack_0n[22], wack_0n[23]);
  C3 I220 (internal_0n[8], wack_0n[24], wack_0n[25], wack_0n[26]);
  C3 I221 (internal_0n[9], wack_0n[27], wack_0n[28], wack_0n[29]);
  C3 I222 (internal_0n[10], wack_0n[30], wack_0n[31], wack_0n[32]);
  C2 I223 (internal_0n[11], wack_0n[33], wack_0n[34]);
  C3 I224 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I225 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I226 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I227 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I228 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I229 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I230 (write_0a, internal_0n[16], internal_0n[17]);
  DRLATCH I231 (write_0r0d[0], write_0r1d[0], wack_0n[0], ldata_0n[0], ldata_1n[0]);
  DRLATCH I232 (write_0r0d[1], write_0r1d[1], wack_0n[1], ldata_0n[1], ldata_1n[1]);
  DRLATCH I233 (write_0r0d[2], write_0r1d[2], wack_0n[2], ldata_0n[2], ldata_1n[2]);
  DRLATCH I234 (write_0r0d[3], write_0r1d[3], wack_0n[3], ldata_0n[3], ldata_1n[3]);
  DRLATCH I235 (write_0r0d[4], write_0r1d[4], wack_0n[4], ldata_0n[4], ldata_1n[4]);
  DRLATCH I236 (write_0r0d[5], write_0r1d[5], wack_0n[5], ldata_0n[5], ldata_1n[5]);
  DRLATCH I237 (write_0r0d[6], write_0r1d[6], wack_0n[6], ldata_0n[6], ldata_1n[6]);
  DRLATCH I238 (write_0r0d[7], write_0r1d[7], wack_0n[7], ldata_0n[7], ldata_1n[7]);
  DRLATCH I239 (write_0r0d[8], write_0r1d[8], wack_0n[8], ldata_0n[8], ldata_1n[8]);
  DRLATCH I240 (write_0r0d[9], write_0r1d[9], wack_0n[9], ldata_0n[9], ldata_1n[9]);
  DRLATCH I241 (write_0r0d[10], write_0r1d[10], wack_0n[10], ldata_0n[10], ldata_1n[10]);
  DRLATCH I242 (write_0r0d[11], write_0r1d[11], wack_0n[11], ldata_0n[11], ldata_1n[11]);
  DRLATCH I243 (write_0r0d[12], write_0r1d[12], wack_0n[12], ldata_0n[12], ldata_1n[12]);
  DRLATCH I244 (write_0r0d[13], write_0r1d[13], wack_0n[13], ldata_0n[13], ldata_1n[13]);
  DRLATCH I245 (write_0r0d[14], write_0r1d[14], wack_0n[14], ldata_0n[14], ldata_1n[14]);
  DRLATCH I246 (write_0r0d[15], write_0r1d[15], wack_0n[15], ldata_0n[15], ldata_1n[15]);
  DRLATCH I247 (write_0r0d[16], write_0r1d[16], wack_0n[16], ldata_0n[16], ldata_1n[16]);
  DRLATCH I248 (write_0r0d[17], write_0r1d[17], wack_0n[17], ldata_0n[17], ldata_1n[17]);
  DRLATCH I249 (write_0r0d[18], write_0r1d[18], wack_0n[18], ldata_0n[18], ldata_1n[18]);
  DRLATCH I250 (write_0r0d[19], write_0r1d[19], wack_0n[19], ldata_0n[19], ldata_1n[19]);
  DRLATCH I251 (write_0r0d[20], write_0r1d[20], wack_0n[20], ldata_0n[20], ldata_1n[20]);
  DRLATCH I252 (write_0r0d[21], write_0r1d[21], wack_0n[21], ldata_0n[21], ldata_1n[21]);
  DRLATCH I253 (write_0r0d[22], write_0r1d[22], wack_0n[22], ldata_0n[22], ldata_1n[22]);
  DRLATCH I254 (write_0r0d[23], write_0r1d[23], wack_0n[23], ldata_0n[23], ldata_1n[23]);
  DRLATCH I255 (write_0r0d[24], write_0r1d[24], wack_0n[24], ldata_0n[24], ldata_1n[24]);
  DRLATCH I256 (write_0r0d[25], write_0r1d[25], wack_0n[25], ldata_0n[25], ldata_1n[25]);
  DRLATCH I257 (write_0r0d[26], write_0r1d[26], wack_0n[26], ldata_0n[26], ldata_1n[26]);
  DRLATCH I258 (write_0r0d[27], write_0r1d[27], wack_0n[27], ldata_0n[27], ldata_1n[27]);
  DRLATCH I259 (write_0r0d[28], write_0r1d[28], wack_0n[28], ldata_0n[28], ldata_1n[28]);
  DRLATCH I260 (write_0r0d[29], write_0r1d[29], wack_0n[29], ldata_0n[29], ldata_1n[29]);
  DRLATCH I261 (write_0r0d[30], write_0r1d[30], wack_0n[30], ldata_0n[30], ldata_1n[30]);
  DRLATCH I262 (write_0r0d[31], write_0r1d[31], wack_0n[31], ldata_0n[31], ldata_1n[31]);
  DRLATCH I263 (write_0r0d[32], write_0r1d[32], wack_0n[32], ldata_0n[32], ldata_1n[32]);
  DRLATCH I264 (write_0r0d[33], write_0r1d[33], wack_0n[33], ldata_0n[33], ldata_1n[33]);
  DRLATCH I265 (write_0r0d[34], write_0r1d[34], wack_0n[34], ldata_0n[34], ldata_1n[34]);
endmodule

module BrzVariable_35_2_s12__3b0_2e_2e30 (
  write_0r0d, write_0r1d, write_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d
);
  input [34:0] write_0r0d;
  input [34:0] write_0r1d;
  output write_0a;
  input read_0r;
  output [34:0] read_0a0d;
  output [34:0] read_0a1d;
  input read_1r;
  output [30:0] read_1a0d;
  output [30:0] read_1a1d;
  wire [17:0] internal_0n;
  wire [34:0] store_0n;
  wire [34:0] store_1n;
  wire [34:0] ldata_0n;
  wire [34:0] ldata_1n;
  wire [34:0] wack_0n;
  wire readReq_0n;
  wire readReq_1n;
  AND2 I0 (read_1a1d[0], store_1n[0], readReq_1n);
  AND2 I1 (read_1a1d[1], store_1n[1], readReq_1n);
  AND2 I2 (read_1a1d[2], store_1n[2], readReq_1n);
  AND2 I3 (read_1a1d[3], store_1n[3], readReq_1n);
  AND2 I4 (read_1a1d[4], store_1n[4], readReq_1n);
  AND2 I5 (read_1a1d[5], store_1n[5], readReq_1n);
  AND2 I6 (read_1a1d[6], store_1n[6], readReq_1n);
  AND2 I7 (read_1a1d[7], store_1n[7], readReq_1n);
  AND2 I8 (read_1a1d[8], store_1n[8], readReq_1n);
  AND2 I9 (read_1a1d[9], store_1n[9], readReq_1n);
  AND2 I10 (read_1a1d[10], store_1n[10], readReq_1n);
  AND2 I11 (read_1a1d[11], store_1n[11], readReq_1n);
  AND2 I12 (read_1a1d[12], store_1n[12], readReq_1n);
  AND2 I13 (read_1a1d[13], store_1n[13], readReq_1n);
  AND2 I14 (read_1a1d[14], store_1n[14], readReq_1n);
  AND2 I15 (read_1a1d[15], store_1n[15], readReq_1n);
  AND2 I16 (read_1a1d[16], store_1n[16], readReq_1n);
  AND2 I17 (read_1a1d[17], store_1n[17], readReq_1n);
  AND2 I18 (read_1a1d[18], store_1n[18], readReq_1n);
  AND2 I19 (read_1a1d[19], store_1n[19], readReq_1n);
  AND2 I20 (read_1a1d[20], store_1n[20], readReq_1n);
  AND2 I21 (read_1a1d[21], store_1n[21], readReq_1n);
  AND2 I22 (read_1a1d[22], store_1n[22], readReq_1n);
  AND2 I23 (read_1a1d[23], store_1n[23], readReq_1n);
  AND2 I24 (read_1a1d[24], store_1n[24], readReq_1n);
  AND2 I25 (read_1a1d[25], store_1n[25], readReq_1n);
  AND2 I26 (read_1a1d[26], store_1n[26], readReq_1n);
  AND2 I27 (read_1a1d[27], store_1n[27], readReq_1n);
  AND2 I28 (read_1a1d[28], store_1n[28], readReq_1n);
  AND2 I29 (read_1a1d[29], store_1n[29], readReq_1n);
  AND2 I30 (read_1a1d[30], store_1n[30], readReq_1n);
  AND2 I31 (read_1a0d[0], store_0n[0], readReq_1n);
  AND2 I32 (read_1a0d[1], store_0n[1], readReq_1n);
  AND2 I33 (read_1a0d[2], store_0n[2], readReq_1n);
  AND2 I34 (read_1a0d[3], store_0n[3], readReq_1n);
  AND2 I35 (read_1a0d[4], store_0n[4], readReq_1n);
  AND2 I36 (read_1a0d[5], store_0n[5], readReq_1n);
  AND2 I37 (read_1a0d[6], store_0n[6], readReq_1n);
  AND2 I38 (read_1a0d[7], store_0n[7], readReq_1n);
  AND2 I39 (read_1a0d[8], store_0n[8], readReq_1n);
  AND2 I40 (read_1a0d[9], store_0n[9], readReq_1n);
  AND2 I41 (read_1a0d[10], store_0n[10], readReq_1n);
  AND2 I42 (read_1a0d[11], store_0n[11], readReq_1n);
  AND2 I43 (read_1a0d[12], store_0n[12], readReq_1n);
  AND2 I44 (read_1a0d[13], store_0n[13], readReq_1n);
  AND2 I45 (read_1a0d[14], store_0n[14], readReq_1n);
  AND2 I46 (read_1a0d[15], store_0n[15], readReq_1n);
  AND2 I47 (read_1a0d[16], store_0n[16], readReq_1n);
  AND2 I48 (read_1a0d[17], store_0n[17], readReq_1n);
  AND2 I49 (read_1a0d[18], store_0n[18], readReq_1n);
  AND2 I50 (read_1a0d[19], store_0n[19], readReq_1n);
  AND2 I51 (read_1a0d[20], store_0n[20], readReq_1n);
  AND2 I52 (read_1a0d[21], store_0n[21], readReq_1n);
  AND2 I53 (read_1a0d[22], store_0n[22], readReq_1n);
  AND2 I54 (read_1a0d[23], store_0n[23], readReq_1n);
  AND2 I55 (read_1a0d[24], store_0n[24], readReq_1n);
  AND2 I56 (read_1a0d[25], store_0n[25], readReq_1n);
  AND2 I57 (read_1a0d[26], store_0n[26], readReq_1n);
  AND2 I58 (read_1a0d[27], store_0n[27], readReq_1n);
  AND2 I59 (read_1a0d[28], store_0n[28], readReq_1n);
  AND2 I60 (read_1a0d[29], store_0n[29], readReq_1n);
  AND2 I61 (read_1a0d[30], store_0n[30], readReq_1n);
  AND2 I62 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I63 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I64 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I65 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I66 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I67 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I68 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I69 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I70 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I71 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I72 (read_0a1d[10], store_1n[10], readReq_0n);
  AND2 I73 (read_0a1d[11], store_1n[11], readReq_0n);
  AND2 I74 (read_0a1d[12], store_1n[12], readReq_0n);
  AND2 I75 (read_0a1d[13], store_1n[13], readReq_0n);
  AND2 I76 (read_0a1d[14], store_1n[14], readReq_0n);
  AND2 I77 (read_0a1d[15], store_1n[15], readReq_0n);
  AND2 I78 (read_0a1d[16], store_1n[16], readReq_0n);
  AND2 I79 (read_0a1d[17], store_1n[17], readReq_0n);
  AND2 I80 (read_0a1d[18], store_1n[18], readReq_0n);
  AND2 I81 (read_0a1d[19], store_1n[19], readReq_0n);
  AND2 I82 (read_0a1d[20], store_1n[20], readReq_0n);
  AND2 I83 (read_0a1d[21], store_1n[21], readReq_0n);
  AND2 I84 (read_0a1d[22], store_1n[22], readReq_0n);
  AND2 I85 (read_0a1d[23], store_1n[23], readReq_0n);
  AND2 I86 (read_0a1d[24], store_1n[24], readReq_0n);
  AND2 I87 (read_0a1d[25], store_1n[25], readReq_0n);
  AND2 I88 (read_0a1d[26], store_1n[26], readReq_0n);
  AND2 I89 (read_0a1d[27], store_1n[27], readReq_0n);
  AND2 I90 (read_0a1d[28], store_1n[28], readReq_0n);
  AND2 I91 (read_0a1d[29], store_1n[29], readReq_0n);
  AND2 I92 (read_0a1d[30], store_1n[30], readReq_0n);
  AND2 I93 (read_0a1d[31], store_1n[31], readReq_0n);
  AND2 I94 (read_0a1d[32], store_1n[32], readReq_0n);
  AND2 I95 (read_0a1d[33], store_1n[33], readReq_0n);
  AND2 I96 (read_0a1d[34], store_1n[34], readReq_0n);
  AND2 I97 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I98 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I99 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I100 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I101 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I102 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I103 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I104 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I105 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I106 (read_0a0d[9], store_0n[9], readReq_0n);
  AND2 I107 (read_0a0d[10], store_0n[10], readReq_0n);
  AND2 I108 (read_0a0d[11], store_0n[11], readReq_0n);
  AND2 I109 (read_0a0d[12], store_0n[12], readReq_0n);
  AND2 I110 (read_0a0d[13], store_0n[13], readReq_0n);
  AND2 I111 (read_0a0d[14], store_0n[14], readReq_0n);
  AND2 I112 (read_0a0d[15], store_0n[15], readReq_0n);
  AND2 I113 (read_0a0d[16], store_0n[16], readReq_0n);
  AND2 I114 (read_0a0d[17], store_0n[17], readReq_0n);
  AND2 I115 (read_0a0d[18], store_0n[18], readReq_0n);
  AND2 I116 (read_0a0d[19], store_0n[19], readReq_0n);
  AND2 I117 (read_0a0d[20], store_0n[20], readReq_0n);
  AND2 I118 (read_0a0d[21], store_0n[21], readReq_0n);
  AND2 I119 (read_0a0d[22], store_0n[22], readReq_0n);
  AND2 I120 (read_0a0d[23], store_0n[23], readReq_0n);
  AND2 I121 (read_0a0d[24], store_0n[24], readReq_0n);
  AND2 I122 (read_0a0d[25], store_0n[25], readReq_0n);
  AND2 I123 (read_0a0d[26], store_0n[26], readReq_0n);
  AND2 I124 (read_0a0d[27], store_0n[27], readReq_0n);
  AND2 I125 (read_0a0d[28], store_0n[28], readReq_0n);
  AND2 I126 (read_0a0d[29], store_0n[29], readReq_0n);
  AND2 I127 (read_0a0d[30], store_0n[30], readReq_0n);
  AND2 I128 (read_0a0d[31], store_0n[31], readReq_0n);
  AND2 I129 (read_0a0d[32], store_0n[32], readReq_0n);
  AND2 I130 (read_0a0d[33], store_0n[33], readReq_0n);
  AND2 I131 (read_0a0d[34], store_0n[34], readReq_0n);
  BUFF I132 (readReq_0n, read_0r);
  BUFF I133 (readReq_1n, read_1r);
  BUFF I134 (store_0n[0], ldata_0n[0]);
  BUFF I135 (store_0n[1], ldata_0n[1]);
  BUFF I136 (store_0n[2], ldata_0n[2]);
  BUFF I137 (store_0n[3], ldata_0n[3]);
  BUFF I138 (store_0n[4], ldata_0n[4]);
  BUFF I139 (store_0n[5], ldata_0n[5]);
  BUFF I140 (store_0n[6], ldata_0n[6]);
  BUFF I141 (store_0n[7], ldata_0n[7]);
  BUFF I142 (store_0n[8], ldata_0n[8]);
  BUFF I143 (store_0n[9], ldata_0n[9]);
  BUFF I144 (store_0n[10], ldata_0n[10]);
  BUFF I145 (store_0n[11], ldata_0n[11]);
  BUFF I146 (store_0n[12], ldata_0n[12]);
  BUFF I147 (store_0n[13], ldata_0n[13]);
  BUFF I148 (store_0n[14], ldata_0n[14]);
  BUFF I149 (store_0n[15], ldata_0n[15]);
  BUFF I150 (store_0n[16], ldata_0n[16]);
  BUFF I151 (store_0n[17], ldata_0n[17]);
  BUFF I152 (store_0n[18], ldata_0n[18]);
  BUFF I153 (store_0n[19], ldata_0n[19]);
  BUFF I154 (store_0n[20], ldata_0n[20]);
  BUFF I155 (store_0n[21], ldata_0n[21]);
  BUFF I156 (store_0n[22], ldata_0n[22]);
  BUFF I157 (store_0n[23], ldata_0n[23]);
  BUFF I158 (store_0n[24], ldata_0n[24]);
  BUFF I159 (store_0n[25], ldata_0n[25]);
  BUFF I160 (store_0n[26], ldata_0n[26]);
  BUFF I161 (store_0n[27], ldata_0n[27]);
  BUFF I162 (store_0n[28], ldata_0n[28]);
  BUFF I163 (store_0n[29], ldata_0n[29]);
  BUFF I164 (store_0n[30], ldata_0n[30]);
  BUFF I165 (store_0n[31], ldata_0n[31]);
  BUFF I166 (store_0n[32], ldata_0n[32]);
  BUFF I167 (store_0n[33], ldata_0n[33]);
  BUFF I168 (store_0n[34], ldata_0n[34]);
  BUFF I169 (store_1n[0], ldata_1n[0]);
  BUFF I170 (store_1n[1], ldata_1n[1]);
  BUFF I171 (store_1n[2], ldata_1n[2]);
  BUFF I172 (store_1n[3], ldata_1n[3]);
  BUFF I173 (store_1n[4], ldata_1n[4]);
  BUFF I174 (store_1n[5], ldata_1n[5]);
  BUFF I175 (store_1n[6], ldata_1n[6]);
  BUFF I176 (store_1n[7], ldata_1n[7]);
  BUFF I177 (store_1n[8], ldata_1n[8]);
  BUFF I178 (store_1n[9], ldata_1n[9]);
  BUFF I179 (store_1n[10], ldata_1n[10]);
  BUFF I180 (store_1n[11], ldata_1n[11]);
  BUFF I181 (store_1n[12], ldata_1n[12]);
  BUFF I182 (store_1n[13], ldata_1n[13]);
  BUFF I183 (store_1n[14], ldata_1n[14]);
  BUFF I184 (store_1n[15], ldata_1n[15]);
  BUFF I185 (store_1n[16], ldata_1n[16]);
  BUFF I186 (store_1n[17], ldata_1n[17]);
  BUFF I187 (store_1n[18], ldata_1n[18]);
  BUFF I188 (store_1n[19], ldata_1n[19]);
  BUFF I189 (store_1n[20], ldata_1n[20]);
  BUFF I190 (store_1n[21], ldata_1n[21]);
  BUFF I191 (store_1n[22], ldata_1n[22]);
  BUFF I192 (store_1n[23], ldata_1n[23]);
  BUFF I193 (store_1n[24], ldata_1n[24]);
  BUFF I194 (store_1n[25], ldata_1n[25]);
  BUFF I195 (store_1n[26], ldata_1n[26]);
  BUFF I196 (store_1n[27], ldata_1n[27]);
  BUFF I197 (store_1n[28], ldata_1n[28]);
  BUFF I198 (store_1n[29], ldata_1n[29]);
  BUFF I199 (store_1n[30], ldata_1n[30]);
  BUFF I200 (store_1n[31], ldata_1n[31]);
  BUFF I201 (store_1n[32], ldata_1n[32]);
  BUFF I202 (store_1n[33], ldata_1n[33]);
  BUFF I203 (store_1n[34], ldata_1n[34]);
  C3 I204 (internal_0n[0], wack_0n[0], wack_0n[1], wack_0n[2]);
  C3 I205 (internal_0n[1], wack_0n[3], wack_0n[4], wack_0n[5]);
  C3 I206 (internal_0n[2], wack_0n[6], wack_0n[7], wack_0n[8]);
  C3 I207 (internal_0n[3], wack_0n[9], wack_0n[10], wack_0n[11]);
  C3 I208 (internal_0n[4], wack_0n[12], wack_0n[13], wack_0n[14]);
  C3 I209 (internal_0n[5], wack_0n[15], wack_0n[16], wack_0n[17]);
  C3 I210 (internal_0n[6], wack_0n[18], wack_0n[19], wack_0n[20]);
  C3 I211 (internal_0n[7], wack_0n[21], wack_0n[22], wack_0n[23]);
  C3 I212 (internal_0n[8], wack_0n[24], wack_0n[25], wack_0n[26]);
  C3 I213 (internal_0n[9], wack_0n[27], wack_0n[28], wack_0n[29]);
  C3 I214 (internal_0n[10], wack_0n[30], wack_0n[31], wack_0n[32]);
  C2 I215 (internal_0n[11], wack_0n[33], wack_0n[34]);
  C3 I216 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I217 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I218 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I219 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I220 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I221 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I222 (write_0a, internal_0n[16], internal_0n[17]);
  DRLATCH I223 (write_0r0d[0], write_0r1d[0], wack_0n[0], ldata_0n[0], ldata_1n[0]);
  DRLATCH I224 (write_0r0d[1], write_0r1d[1], wack_0n[1], ldata_0n[1], ldata_1n[1]);
  DRLATCH I225 (write_0r0d[2], write_0r1d[2], wack_0n[2], ldata_0n[2], ldata_1n[2]);
  DRLATCH I226 (write_0r0d[3], write_0r1d[3], wack_0n[3], ldata_0n[3], ldata_1n[3]);
  DRLATCH I227 (write_0r0d[4], write_0r1d[4], wack_0n[4], ldata_0n[4], ldata_1n[4]);
  DRLATCH I228 (write_0r0d[5], write_0r1d[5], wack_0n[5], ldata_0n[5], ldata_1n[5]);
  DRLATCH I229 (write_0r0d[6], write_0r1d[6], wack_0n[6], ldata_0n[6], ldata_1n[6]);
  DRLATCH I230 (write_0r0d[7], write_0r1d[7], wack_0n[7], ldata_0n[7], ldata_1n[7]);
  DRLATCH I231 (write_0r0d[8], write_0r1d[8], wack_0n[8], ldata_0n[8], ldata_1n[8]);
  DRLATCH I232 (write_0r0d[9], write_0r1d[9], wack_0n[9], ldata_0n[9], ldata_1n[9]);
  DRLATCH I233 (write_0r0d[10], write_0r1d[10], wack_0n[10], ldata_0n[10], ldata_1n[10]);
  DRLATCH I234 (write_0r0d[11], write_0r1d[11], wack_0n[11], ldata_0n[11], ldata_1n[11]);
  DRLATCH I235 (write_0r0d[12], write_0r1d[12], wack_0n[12], ldata_0n[12], ldata_1n[12]);
  DRLATCH I236 (write_0r0d[13], write_0r1d[13], wack_0n[13], ldata_0n[13], ldata_1n[13]);
  DRLATCH I237 (write_0r0d[14], write_0r1d[14], wack_0n[14], ldata_0n[14], ldata_1n[14]);
  DRLATCH I238 (write_0r0d[15], write_0r1d[15], wack_0n[15], ldata_0n[15], ldata_1n[15]);
  DRLATCH I239 (write_0r0d[16], write_0r1d[16], wack_0n[16], ldata_0n[16], ldata_1n[16]);
  DRLATCH I240 (write_0r0d[17], write_0r1d[17], wack_0n[17], ldata_0n[17], ldata_1n[17]);
  DRLATCH I241 (write_0r0d[18], write_0r1d[18], wack_0n[18], ldata_0n[18], ldata_1n[18]);
  DRLATCH I242 (write_0r0d[19], write_0r1d[19], wack_0n[19], ldata_0n[19], ldata_1n[19]);
  DRLATCH I243 (write_0r0d[20], write_0r1d[20], wack_0n[20], ldata_0n[20], ldata_1n[20]);
  DRLATCH I244 (write_0r0d[21], write_0r1d[21], wack_0n[21], ldata_0n[21], ldata_1n[21]);
  DRLATCH I245 (write_0r0d[22], write_0r1d[22], wack_0n[22], ldata_0n[22], ldata_1n[22]);
  DRLATCH I246 (write_0r0d[23], write_0r1d[23], wack_0n[23], ldata_0n[23], ldata_1n[23]);
  DRLATCH I247 (write_0r0d[24], write_0r1d[24], wack_0n[24], ldata_0n[24], ldata_1n[24]);
  DRLATCH I248 (write_0r0d[25], write_0r1d[25], wack_0n[25], ldata_0n[25], ldata_1n[25]);
  DRLATCH I249 (write_0r0d[26], write_0r1d[26], wack_0n[26], ldata_0n[26], ldata_1n[26]);
  DRLATCH I250 (write_0r0d[27], write_0r1d[27], wack_0n[27], ldata_0n[27], ldata_1n[27]);
  DRLATCH I251 (write_0r0d[28], write_0r1d[28], wack_0n[28], ldata_0n[28], ldata_1n[28]);
  DRLATCH I252 (write_0r0d[29], write_0r1d[29], wack_0n[29], ldata_0n[29], ldata_1n[29]);
  DRLATCH I253 (write_0r0d[30], write_0r1d[30], wack_0n[30], ldata_0n[30], ldata_1n[30]);
  DRLATCH I254 (write_0r0d[31], write_0r1d[31], wack_0n[31], ldata_0n[31], ldata_1n[31]);
  DRLATCH I255 (write_0r0d[32], write_0r1d[32], wack_0n[32], ldata_0n[32], ldata_1n[32]);
  DRLATCH I256 (write_0r0d[33], write_0r1d[33], wack_0n[33], ldata_0n[33], ldata_1n[33]);
  DRLATCH I257 (write_0r0d[34], write_0r1d[34], wack_0n[34], ldata_0n[34], ldata_1n[34]);
endmodule

module BrzVariable_35_4_s47_2_2e_2e34_3b34_2e_2e3_m29m (
  write_0r0d, write_0r1d, write_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d,
  read_2r, read_2a0d, read_2a1d,
  read_3r, read_3a0d, read_3a1d
);
  input [34:0] write_0r0d;
  input [34:0] write_0r1d;
  output write_0a;
  input read_0r;
  output [32:0] read_0a0d;
  output [32:0] read_0a1d;
  input read_1r;
  output read_1a0d;
  output read_1a1d;
  input read_2r;
  output read_2a0d;
  output read_2a1d;
  input read_3r;
  output [31:0] read_3a0d;
  output [31:0] read_3a1d;
  wire [17:0] internal_0n;
  wire [34:0] store_0n;
  wire [34:0] store_1n;
  wire [34:0] ldata_0n;
  wire [34:0] ldata_1n;
  wire [34:0] wack_0n;
  wire readReq_0n;
  wire readReq_1n;
  wire readReq_2n;
  wire readReq_3n;
  AND2 I0 (read_3a1d[0], store_1n[1], readReq_3n);
  AND2 I1 (read_3a1d[1], store_1n[2], readReq_3n);
  AND2 I2 (read_3a1d[2], store_1n[3], readReq_3n);
  AND2 I3 (read_3a1d[3], store_1n[4], readReq_3n);
  AND2 I4 (read_3a1d[4], store_1n[5], readReq_3n);
  AND2 I5 (read_3a1d[5], store_1n[6], readReq_3n);
  AND2 I6 (read_3a1d[6], store_1n[7], readReq_3n);
  AND2 I7 (read_3a1d[7], store_1n[8], readReq_3n);
  AND2 I8 (read_3a1d[8], store_1n[9], readReq_3n);
  AND2 I9 (read_3a1d[9], store_1n[10], readReq_3n);
  AND2 I10 (read_3a1d[10], store_1n[11], readReq_3n);
  AND2 I11 (read_3a1d[11], store_1n[12], readReq_3n);
  AND2 I12 (read_3a1d[12], store_1n[13], readReq_3n);
  AND2 I13 (read_3a1d[13], store_1n[14], readReq_3n);
  AND2 I14 (read_3a1d[14], store_1n[15], readReq_3n);
  AND2 I15 (read_3a1d[15], store_1n[16], readReq_3n);
  AND2 I16 (read_3a1d[16], store_1n[17], readReq_3n);
  AND2 I17 (read_3a1d[17], store_1n[18], readReq_3n);
  AND2 I18 (read_3a1d[18], store_1n[19], readReq_3n);
  AND2 I19 (read_3a1d[19], store_1n[20], readReq_3n);
  AND2 I20 (read_3a1d[20], store_1n[21], readReq_3n);
  AND2 I21 (read_3a1d[21], store_1n[22], readReq_3n);
  AND2 I22 (read_3a1d[22], store_1n[23], readReq_3n);
  AND2 I23 (read_3a1d[23], store_1n[24], readReq_3n);
  AND2 I24 (read_3a1d[24], store_1n[25], readReq_3n);
  AND2 I25 (read_3a1d[25], store_1n[26], readReq_3n);
  AND2 I26 (read_3a1d[26], store_1n[27], readReq_3n);
  AND2 I27 (read_3a1d[27], store_1n[28], readReq_3n);
  AND2 I28 (read_3a1d[28], store_1n[29], readReq_3n);
  AND2 I29 (read_3a1d[29], store_1n[30], readReq_3n);
  AND2 I30 (read_3a1d[30], store_1n[31], readReq_3n);
  AND2 I31 (read_3a1d[31], store_1n[32], readReq_3n);
  AND2 I32 (read_3a0d[0], store_0n[1], readReq_3n);
  AND2 I33 (read_3a0d[1], store_0n[2], readReq_3n);
  AND2 I34 (read_3a0d[2], store_0n[3], readReq_3n);
  AND2 I35 (read_3a0d[3], store_0n[4], readReq_3n);
  AND2 I36 (read_3a0d[4], store_0n[5], readReq_3n);
  AND2 I37 (read_3a0d[5], store_0n[6], readReq_3n);
  AND2 I38 (read_3a0d[6], store_0n[7], readReq_3n);
  AND2 I39 (read_3a0d[7], store_0n[8], readReq_3n);
  AND2 I40 (read_3a0d[8], store_0n[9], readReq_3n);
  AND2 I41 (read_3a0d[9], store_0n[10], readReq_3n);
  AND2 I42 (read_3a0d[10], store_0n[11], readReq_3n);
  AND2 I43 (read_3a0d[11], store_0n[12], readReq_3n);
  AND2 I44 (read_3a0d[12], store_0n[13], readReq_3n);
  AND2 I45 (read_3a0d[13], store_0n[14], readReq_3n);
  AND2 I46 (read_3a0d[14], store_0n[15], readReq_3n);
  AND2 I47 (read_3a0d[15], store_0n[16], readReq_3n);
  AND2 I48 (read_3a0d[16], store_0n[17], readReq_3n);
  AND2 I49 (read_3a0d[17], store_0n[18], readReq_3n);
  AND2 I50 (read_3a0d[18], store_0n[19], readReq_3n);
  AND2 I51 (read_3a0d[19], store_0n[20], readReq_3n);
  AND2 I52 (read_3a0d[20], store_0n[21], readReq_3n);
  AND2 I53 (read_3a0d[21], store_0n[22], readReq_3n);
  AND2 I54 (read_3a0d[22], store_0n[23], readReq_3n);
  AND2 I55 (read_3a0d[23], store_0n[24], readReq_3n);
  AND2 I56 (read_3a0d[24], store_0n[25], readReq_3n);
  AND2 I57 (read_3a0d[25], store_0n[26], readReq_3n);
  AND2 I58 (read_3a0d[26], store_0n[27], readReq_3n);
  AND2 I59 (read_3a0d[27], store_0n[28], readReq_3n);
  AND2 I60 (read_3a0d[28], store_0n[29], readReq_3n);
  AND2 I61 (read_3a0d[29], store_0n[30], readReq_3n);
  AND2 I62 (read_3a0d[30], store_0n[31], readReq_3n);
  AND2 I63 (read_3a0d[31], store_0n[32], readReq_3n);
  AND2 I64 (read_2a1d, store_1n[34], readReq_2n);
  AND2 I65 (read_2a0d, store_0n[34], readReq_2n);
  AND2 I66 (read_1a1d, store_1n[34], readReq_1n);
  AND2 I67 (read_1a0d, store_0n[34], readReq_1n);
  AND2 I68 (read_0a1d[0], store_1n[2], readReq_0n);
  AND2 I69 (read_0a1d[1], store_1n[3], readReq_0n);
  AND2 I70 (read_0a1d[2], store_1n[4], readReq_0n);
  AND2 I71 (read_0a1d[3], store_1n[5], readReq_0n);
  AND2 I72 (read_0a1d[4], store_1n[6], readReq_0n);
  AND2 I73 (read_0a1d[5], store_1n[7], readReq_0n);
  AND2 I74 (read_0a1d[6], store_1n[8], readReq_0n);
  AND2 I75 (read_0a1d[7], store_1n[9], readReq_0n);
  AND2 I76 (read_0a1d[8], store_1n[10], readReq_0n);
  AND2 I77 (read_0a1d[9], store_1n[11], readReq_0n);
  AND2 I78 (read_0a1d[10], store_1n[12], readReq_0n);
  AND2 I79 (read_0a1d[11], store_1n[13], readReq_0n);
  AND2 I80 (read_0a1d[12], store_1n[14], readReq_0n);
  AND2 I81 (read_0a1d[13], store_1n[15], readReq_0n);
  AND2 I82 (read_0a1d[14], store_1n[16], readReq_0n);
  AND2 I83 (read_0a1d[15], store_1n[17], readReq_0n);
  AND2 I84 (read_0a1d[16], store_1n[18], readReq_0n);
  AND2 I85 (read_0a1d[17], store_1n[19], readReq_0n);
  AND2 I86 (read_0a1d[18], store_1n[20], readReq_0n);
  AND2 I87 (read_0a1d[19], store_1n[21], readReq_0n);
  AND2 I88 (read_0a1d[20], store_1n[22], readReq_0n);
  AND2 I89 (read_0a1d[21], store_1n[23], readReq_0n);
  AND2 I90 (read_0a1d[22], store_1n[24], readReq_0n);
  AND2 I91 (read_0a1d[23], store_1n[25], readReq_0n);
  AND2 I92 (read_0a1d[24], store_1n[26], readReq_0n);
  AND2 I93 (read_0a1d[25], store_1n[27], readReq_0n);
  AND2 I94 (read_0a1d[26], store_1n[28], readReq_0n);
  AND2 I95 (read_0a1d[27], store_1n[29], readReq_0n);
  AND2 I96 (read_0a1d[28], store_1n[30], readReq_0n);
  AND2 I97 (read_0a1d[29], store_1n[31], readReq_0n);
  AND2 I98 (read_0a1d[30], store_1n[32], readReq_0n);
  AND2 I99 (read_0a1d[31], store_1n[33], readReq_0n);
  AND2 I100 (read_0a1d[32], store_1n[34], readReq_0n);
  AND2 I101 (read_0a0d[0], store_0n[2], readReq_0n);
  AND2 I102 (read_0a0d[1], store_0n[3], readReq_0n);
  AND2 I103 (read_0a0d[2], store_0n[4], readReq_0n);
  AND2 I104 (read_0a0d[3], store_0n[5], readReq_0n);
  AND2 I105 (read_0a0d[4], store_0n[6], readReq_0n);
  AND2 I106 (read_0a0d[5], store_0n[7], readReq_0n);
  AND2 I107 (read_0a0d[6], store_0n[8], readReq_0n);
  AND2 I108 (read_0a0d[7], store_0n[9], readReq_0n);
  AND2 I109 (read_0a0d[8], store_0n[10], readReq_0n);
  AND2 I110 (read_0a0d[9], store_0n[11], readReq_0n);
  AND2 I111 (read_0a0d[10], store_0n[12], readReq_0n);
  AND2 I112 (read_0a0d[11], store_0n[13], readReq_0n);
  AND2 I113 (read_0a0d[12], store_0n[14], readReq_0n);
  AND2 I114 (read_0a0d[13], store_0n[15], readReq_0n);
  AND2 I115 (read_0a0d[14], store_0n[16], readReq_0n);
  AND2 I116 (read_0a0d[15], store_0n[17], readReq_0n);
  AND2 I117 (read_0a0d[16], store_0n[18], readReq_0n);
  AND2 I118 (read_0a0d[17], store_0n[19], readReq_0n);
  AND2 I119 (read_0a0d[18], store_0n[20], readReq_0n);
  AND2 I120 (read_0a0d[19], store_0n[21], readReq_0n);
  AND2 I121 (read_0a0d[20], store_0n[22], readReq_0n);
  AND2 I122 (read_0a0d[21], store_0n[23], readReq_0n);
  AND2 I123 (read_0a0d[22], store_0n[24], readReq_0n);
  AND2 I124 (read_0a0d[23], store_0n[25], readReq_0n);
  AND2 I125 (read_0a0d[24], store_0n[26], readReq_0n);
  AND2 I126 (read_0a0d[25], store_0n[27], readReq_0n);
  AND2 I127 (read_0a0d[26], store_0n[28], readReq_0n);
  AND2 I128 (read_0a0d[27], store_0n[29], readReq_0n);
  AND2 I129 (read_0a0d[28], store_0n[30], readReq_0n);
  AND2 I130 (read_0a0d[29], store_0n[31], readReq_0n);
  AND2 I131 (read_0a0d[30], store_0n[32], readReq_0n);
  AND2 I132 (read_0a0d[31], store_0n[33], readReq_0n);
  AND2 I133 (read_0a0d[32], store_0n[34], readReq_0n);
  BUFF I134 (readReq_0n, read_0r);
  BUFF I135 (readReq_1n, read_1r);
  BUFF I136 (readReq_2n, read_2r);
  BUFF I137 (readReq_3n, read_3r);
  BUFF I138 (store_0n[0], ldata_0n[0]);
  BUFF I139 (store_0n[1], ldata_0n[1]);
  BUFF I140 (store_0n[2], ldata_0n[2]);
  BUFF I141 (store_0n[3], ldata_0n[3]);
  BUFF I142 (store_0n[4], ldata_0n[4]);
  BUFF I143 (store_0n[5], ldata_0n[5]);
  BUFF I144 (store_0n[6], ldata_0n[6]);
  BUFF I145 (store_0n[7], ldata_0n[7]);
  BUFF I146 (store_0n[8], ldata_0n[8]);
  BUFF I147 (store_0n[9], ldata_0n[9]);
  BUFF I148 (store_0n[10], ldata_0n[10]);
  BUFF I149 (store_0n[11], ldata_0n[11]);
  BUFF I150 (store_0n[12], ldata_0n[12]);
  BUFF I151 (store_0n[13], ldata_0n[13]);
  BUFF I152 (store_0n[14], ldata_0n[14]);
  BUFF I153 (store_0n[15], ldata_0n[15]);
  BUFF I154 (store_0n[16], ldata_0n[16]);
  BUFF I155 (store_0n[17], ldata_0n[17]);
  BUFF I156 (store_0n[18], ldata_0n[18]);
  BUFF I157 (store_0n[19], ldata_0n[19]);
  BUFF I158 (store_0n[20], ldata_0n[20]);
  BUFF I159 (store_0n[21], ldata_0n[21]);
  BUFF I160 (store_0n[22], ldata_0n[22]);
  BUFF I161 (store_0n[23], ldata_0n[23]);
  BUFF I162 (store_0n[24], ldata_0n[24]);
  BUFF I163 (store_0n[25], ldata_0n[25]);
  BUFF I164 (store_0n[26], ldata_0n[26]);
  BUFF I165 (store_0n[27], ldata_0n[27]);
  BUFF I166 (store_0n[28], ldata_0n[28]);
  BUFF I167 (store_0n[29], ldata_0n[29]);
  BUFF I168 (store_0n[30], ldata_0n[30]);
  BUFF I169 (store_0n[31], ldata_0n[31]);
  BUFF I170 (store_0n[32], ldata_0n[32]);
  BUFF I171 (store_0n[33], ldata_0n[33]);
  BUFF I172 (store_0n[34], ldata_0n[34]);
  BUFF I173 (store_1n[0], ldata_1n[0]);
  BUFF I174 (store_1n[1], ldata_1n[1]);
  BUFF I175 (store_1n[2], ldata_1n[2]);
  BUFF I176 (store_1n[3], ldata_1n[3]);
  BUFF I177 (store_1n[4], ldata_1n[4]);
  BUFF I178 (store_1n[5], ldata_1n[5]);
  BUFF I179 (store_1n[6], ldata_1n[6]);
  BUFF I180 (store_1n[7], ldata_1n[7]);
  BUFF I181 (store_1n[8], ldata_1n[8]);
  BUFF I182 (store_1n[9], ldata_1n[9]);
  BUFF I183 (store_1n[10], ldata_1n[10]);
  BUFF I184 (store_1n[11], ldata_1n[11]);
  BUFF I185 (store_1n[12], ldata_1n[12]);
  BUFF I186 (store_1n[13], ldata_1n[13]);
  BUFF I187 (store_1n[14], ldata_1n[14]);
  BUFF I188 (store_1n[15], ldata_1n[15]);
  BUFF I189 (store_1n[16], ldata_1n[16]);
  BUFF I190 (store_1n[17], ldata_1n[17]);
  BUFF I191 (store_1n[18], ldata_1n[18]);
  BUFF I192 (store_1n[19], ldata_1n[19]);
  BUFF I193 (store_1n[20], ldata_1n[20]);
  BUFF I194 (store_1n[21], ldata_1n[21]);
  BUFF I195 (store_1n[22], ldata_1n[22]);
  BUFF I196 (store_1n[23], ldata_1n[23]);
  BUFF I197 (store_1n[24], ldata_1n[24]);
  BUFF I198 (store_1n[25], ldata_1n[25]);
  BUFF I199 (store_1n[26], ldata_1n[26]);
  BUFF I200 (store_1n[27], ldata_1n[27]);
  BUFF I201 (store_1n[28], ldata_1n[28]);
  BUFF I202 (store_1n[29], ldata_1n[29]);
  BUFF I203 (store_1n[30], ldata_1n[30]);
  BUFF I204 (store_1n[31], ldata_1n[31]);
  BUFF I205 (store_1n[32], ldata_1n[32]);
  BUFF I206 (store_1n[33], ldata_1n[33]);
  BUFF I207 (store_1n[34], ldata_1n[34]);
  C3 I208 (internal_0n[0], wack_0n[0], wack_0n[1], wack_0n[2]);
  C3 I209 (internal_0n[1], wack_0n[3], wack_0n[4], wack_0n[5]);
  C3 I210 (internal_0n[2], wack_0n[6], wack_0n[7], wack_0n[8]);
  C3 I211 (internal_0n[3], wack_0n[9], wack_0n[10], wack_0n[11]);
  C3 I212 (internal_0n[4], wack_0n[12], wack_0n[13], wack_0n[14]);
  C3 I213 (internal_0n[5], wack_0n[15], wack_0n[16], wack_0n[17]);
  C3 I214 (internal_0n[6], wack_0n[18], wack_0n[19], wack_0n[20]);
  C3 I215 (internal_0n[7], wack_0n[21], wack_0n[22], wack_0n[23]);
  C3 I216 (internal_0n[8], wack_0n[24], wack_0n[25], wack_0n[26]);
  C3 I217 (internal_0n[9], wack_0n[27], wack_0n[28], wack_0n[29]);
  C3 I218 (internal_0n[10], wack_0n[30], wack_0n[31], wack_0n[32]);
  C2 I219 (internal_0n[11], wack_0n[33], wack_0n[34]);
  C3 I220 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I221 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I222 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I223 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I224 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I225 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I226 (write_0a, internal_0n[16], internal_0n[17]);
  DRLATCH I227 (write_0r0d[0], write_0r1d[0], wack_0n[0], ldata_0n[0], ldata_1n[0]);
  DRLATCH I228 (write_0r0d[1], write_0r1d[1], wack_0n[1], ldata_0n[1], ldata_1n[1]);
  DRLATCH I229 (write_0r0d[2], write_0r1d[2], wack_0n[2], ldata_0n[2], ldata_1n[2]);
  DRLATCH I230 (write_0r0d[3], write_0r1d[3], wack_0n[3], ldata_0n[3], ldata_1n[3]);
  DRLATCH I231 (write_0r0d[4], write_0r1d[4], wack_0n[4], ldata_0n[4], ldata_1n[4]);
  DRLATCH I232 (write_0r0d[5], write_0r1d[5], wack_0n[5], ldata_0n[5], ldata_1n[5]);
  DRLATCH I233 (write_0r0d[6], write_0r1d[6], wack_0n[6], ldata_0n[6], ldata_1n[6]);
  DRLATCH I234 (write_0r0d[7], write_0r1d[7], wack_0n[7], ldata_0n[7], ldata_1n[7]);
  DRLATCH I235 (write_0r0d[8], write_0r1d[8], wack_0n[8], ldata_0n[8], ldata_1n[8]);
  DRLATCH I236 (write_0r0d[9], write_0r1d[9], wack_0n[9], ldata_0n[9], ldata_1n[9]);
  DRLATCH I237 (write_0r0d[10], write_0r1d[10], wack_0n[10], ldata_0n[10], ldata_1n[10]);
  DRLATCH I238 (write_0r0d[11], write_0r1d[11], wack_0n[11], ldata_0n[11], ldata_1n[11]);
  DRLATCH I239 (write_0r0d[12], write_0r1d[12], wack_0n[12], ldata_0n[12], ldata_1n[12]);
  DRLATCH I240 (write_0r0d[13], write_0r1d[13], wack_0n[13], ldata_0n[13], ldata_1n[13]);
  DRLATCH I241 (write_0r0d[14], write_0r1d[14], wack_0n[14], ldata_0n[14], ldata_1n[14]);
  DRLATCH I242 (write_0r0d[15], write_0r1d[15], wack_0n[15], ldata_0n[15], ldata_1n[15]);
  DRLATCH I243 (write_0r0d[16], write_0r1d[16], wack_0n[16], ldata_0n[16], ldata_1n[16]);
  DRLATCH I244 (write_0r0d[17], write_0r1d[17], wack_0n[17], ldata_0n[17], ldata_1n[17]);
  DRLATCH I245 (write_0r0d[18], write_0r1d[18], wack_0n[18], ldata_0n[18], ldata_1n[18]);
  DRLATCH I246 (write_0r0d[19], write_0r1d[19], wack_0n[19], ldata_0n[19], ldata_1n[19]);
  DRLATCH I247 (write_0r0d[20], write_0r1d[20], wack_0n[20], ldata_0n[20], ldata_1n[20]);
  DRLATCH I248 (write_0r0d[21], write_0r1d[21], wack_0n[21], ldata_0n[21], ldata_1n[21]);
  DRLATCH I249 (write_0r0d[22], write_0r1d[22], wack_0n[22], ldata_0n[22], ldata_1n[22]);
  DRLATCH I250 (write_0r0d[23], write_0r1d[23], wack_0n[23], ldata_0n[23], ldata_1n[23]);
  DRLATCH I251 (write_0r0d[24], write_0r1d[24], wack_0n[24], ldata_0n[24], ldata_1n[24]);
  DRLATCH I252 (write_0r0d[25], write_0r1d[25], wack_0n[25], ldata_0n[25], ldata_1n[25]);
  DRLATCH I253 (write_0r0d[26], write_0r1d[26], wack_0n[26], ldata_0n[26], ldata_1n[26]);
  DRLATCH I254 (write_0r0d[27], write_0r1d[27], wack_0n[27], ldata_0n[27], ldata_1n[27]);
  DRLATCH I255 (write_0r0d[28], write_0r1d[28], wack_0n[28], ldata_0n[28], ldata_1n[28]);
  DRLATCH I256 (write_0r0d[29], write_0r1d[29], wack_0n[29], ldata_0n[29], ldata_1n[29]);
  DRLATCH I257 (write_0r0d[30], write_0r1d[30], wack_0n[30], ldata_0n[30], ldata_1n[30]);
  DRLATCH I258 (write_0r0d[31], write_0r1d[31], wack_0n[31], ldata_0n[31], ldata_1n[31]);
  DRLATCH I259 (write_0r0d[32], write_0r1d[32], wack_0n[32], ldata_0n[32], ldata_1n[32]);
  DRLATCH I260 (write_0r0d[33], write_0r1d[33], wack_0n[33], ldata_0n[33], ldata_1n[33]);
  DRLATCH I261 (write_0r0d[34], write_0r1d[34], wack_0n[34], ldata_0n[34], ldata_1n[34]);
endmodule

module BrzVariable_36_1_s9_3_2e_2e34 (
  write_0r0d, write_0r1d, write_0a,
  read_0r, read_0a0d, read_0a1d
);
  input [35:0] write_0r0d;
  input [35:0] write_0r1d;
  output write_0a;
  input read_0r;
  output [31:0] read_0a0d;
  output [31:0] read_0a1d;
  wire [17:0] internal_0n;
  wire [35:0] store_0n;
  wire [35:0] store_1n;
  wire [35:0] ldata_0n;
  wire [35:0] ldata_1n;
  wire [35:0] wack_0n;
  wire readReq_0n;
  AND2 I0 (read_0a1d[0], store_1n[3], readReq_0n);
  AND2 I1 (read_0a1d[1], store_1n[4], readReq_0n);
  AND2 I2 (read_0a1d[2], store_1n[5], readReq_0n);
  AND2 I3 (read_0a1d[3], store_1n[6], readReq_0n);
  AND2 I4 (read_0a1d[4], store_1n[7], readReq_0n);
  AND2 I5 (read_0a1d[5], store_1n[8], readReq_0n);
  AND2 I6 (read_0a1d[6], store_1n[9], readReq_0n);
  AND2 I7 (read_0a1d[7], store_1n[10], readReq_0n);
  AND2 I8 (read_0a1d[8], store_1n[11], readReq_0n);
  AND2 I9 (read_0a1d[9], store_1n[12], readReq_0n);
  AND2 I10 (read_0a1d[10], store_1n[13], readReq_0n);
  AND2 I11 (read_0a1d[11], store_1n[14], readReq_0n);
  AND2 I12 (read_0a1d[12], store_1n[15], readReq_0n);
  AND2 I13 (read_0a1d[13], store_1n[16], readReq_0n);
  AND2 I14 (read_0a1d[14], store_1n[17], readReq_0n);
  AND2 I15 (read_0a1d[15], store_1n[18], readReq_0n);
  AND2 I16 (read_0a1d[16], store_1n[19], readReq_0n);
  AND2 I17 (read_0a1d[17], store_1n[20], readReq_0n);
  AND2 I18 (read_0a1d[18], store_1n[21], readReq_0n);
  AND2 I19 (read_0a1d[19], store_1n[22], readReq_0n);
  AND2 I20 (read_0a1d[20], store_1n[23], readReq_0n);
  AND2 I21 (read_0a1d[21], store_1n[24], readReq_0n);
  AND2 I22 (read_0a1d[22], store_1n[25], readReq_0n);
  AND2 I23 (read_0a1d[23], store_1n[26], readReq_0n);
  AND2 I24 (read_0a1d[24], store_1n[27], readReq_0n);
  AND2 I25 (read_0a1d[25], store_1n[28], readReq_0n);
  AND2 I26 (read_0a1d[26], store_1n[29], readReq_0n);
  AND2 I27 (read_0a1d[27], store_1n[30], readReq_0n);
  AND2 I28 (read_0a1d[28], store_1n[31], readReq_0n);
  AND2 I29 (read_0a1d[29], store_1n[32], readReq_0n);
  AND2 I30 (read_0a1d[30], store_1n[33], readReq_0n);
  AND2 I31 (read_0a1d[31], store_1n[34], readReq_0n);
  AND2 I32 (read_0a0d[0], store_0n[3], readReq_0n);
  AND2 I33 (read_0a0d[1], store_0n[4], readReq_0n);
  AND2 I34 (read_0a0d[2], store_0n[5], readReq_0n);
  AND2 I35 (read_0a0d[3], store_0n[6], readReq_0n);
  AND2 I36 (read_0a0d[4], store_0n[7], readReq_0n);
  AND2 I37 (read_0a0d[5], store_0n[8], readReq_0n);
  AND2 I38 (read_0a0d[6], store_0n[9], readReq_0n);
  AND2 I39 (read_0a0d[7], store_0n[10], readReq_0n);
  AND2 I40 (read_0a0d[8], store_0n[11], readReq_0n);
  AND2 I41 (read_0a0d[9], store_0n[12], readReq_0n);
  AND2 I42 (read_0a0d[10], store_0n[13], readReq_0n);
  AND2 I43 (read_0a0d[11], store_0n[14], readReq_0n);
  AND2 I44 (read_0a0d[12], store_0n[15], readReq_0n);
  AND2 I45 (read_0a0d[13], store_0n[16], readReq_0n);
  AND2 I46 (read_0a0d[14], store_0n[17], readReq_0n);
  AND2 I47 (read_0a0d[15], store_0n[18], readReq_0n);
  AND2 I48 (read_0a0d[16], store_0n[19], readReq_0n);
  AND2 I49 (read_0a0d[17], store_0n[20], readReq_0n);
  AND2 I50 (read_0a0d[18], store_0n[21], readReq_0n);
  AND2 I51 (read_0a0d[19], store_0n[22], readReq_0n);
  AND2 I52 (read_0a0d[20], store_0n[23], readReq_0n);
  AND2 I53 (read_0a0d[21], store_0n[24], readReq_0n);
  AND2 I54 (read_0a0d[22], store_0n[25], readReq_0n);
  AND2 I55 (read_0a0d[23], store_0n[26], readReq_0n);
  AND2 I56 (read_0a0d[24], store_0n[27], readReq_0n);
  AND2 I57 (read_0a0d[25], store_0n[28], readReq_0n);
  AND2 I58 (read_0a0d[26], store_0n[29], readReq_0n);
  AND2 I59 (read_0a0d[27], store_0n[30], readReq_0n);
  AND2 I60 (read_0a0d[28], store_0n[31], readReq_0n);
  AND2 I61 (read_0a0d[29], store_0n[32], readReq_0n);
  AND2 I62 (read_0a0d[30], store_0n[33], readReq_0n);
  AND2 I63 (read_0a0d[31], store_0n[34], readReq_0n);
  BUFF I64 (readReq_0n, read_0r);
  BUFF I65 (store_0n[0], ldata_0n[0]);
  BUFF I66 (store_0n[1], ldata_0n[1]);
  BUFF I67 (store_0n[2], ldata_0n[2]);
  BUFF I68 (store_0n[3], ldata_0n[3]);
  BUFF I69 (store_0n[4], ldata_0n[4]);
  BUFF I70 (store_0n[5], ldata_0n[5]);
  BUFF I71 (store_0n[6], ldata_0n[6]);
  BUFF I72 (store_0n[7], ldata_0n[7]);
  BUFF I73 (store_0n[8], ldata_0n[8]);
  BUFF I74 (store_0n[9], ldata_0n[9]);
  BUFF I75 (store_0n[10], ldata_0n[10]);
  BUFF I76 (store_0n[11], ldata_0n[11]);
  BUFF I77 (store_0n[12], ldata_0n[12]);
  BUFF I78 (store_0n[13], ldata_0n[13]);
  BUFF I79 (store_0n[14], ldata_0n[14]);
  BUFF I80 (store_0n[15], ldata_0n[15]);
  BUFF I81 (store_0n[16], ldata_0n[16]);
  BUFF I82 (store_0n[17], ldata_0n[17]);
  BUFF I83 (store_0n[18], ldata_0n[18]);
  BUFF I84 (store_0n[19], ldata_0n[19]);
  BUFF I85 (store_0n[20], ldata_0n[20]);
  BUFF I86 (store_0n[21], ldata_0n[21]);
  BUFF I87 (store_0n[22], ldata_0n[22]);
  BUFF I88 (store_0n[23], ldata_0n[23]);
  BUFF I89 (store_0n[24], ldata_0n[24]);
  BUFF I90 (store_0n[25], ldata_0n[25]);
  BUFF I91 (store_0n[26], ldata_0n[26]);
  BUFF I92 (store_0n[27], ldata_0n[27]);
  BUFF I93 (store_0n[28], ldata_0n[28]);
  BUFF I94 (store_0n[29], ldata_0n[29]);
  BUFF I95 (store_0n[30], ldata_0n[30]);
  BUFF I96 (store_0n[31], ldata_0n[31]);
  BUFF I97 (store_0n[32], ldata_0n[32]);
  BUFF I98 (store_0n[33], ldata_0n[33]);
  BUFF I99 (store_0n[34], ldata_0n[34]);
  BUFF I100 (store_0n[35], ldata_0n[35]);
  BUFF I101 (store_1n[0], ldata_1n[0]);
  BUFF I102 (store_1n[1], ldata_1n[1]);
  BUFF I103 (store_1n[2], ldata_1n[2]);
  BUFF I104 (store_1n[3], ldata_1n[3]);
  BUFF I105 (store_1n[4], ldata_1n[4]);
  BUFF I106 (store_1n[5], ldata_1n[5]);
  BUFF I107 (store_1n[6], ldata_1n[6]);
  BUFF I108 (store_1n[7], ldata_1n[7]);
  BUFF I109 (store_1n[8], ldata_1n[8]);
  BUFF I110 (store_1n[9], ldata_1n[9]);
  BUFF I111 (store_1n[10], ldata_1n[10]);
  BUFF I112 (store_1n[11], ldata_1n[11]);
  BUFF I113 (store_1n[12], ldata_1n[12]);
  BUFF I114 (store_1n[13], ldata_1n[13]);
  BUFF I115 (store_1n[14], ldata_1n[14]);
  BUFF I116 (store_1n[15], ldata_1n[15]);
  BUFF I117 (store_1n[16], ldata_1n[16]);
  BUFF I118 (store_1n[17], ldata_1n[17]);
  BUFF I119 (store_1n[18], ldata_1n[18]);
  BUFF I120 (store_1n[19], ldata_1n[19]);
  BUFF I121 (store_1n[20], ldata_1n[20]);
  BUFF I122 (store_1n[21], ldata_1n[21]);
  BUFF I123 (store_1n[22], ldata_1n[22]);
  BUFF I124 (store_1n[23], ldata_1n[23]);
  BUFF I125 (store_1n[24], ldata_1n[24]);
  BUFF I126 (store_1n[25], ldata_1n[25]);
  BUFF I127 (store_1n[26], ldata_1n[26]);
  BUFF I128 (store_1n[27], ldata_1n[27]);
  BUFF I129 (store_1n[28], ldata_1n[28]);
  BUFF I130 (store_1n[29], ldata_1n[29]);
  BUFF I131 (store_1n[30], ldata_1n[30]);
  BUFF I132 (store_1n[31], ldata_1n[31]);
  BUFF I133 (store_1n[32], ldata_1n[32]);
  BUFF I134 (store_1n[33], ldata_1n[33]);
  BUFF I135 (store_1n[34], ldata_1n[34]);
  BUFF I136 (store_1n[35], ldata_1n[35]);
  C3 I137 (internal_0n[0], wack_0n[0], wack_0n[1], wack_0n[2]);
  C3 I138 (internal_0n[1], wack_0n[3], wack_0n[4], wack_0n[5]);
  C3 I139 (internal_0n[2], wack_0n[6], wack_0n[7], wack_0n[8]);
  C3 I140 (internal_0n[3], wack_0n[9], wack_0n[10], wack_0n[11]);
  C3 I141 (internal_0n[4], wack_0n[12], wack_0n[13], wack_0n[14]);
  C3 I142 (internal_0n[5], wack_0n[15], wack_0n[16], wack_0n[17]);
  C3 I143 (internal_0n[6], wack_0n[18], wack_0n[19], wack_0n[20]);
  C3 I144 (internal_0n[7], wack_0n[21], wack_0n[22], wack_0n[23]);
  C3 I145 (internal_0n[8], wack_0n[24], wack_0n[25], wack_0n[26]);
  C3 I146 (internal_0n[9], wack_0n[27], wack_0n[28], wack_0n[29]);
  C3 I147 (internal_0n[10], wack_0n[30], wack_0n[31], wack_0n[32]);
  C3 I148 (internal_0n[11], wack_0n[33], wack_0n[34], wack_0n[35]);
  C3 I149 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I150 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I151 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I152 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I153 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I154 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I155 (write_0a, internal_0n[16], internal_0n[17]);
  DRLATCH I156 (write_0r0d[0], write_0r1d[0], wack_0n[0], ldata_0n[0], ldata_1n[0]);
  DRLATCH I157 (write_0r0d[1], write_0r1d[1], wack_0n[1], ldata_0n[1], ldata_1n[1]);
  DRLATCH I158 (write_0r0d[2], write_0r1d[2], wack_0n[2], ldata_0n[2], ldata_1n[2]);
  DRLATCH I159 (write_0r0d[3], write_0r1d[3], wack_0n[3], ldata_0n[3], ldata_1n[3]);
  DRLATCH I160 (write_0r0d[4], write_0r1d[4], wack_0n[4], ldata_0n[4], ldata_1n[4]);
  DRLATCH I161 (write_0r0d[5], write_0r1d[5], wack_0n[5], ldata_0n[5], ldata_1n[5]);
  DRLATCH I162 (write_0r0d[6], write_0r1d[6], wack_0n[6], ldata_0n[6], ldata_1n[6]);
  DRLATCH I163 (write_0r0d[7], write_0r1d[7], wack_0n[7], ldata_0n[7], ldata_1n[7]);
  DRLATCH I164 (write_0r0d[8], write_0r1d[8], wack_0n[8], ldata_0n[8], ldata_1n[8]);
  DRLATCH I165 (write_0r0d[9], write_0r1d[9], wack_0n[9], ldata_0n[9], ldata_1n[9]);
  DRLATCH I166 (write_0r0d[10], write_0r1d[10], wack_0n[10], ldata_0n[10], ldata_1n[10]);
  DRLATCH I167 (write_0r0d[11], write_0r1d[11], wack_0n[11], ldata_0n[11], ldata_1n[11]);
  DRLATCH I168 (write_0r0d[12], write_0r1d[12], wack_0n[12], ldata_0n[12], ldata_1n[12]);
  DRLATCH I169 (write_0r0d[13], write_0r1d[13], wack_0n[13], ldata_0n[13], ldata_1n[13]);
  DRLATCH I170 (write_0r0d[14], write_0r1d[14], wack_0n[14], ldata_0n[14], ldata_1n[14]);
  DRLATCH I171 (write_0r0d[15], write_0r1d[15], wack_0n[15], ldata_0n[15], ldata_1n[15]);
  DRLATCH I172 (write_0r0d[16], write_0r1d[16], wack_0n[16], ldata_0n[16], ldata_1n[16]);
  DRLATCH I173 (write_0r0d[17], write_0r1d[17], wack_0n[17], ldata_0n[17], ldata_1n[17]);
  DRLATCH I174 (write_0r0d[18], write_0r1d[18], wack_0n[18], ldata_0n[18], ldata_1n[18]);
  DRLATCH I175 (write_0r0d[19], write_0r1d[19], wack_0n[19], ldata_0n[19], ldata_1n[19]);
  DRLATCH I176 (write_0r0d[20], write_0r1d[20], wack_0n[20], ldata_0n[20], ldata_1n[20]);
  DRLATCH I177 (write_0r0d[21], write_0r1d[21], wack_0n[21], ldata_0n[21], ldata_1n[21]);
  DRLATCH I178 (write_0r0d[22], write_0r1d[22], wack_0n[22], ldata_0n[22], ldata_1n[22]);
  DRLATCH I179 (write_0r0d[23], write_0r1d[23], wack_0n[23], ldata_0n[23], ldata_1n[23]);
  DRLATCH I180 (write_0r0d[24], write_0r1d[24], wack_0n[24], ldata_0n[24], ldata_1n[24]);
  DRLATCH I181 (write_0r0d[25], write_0r1d[25], wack_0n[25], ldata_0n[25], ldata_1n[25]);
  DRLATCH I182 (write_0r0d[26], write_0r1d[26], wack_0n[26], ldata_0n[26], ldata_1n[26]);
  DRLATCH I183 (write_0r0d[27], write_0r1d[27], wack_0n[27], ldata_0n[27], ldata_1n[27]);
  DRLATCH I184 (write_0r0d[28], write_0r1d[28], wack_0n[28], ldata_0n[28], ldata_1n[28]);
  DRLATCH I185 (write_0r0d[29], write_0r1d[29], wack_0n[29], ldata_0n[29], ldata_1n[29]);
  DRLATCH I186 (write_0r0d[30], write_0r1d[30], wack_0n[30], ldata_0n[30], ldata_1n[30]);
  DRLATCH I187 (write_0r0d[31], write_0r1d[31], wack_0n[31], ldata_0n[31], ldata_1n[31]);
  DRLATCH I188 (write_0r0d[32], write_0r1d[32], wack_0n[32], ldata_0n[32], ldata_1n[32]);
  DRLATCH I189 (write_0r0d[33], write_0r1d[33], wack_0n[33], ldata_0n[33], ldata_1n[33]);
  DRLATCH I190 (write_0r0d[34], write_0r1d[34], wack_0n[34], ldata_0n[34], ldata_1n[34]);
  DRLATCH I191 (write_0r0d[35], write_0r1d[35], wack_0n[35], ldata_0n[35], ldata_1n[35]);
endmodule

module BrzVariable_36_2_s12__3b2_2e_2e33 (
  write_0r0d, write_0r1d, write_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d
);
  input [35:0] write_0r0d;
  input [35:0] write_0r1d;
  output write_0a;
  input read_0r;
  output [35:0] read_0a0d;
  output [35:0] read_0a1d;
  input read_1r;
  output [31:0] read_1a0d;
  output [31:0] read_1a1d;
  wire [17:0] internal_0n;
  wire [35:0] store_0n;
  wire [35:0] store_1n;
  wire [35:0] ldata_0n;
  wire [35:0] ldata_1n;
  wire [35:0] wack_0n;
  wire readReq_0n;
  wire readReq_1n;
  AND2 I0 (read_1a1d[0], store_1n[2], readReq_1n);
  AND2 I1 (read_1a1d[1], store_1n[3], readReq_1n);
  AND2 I2 (read_1a1d[2], store_1n[4], readReq_1n);
  AND2 I3 (read_1a1d[3], store_1n[5], readReq_1n);
  AND2 I4 (read_1a1d[4], store_1n[6], readReq_1n);
  AND2 I5 (read_1a1d[5], store_1n[7], readReq_1n);
  AND2 I6 (read_1a1d[6], store_1n[8], readReq_1n);
  AND2 I7 (read_1a1d[7], store_1n[9], readReq_1n);
  AND2 I8 (read_1a1d[8], store_1n[10], readReq_1n);
  AND2 I9 (read_1a1d[9], store_1n[11], readReq_1n);
  AND2 I10 (read_1a1d[10], store_1n[12], readReq_1n);
  AND2 I11 (read_1a1d[11], store_1n[13], readReq_1n);
  AND2 I12 (read_1a1d[12], store_1n[14], readReq_1n);
  AND2 I13 (read_1a1d[13], store_1n[15], readReq_1n);
  AND2 I14 (read_1a1d[14], store_1n[16], readReq_1n);
  AND2 I15 (read_1a1d[15], store_1n[17], readReq_1n);
  AND2 I16 (read_1a1d[16], store_1n[18], readReq_1n);
  AND2 I17 (read_1a1d[17], store_1n[19], readReq_1n);
  AND2 I18 (read_1a1d[18], store_1n[20], readReq_1n);
  AND2 I19 (read_1a1d[19], store_1n[21], readReq_1n);
  AND2 I20 (read_1a1d[20], store_1n[22], readReq_1n);
  AND2 I21 (read_1a1d[21], store_1n[23], readReq_1n);
  AND2 I22 (read_1a1d[22], store_1n[24], readReq_1n);
  AND2 I23 (read_1a1d[23], store_1n[25], readReq_1n);
  AND2 I24 (read_1a1d[24], store_1n[26], readReq_1n);
  AND2 I25 (read_1a1d[25], store_1n[27], readReq_1n);
  AND2 I26 (read_1a1d[26], store_1n[28], readReq_1n);
  AND2 I27 (read_1a1d[27], store_1n[29], readReq_1n);
  AND2 I28 (read_1a1d[28], store_1n[30], readReq_1n);
  AND2 I29 (read_1a1d[29], store_1n[31], readReq_1n);
  AND2 I30 (read_1a1d[30], store_1n[32], readReq_1n);
  AND2 I31 (read_1a1d[31], store_1n[33], readReq_1n);
  AND2 I32 (read_1a0d[0], store_0n[2], readReq_1n);
  AND2 I33 (read_1a0d[1], store_0n[3], readReq_1n);
  AND2 I34 (read_1a0d[2], store_0n[4], readReq_1n);
  AND2 I35 (read_1a0d[3], store_0n[5], readReq_1n);
  AND2 I36 (read_1a0d[4], store_0n[6], readReq_1n);
  AND2 I37 (read_1a0d[5], store_0n[7], readReq_1n);
  AND2 I38 (read_1a0d[6], store_0n[8], readReq_1n);
  AND2 I39 (read_1a0d[7], store_0n[9], readReq_1n);
  AND2 I40 (read_1a0d[8], store_0n[10], readReq_1n);
  AND2 I41 (read_1a0d[9], store_0n[11], readReq_1n);
  AND2 I42 (read_1a0d[10], store_0n[12], readReq_1n);
  AND2 I43 (read_1a0d[11], store_0n[13], readReq_1n);
  AND2 I44 (read_1a0d[12], store_0n[14], readReq_1n);
  AND2 I45 (read_1a0d[13], store_0n[15], readReq_1n);
  AND2 I46 (read_1a0d[14], store_0n[16], readReq_1n);
  AND2 I47 (read_1a0d[15], store_0n[17], readReq_1n);
  AND2 I48 (read_1a0d[16], store_0n[18], readReq_1n);
  AND2 I49 (read_1a0d[17], store_0n[19], readReq_1n);
  AND2 I50 (read_1a0d[18], store_0n[20], readReq_1n);
  AND2 I51 (read_1a0d[19], store_0n[21], readReq_1n);
  AND2 I52 (read_1a0d[20], store_0n[22], readReq_1n);
  AND2 I53 (read_1a0d[21], store_0n[23], readReq_1n);
  AND2 I54 (read_1a0d[22], store_0n[24], readReq_1n);
  AND2 I55 (read_1a0d[23], store_0n[25], readReq_1n);
  AND2 I56 (read_1a0d[24], store_0n[26], readReq_1n);
  AND2 I57 (read_1a0d[25], store_0n[27], readReq_1n);
  AND2 I58 (read_1a0d[26], store_0n[28], readReq_1n);
  AND2 I59 (read_1a0d[27], store_0n[29], readReq_1n);
  AND2 I60 (read_1a0d[28], store_0n[30], readReq_1n);
  AND2 I61 (read_1a0d[29], store_0n[31], readReq_1n);
  AND2 I62 (read_1a0d[30], store_0n[32], readReq_1n);
  AND2 I63 (read_1a0d[31], store_0n[33], readReq_1n);
  AND2 I64 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I65 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I66 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I67 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I68 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I69 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I70 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I71 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I72 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I73 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I74 (read_0a1d[10], store_1n[10], readReq_0n);
  AND2 I75 (read_0a1d[11], store_1n[11], readReq_0n);
  AND2 I76 (read_0a1d[12], store_1n[12], readReq_0n);
  AND2 I77 (read_0a1d[13], store_1n[13], readReq_0n);
  AND2 I78 (read_0a1d[14], store_1n[14], readReq_0n);
  AND2 I79 (read_0a1d[15], store_1n[15], readReq_0n);
  AND2 I80 (read_0a1d[16], store_1n[16], readReq_0n);
  AND2 I81 (read_0a1d[17], store_1n[17], readReq_0n);
  AND2 I82 (read_0a1d[18], store_1n[18], readReq_0n);
  AND2 I83 (read_0a1d[19], store_1n[19], readReq_0n);
  AND2 I84 (read_0a1d[20], store_1n[20], readReq_0n);
  AND2 I85 (read_0a1d[21], store_1n[21], readReq_0n);
  AND2 I86 (read_0a1d[22], store_1n[22], readReq_0n);
  AND2 I87 (read_0a1d[23], store_1n[23], readReq_0n);
  AND2 I88 (read_0a1d[24], store_1n[24], readReq_0n);
  AND2 I89 (read_0a1d[25], store_1n[25], readReq_0n);
  AND2 I90 (read_0a1d[26], store_1n[26], readReq_0n);
  AND2 I91 (read_0a1d[27], store_1n[27], readReq_0n);
  AND2 I92 (read_0a1d[28], store_1n[28], readReq_0n);
  AND2 I93 (read_0a1d[29], store_1n[29], readReq_0n);
  AND2 I94 (read_0a1d[30], store_1n[30], readReq_0n);
  AND2 I95 (read_0a1d[31], store_1n[31], readReq_0n);
  AND2 I96 (read_0a1d[32], store_1n[32], readReq_0n);
  AND2 I97 (read_0a1d[33], store_1n[33], readReq_0n);
  AND2 I98 (read_0a1d[34], store_1n[34], readReq_0n);
  AND2 I99 (read_0a1d[35], store_1n[35], readReq_0n);
  AND2 I100 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I101 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I102 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I103 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I104 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I105 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I106 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I107 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I108 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I109 (read_0a0d[9], store_0n[9], readReq_0n);
  AND2 I110 (read_0a0d[10], store_0n[10], readReq_0n);
  AND2 I111 (read_0a0d[11], store_0n[11], readReq_0n);
  AND2 I112 (read_0a0d[12], store_0n[12], readReq_0n);
  AND2 I113 (read_0a0d[13], store_0n[13], readReq_0n);
  AND2 I114 (read_0a0d[14], store_0n[14], readReq_0n);
  AND2 I115 (read_0a0d[15], store_0n[15], readReq_0n);
  AND2 I116 (read_0a0d[16], store_0n[16], readReq_0n);
  AND2 I117 (read_0a0d[17], store_0n[17], readReq_0n);
  AND2 I118 (read_0a0d[18], store_0n[18], readReq_0n);
  AND2 I119 (read_0a0d[19], store_0n[19], readReq_0n);
  AND2 I120 (read_0a0d[20], store_0n[20], readReq_0n);
  AND2 I121 (read_0a0d[21], store_0n[21], readReq_0n);
  AND2 I122 (read_0a0d[22], store_0n[22], readReq_0n);
  AND2 I123 (read_0a0d[23], store_0n[23], readReq_0n);
  AND2 I124 (read_0a0d[24], store_0n[24], readReq_0n);
  AND2 I125 (read_0a0d[25], store_0n[25], readReq_0n);
  AND2 I126 (read_0a0d[26], store_0n[26], readReq_0n);
  AND2 I127 (read_0a0d[27], store_0n[27], readReq_0n);
  AND2 I128 (read_0a0d[28], store_0n[28], readReq_0n);
  AND2 I129 (read_0a0d[29], store_0n[29], readReq_0n);
  AND2 I130 (read_0a0d[30], store_0n[30], readReq_0n);
  AND2 I131 (read_0a0d[31], store_0n[31], readReq_0n);
  AND2 I132 (read_0a0d[32], store_0n[32], readReq_0n);
  AND2 I133 (read_0a0d[33], store_0n[33], readReq_0n);
  AND2 I134 (read_0a0d[34], store_0n[34], readReq_0n);
  AND2 I135 (read_0a0d[35], store_0n[35], readReq_0n);
  BUFF I136 (readReq_0n, read_0r);
  BUFF I137 (readReq_1n, read_1r);
  BUFF I138 (store_0n[0], ldata_0n[0]);
  BUFF I139 (store_0n[1], ldata_0n[1]);
  BUFF I140 (store_0n[2], ldata_0n[2]);
  BUFF I141 (store_0n[3], ldata_0n[3]);
  BUFF I142 (store_0n[4], ldata_0n[4]);
  BUFF I143 (store_0n[5], ldata_0n[5]);
  BUFF I144 (store_0n[6], ldata_0n[6]);
  BUFF I145 (store_0n[7], ldata_0n[7]);
  BUFF I146 (store_0n[8], ldata_0n[8]);
  BUFF I147 (store_0n[9], ldata_0n[9]);
  BUFF I148 (store_0n[10], ldata_0n[10]);
  BUFF I149 (store_0n[11], ldata_0n[11]);
  BUFF I150 (store_0n[12], ldata_0n[12]);
  BUFF I151 (store_0n[13], ldata_0n[13]);
  BUFF I152 (store_0n[14], ldata_0n[14]);
  BUFF I153 (store_0n[15], ldata_0n[15]);
  BUFF I154 (store_0n[16], ldata_0n[16]);
  BUFF I155 (store_0n[17], ldata_0n[17]);
  BUFF I156 (store_0n[18], ldata_0n[18]);
  BUFF I157 (store_0n[19], ldata_0n[19]);
  BUFF I158 (store_0n[20], ldata_0n[20]);
  BUFF I159 (store_0n[21], ldata_0n[21]);
  BUFF I160 (store_0n[22], ldata_0n[22]);
  BUFF I161 (store_0n[23], ldata_0n[23]);
  BUFF I162 (store_0n[24], ldata_0n[24]);
  BUFF I163 (store_0n[25], ldata_0n[25]);
  BUFF I164 (store_0n[26], ldata_0n[26]);
  BUFF I165 (store_0n[27], ldata_0n[27]);
  BUFF I166 (store_0n[28], ldata_0n[28]);
  BUFF I167 (store_0n[29], ldata_0n[29]);
  BUFF I168 (store_0n[30], ldata_0n[30]);
  BUFF I169 (store_0n[31], ldata_0n[31]);
  BUFF I170 (store_0n[32], ldata_0n[32]);
  BUFF I171 (store_0n[33], ldata_0n[33]);
  BUFF I172 (store_0n[34], ldata_0n[34]);
  BUFF I173 (store_0n[35], ldata_0n[35]);
  BUFF I174 (store_1n[0], ldata_1n[0]);
  BUFF I175 (store_1n[1], ldata_1n[1]);
  BUFF I176 (store_1n[2], ldata_1n[2]);
  BUFF I177 (store_1n[3], ldata_1n[3]);
  BUFF I178 (store_1n[4], ldata_1n[4]);
  BUFF I179 (store_1n[5], ldata_1n[5]);
  BUFF I180 (store_1n[6], ldata_1n[6]);
  BUFF I181 (store_1n[7], ldata_1n[7]);
  BUFF I182 (store_1n[8], ldata_1n[8]);
  BUFF I183 (store_1n[9], ldata_1n[9]);
  BUFF I184 (store_1n[10], ldata_1n[10]);
  BUFF I185 (store_1n[11], ldata_1n[11]);
  BUFF I186 (store_1n[12], ldata_1n[12]);
  BUFF I187 (store_1n[13], ldata_1n[13]);
  BUFF I188 (store_1n[14], ldata_1n[14]);
  BUFF I189 (store_1n[15], ldata_1n[15]);
  BUFF I190 (store_1n[16], ldata_1n[16]);
  BUFF I191 (store_1n[17], ldata_1n[17]);
  BUFF I192 (store_1n[18], ldata_1n[18]);
  BUFF I193 (store_1n[19], ldata_1n[19]);
  BUFF I194 (store_1n[20], ldata_1n[20]);
  BUFF I195 (store_1n[21], ldata_1n[21]);
  BUFF I196 (store_1n[22], ldata_1n[22]);
  BUFF I197 (store_1n[23], ldata_1n[23]);
  BUFF I198 (store_1n[24], ldata_1n[24]);
  BUFF I199 (store_1n[25], ldata_1n[25]);
  BUFF I200 (store_1n[26], ldata_1n[26]);
  BUFF I201 (store_1n[27], ldata_1n[27]);
  BUFF I202 (store_1n[28], ldata_1n[28]);
  BUFF I203 (store_1n[29], ldata_1n[29]);
  BUFF I204 (store_1n[30], ldata_1n[30]);
  BUFF I205 (store_1n[31], ldata_1n[31]);
  BUFF I206 (store_1n[32], ldata_1n[32]);
  BUFF I207 (store_1n[33], ldata_1n[33]);
  BUFF I208 (store_1n[34], ldata_1n[34]);
  BUFF I209 (store_1n[35], ldata_1n[35]);
  C3 I210 (internal_0n[0], wack_0n[0], wack_0n[1], wack_0n[2]);
  C3 I211 (internal_0n[1], wack_0n[3], wack_0n[4], wack_0n[5]);
  C3 I212 (internal_0n[2], wack_0n[6], wack_0n[7], wack_0n[8]);
  C3 I213 (internal_0n[3], wack_0n[9], wack_0n[10], wack_0n[11]);
  C3 I214 (internal_0n[4], wack_0n[12], wack_0n[13], wack_0n[14]);
  C3 I215 (internal_0n[5], wack_0n[15], wack_0n[16], wack_0n[17]);
  C3 I216 (internal_0n[6], wack_0n[18], wack_0n[19], wack_0n[20]);
  C3 I217 (internal_0n[7], wack_0n[21], wack_0n[22], wack_0n[23]);
  C3 I218 (internal_0n[8], wack_0n[24], wack_0n[25], wack_0n[26]);
  C3 I219 (internal_0n[9], wack_0n[27], wack_0n[28], wack_0n[29]);
  C3 I220 (internal_0n[10], wack_0n[30], wack_0n[31], wack_0n[32]);
  C3 I221 (internal_0n[11], wack_0n[33], wack_0n[34], wack_0n[35]);
  C3 I222 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I223 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I224 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I225 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I226 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I227 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I228 (write_0a, internal_0n[16], internal_0n[17]);
  DRLATCH I229 (write_0r0d[0], write_0r1d[0], wack_0n[0], ldata_0n[0], ldata_1n[0]);
  DRLATCH I230 (write_0r0d[1], write_0r1d[1], wack_0n[1], ldata_0n[1], ldata_1n[1]);
  DRLATCH I231 (write_0r0d[2], write_0r1d[2], wack_0n[2], ldata_0n[2], ldata_1n[2]);
  DRLATCH I232 (write_0r0d[3], write_0r1d[3], wack_0n[3], ldata_0n[3], ldata_1n[3]);
  DRLATCH I233 (write_0r0d[4], write_0r1d[4], wack_0n[4], ldata_0n[4], ldata_1n[4]);
  DRLATCH I234 (write_0r0d[5], write_0r1d[5], wack_0n[5], ldata_0n[5], ldata_1n[5]);
  DRLATCH I235 (write_0r0d[6], write_0r1d[6], wack_0n[6], ldata_0n[6], ldata_1n[6]);
  DRLATCH I236 (write_0r0d[7], write_0r1d[7], wack_0n[7], ldata_0n[7], ldata_1n[7]);
  DRLATCH I237 (write_0r0d[8], write_0r1d[8], wack_0n[8], ldata_0n[8], ldata_1n[8]);
  DRLATCH I238 (write_0r0d[9], write_0r1d[9], wack_0n[9], ldata_0n[9], ldata_1n[9]);
  DRLATCH I239 (write_0r0d[10], write_0r1d[10], wack_0n[10], ldata_0n[10], ldata_1n[10]);
  DRLATCH I240 (write_0r0d[11], write_0r1d[11], wack_0n[11], ldata_0n[11], ldata_1n[11]);
  DRLATCH I241 (write_0r0d[12], write_0r1d[12], wack_0n[12], ldata_0n[12], ldata_1n[12]);
  DRLATCH I242 (write_0r0d[13], write_0r1d[13], wack_0n[13], ldata_0n[13], ldata_1n[13]);
  DRLATCH I243 (write_0r0d[14], write_0r1d[14], wack_0n[14], ldata_0n[14], ldata_1n[14]);
  DRLATCH I244 (write_0r0d[15], write_0r1d[15], wack_0n[15], ldata_0n[15], ldata_1n[15]);
  DRLATCH I245 (write_0r0d[16], write_0r1d[16], wack_0n[16], ldata_0n[16], ldata_1n[16]);
  DRLATCH I246 (write_0r0d[17], write_0r1d[17], wack_0n[17], ldata_0n[17], ldata_1n[17]);
  DRLATCH I247 (write_0r0d[18], write_0r1d[18], wack_0n[18], ldata_0n[18], ldata_1n[18]);
  DRLATCH I248 (write_0r0d[19], write_0r1d[19], wack_0n[19], ldata_0n[19], ldata_1n[19]);
  DRLATCH I249 (write_0r0d[20], write_0r1d[20], wack_0n[20], ldata_0n[20], ldata_1n[20]);
  DRLATCH I250 (write_0r0d[21], write_0r1d[21], wack_0n[21], ldata_0n[21], ldata_1n[21]);
  DRLATCH I251 (write_0r0d[22], write_0r1d[22], wack_0n[22], ldata_0n[22], ldata_1n[22]);
  DRLATCH I252 (write_0r0d[23], write_0r1d[23], wack_0n[23], ldata_0n[23], ldata_1n[23]);
  DRLATCH I253 (write_0r0d[24], write_0r1d[24], wack_0n[24], ldata_0n[24], ldata_1n[24]);
  DRLATCH I254 (write_0r0d[25], write_0r1d[25], wack_0n[25], ldata_0n[25], ldata_1n[25]);
  DRLATCH I255 (write_0r0d[26], write_0r1d[26], wack_0n[26], ldata_0n[26], ldata_1n[26]);
  DRLATCH I256 (write_0r0d[27], write_0r1d[27], wack_0n[27], ldata_0n[27], ldata_1n[27]);
  DRLATCH I257 (write_0r0d[28], write_0r1d[28], wack_0n[28], ldata_0n[28], ldata_1n[28]);
  DRLATCH I258 (write_0r0d[29], write_0r1d[29], wack_0n[29], ldata_0n[29], ldata_1n[29]);
  DRLATCH I259 (write_0r0d[30], write_0r1d[30], wack_0n[30], ldata_0n[30], ldata_1n[30]);
  DRLATCH I260 (write_0r0d[31], write_0r1d[31], wack_0n[31], ldata_0n[31], ldata_1n[31]);
  DRLATCH I261 (write_0r0d[32], write_0r1d[32], wack_0n[32], ldata_0n[32], ldata_1n[32]);
  DRLATCH I262 (write_0r0d[33], write_0r1d[33], wack_0n[33], ldata_0n[33], ldata_1n[33]);
  DRLATCH I263 (write_0r0d[34], write_0r1d[34], wack_0n[34], ldata_0n[34], ldata_1n[34]);
  DRLATCH I264 (write_0r0d[35], write_0r1d[35], wack_0n[35], ldata_0n[35], ldata_1n[35]);
endmodule

module BrzVariable_36_4_s36__3b0_2e_2e3_3b2_2e_2e_m31m (
  write_0r0d, write_0r1d, write_0a,
  read_0r, read_0a0d, read_0a1d,
  read_1r, read_1a0d, read_1a1d,
  read_2r, read_2a0d, read_2a1d,
  read_3r, read_3a0d, read_3a1d
);
  input [35:0] write_0r0d;
  input [35:0] write_0r1d;
  output write_0a;
  input read_0r;
  output [35:0] read_0a0d;
  output [35:0] read_0a1d;
  input read_1r;
  output [3:0] read_1a0d;
  output [3:0] read_1a1d;
  input read_2r;
  output [31:0] read_2a0d;
  output [31:0] read_2a1d;
  input read_3r;
  output read_3a0d;
  output read_3a1d;
  wire [17:0] internal_0n;
  wire [35:0] store_0n;
  wire [35:0] store_1n;
  wire [35:0] ldata_0n;
  wire [35:0] ldata_1n;
  wire [35:0] wack_0n;
  wire readReq_0n;
  wire readReq_1n;
  wire readReq_2n;
  wire readReq_3n;
  AND2 I0 (read_3a1d, store_1n[34], readReq_3n);
  AND2 I1 (read_3a0d, store_0n[34], readReq_3n);
  AND2 I2 (read_2a1d[0], store_1n[2], readReq_2n);
  AND2 I3 (read_2a1d[1], store_1n[3], readReq_2n);
  AND2 I4 (read_2a1d[2], store_1n[4], readReq_2n);
  AND2 I5 (read_2a1d[3], store_1n[5], readReq_2n);
  AND2 I6 (read_2a1d[4], store_1n[6], readReq_2n);
  AND2 I7 (read_2a1d[5], store_1n[7], readReq_2n);
  AND2 I8 (read_2a1d[6], store_1n[8], readReq_2n);
  AND2 I9 (read_2a1d[7], store_1n[9], readReq_2n);
  AND2 I10 (read_2a1d[8], store_1n[10], readReq_2n);
  AND2 I11 (read_2a1d[9], store_1n[11], readReq_2n);
  AND2 I12 (read_2a1d[10], store_1n[12], readReq_2n);
  AND2 I13 (read_2a1d[11], store_1n[13], readReq_2n);
  AND2 I14 (read_2a1d[12], store_1n[14], readReq_2n);
  AND2 I15 (read_2a1d[13], store_1n[15], readReq_2n);
  AND2 I16 (read_2a1d[14], store_1n[16], readReq_2n);
  AND2 I17 (read_2a1d[15], store_1n[17], readReq_2n);
  AND2 I18 (read_2a1d[16], store_1n[18], readReq_2n);
  AND2 I19 (read_2a1d[17], store_1n[19], readReq_2n);
  AND2 I20 (read_2a1d[18], store_1n[20], readReq_2n);
  AND2 I21 (read_2a1d[19], store_1n[21], readReq_2n);
  AND2 I22 (read_2a1d[20], store_1n[22], readReq_2n);
  AND2 I23 (read_2a1d[21], store_1n[23], readReq_2n);
  AND2 I24 (read_2a1d[22], store_1n[24], readReq_2n);
  AND2 I25 (read_2a1d[23], store_1n[25], readReq_2n);
  AND2 I26 (read_2a1d[24], store_1n[26], readReq_2n);
  AND2 I27 (read_2a1d[25], store_1n[27], readReq_2n);
  AND2 I28 (read_2a1d[26], store_1n[28], readReq_2n);
  AND2 I29 (read_2a1d[27], store_1n[29], readReq_2n);
  AND2 I30 (read_2a1d[28], store_1n[30], readReq_2n);
  AND2 I31 (read_2a1d[29], store_1n[31], readReq_2n);
  AND2 I32 (read_2a1d[30], store_1n[32], readReq_2n);
  AND2 I33 (read_2a1d[31], store_1n[33], readReq_2n);
  AND2 I34 (read_2a0d[0], store_0n[2], readReq_2n);
  AND2 I35 (read_2a0d[1], store_0n[3], readReq_2n);
  AND2 I36 (read_2a0d[2], store_0n[4], readReq_2n);
  AND2 I37 (read_2a0d[3], store_0n[5], readReq_2n);
  AND2 I38 (read_2a0d[4], store_0n[6], readReq_2n);
  AND2 I39 (read_2a0d[5], store_0n[7], readReq_2n);
  AND2 I40 (read_2a0d[6], store_0n[8], readReq_2n);
  AND2 I41 (read_2a0d[7], store_0n[9], readReq_2n);
  AND2 I42 (read_2a0d[8], store_0n[10], readReq_2n);
  AND2 I43 (read_2a0d[9], store_0n[11], readReq_2n);
  AND2 I44 (read_2a0d[10], store_0n[12], readReq_2n);
  AND2 I45 (read_2a0d[11], store_0n[13], readReq_2n);
  AND2 I46 (read_2a0d[12], store_0n[14], readReq_2n);
  AND2 I47 (read_2a0d[13], store_0n[15], readReq_2n);
  AND2 I48 (read_2a0d[14], store_0n[16], readReq_2n);
  AND2 I49 (read_2a0d[15], store_0n[17], readReq_2n);
  AND2 I50 (read_2a0d[16], store_0n[18], readReq_2n);
  AND2 I51 (read_2a0d[17], store_0n[19], readReq_2n);
  AND2 I52 (read_2a0d[18], store_0n[20], readReq_2n);
  AND2 I53 (read_2a0d[19], store_0n[21], readReq_2n);
  AND2 I54 (read_2a0d[20], store_0n[22], readReq_2n);
  AND2 I55 (read_2a0d[21], store_0n[23], readReq_2n);
  AND2 I56 (read_2a0d[22], store_0n[24], readReq_2n);
  AND2 I57 (read_2a0d[23], store_0n[25], readReq_2n);
  AND2 I58 (read_2a0d[24], store_0n[26], readReq_2n);
  AND2 I59 (read_2a0d[25], store_0n[27], readReq_2n);
  AND2 I60 (read_2a0d[26], store_0n[28], readReq_2n);
  AND2 I61 (read_2a0d[27], store_0n[29], readReq_2n);
  AND2 I62 (read_2a0d[28], store_0n[30], readReq_2n);
  AND2 I63 (read_2a0d[29], store_0n[31], readReq_2n);
  AND2 I64 (read_2a0d[30], store_0n[32], readReq_2n);
  AND2 I65 (read_2a0d[31], store_0n[33], readReq_2n);
  AND2 I66 (read_1a1d[0], store_1n[0], readReq_1n);
  AND2 I67 (read_1a1d[1], store_1n[1], readReq_1n);
  AND2 I68 (read_1a1d[2], store_1n[2], readReq_1n);
  AND2 I69 (read_1a1d[3], store_1n[3], readReq_1n);
  AND2 I70 (read_1a0d[0], store_0n[0], readReq_1n);
  AND2 I71 (read_1a0d[1], store_0n[1], readReq_1n);
  AND2 I72 (read_1a0d[2], store_0n[2], readReq_1n);
  AND2 I73 (read_1a0d[3], store_0n[3], readReq_1n);
  AND2 I74 (read_0a1d[0], store_1n[0], readReq_0n);
  AND2 I75 (read_0a1d[1], store_1n[1], readReq_0n);
  AND2 I76 (read_0a1d[2], store_1n[2], readReq_0n);
  AND2 I77 (read_0a1d[3], store_1n[3], readReq_0n);
  AND2 I78 (read_0a1d[4], store_1n[4], readReq_0n);
  AND2 I79 (read_0a1d[5], store_1n[5], readReq_0n);
  AND2 I80 (read_0a1d[6], store_1n[6], readReq_0n);
  AND2 I81 (read_0a1d[7], store_1n[7], readReq_0n);
  AND2 I82 (read_0a1d[8], store_1n[8], readReq_0n);
  AND2 I83 (read_0a1d[9], store_1n[9], readReq_0n);
  AND2 I84 (read_0a1d[10], store_1n[10], readReq_0n);
  AND2 I85 (read_0a1d[11], store_1n[11], readReq_0n);
  AND2 I86 (read_0a1d[12], store_1n[12], readReq_0n);
  AND2 I87 (read_0a1d[13], store_1n[13], readReq_0n);
  AND2 I88 (read_0a1d[14], store_1n[14], readReq_0n);
  AND2 I89 (read_0a1d[15], store_1n[15], readReq_0n);
  AND2 I90 (read_0a1d[16], store_1n[16], readReq_0n);
  AND2 I91 (read_0a1d[17], store_1n[17], readReq_0n);
  AND2 I92 (read_0a1d[18], store_1n[18], readReq_0n);
  AND2 I93 (read_0a1d[19], store_1n[19], readReq_0n);
  AND2 I94 (read_0a1d[20], store_1n[20], readReq_0n);
  AND2 I95 (read_0a1d[21], store_1n[21], readReq_0n);
  AND2 I96 (read_0a1d[22], store_1n[22], readReq_0n);
  AND2 I97 (read_0a1d[23], store_1n[23], readReq_0n);
  AND2 I98 (read_0a1d[24], store_1n[24], readReq_0n);
  AND2 I99 (read_0a1d[25], store_1n[25], readReq_0n);
  AND2 I100 (read_0a1d[26], store_1n[26], readReq_0n);
  AND2 I101 (read_0a1d[27], store_1n[27], readReq_0n);
  AND2 I102 (read_0a1d[28], store_1n[28], readReq_0n);
  AND2 I103 (read_0a1d[29], store_1n[29], readReq_0n);
  AND2 I104 (read_0a1d[30], store_1n[30], readReq_0n);
  AND2 I105 (read_0a1d[31], store_1n[31], readReq_0n);
  AND2 I106 (read_0a1d[32], store_1n[32], readReq_0n);
  AND2 I107 (read_0a1d[33], store_1n[33], readReq_0n);
  AND2 I108 (read_0a1d[34], store_1n[34], readReq_0n);
  AND2 I109 (read_0a1d[35], store_1n[35], readReq_0n);
  AND2 I110 (read_0a0d[0], store_0n[0], readReq_0n);
  AND2 I111 (read_0a0d[1], store_0n[1], readReq_0n);
  AND2 I112 (read_0a0d[2], store_0n[2], readReq_0n);
  AND2 I113 (read_0a0d[3], store_0n[3], readReq_0n);
  AND2 I114 (read_0a0d[4], store_0n[4], readReq_0n);
  AND2 I115 (read_0a0d[5], store_0n[5], readReq_0n);
  AND2 I116 (read_0a0d[6], store_0n[6], readReq_0n);
  AND2 I117 (read_0a0d[7], store_0n[7], readReq_0n);
  AND2 I118 (read_0a0d[8], store_0n[8], readReq_0n);
  AND2 I119 (read_0a0d[9], store_0n[9], readReq_0n);
  AND2 I120 (read_0a0d[10], store_0n[10], readReq_0n);
  AND2 I121 (read_0a0d[11], store_0n[11], readReq_0n);
  AND2 I122 (read_0a0d[12], store_0n[12], readReq_0n);
  AND2 I123 (read_0a0d[13], store_0n[13], readReq_0n);
  AND2 I124 (read_0a0d[14], store_0n[14], readReq_0n);
  AND2 I125 (read_0a0d[15], store_0n[15], readReq_0n);
  AND2 I126 (read_0a0d[16], store_0n[16], readReq_0n);
  AND2 I127 (read_0a0d[17], store_0n[17], readReq_0n);
  AND2 I128 (read_0a0d[18], store_0n[18], readReq_0n);
  AND2 I129 (read_0a0d[19], store_0n[19], readReq_0n);
  AND2 I130 (read_0a0d[20], store_0n[20], readReq_0n);
  AND2 I131 (read_0a0d[21], store_0n[21], readReq_0n);
  AND2 I132 (read_0a0d[22], store_0n[22], readReq_0n);
  AND2 I133 (read_0a0d[23], store_0n[23], readReq_0n);
  AND2 I134 (read_0a0d[24], store_0n[24], readReq_0n);
  AND2 I135 (read_0a0d[25], store_0n[25], readReq_0n);
  AND2 I136 (read_0a0d[26], store_0n[26], readReq_0n);
  AND2 I137 (read_0a0d[27], store_0n[27], readReq_0n);
  AND2 I138 (read_0a0d[28], store_0n[28], readReq_0n);
  AND2 I139 (read_0a0d[29], store_0n[29], readReq_0n);
  AND2 I140 (read_0a0d[30], store_0n[30], readReq_0n);
  AND2 I141 (read_0a0d[31], store_0n[31], readReq_0n);
  AND2 I142 (read_0a0d[32], store_0n[32], readReq_0n);
  AND2 I143 (read_0a0d[33], store_0n[33], readReq_0n);
  AND2 I144 (read_0a0d[34], store_0n[34], readReq_0n);
  AND2 I145 (read_0a0d[35], store_0n[35], readReq_0n);
  BUFF I146 (readReq_0n, read_0r);
  BUFF I147 (readReq_1n, read_1r);
  BUFF I148 (readReq_2n, read_2r);
  BUFF I149 (readReq_3n, read_3r);
  BUFF I150 (store_0n[0], ldata_0n[0]);
  BUFF I151 (store_0n[1], ldata_0n[1]);
  BUFF I152 (store_0n[2], ldata_0n[2]);
  BUFF I153 (store_0n[3], ldata_0n[3]);
  BUFF I154 (store_0n[4], ldata_0n[4]);
  BUFF I155 (store_0n[5], ldata_0n[5]);
  BUFF I156 (store_0n[6], ldata_0n[6]);
  BUFF I157 (store_0n[7], ldata_0n[7]);
  BUFF I158 (store_0n[8], ldata_0n[8]);
  BUFF I159 (store_0n[9], ldata_0n[9]);
  BUFF I160 (store_0n[10], ldata_0n[10]);
  BUFF I161 (store_0n[11], ldata_0n[11]);
  BUFF I162 (store_0n[12], ldata_0n[12]);
  BUFF I163 (store_0n[13], ldata_0n[13]);
  BUFF I164 (store_0n[14], ldata_0n[14]);
  BUFF I165 (store_0n[15], ldata_0n[15]);
  BUFF I166 (store_0n[16], ldata_0n[16]);
  BUFF I167 (store_0n[17], ldata_0n[17]);
  BUFF I168 (store_0n[18], ldata_0n[18]);
  BUFF I169 (store_0n[19], ldata_0n[19]);
  BUFF I170 (store_0n[20], ldata_0n[20]);
  BUFF I171 (store_0n[21], ldata_0n[21]);
  BUFF I172 (store_0n[22], ldata_0n[22]);
  BUFF I173 (store_0n[23], ldata_0n[23]);
  BUFF I174 (store_0n[24], ldata_0n[24]);
  BUFF I175 (store_0n[25], ldata_0n[25]);
  BUFF I176 (store_0n[26], ldata_0n[26]);
  BUFF I177 (store_0n[27], ldata_0n[27]);
  BUFF I178 (store_0n[28], ldata_0n[28]);
  BUFF I179 (store_0n[29], ldata_0n[29]);
  BUFF I180 (store_0n[30], ldata_0n[30]);
  BUFF I181 (store_0n[31], ldata_0n[31]);
  BUFF I182 (store_0n[32], ldata_0n[32]);
  BUFF I183 (store_0n[33], ldata_0n[33]);
  BUFF I184 (store_0n[34], ldata_0n[34]);
  BUFF I185 (store_0n[35], ldata_0n[35]);
  BUFF I186 (store_1n[0], ldata_1n[0]);
  BUFF I187 (store_1n[1], ldata_1n[1]);
  BUFF I188 (store_1n[2], ldata_1n[2]);
  BUFF I189 (store_1n[3], ldata_1n[3]);
  BUFF I190 (store_1n[4], ldata_1n[4]);
  BUFF I191 (store_1n[5], ldata_1n[5]);
  BUFF I192 (store_1n[6], ldata_1n[6]);
  BUFF I193 (store_1n[7], ldata_1n[7]);
  BUFF I194 (store_1n[8], ldata_1n[8]);
  BUFF I195 (store_1n[9], ldata_1n[9]);
  BUFF I196 (store_1n[10], ldata_1n[10]);
  BUFF I197 (store_1n[11], ldata_1n[11]);
  BUFF I198 (store_1n[12], ldata_1n[12]);
  BUFF I199 (store_1n[13], ldata_1n[13]);
  BUFF I200 (store_1n[14], ldata_1n[14]);
  BUFF I201 (store_1n[15], ldata_1n[15]);
  BUFF I202 (store_1n[16], ldata_1n[16]);
  BUFF I203 (store_1n[17], ldata_1n[17]);
  BUFF I204 (store_1n[18], ldata_1n[18]);
  BUFF I205 (store_1n[19], ldata_1n[19]);
  BUFF I206 (store_1n[20], ldata_1n[20]);
  BUFF I207 (store_1n[21], ldata_1n[21]);
  BUFF I208 (store_1n[22], ldata_1n[22]);
  BUFF I209 (store_1n[23], ldata_1n[23]);
  BUFF I210 (store_1n[24], ldata_1n[24]);
  BUFF I211 (store_1n[25], ldata_1n[25]);
  BUFF I212 (store_1n[26], ldata_1n[26]);
  BUFF I213 (store_1n[27], ldata_1n[27]);
  BUFF I214 (store_1n[28], ldata_1n[28]);
  BUFF I215 (store_1n[29], ldata_1n[29]);
  BUFF I216 (store_1n[30], ldata_1n[30]);
  BUFF I217 (store_1n[31], ldata_1n[31]);
  BUFF I218 (store_1n[32], ldata_1n[32]);
  BUFF I219 (store_1n[33], ldata_1n[33]);
  BUFF I220 (store_1n[34], ldata_1n[34]);
  BUFF I221 (store_1n[35], ldata_1n[35]);
  C3 I222 (internal_0n[0], wack_0n[0], wack_0n[1], wack_0n[2]);
  C3 I223 (internal_0n[1], wack_0n[3], wack_0n[4], wack_0n[5]);
  C3 I224 (internal_0n[2], wack_0n[6], wack_0n[7], wack_0n[8]);
  C3 I225 (internal_0n[3], wack_0n[9], wack_0n[10], wack_0n[11]);
  C3 I226 (internal_0n[4], wack_0n[12], wack_0n[13], wack_0n[14]);
  C3 I227 (internal_0n[5], wack_0n[15], wack_0n[16], wack_0n[17]);
  C3 I228 (internal_0n[6], wack_0n[18], wack_0n[19], wack_0n[20]);
  C3 I229 (internal_0n[7], wack_0n[21], wack_0n[22], wack_0n[23]);
  C3 I230 (internal_0n[8], wack_0n[24], wack_0n[25], wack_0n[26]);
  C3 I231 (internal_0n[9], wack_0n[27], wack_0n[28], wack_0n[29]);
  C3 I232 (internal_0n[10], wack_0n[30], wack_0n[31], wack_0n[32]);
  C3 I233 (internal_0n[11], wack_0n[33], wack_0n[34], wack_0n[35]);
  C3 I234 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I235 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I236 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I237 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I238 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I239 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I240 (write_0a, internal_0n[16], internal_0n[17]);
  DRLATCH I241 (write_0r0d[0], write_0r1d[0], wack_0n[0], ldata_0n[0], ldata_1n[0]);
  DRLATCH I242 (write_0r0d[1], write_0r1d[1], wack_0n[1], ldata_0n[1], ldata_1n[1]);
  DRLATCH I243 (write_0r0d[2], write_0r1d[2], wack_0n[2], ldata_0n[2], ldata_1n[2]);
  DRLATCH I244 (write_0r0d[3], write_0r1d[3], wack_0n[3], ldata_0n[3], ldata_1n[3]);
  DRLATCH I245 (write_0r0d[4], write_0r1d[4], wack_0n[4], ldata_0n[4], ldata_1n[4]);
  DRLATCH I246 (write_0r0d[5], write_0r1d[5], wack_0n[5], ldata_0n[5], ldata_1n[5]);
  DRLATCH I247 (write_0r0d[6], write_0r1d[6], wack_0n[6], ldata_0n[6], ldata_1n[6]);
  DRLATCH I248 (write_0r0d[7], write_0r1d[7], wack_0n[7], ldata_0n[7], ldata_1n[7]);
  DRLATCH I249 (write_0r0d[8], write_0r1d[8], wack_0n[8], ldata_0n[8], ldata_1n[8]);
  DRLATCH I250 (write_0r0d[9], write_0r1d[9], wack_0n[9], ldata_0n[9], ldata_1n[9]);
  DRLATCH I251 (write_0r0d[10], write_0r1d[10], wack_0n[10], ldata_0n[10], ldata_1n[10]);
  DRLATCH I252 (write_0r0d[11], write_0r1d[11], wack_0n[11], ldata_0n[11], ldata_1n[11]);
  DRLATCH I253 (write_0r0d[12], write_0r1d[12], wack_0n[12], ldata_0n[12], ldata_1n[12]);
  DRLATCH I254 (write_0r0d[13], write_0r1d[13], wack_0n[13], ldata_0n[13], ldata_1n[13]);
  DRLATCH I255 (write_0r0d[14], write_0r1d[14], wack_0n[14], ldata_0n[14], ldata_1n[14]);
  DRLATCH I256 (write_0r0d[15], write_0r1d[15], wack_0n[15], ldata_0n[15], ldata_1n[15]);
  DRLATCH I257 (write_0r0d[16], write_0r1d[16], wack_0n[16], ldata_0n[16], ldata_1n[16]);
  DRLATCH I258 (write_0r0d[17], write_0r1d[17], wack_0n[17], ldata_0n[17], ldata_1n[17]);
  DRLATCH I259 (write_0r0d[18], write_0r1d[18], wack_0n[18], ldata_0n[18], ldata_1n[18]);
  DRLATCH I260 (write_0r0d[19], write_0r1d[19], wack_0n[19], ldata_0n[19], ldata_1n[19]);
  DRLATCH I261 (write_0r0d[20], write_0r1d[20], wack_0n[20], ldata_0n[20], ldata_1n[20]);
  DRLATCH I262 (write_0r0d[21], write_0r1d[21], wack_0n[21], ldata_0n[21], ldata_1n[21]);
  DRLATCH I263 (write_0r0d[22], write_0r1d[22], wack_0n[22], ldata_0n[22], ldata_1n[22]);
  DRLATCH I264 (write_0r0d[23], write_0r1d[23], wack_0n[23], ldata_0n[23], ldata_1n[23]);
  DRLATCH I265 (write_0r0d[24], write_0r1d[24], wack_0n[24], ldata_0n[24], ldata_1n[24]);
  DRLATCH I266 (write_0r0d[25], write_0r1d[25], wack_0n[25], ldata_0n[25], ldata_1n[25]);
  DRLATCH I267 (write_0r0d[26], write_0r1d[26], wack_0n[26], ldata_0n[26], ldata_1n[26]);
  DRLATCH I268 (write_0r0d[27], write_0r1d[27], wack_0n[27], ldata_0n[27], ldata_1n[27]);
  DRLATCH I269 (write_0r0d[28], write_0r1d[28], wack_0n[28], ldata_0n[28], ldata_1n[28]);
  DRLATCH I270 (write_0r0d[29], write_0r1d[29], wack_0n[29], ldata_0n[29], ldata_1n[29]);
  DRLATCH I271 (write_0r0d[30], write_0r1d[30], wack_0n[30], ldata_0n[30], ldata_1n[30]);
  DRLATCH I272 (write_0r0d[31], write_0r1d[31], wack_0n[31], ldata_0n[31], ldata_1n[31]);
  DRLATCH I273 (write_0r0d[32], write_0r1d[32], wack_0n[32], ldata_0n[32], ldata_1n[32]);
  DRLATCH I274 (write_0r0d[33], write_0r1d[33], wack_0n[33], ldata_0n[33], ldata_1n[33]);
  DRLATCH I275 (write_0r0d[34], write_0r1d[34], wack_0n[34], ldata_0n[34], ldata_1n[34]);
  DRLATCH I276 (write_0r0d[35], write_0r1d[35], wack_0n[35], ldata_0n[35], ldata_1n[35]);
endmodule

module BrzWhile (
  activate_0r, activate_0a,
  guard_0r, guard_0a0d, guard_0a1d,
  activateOut_0r, activateOut_0a
);
  input activate_0r;
  output activate_0a;
  output guard_0r;
  input guard_0a0d;
  input guard_0a1d;
  output activateOut_0r;
  input activateOut_0a;
  wire guardReq_0n;
  wire nReq_0n;
  BALSA_SELEM I0 (guardReq_0n, activateOut_0r, guard_0r, guard_0a1d);
  INV I1 (nReq_0n, activate_0r);
  NOR2 I2 (guardReq_0n, nReq_0n, activateOut_0a);
  BUFF I3 (activate_0a, guard_0a0d);
endmodule

module BrzWireFork_13 (
  inp_0r, inp_0a,
  out_0r, out_0a,
  out_1r, out_1a,
  out_2r, out_2a,
  out_3r, out_3a,
  out_4r, out_4a,
  out_5r, out_5a,
  out_6r, out_6a,
  out_7r, out_7a,
  out_8r, out_8a,
  out_9r, out_9a,
  out_10r, out_10a,
  out_11r, out_11a,
  out_12r, out_12a
);
  input inp_0r;
  output inp_0a;
  output out_0r;
  input out_0a;
  output out_1r;
  input out_1a;
  output out_2r;
  input out_2a;
  output out_3r;
  input out_3a;
  output out_4r;
  input out_4a;
  output out_5r;
  input out_5a;
  output out_6r;
  input out_6a;
  output out_7r;
  input out_7a;
  output out_8r;
  input out_8a;
  output out_9r;
  input out_9a;
  output out_10r;
  input out_10a;
  output out_11r;
  input out_11a;
  output out_12r;
  input out_12a;
  supply0 gnd;
  BUFF I0 (inp_0a, gnd);
  BUFF I1 (out_0r, inp_0r);
  BUFF I2 (out_1r, inp_0r);
  BUFF I3 (out_2r, inp_0r);
  BUFF I4 (out_3r, inp_0r);
  BUFF I5 (out_4r, inp_0r);
  BUFF I6 (out_5r, inp_0r);
  BUFF I7 (out_6r, inp_0r);
  BUFF I8 (out_7r, inp_0r);
  BUFF I9 (out_8r, inp_0r);
  BUFF I10 (out_9r, inp_0r);
  BUFF I11 (out_10r, inp_0r);
  BUFF I12 (out_11r, inp_0r);
  BUFF I13 (out_12r, inp_0r);
endmodule

module Balsa_CSAdder__DP2 (
  activate_0r, activate_0a,
  a_0r, a_0a0d, a_0a1d,
  b_0r, b_0a0d, b_0a1d,
  cs_0r, cs_0a0d, cs_0a1d,
  cout_0r0d, cout_0r1d, cout_0a,
  s_0r0d, s_0r1d, s_0a
);
  input activate_0r;
  output activate_0a;
  output a_0r;
  input [34:0] a_0a0d;
  input [34:0] a_0a1d;
  output b_0r;
  input [34:0] b_0a0d;
  input [34:0] b_0a1d;
  output cs_0r;
  input [34:0] cs_0a0d;
  input [34:0] cs_0a1d;
  output [34:0] cout_0r0d;
  output [34:0] cout_0r1d;
  input cout_0a;
  output [34:0] s_0r0d;
  output [34:0] s_0r1d;
  input s_0a;
  wire c32_r;
  wire c32_a;
  wire c31_r;
  wire c31_a;
  wire c30_r;
  wire c30_a;
  wire c29_r;
  wire c29_a;
  wire c28_r;
  wire c28_a;
  wire c27_r;
  wire c27_a;
  wire c26_r;
  wire c26_a;
  wire c25_r;
  wire c25_a;
  wire c24_r;
  wire c24_a;
  wire c23_r;
  wire [34:0] c23_a0d;
  wire [34:0] c23_a1d;
  wire c22_r;
  wire [34:0] c22_a0d;
  wire [34:0] c22_a1d;
  wire c21_r;
  wire [34:0] c21_a0d;
  wire [34:0] c21_a1d;
  wire c20_r;
  wire [34:0] c20_a0d;
  wire [34:0] c20_a1d;
  wire c19_r;
  wire [34:0] c19_a0d;
  wire [34:0] c19_a1d;
  wire c18_r;
  wire c18_a;
  wire c17_r;
  wire [34:0] c17_a0d;
  wire [34:0] c17_a1d;
  wire c16_r;
  wire [34:0] c16_a0d;
  wire [34:0] c16_a1d;
  wire c15_r;
  wire [34:0] c15_a0d;
  wire [34:0] c15_a1d;
  wire c14_r;
  wire [34:0] c14_a0d;
  wire [34:0] c14_a1d;
  wire c13_r;
  wire [34:0] c13_a0d;
  wire [34:0] c13_a1d;
  wire c12_r;
  wire [34:0] c12_a0d;
  wire [34:0] c12_a1d;
  wire c11_r;
  wire [34:0] c11_a0d;
  wire [34:0] c11_a1d;
  wire c10_r;
  wire [34:0] c10_a0d;
  wire [34:0] c10_a1d;
  wire c9_r;
  wire [34:0] c9_a0d;
  wire [34:0] c9_a1d;
  wire c8_r;
  wire [34:0] c8_a0d;
  wire [34:0] c8_a1d;
  wire c7_r;
  wire [34:0] c7_a0d;
  wire [34:0] c7_a1d;
  BrzBinaryFunc_35_35_35_s3_And_s5_false_s5__m19m I0 (c9_r, c9_a0d[34:0], c9_a1d[34:0], c8_r, c8_a0d[34:0], c8_a1d[34:0], c7_r, c7_a0d[34:0], c7_a1d[34:0]);
  BrzBinaryFunc_35_35_35_s3_And_s5_false_s5__m19m I1 (c12_r, c12_a0d[34:0], c12_a1d[34:0], c11_r, c11_a0d[34:0], c11_a1d[34:0], c10_r, c10_a0d[34:0], c10_a1d[34:0]);
  BrzBinaryFunc_35_35_35_s3_And_s5_false_s5__m19m I2 (c15_r, c15_a0d[34:0], c15_a1d[34:0], c14_r, c14_a0d[34:0], c14_a1d[34:0], c13_r, c13_a0d[34:0], c13_a1d[34:0]);
  BrzBinaryFunc_35_35_35_s2_Or_s5_false_s5_f_m21m I3 (c16_r, c16_a0d[34:0], c16_a1d[34:0], c15_r, c15_a0d[34:0], c15_a1d[34:0], c12_r, c12_a0d[34:0], c12_a1d[34:0]);
  BrzBinaryFunc_35_35_35_s2_Or_s5_false_s5_f_m21m I4 (c17_r, c17_a0d[34:0], c17_a1d[34:0], c16_r, c16_a0d[34:0], c16_a1d[34:0], c9_r, c9_a0d[34:0], c9_a1d[34:0]);
  BrzFetch_35_s5_false I5 (c18_r, c18_a, c17_r, c17_a0d[34:0], c17_a1d[34:0], cout_0r0d[34:0], cout_0r1d[34:0], cout_0a);
  BrzBinaryFunc_35_35_35_s3_Xor_s5_false_s5__m23m I6 (c22_r, c22_a0d[34:0], c22_a1d[34:0], c21_r, c21_a0d[34:0], c21_a1d[34:0], c20_r, c20_a0d[34:0], c20_a1d[34:0]);
  BrzBinaryFunc_35_35_35_s3_Xor_s5_false_s5__m23m I7 (c23_r, c23_a0d[34:0], c23_a1d[34:0], c22_r, c22_a0d[34:0], c22_a1d[34:0], c19_r, c19_a0d[34:0], c19_a1d[34:0]);
  BrzFetch_35_s5_false I8 (c24_r, c24_a, c23_r, c23_a0d[34:0], c23_a1d[34:0], s_0r0d[34:0], s_0r1d[34:0], s_0a);
  BrzConcur_2 I9 (c32_r, c32_a, c24_r, c24_a, c18_r, c18_a);
  BrzActiveEagerFalseVariable_35_3_s0_ I10 (c26_r, c26_a, a_0r, a_0a0d[34:0], a_0a1d[34:0], c25_r, c25_a, c21_r, c21_a0d[34:0], c21_a1d[34:0], c14_r, c14_a0d[34:0], c14_a1d[34:0], c10_r, c10_a0d[34:0], c10_a1d[34:0]);
  BrzActiveEagerFalseVariable_35_3_s0_ I11 (c28_r, c28_a, b_0r, b_0a0d[34:0], b_0a1d[34:0], c27_r, c27_a, c20_r, c20_a0d[34:0], c20_a1d[34:0], c13_r, c13_a0d[34:0], c13_a1d[34:0], c7_r, c7_a0d[34:0], c7_a1d[34:0]);
  BrzActiveEagerFalseVariable_35_3_s0_ I12 (c30_r, c30_a, cs_0r, cs_0a0d[34:0], cs_0a1d[34:0], c29_r, c29_a, c19_r, c19_a0d[34:0], c19_a1d[34:0], c11_r, c11_a0d[34:0], c11_a1d[34:0], c8_r, c8_a0d[34:0], c8_a1d[34:0]);
  BrzFork_3 I13 (c31_r, c31_a, c30_r, c30_a, c28_r, c28_a, c26_r, c26_a);
  BrzSynch_3 I14 (c29_r, c29_a, c27_r, c27_a, c25_r, c25_a, c32_r, c32_a);
  BrzLoop I15 (activate_0r, activate_0a, c31_r, c31_a);
endmodule

module Balsa_CPadder (
  activate_0r, activate_0a,
  a_0r, a_0a0d, a_0a1d,
  b_0r, b_0a0d, b_0a1d,
  c0_0r, c0_0a0d, c0_0a1d,
  s_0r0d, s_0r1d, s_0a,
  cN_0r0d, cN_0r1d, cN_0a
);
  input activate_0r;
  output activate_0a;
  output a_0r;
  input [31:0] a_0a0d;
  input [31:0] a_0a1d;
  output b_0r;
  input [31:0] b_0a0d;
  input [31:0] b_0a1d;
  output c0_0r;
  input c0_0a0d;
  input c0_0a1d;
  output [31:0] s_0r0d;
  output [31:0] s_0r1d;
  input s_0a;
  output cN_0r0d;
  output cN_0r1d;
  input cN_0a;
  wire c44_r;
  wire c44_a;
  wire c43_r;
  wire c43_a;
  wire c42_r;
  wire c42_a;
  wire c41_r;
  wire c41_a;
  wire c40_r;
  wire c40_a;
  wire c39_r;
  wire c39_a;
  wire c38_r;
  wire c38_a;
  wire c37_r;
  wire c37_a;
  wire c36_r;
  wire c36_a;
  wire c35_r;
  wire c35_a;
  wire [32:0] c34_r0d;
  wire [32:0] c34_r1d;
  wire c34_a;
  wire c33_r;
  wire [32:0] c33_a0d;
  wire [32:0] c33_a1d;
  wire c32_r;
  wire c32_a0d;
  wire c32_a1d;
  wire c31_r;
  wire [31:0] c31_a0d;
  wire [31:0] c31_a1d;
  wire c30_r;
  wire c30_a;
  wire [32:0] c29_r0d;
  wire [32:0] c29_r1d;
  wire c29_a;
  wire c28_r;
  wire [32:0] c28_a0d;
  wire [32:0] c28_a1d;
  wire c27_r;
  wire c27_a0d;
  wire c27_a1d;
  wire c26_r;
  wire [31:0] c26_a0d;
  wire [31:0] c26_a1d;
  wire c25_r;
  wire c25_a;
  wire c24_r;
  wire c24_a;
  wire c23_r;
  wire c23_a;
  wire c22_r;
  wire c22_a;
  wire c21_r;
  wire c21_a;
  wire c20_r;
  wire c20_a;
  wire [33:0] c19_r0d;
  wire [33:0] c19_r1d;
  wire c19_a;
  wire c18_r;
  wire [33:0] c18_a0d;
  wire [33:0] c18_a1d;
  wire c17_r;
  wire [32:0] c17_a0d;
  wire [32:0] c17_a1d;
  wire c16_r;
  wire [32:0] c16_a0d;
  wire [32:0] c16_a1d;
  wire c15_r;
  wire [32:0] c15_a0d;
  wire [32:0] c15_a1d;
  wire c14_r;
  wire [32:0] c14_a0d;
  wire [32:0] c14_a1d;
  wire c13_r;
  wire c13_a;
  wire c12_r;
  wire c12_a;
  wire c11_r;
  wire c11_a;
  wire c10_r;
  wire [31:0] c10_a0d;
  wire [31:0] c10_a1d;
  wire c9_r;
  wire c9_a;
  wire c8_r;
  wire c8_a0d;
  wire c8_a1d;
  wire c7_r;
  wire [33:0] c7_a0d;
  wire [33:0] c7_a1d;
  BrzFetch_1_s5_false I0 (c9_r, c9_a, c8_r, c8_a0d, c8_a1d, cN_0r0d, cN_0r1d, cN_0a);
  BrzFetch_32_s5_false I1 (c11_r, c11_a, c10_r, c10_a0d[31:0], c10_a1d[31:0], s_0r0d[31:0], s_0r1d[31:0], s_0a);
  BrzConcur_2 I2 (c12_r, c12_a, c11_r, c11_a, c9_r, c9_a);
  BrzActiveEagerFalseVariable_34_2_s22_1_2e__m5m I3 (c13_r, c13_a, c7_r, c7_a0d[33:0], c7_a1d[33:0], c12_r, c12_a, c10_r, c10_a0d[31:0], c10_a1d[31:0], c8_r, c8_a0d, c8_a1d);
  BrzBinaryFunc_34_33_33_s3_Add_s5_false_s5__m17m I4 (c18_r, c18_a0d[33:0], c18_a1d[33:0], c17_r, c17_a0d[32:0], c17_a1d[32:0], c16_r, c16_a0d[32:0], c16_a1d[32:0]);
  BrzFetch_34_s5_false I5 (c25_r, c25_a, c18_r, c18_a0d[33:0], c18_a1d[33:0], c19_r0d[33:0], c19_r1d[33:0], c19_a);
  BrzActiveEagerFalseVariable_33_1_s0_ I6 (c21_r, c21_a, c15_r, c15_a0d[32:0], c15_a1d[32:0], c20_r, c20_a, c16_r, c16_a0d[32:0], c16_a1d[32:0]);
  BrzActiveEagerFalseVariable_33_1_s0_ I7 (c23_r, c23_a, c14_r, c14_a0d[32:0], c14_a1d[32:0], c22_r, c22_a, c17_r, c17_a0d[32:0], c17_a1d[32:0]);
  BrzFork_2 I8 (c24_r, c24_a, c23_r, c23_a, c21_r, c21_a);
  BrzSynch_2 I9 (c22_r, c22_a, c20_r, c20_a, c25_r, c25_a);
  BrzCombine_33_1_32 I10 (c28_r, c28_a0d[32:0], c28_a1d[32:0], c27_r, c27_a0d, c27_a1d, c26_r, c26_a0d[31:0], c26_a1d[31:0]);
  BrzFetch_33_s5_false I11 (c30_r, c30_a, c28_r, c28_a0d[32:0], c28_a1d[32:0], c29_r0d[32:0], c29_r1d[32:0], c29_a);
  BrzCombine_33_1_32 I12 (c33_r, c33_a0d[32:0], c33_a1d[32:0], c32_r, c32_a0d, c32_a1d, c31_r, c31_a0d[31:0], c31_a1d[31:0]);
  BrzFetch_33_s5_false I13 (c35_r, c35_a, c33_r, c33_a0d[32:0], c33_a1d[32:0], c34_r0d[32:0], c34_r1d[32:0], c34_a);
  BrzConcur_2 I14 (c43_r, c43_a, c35_r, c35_a, c30_r, c30_a);
  BrzActiveEagerFalseVariable_32_1_s0_ I15 (c37_r, c37_a, a_0r, a_0a0d[31:0], a_0a1d[31:0], c36_r, c36_a, c31_r, c31_a0d[31:0], c31_a1d[31:0]);
  BrzActiveEagerFalseVariable_32_1_s0_ I16 (c39_r, c39_a, b_0r, b_0a0d[31:0], b_0a1d[31:0], c38_r, c38_a, c26_r, c26_a0d[31:0], c26_a1d[31:0]);
  BrzActiveEagerFalseVariable_1_2_s0_ I17 (c41_r, c41_a, c0_0r, c0_0a0d, c0_0a1d, c40_r, c40_a, c32_r, c32_a0d, c32_a1d, c27_r, c27_a0d, c27_a1d);
  BrzFork_3 I18 (c42_r, c42_a, c41_r, c41_a, c39_r, c39_a, c37_r, c37_a);
  BrzSynch_3 I19 (c40_r, c40_a, c38_r, c38_a, c36_r, c36_a, c43_r, c43_a);
  BrzPassivatorPush_33_1 I20 (c15_r, c15_a0d[32:0], c15_a1d[32:0], c29_r0d[32:0], c29_r1d[32:0], c29_a);
  BrzPassivatorPush_33_1 I21 (c14_r, c14_a0d[32:0], c14_a1d[32:0], c34_r0d[32:0], c34_r1d[32:0], c34_a);
  BrzConcur_3 I22 (c44_r, c44_a, c42_r, c42_a, c24_r, c24_a, c13_r, c13_a);
  BrzPassivatorPush_34_1 I23 (c7_r, c7_a0d[33:0], c7_a1d[33:0], c19_r0d[33:0], c19_r1d[33:0], c19_a);
  BrzLoop I24 (activate_0r, activate_0a, c44_r, c44_a);
endmodule

module Balsa_doByPass (
  activate_0r, activate_0a,
  bH_0r, bH_0a0d, bH_0a1d,
  bL_0r, bL_0a0d, bL_0a1d,
  bpH_0r, bpH_0a0d, bpH_0a1d,
  bpL_0r, bpL_0a0d, bpL_0a1d,
  bmZ_0r, bmZ_0a0d, bmZ_0a1d,
  bmN_0r, bmN_0a0d, bmN_0a1d,
  mpH_0r0d, mpH_0r1d, mpH_0a,
  mpL_0r0d, mpL_0r1d, mpL_0a,
  mZ_0r0d, mZ_0r1d, mZ_0a,
  mN_0r0d, mN_0r1d, mN_0a
);
  input activate_0r;
  output activate_0a;
  output bH_0r;
  input bH_0a0d;
  input bH_0a1d;
  output bL_0r;
  input bL_0a0d;
  input bL_0a1d;
  output bpH_0r;
  input [31:0] bpH_0a0d;
  input [31:0] bpH_0a1d;
  output bpL_0r;
  input [31:0] bpL_0a0d;
  input [31:0] bpL_0a1d;
  output bmZ_0r;
  input bmZ_0a0d;
  input bmZ_0a1d;
  output bmN_0r;
  input bmN_0a0d;
  input bmN_0a1d;
  output [31:0] mpH_0r0d;
  output [31:0] mpH_0r1d;
  input mpH_0a;
  output [31:0] mpL_0r0d;
  output [31:0] mpL_0r1d;
  input mpL_0a;
  output mZ_0r0d;
  output mZ_0r1d;
  input mZ_0a;
  output mN_0r0d;
  output mN_0r1d;
  input mN_0a;
  wire c47_r;
  wire c47_a;
  wire c46_r;
  wire c46_a;
  wire c45_r;
  wire c45_a;
  wire c44_r;
  wire c44_a;
  wire c43_r;
  wire c43_a;
  wire c42_r;
  wire c42_a;
  wire c41_r0d;
  wire c41_r1d;
  wire c41_a;
  wire c40_r;
  wire c40_a0d;
  wire c40_a1d;
  wire c39_r;
  wire c39_a;
  wire c38_r;
  wire c38_a;
  wire [31:0] c37_r0d;
  wire [31:0] c37_r1d;
  wire c37_a;
  wire c36_r;
  wire [31:0] c36_a0d;
  wire [31:0] c36_a1d;
  wire c35_r;
  wire c35_a;
  wire c34_r0d;
  wire c34_r1d;
  wire c34_a;
  wire c33_r;
  wire c33_a0d;
  wire c33_a1d;
  wire c32_r;
  wire c32_a;
  wire c31_r0d;
  wire c31_r1d;
  wire c31_a;
  wire c30_r;
  wire c30_a0d;
  wire c30_a1d;
  wire c29_r0d;
  wire c29_r1d;
  wire c29_a;
  wire c28_r;
  wire c28_a;
  wire c27_r;
  wire c27_a0d;
  wire c27_a1d;
  wire c26_r;
  wire c26_a;
  wire [31:0] c25_r0d;
  wire [31:0] c25_r1d;
  wire c25_a;
  wire c24_r;
  wire [31:0] c24_a0d;
  wire [31:0] c24_a1d;
  wire c23_r;
  wire c23_a;
  wire c22_r;
  wire c22_a;
  wire [31:0] c21_r0d;
  wire [31:0] c21_r1d;
  wire c21_a;
  wire c20_r;
  wire c20_a;
  wire c19_r0d;
  wire c19_r1d;
  wire c19_a;
  wire c18_r;
  wire c18_a;
  wire c17_r0d;
  wire c17_r1d;
  wire c17_a;
  wire c16_r0d;
  wire c16_r1d;
  wire c16_a;
  wire c15_r;
  wire c15_a;
  wire c14_r;
  wire c14_a0d;
  wire c14_a1d;
  wire c13_r;
  wire c13_a;
  wire [31:0] c12_r0d;
  wire [31:0] c12_r1d;
  wire c12_a;
  BrzFetch_32_s4_true I0 (c13_r, c13_a, bpH_0r, bpH_0a0d[31:0], bpH_0a1d[31:0], c12_r0d[31:0], c12_r1d[31:0], c12_a);
  BrzFetch_1_s5_false I1 (c15_r, c15_a, c14_r, c14_a0d, c14_a1d, c16_r0d, c16_r1d, c16_a);
  BrzCase_1_1_s1_1 I2 (c16_r0d, c16_r1d, c16_a, c13_r, c13_a);
  BrzFetch_1_s4_true I3 (c18_r, c18_a, bmN_0r, bmN_0a0d, bmN_0a1d, c17_r0d, c17_r1d, c17_a);
  BrzFetch_1_s4_true I4 (c20_r, c20_a, bmZ_0r, bmZ_0a0d, bmZ_0a1d, c19_r0d, c19_r1d, c19_a);
  BrzFetch_32_s4_true I5 (c22_r, c22_a, bpL_0r, bpL_0a0d[31:0], bpL_0a1d[31:0], c21_r0d[31:0], c21_r1d[31:0], c21_a);
  BrzConcur_4 I6 (c23_r, c23_a, c22_r, c22_a, c20_r, c20_a, c18_r, c18_a, c15_r, c15_a);
  BrzConstant_32_0 I7 (c24_r, c24_a0d[31:0], c24_a1d[31:0]);
  BrzFetch_32_s5_false I8 (c26_r, c26_a, c24_r, c24_a0d[31:0], c24_a1d[31:0], c25_r0d[31:0], c25_r1d[31:0], c25_a);
  BrzFetch_1_s5_false I9 (c28_r, c28_a, c27_r, c27_a0d, c27_a1d, c29_r0d, c29_r1d, c29_a);
  BrzCase_1_1_s1_1 I10 (c29_r0d, c29_r1d, c29_a, c26_r, c26_a);
  BrzConstant_1_0 I11 (c30_r, c30_a0d, c30_a1d);
  BrzFetch_1_s5_false I12 (c32_r, c32_a, c30_r, c30_a0d, c30_a1d, c31_r0d, c31_r1d, c31_a);
  BrzConstant_1_0 I13 (c33_r, c33_a0d, c33_a1d);
  BrzFetch_1_s5_false I14 (c35_r, c35_a, c33_r, c33_a0d, c33_a1d, c34_r0d, c34_r1d, c34_a);
  BrzConstant_32_0 I15 (c36_r, c36_a0d[31:0], c36_a1d[31:0]);
  BrzFetch_32_s5_false I16 (c38_r, c38_a, c36_r, c36_a0d[31:0], c36_a1d[31:0], c37_r0d[31:0], c37_r1d[31:0], c37_a);
  BrzConcur_4 I17 (c39_r, c39_a, c38_r, c38_a, c35_r, c35_a, c32_r, c32_a, c28_r, c28_a);
  BrzCallMux_32_2 I18 (c25_r0d[31:0], c25_r1d[31:0], c25_a, c12_r0d[31:0], c12_r1d[31:0], c12_a, mpH_0r0d[31:0], mpH_0r1d[31:0], mpH_0a);
  BrzCallMux_32_2 I19 (c37_r0d[31:0], c37_r1d[31:0], c37_a, c21_r0d[31:0], c21_r1d[31:0], c21_a, mpL_0r0d[31:0], mpL_0r1d[31:0], mpL_0a);
  BrzCallMux_1_2 I20 (c34_r0d, c34_r1d, c34_a, c19_r0d, c19_r1d, c19_a, mZ_0r0d, mZ_0r1d, mZ_0a);
  BrzCallMux_1_2 I21 (c31_r0d, c31_r1d, c31_a, c17_r0d, c17_r1d, c17_a, mN_0r0d, mN_0r1d, mN_0a);
  BrzFetch_1_s5_false I22 (c47_r, c47_a, c40_r, c40_a0d, c40_a1d, c41_r0d, c41_r1d, c41_a);
  BrzCase_1_2_s5_0_3b1 I23 (c41_r0d, c41_r1d, c41_a, c23_r, c23_a, c39_r, c39_a);
  BrzActiveEagerFalseVariable_1_2_s0_ I24 (c43_r, c43_a, bH_0r, bH_0a0d, bH_0a1d, c42_r, c42_a, c27_r, c27_a0d, c27_a1d, c14_r, c14_a0d, c14_a1d);
  BrzActiveEagerFalseVariable_1_1_s0_ I25 (c45_r, c45_a, bL_0r, bL_0a0d, bL_0a1d, c44_r, c44_a, c40_r, c40_a0d, c40_a1d);
  BrzFork_2 I26 (c46_r, c46_a, c45_r, c45_a, c43_r, c43_a);
  BrzSynch_2 I27 (c44_r, c44_a, c42_r, c42_a, c47_r, c47_a);
  BrzLoop I28 (activate_0r, activate_0a, c46_r, c46_a);
endmodule

module Balsa_bypassMul (
  activate_0r, activate_0a,
  bypass_0r, bypass_0a0d, bypass_0a1d,
  bypassH_0r, bypassH_0a0d, bypassH_0a1d,
  mulOpA_0r, mulOpA_0a0d, mulOpA_0a1d,
  mulOpB_0r, mulOpB_0a0d, mulOpB_0a1d,
  mulOpC_0r, mulOpC_0a0d, mulOpC_0a1d,
  mulType_0r, mulType_0a0d, mulType_0a1d,
  mulOpAo_0r0d, mulOpAo_0r1d, mulOpAo_0a,
  mulOpBo_0r0d, mulOpBo_0r1d, mulOpBo_0a,
  mulOpCo_0r0d, mulOpCo_0r1d, mulOpCo_0a,
  mulTypeo_0r0d, mulTypeo_0r1d, mulTypeo_0a,
  bH_0r0d, bH_0r1d, bH_0a,
  bL_0r0d, bL_0r1d, bL_0a
);
  input activate_0r;
  output activate_0a;
  output bypass_0r;
  input bypass_0a0d;
  input bypass_0a1d;
  output bypassH_0r;
  input bypassH_0a0d;
  input bypassH_0a1d;
  output mulOpA_0r;
  input [31:0] mulOpA_0a0d;
  input [31:0] mulOpA_0a1d;
  output mulOpB_0r;
  input [31:0] mulOpB_0a0d;
  input [31:0] mulOpB_0a1d;
  output mulOpC_0r;
  input [31:0] mulOpC_0a0d;
  input [31:0] mulOpC_0a1d;
  output mulType_0r;
  input [2:0] mulType_0a0d;
  input [2:0] mulType_0a1d;
  output [31:0] mulOpAo_0r0d;
  output [31:0] mulOpAo_0r1d;
  input mulOpAo_0a;
  output [31:0] mulOpBo_0r0d;
  output [31:0] mulOpBo_0r1d;
  input mulOpBo_0a;
  output [31:0] mulOpCo_0r0d;
  output [31:0] mulOpCo_0r1d;
  input mulOpCo_0a;
  output [2:0] mulTypeo_0r0d;
  output [2:0] mulTypeo_0r1d;
  input mulTypeo_0a;
  output bH_0r0d;
  output bH_0r1d;
  input bH_0a;
  output bL_0r0d;
  output bL_0r1d;
  input bL_0a;
  wire c58_r;
  wire c58_a;
  wire c57_r;
  wire c57_a;
  wire c56_r;
  wire c56_a;
  wire c55_r;
  wire c55_a;
  wire c54_r;
  wire c54_a;
  wire c53_r;
  wire c53_a;
  wire c52_r;
  wire c52_a;
  wire c51_r;
  wire c51_a;
  wire c50_r;
  wire c50_a;
  wire c49_r;
  wire c49_a;
  wire c48_r;
  wire c48_a;
  wire c47_r;
  wire c47_a;
  wire c46_r;
  wire c46_a;
  wire c45_r;
  wire c45_a;
  wire c44_r0d;
  wire c44_r1d;
  wire c44_a;
  wire c43_r;
  wire c43_a0d;
  wire c43_a1d;
  wire [2:0] c42_r0d;
  wire [2:0] c42_r1d;
  wire c42_a;
  wire c41_r;
  wire c41_a;
  wire c40_r;
  wire [2:0] c40_a0d;
  wire [2:0] c40_a1d;
  wire c39_r;
  wire c39_a;
  wire c38_r;
  wire c38_a;
  wire c37_r;
  wire [31:0] c37_a0d;
  wire [31:0] c37_a1d;
  wire c36_r;
  wire c36_a;
  wire c35_r;
  wire c35_a;
  wire c34_r;
  wire c34_a;
  wire c33_r;
  wire [31:0] c33_a0d;
  wire [31:0] c33_a1d;
  wire c32_r;
  wire c32_a;
  wire c31_r;
  wire [31:0] c31_a0d;
  wire [31:0] c31_a1d;
  wire c30_r;
  wire c30_a;
  wire c29_r;
  wire [2:0] c29_a0d;
  wire [2:0] c29_a1d;
  wire [2:0] c28_r0d;
  wire [2:0] c28_r1d;
  wire c28_a;
  wire c27_r;
  wire c27_a;
  wire c26_r;
  wire [2:0] c26_a0d;
  wire [2:0] c26_a1d;
  wire c25_r;
  wire c25_a;
  wire c24_r;
  wire c24_a;
  wire [31:0] c23_r0d;
  wire [31:0] c23_r1d;
  wire c23_a;
  wire c22_r;
  wire [31:0] c22_a0d;
  wire [31:0] c22_a1d;
  wire c21_r;
  wire [31:0] c21_a0d;
  wire [31:0] c21_a1d;
  wire c20_r;
  wire c20_a;
  wire [31:0] c19_r0d;
  wire [31:0] c19_r1d;
  wire c19_a;
  wire c18_r;
  wire [31:0] c18_a0d;
  wire [31:0] c18_a1d;
  wire c17_r;
  wire c17_a;
  wire c16_r;
  wire c16_a0d;
  wire c16_a1d;
  wire c15_r;
  wire c15_a;
  wire c14_r;
  wire c14_a0d;
  wire c14_a1d;
  BrzFetch_1_s5_false I0 (c15_r, c15_a, c14_r, c14_a0d, c14_a1d, bH_0r0d, bH_0r1d, bH_0a);
  BrzFetch_1_s5_false I1 (c17_r, c17_a, c16_r, c16_a0d, c16_a1d, bL_0r0d, bL_0r1d, bL_0a);
  BrzConstant_32_0 I2 (c18_r, c18_a0d[31:0], c18_a1d[31:0]);
  BrzFetch_32_s5_false I3 (c20_r, c20_a, c18_r, c18_a0d[31:0], c18_a1d[31:0], c19_r0d[31:0], c19_r1d[31:0], c19_a);
  BrzFetch_32_s5_false I4 (c24_r, c24_a, c22_r, c22_a0d[31:0], c22_a1d[31:0], c23_r0d[31:0], c23_r1d[31:0], c23_a);
  BrzActiveEagerFalseVariable_32_1_s0_ I5 (c25_r, c25_a, c21_r, c21_a0d[31:0], c21_a1d[31:0], c24_r, c24_a, c22_r, c22_a0d[31:0], c22_a1d[31:0]);
  BrzCallMux_32_2 I6 (c23_r0d[31:0], c23_r1d[31:0], c23_a, c19_r0d[31:0], c19_r1d[31:0], c19_a, mulOpCo_0r0d[31:0], mulOpCo_0r1d[31:0], mulOpCo_0a);
  BrzFetch_3_s5_false I7 (c27_r, c27_a, c26_r, c26_a0d[2:0], c26_a1d[2:0], c28_r0d[2:0], c28_r1d[2:0], c28_a);
  BrzCase_3_2_s19_3_2c0m6_3b7_2c5_2c1 I8 (c28_r0d[2:0], c28_r1d[2:0], c28_a, c20_r, c20_a, c25_r, c25_a);
  BrzFetch_3_s5_false I9 (c30_r, c30_a, c29_r, c29_a0d[2:0], c29_a1d[2:0], mulTypeo_0r0d[2:0], mulTypeo_0r1d[2:0], mulTypeo_0a);
  BrzFetch_32_s5_false I10 (c32_r, c32_a, c31_r, c31_a0d[31:0], c31_a1d[31:0], mulOpBo_0r0d[31:0], mulOpBo_0r1d[31:0], mulOpBo_0a);
  BrzFetch_32_s5_false I11 (c34_r, c34_a, c33_r, c33_a0d[31:0], c33_a1d[31:0], mulOpAo_0r0d[31:0], mulOpAo_0r1d[31:0], mulOpAo_0a);
  BrzConcur_4 I12 (c35_r, c35_a, c34_r, c34_a, c32_r, c32_a, c30_r, c30_a, c27_r, c27_a);
  BrzContinue I13 (c36_r, c36_a);
  BrzContinue I14 (c39_r, c39_a);
  BrzActiveEagerNullAdapt_32 I15 (c38_r, c38_a, c37_r, c37_a0d[31:0], c37_a1d[31:0], c39_r, c39_a);
  BrzFetch_3_s5_false I16 (c41_r, c41_a, c40_r, c40_a0d[2:0], c40_a1d[2:0], c42_r0d[2:0], c42_r1d[2:0], c42_a);
  BrzCase_3_2_s19_3_2c0m6_3b7_2c5_2c1 I17 (c42_r0d[2:0], c42_r1d[2:0], c42_a, c36_r, c36_a, c38_r, c38_a);
  BrzCallDemux_32_2 I18 (c37_r, c37_a0d[31:0], c37_a1d[31:0], c21_r, c21_a0d[31:0], c21_a1d[31:0], mulOpC_0r, mulOpC_0a0d[31:0], mulOpC_0a1d[31:0]);
  BrzFetch_1_s5_false I19 (c50_r, c50_a, c43_r, c43_a0d, c43_a1d, c44_r0d, c44_r1d, c44_a);
  BrzCase_1_2_s5_0_3b1 I20 (c44_r0d, c44_r1d, c44_a, c35_r, c35_a, c41_r, c41_a);
  BrzActiveEagerFalseVariable_32_1_s0_ I21 (c46_r, c46_a, mulOpA_0r, mulOpA_0a0d[31:0], mulOpA_0a1d[31:0], c45_r, c45_a, c33_r, c33_a0d[31:0], c33_a1d[31:0]);
  BrzActiveEagerFalseVariable_32_1_s0_ I22 (c48_r, c48_a, mulOpB_0r, mulOpB_0a0d[31:0], mulOpB_0a1d[31:0], c47_r, c47_a, c31_r, c31_a0d[31:0], c31_a1d[31:0]);
  BrzFork_2 I23 (c49_r, c49_a, c48_r, c48_a, c46_r, c46_a);
  BrzSynch_2 I24 (c47_r, c47_a, c45_r, c45_a, c50_r, c50_a);
  BrzConcur_3 I25 (c58_r, c58_a, c49_r, c49_a, c17_r, c17_a, c15_r, c15_a);
  BrzActiveEagerFalseVariable_1_2_s0_ I26 (c52_r, c52_a, bypass_0r, bypass_0a0d, bypass_0a1d, c51_r, c51_a, c43_r, c43_a0d, c43_a1d, c16_r, c16_a0d, c16_a1d);
  BrzActiveEagerFalseVariable_1_1_s0_ I27 (c54_r, c54_a, bypassH_0r, bypassH_0a0d, bypassH_0a1d, c53_r, c53_a, c14_r, c14_a0d, c14_a1d);
  BrzActiveEagerFalseVariable_3_3_s0_ I28 (c56_r, c56_a, mulType_0r, mulType_0a0d[2:0], mulType_0a1d[2:0], c55_r, c55_a, c40_r, c40_a0d[2:0], c40_a1d[2:0], c29_r, c29_a0d[2:0], c29_a1d[2:0], c26_r, c26_a0d[2:0], c26_a1d[2:0]);
  BrzFork_3 I29 (c57_r, c57_a, c56_r, c56_a, c54_r, c54_a, c52_r, c52_a);
  BrzSynch_3 I30 (c55_r, c55_a, c53_r, c53_a, c51_r, c51_a, c58_r, c58_a);
  BrzLoop I31 (activate_0r, activate_0a, c57_r, c57_a);
endmodule

module Balsa_signAdj (
  activate_0r, activate_0a,
  mType_0r, mType_0a0d, mType_0a1d,
  a_0r, a_0a0d, a_0a1d,
  b_0r, b_0a0d, b_0a1d,
  c_0r, c_0a0d, c_0a1d,
  aa_0r0d, aa_0r1d, aa_0a,
  ba_0r0d, ba_0r1d, ba_0a,
  ca_0r0d, ca_0r1d, ca_0a,
  mlength_0r0d, mlength_0r1d, mlength_0a,
  macc_0r0d, macc_0r1d, macc_0a
);
  input activate_0r;
  output activate_0a;
  output mType_0r;
  input [2:0] mType_0a0d;
  input [2:0] mType_0a1d;
  output a_0r;
  input [31:0] a_0a0d;
  input [31:0] a_0a1d;
  output b_0r;
  input [31:0] b_0a0d;
  input [31:0] b_0a1d;
  output c_0r;
  input [31:0] c_0a0d;
  input [31:0] c_0a1d;
  output [34:0] aa_0r0d;
  output [34:0] aa_0r1d;
  input aa_0a;
  output [35:0] ba_0r0d;
  output [35:0] ba_0r1d;
  input ba_0a;
  output [34:0] ca_0r0d;
  output [34:0] ca_0r1d;
  input ca_0a;
  output mlength_0r0d;
  output mlength_0r1d;
  input mlength_0a;
  output macc_0r0d;
  output macc_0r1d;
  input macc_0a;
  wire c52_r;
  wire c52_a;
  wire c51_r;
  wire c51_a;
  wire c50_r;
  wire c50_a;
  wire c49_r;
  wire c49_a;
  wire c48_r;
  wire c48_a;
  wire c47_r;
  wire c47_a;
  wire c46_r;
  wire c46_a;
  wire c45_r;
  wire c45_a;
  wire c44_r;
  wire c44_a;
  wire c43_r;
  wire c43_a;
  wire [2:0] c42_r0d;
  wire [2:0] c42_r1d;
  wire c42_a;
  wire c41_r;
  wire c41_a;
  wire c40_r;
  wire [2:0] c40_a0d;
  wire [2:0] c40_a1d;
  wire c39_r;
  wire c39_a;
  wire c38_r;
  wire c38_a;
  wire [34:0] c37_r0d;
  wire [34:0] c37_r1d;
  wire c37_a;
  wire c36_r;
  wire [34:0] c36_a0d;
  wire [34:0] c36_a1d;
  wire c35_r;
  wire [31:0] c35_a0d;
  wire [31:0] c35_a1d;
  wire c34_r;
  wire c34_a;
  wire [35:0] c33_r0d;
  wire [35:0] c33_r1d;
  wire c33_a;
  wire c32_r;
  wire [35:0] c32_a0d;
  wire [35:0] c32_a1d;
  wire c31_r;
  wire [32:0] c31_a0d;
  wire [32:0] c31_a1d;
  wire c30_r;
  wire c30_a0d;
  wire c30_a1d;
  wire c29_r;
  wire [31:0] c29_a0d;
  wire [31:0] c29_a1d;
  wire c28_r;
  wire c28_a;
  wire c27_r;
  wire c27_a;
  wire [34:0] c26_r0d;
  wire [34:0] c26_r1d;
  wire c26_a;
  wire c25_r;
  wire [34:0] c25_a0d;
  wire [34:0] c25_a1d;
  wire c24_r;
  wire [31:0] c24_a0d;
  wire [31:0] c24_a1d;
  wire c23_r;
  wire c23_a;
  wire [35:0] c22_r0d;
  wire [35:0] c22_r1d;
  wire c22_a;
  wire c21_r;
  wire [35:0] c21_a0d;
  wire [35:0] c21_a1d;
  wire c20_r;
  wire [32:0] c20_a0d;
  wire [32:0] c20_a1d;
  wire c19_r;
  wire c19_a0d;
  wire c19_a1d;
  wire c18_r;
  wire [31:0] c18_a0d;
  wire [31:0] c18_a1d;
  wire c17_r;
  wire c17_a;
  wire c16_r;
  wire [34:0] c16_a0d;
  wire [34:0] c16_a1d;
  wire c15_r;
  wire [31:0] c15_a0d;
  wire [31:0] c15_a1d;
  wire c14_r;
  wire c14_a;
  wire c13_r;
  wire c13_a0d;
  wire c13_a1d;
  wire c12_r;
  wire c12_a;
  wire c11_r;
  wire c11_a0d;
  wire c11_a1d;
  BrzFetch_1_s5_false I0 (c12_r, c12_a, c11_r, c11_a0d, c11_a1d, macc_0r0d, macc_0r1d, macc_0a);
  BrzFetch_1_s5_false I1 (c14_r, c14_a, c13_r, c13_a0d, c13_a1d, mlength_0r0d, mlength_0r1d, mlength_0a);
  BrzAdapt_35_32_s5_false_s5_false I2 (c16_r, c16_a0d[34:0], c16_a1d[34:0], c15_r, c15_a0d[31:0], c15_a1d[31:0]);
  BrzFetch_35_s5_false I3 (c17_r, c17_a, c16_r, c16_a0d[34:0], c16_a1d[34:0], ca_0r0d[34:0], ca_0r1d[34:0], ca_0a);
  BrzConstant_1_0 I4 (c19_r, c19_a0d, c19_a1d);
  BrzCombine_33_1_32 I5 (c20_r, c20_a0d[32:0], c20_a1d[32:0], c19_r, c19_a0d, c19_a1d, c18_r, c18_a0d[31:0], c18_a1d[31:0]);
  BrzAdapt_36_33_s4_true_s4_true I6 (c21_r, c21_a0d[35:0], c21_a1d[35:0], c20_r, c20_a0d[32:0], c20_a1d[32:0]);
  BrzFetch_36_s5_false I7 (c23_r, c23_a, c21_r, c21_a0d[35:0], c21_a1d[35:0], c22_r0d[35:0], c22_r1d[35:0], c22_a);
  BrzAdapt_35_32_s4_true_s4_true I8 (c25_r, c25_a0d[34:0], c25_a1d[34:0], c24_r, c24_a0d[31:0], c24_a1d[31:0]);
  BrzFetch_35_s5_false I9 (c27_r, c27_a, c25_r, c25_a0d[34:0], c25_a1d[34:0], c26_r0d[34:0], c26_r1d[34:0], c26_a);
  BrzConcur_2 I10 (c28_r, c28_a, c27_r, c27_a, c23_r, c23_a);
  BrzConstant_1_0 I11 (c30_r, c30_a0d, c30_a1d);
  BrzCombine_33_1_32 I12 (c31_r, c31_a0d[32:0], c31_a1d[32:0], c30_r, c30_a0d, c30_a1d, c29_r, c29_a0d[31:0], c29_a1d[31:0]);
  BrzAdapt_36_33_s5_false_s5_false I13 (c32_r, c32_a0d[35:0], c32_a1d[35:0], c31_r, c31_a0d[32:0], c31_a1d[32:0]);
  BrzFetch_36_s5_false I14 (c34_r, c34_a, c32_r, c32_a0d[35:0], c32_a1d[35:0], c33_r0d[35:0], c33_r1d[35:0], c33_a);
  BrzAdapt_35_32_s5_false_s5_false I15 (c36_r, c36_a0d[34:0], c36_a1d[34:0], c35_r, c35_a0d[31:0], c35_a1d[31:0]);
  BrzFetch_35_s5_false I16 (c38_r, c38_a, c36_r, c36_a0d[34:0], c36_a1d[34:0], c37_r0d[34:0], c37_r1d[34:0], c37_a);
  BrzConcur_2 I17 (c39_r, c39_a, c38_r, c38_a, c34_r, c34_a);
  BrzCallMux_35_2 I18 (c37_r0d[34:0], c37_r1d[34:0], c37_a, c26_r0d[34:0], c26_r1d[34:0], c26_a, aa_0r0d[34:0], aa_0r1d[34:0], aa_0a);
  BrzCallMux_36_2 I19 (c33_r0d[35:0], c33_r1d[35:0], c33_a, c22_r0d[35:0], c22_r1d[35:0], c22_a, ba_0r0d[35:0], ba_0r1d[35:0], ba_0a);
  BrzFetch_3_s5_false I20 (c41_r, c41_a, c40_r, c40_a0d[2:0], c40_a1d[2:0], c42_r0d[2:0], c42_r1d[2:0], c42_a);
  BrzCase_3_2_s25_1_2c3m4_2c2m4_3b5_2c4_2c0 I21 (c42_r0d[2:0], c42_r1d[2:0], c42_a, c28_r, c28_a, c39_r, c39_a);
  BrzConcur_4 I22 (c52_r, c52_a, c41_r, c41_a, c17_r, c17_a, c14_r, c14_a, c12_r, c12_a);
  BrzActiveEagerFalseVariable_3_3_s22__3b2_2_m1m I23 (c44_r, c44_a, mType_0r, mType_0a0d[2:0], mType_0a1d[2:0], c43_r, c43_a, c40_r, c40_a0d[2:0], c40_a1d[2:0], c13_r, c13_a0d, c13_a1d, c11_r, c11_a0d, c11_a1d);
  BrzActiveEagerFalseVariable_32_2_s0_ I24 (c46_r, c46_a, a_0r, a_0a0d[31:0], a_0a1d[31:0], c45_r, c45_a, c35_r, c35_a0d[31:0], c35_a1d[31:0], c24_r, c24_a0d[31:0], c24_a1d[31:0]);
  BrzActiveEagerFalseVariable_32_2_s0_ I25 (c48_r, c48_a, b_0r, b_0a0d[31:0], b_0a1d[31:0], c47_r, c47_a, c29_r, c29_a0d[31:0], c29_a1d[31:0], c18_r, c18_a0d[31:0], c18_a1d[31:0]);
  BrzActiveEagerFalseVariable_32_1_s0_ I26 (c50_r, c50_a, c_0r, c_0a0d[31:0], c_0a1d[31:0], c49_r, c49_a, c15_r, c15_a0d[31:0], c15_a1d[31:0]);
  BrzFork_4 I27 (c51_r, c51_a, c50_r, c50_a, c48_r, c48_a, c46_r, c46_a, c44_r, c44_a);
  BrzSynch_4 I28 (c49_r, c49_a, c47_r, c47_a, c45_r, c45_a, c43_r, c43_a, c52_r, c52_a);
  BrzLoop I29 (activate_0r, activate_0a, c51_r, c51_a);
endmodule

module Balsa_mControl10 (
  activate_0r, activate_0a,
  load_0r, load_0a0d, load_0a1d,
  done_0r0d, done_0r1d, done_0a
);
  input activate_0r;
  output activate_0a;
  output load_0r;
  input load_0a0d;
  input load_0a1d;
  output done_0r0d;
  output done_0r1d;
  input done_0a;
  wire [9:0] c31_r0d;
  wire [9:0] c31_r1d;
  wire c31_a;
  wire c30_r;
  wire c30_a;
  wire c29_r;
  wire c29_a;
  wire c28_r;
  wire c28_a;
  wire c27_r0d;
  wire c27_r1d;
  wire c27_a;
  wire c26_r;
  wire c26_a0d;
  wire c26_a1d;
  wire c25_r0d;
  wire c25_r1d;
  wire c25_a;
  wire c24_r;
  wire c24_a;
  wire c23_r;
  wire c23_a0d;
  wire c23_a1d;
  wire c22_r;
  wire c22_a;
  wire c21_r;
  wire c21_a;
  wire [9:0] c20_r0d;
  wire [9:0] c20_r1d;
  wire c20_a;
  wire c19_r;
  wire [9:0] c19_a0d;
  wire [9:0] c19_a1d;
  wire c18_r;
  wire c18_a;
  wire c17_r0d;
  wire c17_r1d;
  wire c17_a;
  wire c16_r;
  wire c16_a0d;
  wire c16_a1d;
  wire c15_r;
  wire c15_a;
  wire c14_r;
  wire c14_a;
  wire c13_r;
  wire c13_a;
  wire c12_r0d;
  wire c12_r1d;
  wire c12_a;
  wire c11_r;
  wire c11_a0d;
  wire c11_a1d;
  wire c10_r;
  wire c10_a;
  wire [9:0] c9_r0d;
  wire [9:0] c9_r1d;
  wire c9_a;
  wire c8_r;
  wire [9:0] c8_a0d;
  wire [9:0] c8_a1d;
  wire c7_r;
  wire [8:0] c7_a0d;
  wire [8:0] c7_a1d;
  wire c6_r;
  wire c6_a;
  wire [9:0] c5_r0d;
  wire [9:0] c5_r1d;
  wire c5_a;
  wire c4_r;
  wire [9:0] c4_a0d;
  wire [9:0] c4_a1d;
  BrzFetch_10_s5_false I0 (c6_r, c6_a, c4_r, c4_a0d[9:0], c4_a1d[9:0], c5_r0d[9:0], c5_r1d[9:0], c5_a);
  BrzAdapt_10_9_s5_false_s5_false I1 (c8_r, c8_a0d[9:0], c8_a1d[9:0], c7_r, c7_a0d[8:0], c7_a1d[8:0]);
  BrzFetch_10_s5_false I2 (c10_r, c10_a, c8_r, c8_a0d[9:0], c8_a1d[9:0], c9_r0d[9:0], c9_r1d[9:0], c9_a);
  BrzFetch_1_s5_false I3 (c13_r, c13_a, c11_r, c11_a0d, c11_a1d, c12_r0d, c12_r1d, c12_a);
  BrzConcur_2 I4 (c14_r, c14_a, c13_r, c13_a, c10_r, c10_a);
  BrzSequenceOptimised_2_s1_S I5 (c15_r, c15_a, c14_r, c14_a, c6_r, c6_a);
  BrzConstant_1_1 I6 (c16_r, c16_a0d, c16_a1d);
  BrzFetch_1_s5_false I7 (c18_r, c18_a, c16_r, c16_a0d, c16_a1d, c17_r0d, c17_r1d, c17_a);
  BrzConstant_10_511 I8 (c19_r, c19_a0d[9:0], c19_a1d[9:0]);
  BrzFetch_10_s5_false I9 (c21_r, c21_a, c19_r, c19_a0d[9:0], c19_a1d[9:0], c20_r0d[9:0], c20_r1d[9:0], c20_a);
  BrzConcur_2 I10 (c22_r, c22_a, c21_r, c21_a, c18_r, c18_a);
  BrzCallMux_1_2 I11 (c17_r0d, c17_r1d, c17_a, c12_r0d, c12_r1d, c12_a, done_0r0d, done_0r1d, done_0a);
  BrzFetch_1_s5_false I12 (c24_r, c24_a, c23_r, c23_a0d, c23_a1d, c25_r0d, c25_r1d, c25_a);
  BrzCase_1_2_s5_0_3b1 I13 (c25_r0d, c25_r1d, c25_a, c15_r, c15_a, c22_r, c22_a);
  BrzFetch_1_s5_false I14 (c28_r, c28_a, c26_r, c26_a0d, c26_a1d, c27_r0d, c27_r1d, c27_a);
  BrzActiveEagerFalseVariable_1_1_s0_ I15 (c29_r, c29_a, load_0r, load_0a0d, load_0a1d, c28_r, c28_a, c26_r, c26_a0d, c26_a1d);
  BrzSequenceOptimised_2_s1_T I16 (c30_r, c30_a, c29_r, c29_a, c24_r, c24_a);
  BrzLoop I17 (activate_0r, activate_0a, c30_r, c30_a);
  BrzVariable_10_1_s0_ I18 (c9_r0d[9:0], c9_r1d[9:0], c9_a, c4_r, c4_a0d[9:0], c4_a1d[9:0]);
  BrzCallMux_10_2 I19 (c5_r0d[9:0], c5_r1d[9:0], c5_a, c20_r0d[9:0], c20_r1d[9:0], c20_a, c31_r0d[9:0], c31_r1d[9:0], c31_a);
  BrzVariable_10_2_s19_0_2e_2e0_3b1_2e_2e9 I20 (c31_r0d[9:0], c31_r1d[9:0], c31_a, c11_r, c11_a0d, c11_a1d, c7_r, c7_a0d[8:0], c7_a1d[8:0]);
  BrzVariable_1_1_s0_ I21 (c27_r0d, c27_r1d, c27_a, c23_r, c23_a0d, c23_a1d);
endmodule

module Balsa_nanoMBoothR3rolled (
  activate_0r, activate_0a,
  cin_0r, cin_0a0d, cin_0a1d,
  res_0r, res_0a0d, res_0a1d,
  a_0r, a_0a0d, a_0a1d,
  b_0r, b_0a0d, b_0a1d,
  c_0r, c_0a0d, c_0a1d,
  mlength_0r, mlength_0a0d, mlength_0a1d,
  macc_0r, macc_0a0d, macc_0a1d,
  load_0r0d, load_0r1d, load_0a,
  done_0r, done_0a0d, done_0a1d,
  opA_0r0d, opA_0r1d, opA_0a,
  opB_0r0d, opB_0r1d, opB_0a,
  cs_0r0d, cs_0r1d, cs_0a,
  raA_0r0d, raA_0r1d, raA_0a,
  raB_0r0d, raB_0r1d, raB_0a,
  rac0_0r0d, rac0_0r1d, rac0_0a,
  raS_0r, raS_0a0d, raS_0a1d,
  racN_0r, racN_0a0d, racN_0a1d,
  pH_0r0d, pH_0r1d, pH_0a,
  pL_0r0d, pL_0r1d, pL_0a,
  z_0r0d, z_0r1d, z_0a,
  n_0r0d, n_0r1d, n_0a
);
  input activate_0r;
  output activate_0a;
  output cin_0r;
  input [34:0] cin_0a0d;
  input [34:0] cin_0a1d;
  output res_0r;
  input [34:0] res_0a0d;
  input [34:0] res_0a1d;
  output a_0r;
  input [34:0] a_0a0d;
  input [34:0] a_0a1d;
  output b_0r;
  input [35:0] b_0a0d;
  input [35:0] b_0a1d;
  output c_0r;
  input [34:0] c_0a0d;
  input [34:0] c_0a1d;
  output mlength_0r;
  input mlength_0a0d;
  input mlength_0a1d;
  output macc_0r;
  input macc_0a0d;
  input macc_0a1d;
  output load_0r0d;
  output load_0r1d;
  input load_0a;
  output done_0r;
  input done_0a0d;
  input done_0a1d;
  output [34:0] opA_0r0d;
  output [34:0] opA_0r1d;
  input opA_0a;
  output [34:0] opB_0r0d;
  output [34:0] opB_0r1d;
  input opB_0a;
  output [34:0] cs_0r0d;
  output [34:0] cs_0r1d;
  input cs_0a;
  output [31:0] raA_0r0d;
  output [31:0] raA_0r1d;
  input raA_0a;
  output [31:0] raB_0r0d;
  output [31:0] raB_0r1d;
  input raB_0a;
  output rac0_0r0d;
  output rac0_0r1d;
  input rac0_0a;
  output raS_0r;
  input [31:0] raS_0a0d;
  input [31:0] raS_0a1d;
  output racN_0r;
  input racN_0a0d;
  input racN_0a1d;
  output [31:0] pH_0r0d;
  output [31:0] pH_0r1d;
  input pH_0a;
  output [31:0] pL_0r0d;
  output [31:0] pL_0r1d;
  input pL_0a;
  output z_0r0d;
  output z_0r1d;
  input z_0a;
  output n_0r0d;
  output n_0r1d;
  input n_0a;
  wire c310_r0d;
  wire c310_r1d;
  wire c310_a;
  wire c309_r;
  wire [32:0] c309_a0d;
  wire [32:0] c309_a1d;
  wire c308_r;
  wire [1:0] c308_a0d;
  wire [1:0] c308_a1d;
  wire c307_r;
  wire [32:0] c307_a0d;
  wire [32:0] c307_a1d;
  wire c306_r;
  wire [1:0] c306_a0d;
  wire [1:0] c306_a1d;
  wire [3:0] c305_r0d;
  wire [3:0] c305_r1d;
  wire c305_a;
  wire [34:0] c304_r0d;
  wire [34:0] c304_r1d;
  wire c304_a;
  wire [34:0] c303_r0d;
  wire [34:0] c303_r1d;
  wire c303_a;
  wire [35:0] c302_r0d;
  wire [35:0] c302_r1d;
  wire c302_a;
  wire [35:0] c301_r0d;
  wire [35:0] c301_r1d;
  wire c301_a;
  wire c300_r0d;
  wire c300_r1d;
  wire c300_a;
  wire c299_r;
  wire c299_a;
  wire c298_r;
  wire c298_a;
  wire c297_r;
  wire c297_a;
  wire c296_r;
  wire c296_a;
  wire c295_r;
  wire c295_a;
  wire c294_r;
  wire c294_a;
  wire c293_r;
  wire c293_a;
  wire c292_r;
  wire c292_a;
  wire c291_r;
  wire c291_a;
  wire c290_r;
  wire c290_a;
  wire c289_r;
  wire c289_a;
  wire c288_r;
  wire c288_a;
  wire c287_r;
  wire c287_a;
  wire c286_r;
  wire c286_a;
  wire c285_r0d;
  wire c285_r1d;
  wire c285_a;
  wire c284_r;
  wire c284_a0d;
  wire c284_a1d;
  wire c283_r;
  wire c283_a;
  wire c282_r0d;
  wire c282_r1d;
  wire c282_a;
  wire c281_r;
  wire c281_a0d;
  wire c281_a1d;
  wire c280_r;
  wire c280_a;
  wire [34:0] c279_r0d;
  wire [34:0] c279_r1d;
  wire c279_a;
  wire c278_r;
  wire [34:0] c278_a0d;
  wire [34:0] c278_a1d;
  wire c277_r;
  wire c277_a;
  wire [34:0] c276_r0d;
  wire [34:0] c276_r1d;
  wire c276_a;
  wire c275_r;
  wire [34:0] c275_a0d;
  wire [34:0] c275_a1d;
  wire c274_r;
  wire c274_a0d;
  wire c274_a1d;
  wire c273_r;
  wire [33:0] c273_a0d;
  wire [33:0] c273_a1d;
  wire c272_r;
  wire c272_a;
  wire [34:0] c271_r0d;
  wire [34:0] c271_r1d;
  wire c271_a;
  wire c270_r;
  wire [34:0] c270_a0d;
  wire [34:0] c270_a1d;
  wire c269_r;
  wire [1:0] c269_a0d;
  wire [1:0] c269_a1d;
  wire c268_r;
  wire [32:0] c268_a0d;
  wire [32:0] c268_a1d;
  wire c267_r;
  wire c267_a;
  wire [31:0] c266_r0d;
  wire [31:0] c266_r1d;
  wire c266_a;
  wire c265_r;
  wire [31:0] c265_a0d;
  wire [31:0] c265_a1d;
  wire c264_r;
  wire c264_a;
  wire [31:0] c263_r0d;
  wire [31:0] c263_r1d;
  wire c263_a;
  wire c262_r;
  wire [31:0] c262_a0d;
  wire [31:0] c262_a1d;
  wire c261_r;
  wire [34:0] c261_a0d;
  wire [34:0] c261_a1d;
  wire c260_r;
  wire c260_a;
  wire c259_r;
  wire c259_a;
  wire c258_r;
  wire c258_a;
  wire c257_r;
  wire c257_a;
  wire c256_r;
  wire c256_a;
  wire c255_r;
  wire c255_a;
  wire c254_r;
  wire c254_a;
  wire [34:0] c253_r0d;
  wire [34:0] c253_r1d;
  wire c253_a;
  wire c252_r;
  wire [34:0] c252_a0d;
  wire [34:0] c252_a1d;
  wire c251_r;
  wire c251_a0d;
  wire c251_a1d;
  wire c250_r;
  wire [31:0] c250_a0d;
  wire [31:0] c250_a1d;
  wire c249_r;
  wire c249_a0d;
  wire c249_a1d;
  wire c248_r;
  wire c248_a0d;
  wire c248_a1d;
  wire c247_r;
  wire [31:0] c247_a0d;
  wire [31:0] c247_a1d;
  wire c246_r;
  wire c246_a0d;
  wire c246_a1d;
  wire c245_r;
  wire c245_a;
  wire [35:0] c244_r0d;
  wire [35:0] c244_r1d;
  wire c244_a;
  wire c243_r;
  wire [35:0] c243_a0d;
  wire [35:0] c243_a1d;
  wire c242_r;
  wire c242_a;
  wire [34:0] c241_r0d;
  wire [34:0] c241_r1d;
  wire c241_a;
  wire c240_r;
  wire [34:0] c240_a0d;
  wire [34:0] c240_a1d;
  wire c239_r;
  wire c239_a;
  wire [3:0] c238_r0d;
  wire [3:0] c238_r1d;
  wire c238_a;
  wire c237_r;
  wire [3:0] c237_a0d;
  wire [3:0] c237_a1d;
  wire c236_r;
  wire c236_a;
  wire [34:0] c235_r0d;
  wire [34:0] c235_r1d;
  wire c235_a;
  wire c234_r;
  wire [34:0] c234_a0d;
  wire [34:0] c234_a1d;
  wire c233_r;
  wire c233_a;
  wire [35:0] c232_r0d;
  wire [35:0] c232_r1d;
  wire c232_a;
  wire c231_r;
  wire [35:0] c231_a0d;
  wire [35:0] c231_a1d;
  wire c230_r;
  wire c230_a;
  wire c229_r;
  wire c229_a;
  wire [34:0] c228_r0d;
  wire [34:0] c228_r1d;
  wire c228_a;
  wire c227_r;
  wire [34:0] c227_a0d;
  wire [34:0] c227_a1d;
  wire c226_r;
  wire [34:0] c226_a0d;
  wire [34:0] c226_a1d;
  wire c225_r;
  wire c225_a;
  wire [34:0] c224_r0d;
  wire [34:0] c224_r1d;
  wire c224_a;
  wire c223_r;
  wire [34:0] c223_a0d;
  wire [34:0] c223_a1d;
  wire c222_r;
  wire [34:0] c222_a0d;
  wire [34:0] c222_a1d;
  wire c221_r;
  wire c221_a;
  wire [34:0] c220_r0d;
  wire [34:0] c220_r1d;
  wire c220_a;
  wire c219_r;
  wire [34:0] c219_a0d;
  wire [34:0] c219_a1d;
  wire c218_r;
  wire [34:0] c218_a0d;
  wire [34:0] c218_a1d;
  wire c217_r;
  wire c217_a;
  wire [34:0] c216_r0d;
  wire [34:0] c216_r1d;
  wire c216_a;
  wire c215_r;
  wire [34:0] c215_a0d;
  wire [34:0] c215_a1d;
  wire c214_r;
  wire [34:0] c214_a0d;
  wire [34:0] c214_a1d;
  wire c213_r;
  wire c213_a;
  wire c212_r;
  wire c212_a;
  wire c211_r;
  wire c211_a;
  wire c210_r;
  wire c210_a;
  wire c209_r;
  wire c209_a;
  wire c208_r;
  wire c208_a;
  wire c207_r;
  wire c207_a0d;
  wire c207_a1d;
  wire c206_r;
  wire c206_a;
  wire c205_r;
  wire c205_a;
  wire [34:0] c204_r0d;
  wire [34:0] c204_r1d;
  wire c204_a;
  wire c203_r;
  wire [34:0] c203_a0d;
  wire [34:0] c203_a1d;
  wire c202_r;
  wire [32:0] c202_a0d;
  wire [32:0] c202_a1d;
  wire c201_r;
  wire c201_a0d;
  wire c201_a1d;
  wire c200_r;
  wire c200_a0d;
  wire c200_a1d;
  wire c199_r;
  wire c199_a;
  wire [35:0] c198_r0d;
  wire [35:0] c198_r1d;
  wire c198_a;
  wire c197_r;
  wire [35:0] c197_a0d;
  wire [35:0] c197_a1d;
  wire c196_r;
  wire c196_a;
  wire [34:0] c195_r0d;
  wire [34:0] c195_r1d;
  wire c195_a;
  wire c194_r;
  wire [34:0] c194_a0d;
  wire [34:0] c194_a1d;
  wire c193_r;
  wire c193_a;
  wire [35:0] c192_r0d;
  wire [35:0] c192_r1d;
  wire c192_a;
  wire c191_r;
  wire [35:0] c191_a0d;
  wire [35:0] c191_a1d;
  wire c190_r;
  wire c190_a;
  wire [3:0] c189_r0d;
  wire [3:0] c189_r1d;
  wire c189_a;
  wire c188_r;
  wire [3:0] c188_a0d;
  wire [3:0] c188_a1d;
  wire c187_r;
  wire c187_a;
  wire c186_r;
  wire c186_a;
  wire c185_r;
  wire c185_a;
  wire c184_r;
  wire [34:0] c184_a0d;
  wire [34:0] c184_a1d;
  wire c183_r;
  wire c183_a;
  wire c182_r;
  wire [34:0] c182_a0d;
  wire [34:0] c182_a1d;
  wire c181_r;
  wire c181_a;
  wire [34:0] c180_r0d;
  wire [34:0] c180_r1d;
  wire c180_a;
  wire c179_r;
  wire c179_a;
  wire [34:0] c178_r0d;
  wire [34:0] c178_r1d;
  wire c178_a;
  wire c177_r;
  wire c177_a;
  wire c176_r0d;
  wire c176_r1d;
  wire c176_a;
  wire c175_r;
  wire c175_a0d;
  wire c175_a1d;
  wire [3:0] c174_r0d;
  wire [3:0] c174_r1d;
  wire c174_a;
  wire c173_r;
  wire c173_a;
  wire c172_r;
  wire [3:0] c172_a0d;
  wire [3:0] c172_a1d;
  wire c171_r;
  wire c171_a;
  wire [34:0] c170_r0d;
  wire [34:0] c170_r1d;
  wire c170_a;
  wire c169_r;
  wire [34:0] c169_a0d;
  wire [34:0] c169_a1d;
  wire c168_r;
  wire c168_a;
  wire [34:0] c167_r0d;
  wire [34:0] c167_r1d;
  wire c167_a;
  wire c166_r;
  wire [34:0] c166_a0d;
  wire [34:0] c166_a1d;
  wire c165_r;
  wire c165_a;
  wire [34:0] c164_r0d;
  wire [34:0] c164_r1d;
  wire c164_a;
  wire c163_r;
  wire [34:0] c163_a0d;
  wire [34:0] c163_a1d;
  wire c162_r;
  wire c162_a;
  wire [34:0] c161_r0d;
  wire [34:0] c161_r1d;
  wire c161_a;
  wire c160_r;
  wire [34:0] c160_a0d;
  wire [34:0] c160_a1d;
  wire c159_r;
  wire c159_a;
  wire [34:0] c158_r0d;
  wire [34:0] c158_r1d;
  wire c158_a;
  wire c157_r;
  wire [34:0] c157_a0d;
  wire [34:0] c157_a1d;
  wire c156_r;
  wire c156_a;
  wire [34:0] c155_r0d;
  wire [34:0] c155_r1d;
  wire c155_a;
  wire c154_r;
  wire [34:0] c154_a0d;
  wire [34:0] c154_a1d;
  wire c153_r;
  wire c153_a;
  wire [34:0] c152_r0d;
  wire [34:0] c152_r1d;
  wire c152_a;
  wire c151_r;
  wire [34:0] c151_a0d;
  wire [34:0] c151_a1d;
  wire c150_r;
  wire c150_a;
  wire [34:0] c149_r0d;
  wire [34:0] c149_r1d;
  wire c149_a;
  wire c148_r;
  wire [34:0] c148_a0d;
  wire [34:0] c148_a1d;
  wire c147_r;
  wire c147_a;
  wire [34:0] c146_r0d;
  wire [34:0] c146_r1d;
  wire c146_a;
  wire c145_r;
  wire [34:0] c145_a0d;
  wire [34:0] c145_a1d;
  wire c144_r;
  wire [3:0] c144_a0d;
  wire [3:0] c144_a1d;
  wire c143_r;
  wire c143_a;
  wire c142_r;
  wire c142_a;
  wire c141_r;
  wire c141_a;
  wire c140_r;
  wire c140_a;
  wire c139_r;
  wire c139_a;
  wire c138_r;
  wire c138_a;
  wire c137_r;
  wire c137_a;
  wire c136_r;
  wire c136_a;
  wire c135_r;
  wire c135_a;
  wire [34:0] c134_r0d;
  wire [34:0] c134_r1d;
  wire c134_a;
  wire c133_r;
  wire [34:0] c133_a0d;
  wire [34:0] c133_a1d;
  wire c132_r;
  wire c132_a;
  wire [35:0] c131_r0d;
  wire [35:0] c131_r1d;
  wire c131_a;
  wire c130_r;
  wire [35:0] c130_a0d;
  wire [35:0] c130_a1d;
  wire c129_r;
  wire [34:0] c129_a0d;
  wire [34:0] c129_a1d;
  wire c128_r;
  wire [31:0] c128_a0d;
  wire [31:0] c128_a1d;
  wire c127_r;
  wire c127_a0d;
  wire c127_a1d;
  wire c126_r;
  wire [1:0] c126_a0d;
  wire [1:0] c126_a1d;
  wire c125_r;
  wire c125_a;
  wire [34:0] c124_r0d;
  wire [34:0] c124_r1d;
  wire c124_a;
  wire c123_r;
  wire [34:0] c123_a0d;
  wire [34:0] c123_a1d;
  wire c122_r;
  wire [31:0] c122_a0d;
  wire [31:0] c122_a1d;
  wire c121_r;
  wire c121_a;
  wire [35:0] c120_r0d;
  wire [35:0] c120_r1d;
  wire c120_a;
  wire c119_r;
  wire [35:0] c119_a0d;
  wire [35:0] c119_a1d;
  wire c118_r;
  wire [34:0] c118_a0d;
  wire [34:0] c118_a1d;
  wire c117_r;
  wire [31:0] c117_a0d;
  wire [31:0] c117_a1d;
  wire c116_r;
  wire [2:0] c116_a0d;
  wire [2:0] c116_a1d;
  wire c115_r;
  wire [34:0] c115_a0d;
  wire [34:0] c115_a1d;
  wire c114_r;
  wire [34:0] c114_a0d;
  wire [34:0] c114_a1d;
  wire c113_r;
  wire c113_a0d;
  wire c113_a1d;
  wire c112_r;
  wire c112_a;
  wire c111_r;
  wire c111_a;
  wire c110_r0d;
  wire c110_r1d;
  wire c110_a;
  wire c109_r;
  wire c109_a0d;
  wire c109_a1d;
  wire c108_r;
  wire c108_a;
  wire c107_r;
  wire c107_a;
  wire [31:0] c106_r0d;
  wire [31:0] c106_r1d;
  wire c106_a;
  wire c105_r;
  wire [31:0] c105_a0d;
  wire [31:0] c105_a1d;
  wire c104_r;
  wire c104_a;
  wire [31:0] c103_r0d;
  wire [31:0] c103_r1d;
  wire c103_a;
  wire c102_r;
  wire [31:0] c102_a0d;
  wire [31:0] c102_a1d;
  wire c101_r;
  wire c101_a;
  wire c100_r;
  wire c100_a;
  wire c99_r;
  wire c99_a;
  wire c98_r;
  wire c98_a;
  wire c97_r;
  wire c97_a;
  wire c96_r;
  wire c96_a;
  wire c95_r;
  wire c95_a;
  wire c94_r;
  wire c94_a;
  wire [31:0] c93_r0d;
  wire [31:0] c93_r1d;
  wire c93_a;
  wire c92_r;
  wire [31:0] c92_a0d;
  wire [31:0] c92_a1d;
  wire c91_r;
  wire c91_a;
  wire c90_r0d;
  wire c90_r1d;
  wire c90_a;
  wire c89_r;
  wire c89_a0d;
  wire c89_a1d;
  wire c88_r;
  wire c88_a;
  wire c87_r0d;
  wire c87_r1d;
  wire c87_a;
  wire c86_r;
  wire c86_a0d;
  wire c86_a1d;
  wire c85_r;
  wire c85_a;
  wire c84_r0d;
  wire c84_r1d;
  wire c84_a;
  wire c83_r;
  wire c83_a0d;
  wire c83_a1d;
  wire c82_r;
  wire [31:0] c82_a0d;
  wire [31:0] c82_a1d;
  wire c81_r;
  wire [31:0] c81_a0d;
  wire [31:0] c81_a1d;
  wire c80_r;
  wire c80_a0d;
  wire c80_a1d;
  wire c79_r0d;
  wire c79_r1d;
  wire c79_a;
  wire c78_r;
  wire c78_a;
  wire c77_r;
  wire c77_a0d;
  wire c77_a1d;
  wire c76_r;
  wire c76_a;
  wire c75_r;
  wire c75_a;
  wire c74_r;
  wire c74_a;
  wire [31:0] c73_r0d;
  wire [31:0] c73_r1d;
  wire c73_a;
  wire c72_r;
  wire [31:0] c72_a0d;
  wire [31:0] c72_a1d;
  wire c71_r;
  wire c71_a0d;
  wire c71_a1d;
  wire c70_r;
  wire [30:0] c70_a0d;
  wire [30:0] c70_a1d;
  wire c69_r;
  wire c69_a;
  wire [31:0] c68_r0d;
  wire [31:0] c68_r1d;
  wire c68_a;
  wire c67_r;
  wire [31:0] c67_a0d;
  wire [31:0] c67_a1d;
  wire c66_r;
  wire c66_a;
  wire c65_r0d;
  wire c65_r1d;
  wire c65_a;
  wire c64_r;
  wire c64_a0d;
  wire c64_a1d;
  wire c63_r;
  wire c63_a;
  wire c62_r;
  wire c62_a;
  wire c61_r;
  wire c61_a;
  wire c60_r;
  wire c60_a;
  wire c59_r;
  wire c59_a;
  wire c58_r;
  wire c58_a;
  wire [31:0] c57_r0d;
  wire [31:0] c57_r1d;
  wire c57_a;
  wire c56_r;
  wire [31:0] c56_a0d;
  wire [31:0] c56_a1d;
  wire c55_r;
  wire [31:0] c55_a0d;
  wire [31:0] c55_a1d;
  wire c54_r;
  wire c54_a0d;
  wire c54_a1d;
  wire c53_r;
  wire c53_a;
  wire c52_r;
  wire c52_a;
  wire c51_r;
  wire [31:0] c51_a0d;
  wire [31:0] c51_a1d;
  wire c50_r;
  wire c50_a;
  wire [31:0] c49_r0d;
  wire [31:0] c49_r1d;
  wire c49_a;
  wire c48_r;
  wire [31:0] c48_a0d;
  wire [31:0] c48_a1d;
  wire c47_r0d;
  wire c47_r1d;
  wire c47_a;
  wire c46_r;
  wire c46_a;
  wire c45_r;
  wire c45_a0d;
  wire c45_a1d;
  wire c44_r;
  wire c44_a;
  wire c43_r0d;
  wire c43_r1d;
  wire c43_a;
  wire c42_r;
  wire c42_a0d;
  wire c42_a1d;
  wire c41_r;
  wire c41_a;
  wire c40_r0d;
  wire c40_r1d;
  wire c40_a;
  wire c39_r;
  wire c39_a0d;
  wire c39_a1d;
  wire c38_r;
  wire c38_a0d;
  wire c38_a1d;
  wire c37_r;
  wire [31:0] c37_a0d;
  wire [31:0] c37_a1d;
  wire c36_r;
  wire c36_a0d;
  wire c36_a1d;
  wire c35_r;
  wire c35_a;
  wire c34_r0d;
  wire c34_r1d;
  wire c34_a;
  wire c33_r;
  wire c33_a0d;
  wire c33_a1d;
  wire c32_r;
  wire c32_a;
  wire c31_r;
  wire c31_a;
  wire [31:0] c30_r0d;
  wire [31:0] c30_r1d;
  wire c30_a;
  wire c29_r;
  wire [31:0] c29_a0d;
  wire [31:0] c29_a1d;
  wire c28_r;
  wire c28_a;
  wire c27_r0d;
  wire c27_r1d;
  wire c27_a;
  wire c26_r;
  wire c26_a0d;
  wire c26_a1d;
  wire c25_r;
  wire c25_a;
  wire c24_r0d;
  wire c24_r1d;
  wire c24_a;
  wire c23_r;
  wire c23_a0d;
  wire c23_a1d;
  BrzEncode_1_2_s5_0_3b0 I0 (c260_r, c260_a, c101_r, c101_a, c310_r0d, c310_r1d, c310_a);
  BrzEncode_1_2_s5_1_3b0 I1 (c213_r, c213_a, c187_r, c187_a, load_0r0d, load_0r1d, load_0a);
  BrzCombineEqual_2_1_2 I2 (c306_r, c306_a0d[1:0], c306_a1d[1:0], c249_r, c249_a0d, c249_a1d, c248_r, c248_a0d, c248_a1d);
  BrzCombine_33_1_32 I3 (c307_r, c307_a0d[32:0], c307_a1d[32:0], c251_r, c251_a0d, c251_a1d, c250_r, c250_a0d[31:0], c250_a1d[31:0]);
  BrzCombine_35_33_2 I4 (c252_r, c252_a0d[34:0], c252_a1d[34:0], c307_r, c307_a0d[32:0], c307_a1d[32:0], c306_r, c306_a0d[1:0], c306_a1d[1:0]);
  BrzCombineEqual_2_1_2 I5 (c308_r, c308_a0d[1:0], c308_a1d[1:0], c201_r, c201_a0d, c201_a1d, c200_r, c200_a0d, c200_a1d);
  BrzCombine_35_33_2 I6 (c203_r, c203_a0d[34:0], c203_a1d[34:0], c202_r, c202_a0d[32:0], c202_a1d[32:0], c308_r, c308_a0d[1:0], c308_a1d[1:0]);
  BrzCombine_33_32_1 I7 (c309_r, c309_a0d[32:0], c309_a1d[32:0], c128_r, c128_a0d[31:0], c128_a1d[31:0], c127_r, c127_a0d, c127_a1d);
  BrzCombine_35_33_2 I8 (c129_r, c129_a0d[34:0], c129_a1d[34:0], c309_r, c309_a0d[32:0], c309_a1d[32:0], c126_r, c126_a0d[1:0], c126_a1d[1:0]);
  BrzFetch_1_s5_false I9 (c25_r, c25_a, c23_r, c23_a0d, c23_a1d, c24_r0d, c24_r1d, c24_a);
  BrzFetch_1_s5_false I10 (c28_r, c28_a, c26_r, c26_a0d, c26_a1d, c27_r0d, c27_r1d, c27_a);
  BrzFetch_32_s5_false I11 (c31_r, c31_a, c29_r, c29_a0d[31:0], c29_a1d[31:0], c30_r0d[31:0], c30_r1d[31:0], c30_a);
  BrzConcur_3 I12 (c32_r, c32_a, c31_r, c31_a, c28_r, c28_a, c25_r, c25_a);
  BrzFetch_1_s5_false I13 (c35_r, c35_a, c33_r, c33_a0d, c33_a1d, c34_r0d, c34_r1d, c34_a);
  BrzBinaryFuncConstR_1_32_1_s6_Equals_s5_fa_m25m I14 (c38_r, c38_a0d, c38_a1d, c37_r, c37_a0d[31:0], c37_a1d[31:0]);
  BrzBinaryFunc_1_1_1_s3_And_s5_false_s5_fal_m15m I15 (c39_r, c39_a0d, c39_a1d, c38_r, c38_a0d, c38_a1d, c36_r, c36_a0d, c36_a1d);
  BrzFetch_1_s5_false I16 (c41_r, c41_a, c39_r, c39_a0d, c39_a1d, c40_r0d, c40_r1d, c40_a);
  BrzFetch_1_s5_false I17 (c44_r, c44_a, c42_r, c42_a0d, c42_a1d, c43_r0d, c43_r1d, c43_a);
  BrzFetch_1_s5_false I18 (c46_r, c46_a, c45_r, c45_a0d, c45_a1d, c47_r0d, c47_r1d, c47_a);
  BrzCase_1_2_s5_0_3b1 I19 (c47_r0d, c47_r1d, c47_a, c41_r, c41_a, c44_r, c44_a);
  BrzFetch_32_s5_false I20 (c50_r, c50_a, c48_r, c48_a0d[31:0], c48_a1d[31:0], c49_r0d[31:0], c49_r1d[31:0], c49_a);
  BrzFetch_32_s5_false I21 (c52_r, c52_a, c51_r, c51_a0d[31:0], c51_a1d[31:0], pH_0r0d[31:0], pH_0r1d[31:0], pH_0a);
  BrzConcur_4 I22 (c53_r, c53_a, c52_r, c52_a, c50_r, c50_a, c46_r, c46_a, c35_r, c35_a);
  BrzFetch_32_s5_false I23 (c63_r, c63_a, c56_r, c56_a0d[31:0], c56_a1d[31:0], c57_r0d[31:0], c57_r1d[31:0], c57_a);
  BrzActiveEagerFalseVariable_32_1_s0_ I24 (c59_r, c59_a, c55_r, c55_a0d[31:0], c55_a1d[31:0], c58_r, c58_a, c56_r, c56_a0d[31:0], c56_a1d[31:0]);
  BrzActiveEagerNullAdapt_1 I25 (c60_r, c60_a, c54_r, c54_a0d, c54_a1d, c61_r, c61_a);
  BrzFork_2 I26 (c62_r, c62_a, c60_r, c60_a, c59_r, c59_a);
  BrzSynch_2 I27 (c61_r, c61_a, c58_r, c58_a, c63_r, c63_a);
  BrzFetch_1_s5_false I28 (c66_r, c66_a, c64_r, c64_a0d, c64_a1d, c65_r0d, c65_r1d, c65_a);
  BrzFetch_32_s5_false I29 (c69_r, c69_a, c67_r, c67_a0d[31:0], c67_a1d[31:0], c68_r0d[31:0], c68_r1d[31:0], c68_a);
  BrzCombine_32_1_31 I30 (c72_r, c72_a0d[31:0], c72_a1d[31:0], c71_r, c71_a0d, c71_a1d, c70_r, c70_a0d[30:0], c70_a1d[30:0]);
  BrzFetch_32_s5_false I31 (c74_r, c74_a, c72_r, c72_a0d[31:0], c72_a1d[31:0], c73_r0d[31:0], c73_r1d[31:0], c73_a);
  BrzConcur_4 I32 (c75_r, c75_a, c74_r, c74_a, c69_r, c69_a, c66_r, c66_a, c62_r, c62_a);
  BrzSequenceOptimised_2_s1_S I33 (c76_r, c76_a, c75_r, c75_a, c53_r, c53_a);
  BrzCallMux_32_2 I34 (c49_r0d[31:0], c49_r1d[31:0], c49_a, c30_r0d[31:0], c30_r1d[31:0], c30_a, pL_0r0d[31:0], pL_0r1d[31:0], pL_0a);
  BrzCallMux_1_3 I35 (c43_r0d, c43_r1d, c43_a, c40_r0d, c40_r1d, c40_a, c27_r0d, c27_r1d, c27_a, z_0r0d, z_0r1d, z_0a);
  BrzCallMux_1_2 I36 (c34_r0d, c34_r1d, c34_a, c24_r0d, c24_r1d, c24_a, n_0r0d, n_0r1d, n_0a);
  BrzFetch_1_s5_false I37 (c78_r, c78_a, c77_r, c77_a0d, c77_a1d, c79_r0d, c79_r1d, c79_a);
  BrzCase_1_2_s5_0_3b1 I38 (c79_r0d, c79_r1d, c79_a, c32_r, c32_a, c76_r, c76_a);
  BrzBinaryFuncConstR_1_32_1_s6_Equals_s5_fa_m25m I39 (c83_r, c83_a0d, c83_a1d, c82_r, c82_a0d[31:0], c82_a1d[31:0]);
  BrzFetch_1_s5_false I40 (c85_r, c85_a, c83_r, c83_a0d, c83_a1d, c84_r0d, c84_r1d, c84_a);
  BrzFetch_1_s5_false I41 (c88_r, c88_a, c86_r, c86_a0d, c86_a1d, c87_r0d, c87_r1d, c87_a);
  BrzFetch_1_s5_false I42 (c91_r, c91_a, c89_r, c89_a0d, c89_a1d, c90_r0d, c90_r1d, c90_a);
  BrzFetch_32_s5_false I43 (c94_r, c94_a, c92_r, c92_a0d[31:0], c92_a1d[31:0], c93_r0d[31:0], c93_r1d[31:0], c93_a);
  BrzConcur_4 I44 (c100_r, c100_a, c94_r, c94_a, c91_r, c91_a, c88_r, c88_a, c85_r, c85_a);
  BrzActiveEagerFalseVariable_32_3_s13__3b31_m3m I45 (c96_r, c96_a, c81_r, c81_a0d[31:0], c81_a1d[31:0], c95_r, c95_a, c92_r, c92_a0d[31:0], c92_a1d[31:0], c86_r, c86_a0d, c86_a1d, c82_r, c82_a0d[31:0], c82_a1d[31:0]);
  BrzActiveEagerFalseVariable_1_1_s0_ I46 (c98_r, c98_a, c80_r, c80_a0d, c80_a1d, c97_r, c97_a, c89_r, c89_a0d, c89_a1d);
  BrzFork_2 I47 (c99_r, c99_a, c98_r, c98_a, c96_r, c96_a);
  BrzSynch_2 I48 (c97_r, c97_a, c95_r, c95_a, c100_r, c100_a);
  BrzFetch_32_s5_false I49 (c104_r, c104_a, c102_r, c102_a0d[31:0], c102_a1d[31:0], c103_r0d[31:0], c103_r1d[31:0], c103_a);
  BrzFetch_32_s5_false I50 (c107_r, c107_a, c105_r, c105_a0d[31:0], c105_a1d[31:0], c106_r0d[31:0], c106_r1d[31:0], c106_a);
  BrzConcur_4 I51 (c108_r, c108_a, c107_r, c107_a, c104_r, c104_a, c101_r, c101_a, c99_r, c99_a);
  BrzFetch_1_s5_false I52 (c111_r, c111_a, c109_r, c109_a0d, c109_a1d, c110_r0d, c110_r1d, c110_a);
  BrzActiveEagerFalseVariable_1_1_s0_ I53 (c112_r, c112_a, done_0r, done_0a0d, done_0a1d, c111_r, c111_a, c109_r, c109_a0d, c109_a1d);
  BrzCombine_35_32_3 I54 (c118_r, c118_a0d[34:0], c118_a1d[34:0], c117_r, c117_a0d[31:0], c117_a1d[31:0], c116_r, c116_a0d[2:0], c116_a1d[2:0]);
  BrzAdapt_36_35_s5_false_s5_false I55 (c119_r, c119_a0d[35:0], c119_a1d[35:0], c118_r, c118_a0d[34:0], c118_a1d[34:0]);
  BrzFetch_36_s5_false I56 (c121_r, c121_a, c119_r, c119_a0d[35:0], c119_a1d[35:0], c120_r0d[35:0], c120_r1d[35:0], c120_a);
  BrzAdapt_35_32_s4_true_s4_true I57 (c123_r, c123_a0d[34:0], c123_a1d[34:0], c122_r, c122_a0d[31:0], c122_a1d[31:0]);
  BrzFetch_35_s5_false I58 (c125_r, c125_a, c123_r, c123_a0d[34:0], c123_a1d[34:0], c124_r0d[34:0], c124_r1d[34:0], c124_a);
  BrzAdapt_36_35_s5_false_s5_false I59 (c130_r, c130_a0d[35:0], c130_a1d[35:0], c129_r, c129_a0d[34:0], c129_a1d[34:0]);
  BrzFetch_36_s5_false I60 (c132_r, c132_a, c130_r, c130_a0d[35:0], c130_a1d[35:0], c131_r0d[35:0], c131_r1d[35:0], c131_a);
  BrzFetch_35_s5_false I61 (c135_r, c135_a, c133_r, c133_a0d[34:0], c133_a1d[34:0], c134_r0d[34:0], c134_r1d[34:0], c134_a);
  BrzConcur_4 I62 (c143_r, c143_a, c135_r, c135_a, c132_r, c132_a, c125_r, c125_a, c121_r, c121_a);
  BrzActiveEagerFalseVariable_1_1_s0_ I63 (c137_r, c137_a, c113_r, c113_a0d, c113_a1d, c136_r, c136_a, c127_r, c127_a0d, c127_a1d);
  BrzActiveEagerFalseVariable_35_2_s11__3b0__m9m I64 (c139_r, c139_a, c114_r, c114_a0d[34:0], c114_a1d[34:0], c138_r, c138_a, c133_r, c133_a0d[34:0], c133_a1d[34:0], c126_r, c126_a0d[1:0], c126_a1d[1:0]);
  BrzActiveEagerFalseVariable_35_2_s20_3_2e__m7m I65 (c141_r, c141_a, c115_r, c115_a0d[34:0], c115_a1d[34:0], c140_r, c140_a, c122_r, c122_a0d[31:0], c122_a1d[31:0], c116_r, c116_a0d[2:0], c116_a1d[2:0]);
  BrzFork_3 I66 (c142_r, c142_a, c141_r, c141_a, c139_r, c139_a, c137_r, c137_a);
  BrzSynch_3 I67 (c140_r, c140_a, c138_r, c138_a, c136_r, c136_a, c143_r, c143_a);
  BrzAdapt_35_4_s4_true_s4_true I68 (c145_r, c145_a0d[34:0], c145_a1d[34:0], c144_r, c144_a0d[3:0], c144_a1d[3:0]);
  BrzFetch_35_s5_false I69 (c147_r, c147_a, c145_r, c145_a0d[34:0], c145_a1d[34:0], c146_r0d[34:0], c146_r1d[34:0], c146_a);
  BrzFetch_35_s5_false I70 (c150_r, c150_a, c148_r, c148_a0d[34:0], c148_a1d[34:0], c149_r0d[34:0], c149_r1d[34:0], c149_a);
  BrzFetch_35_s5_false I71 (c153_r, c153_a, c151_r, c151_a0d[34:0], c151_a1d[34:0], c152_r0d[34:0], c152_r1d[34:0], c152_a);
  BrzFetch_35_s5_false I72 (c156_r, c156_a, c154_r, c154_a0d[34:0], c154_a1d[34:0], c155_r0d[34:0], c155_r1d[34:0], c155_a);
  BrzFetch_35_s5_false I73 (c159_r, c159_a, c157_r, c157_a0d[34:0], c157_a1d[34:0], c158_r0d[34:0], c158_r1d[34:0], c158_a);
  BrzFetch_35_s5_false I74 (c162_r, c162_a, c160_r, c160_a0d[34:0], c160_a1d[34:0], c161_r0d[34:0], c161_r1d[34:0], c161_a);
  BrzFetch_35_s5_false I75 (c165_r, c165_a, c163_r, c163_a0d[34:0], c163_a1d[34:0], c164_r0d[34:0], c164_r1d[34:0], c164_a);
  BrzFetch_35_s5_false I76 (c168_r, c168_a, c166_r, c166_a0d[34:0], c166_a1d[34:0], c167_r0d[34:0], c167_r1d[34:0], c167_a);
  BrzFetch_35_s5_false I77 (c171_r, c171_a, c169_r, c169_a0d[34:0], c169_a1d[34:0], c170_r0d[34:0], c170_r1d[34:0], c170_a);
  BrzCallMux_35_9 I78 (c170_r0d[34:0], c170_r1d[34:0], c170_a, c167_r0d[34:0], c167_r1d[34:0], c167_a, c164_r0d[34:0], c164_r1d[34:0], c164_a, c161_r0d[34:0], c161_r1d[34:0], c161_a, c158_r0d[34:0], c158_r1d[34:0], c158_a, c155_r0d[34:0], c155_r1d[34:0], c155_a, c152_r0d[34:0], c152_r1d[34:0], c152_a, c149_r0d[34:0], c149_r1d[34:0], c149_a, c146_r0d[34:0], c146_r1d[34:0], c146_a, opB_0r0d[34:0], opB_0r1d[34:0], opB_0a);
  BrzFetch_4_s5_false I79 (c173_r, c173_a, c172_r, c172_a0d[3:0], c172_a1d[3:0], c174_r0d[3:0], c174_r1d[3:0], c174_a);
  BrzCase_4_9_s67_15_2c0_3b2_2c1_3b4_2c3_3b6_m27m I80 (c174_r0d[3:0], c174_r1d[3:0], c174_a, c147_r, c147_a, c150_r, c150_a, c153_r, c153_a, c156_r, c156_a, c159_r, c159_a, c162_r, c162_a, c165_r, c165_a, c168_r, c168_a, c171_r, c171_a);
  BrzFetch_1_s5_false I81 (c177_r, c177_a, c175_r, c175_a0d, c175_a1d, c176_r0d, c176_r1d, c176_a);
  BrzFetch_35_s4_true I82 (c179_r, c179_a, cin_0r, cin_0a0d[34:0], cin_0a1d[34:0], c178_r0d[34:0], c178_r1d[34:0], c178_a);
  BrzFetch_35_s4_true I83 (c181_r, c181_a, res_0r, res_0a0d[34:0], res_0a1d[34:0], c180_r0d[34:0], c180_r1d[34:0], c180_a);
  BrzFetch_35_s5_false I84 (c183_r, c183_a, c182_r, c182_a0d[34:0], c182_a1d[34:0], cs_0r0d[34:0], cs_0r1d[34:0], cs_0a);
  BrzFetch_35_s5_false I85 (c185_r, c185_a, c184_r, c184_a0d[34:0], c184_a1d[34:0], opA_0r0d[34:0], opA_0r1d[34:0], opA_0a);
  BrzConcur_8 I86 (c186_r, c186_a, c185_r, c185_a, c183_r, c183_a, c181_r, c181_a, c179_r, c179_a, c177_r, c177_a, c173_r, c173_a, c142_r, c142_a, c112_r, c112_a);
  BrzPassivatorPush_1_1 I87 (c113_r, c113_a0d, c113_a1d, c176_r0d, c176_r1d, c176_a);
  BrzPassivatorPush_35_1 I88 (c114_r, c114_a0d[34:0], c114_a1d[34:0], c178_r0d[34:0], c178_r1d[34:0], c178_a);
  BrzPassivatorPush_35_1 I89 (c115_r, c115_a0d[34:0], c115_a1d[34:0], c180_r0d[34:0], c180_r1d[34:0], c180_a);
  BrzFetch_4_s5_false I90 (c190_r, c190_a, c188_r, c188_a0d[3:0], c188_a1d[3:0], c189_r0d[3:0], c189_r1d[3:0], c189_a);
  BrzFetch_36_s5_false I91 (c193_r, c193_a, c191_r, c191_a0d[35:0], c191_a1d[35:0], c192_r0d[35:0], c192_r1d[35:0], c192_a);
  BrzFetch_35_s5_false I92 (c196_r, c196_a, c194_r, c194_a0d[34:0], c194_a1d[34:0], c195_r0d[34:0], c195_r1d[34:0], c195_a);
  BrzFetch_36_s5_false I93 (c199_r, c199_a, c197_r, c197_a0d[35:0], c197_a1d[35:0], c198_r0d[35:0], c198_r1d[35:0], c198_a);
  BrzFetch_35_s5_false I94 (c205_r, c205_a, c203_r, c203_a0d[34:0], c203_a1d[34:0], c204_r0d[34:0], c204_r1d[34:0], c204_a);
  BrzConcur_6 I95 (c206_r, c206_a, c205_r, c205_a, c199_r, c199_a, c196_r, c196_a, c193_r, c193_a, c190_r, c190_a, c187_r, c187_a);
  BrzWhile I96 (c211_r, c211_a, c207_r, c207_a0d, c207_a1d, c212_r, c212_a);
  BrzCall_2 I97 (c210_r, c210_a, c209_r, c209_a, c186_r, c186_a);
  BrzSequenceOptimised_2_s1_S I98 (c208_r, c208_a, c210_r, c210_a, c211_r, c211_a);
  BrzSequenceOptimised_2_s1_S I99 (c212_r, c212_a, c206_r, c206_a, c209_r, c209_a);
  BrzUnaryFunc_35_35_s6_Invert_s5_false I100 (c215_r, c215_a0d[34:0], c215_a1d[34:0], c214_r, c214_a0d[34:0], c214_a1d[34:0]);
  BrzFetch_35_s5_false I101 (c217_r, c217_a, c215_r, c215_a0d[34:0], c215_a1d[34:0], c216_r0d[34:0], c216_r1d[34:0], c216_a);
  BrzUnaryFunc_35_35_s6_Invert_s5_false I102 (c219_r, c219_a0d[34:0], c219_a1d[34:0], c218_r, c218_a0d[34:0], c218_a1d[34:0]);
  BrzFetch_35_s5_false I103 (c221_r, c221_a, c219_r, c219_a0d[34:0], c219_a1d[34:0], c220_r0d[34:0], c220_r1d[34:0], c220_a);
  BrzUnaryFunc_35_35_s6_Invert_s5_false I104 (c223_r, c223_a0d[34:0], c223_a1d[34:0], c222_r, c222_a0d[34:0], c222_a1d[34:0]);
  BrzFetch_35_s5_false I105 (c225_r, c225_a, c223_r, c223_a0d[34:0], c223_a1d[34:0], c224_r0d[34:0], c224_r1d[34:0], c224_a);
  BrzUnaryFunc_35_35_s6_Invert_s5_false I106 (c227_r, c227_a0d[34:0], c227_a1d[34:0], c226_r, c226_a0d[34:0], c226_a1d[34:0]);
  BrzFetch_35_s5_false I107 (c229_r, c229_a, c227_r, c227_a0d[34:0], c227_a1d[34:0], c228_r0d[34:0], c228_r1d[34:0], c228_a);
  BrzConcur_5 I108 (c230_r, c230_a, c229_r, c229_a, c225_r, c225_a, c221_r, c221_a, c217_r, c217_a, c213_r, c213_a);
  BrzConstant_36_0 I109 (c231_r, c231_a0d[35:0], c231_a1d[35:0]);
  BrzFetch_36_s5_false I110 (c233_r, c233_a, c231_r, c231_a0d[35:0], c231_a1d[35:0], c232_r0d[35:0], c232_r1d[35:0], c232_a);
  BrzConstant_35_0 I111 (c234_r, c234_a0d[34:0], c234_a1d[34:0]);
  BrzFetch_35_s5_false I112 (c236_r, c236_a, c234_r, c234_a0d[34:0], c234_a1d[34:0], c235_r0d[34:0], c235_r1d[34:0], c235_a);
  BrzFetch_4_s5_false I113 (c239_r, c239_a, c237_r, c237_a0d[3:0], c237_a1d[3:0], c238_r0d[3:0], c238_r1d[3:0], c238_a);
  BrzFetch_35_s5_false I114 (c242_r, c242_a, c240_r, c240_a0d[34:0], c240_a1d[34:0], c241_r0d[34:0], c241_r1d[34:0], c241_a);
  BrzFetch_36_s5_false I115 (c245_r, c245_a, c243_r, c243_a0d[35:0], c243_a1d[35:0], c244_r0d[35:0], c244_r1d[35:0], c244_a);
  BrzFetch_35_s5_false I116 (c259_r, c259_a, c252_r, c252_a0d[34:0], c252_a1d[34:0], c253_r0d[34:0], c253_r1d[34:0], c253_a);
  BrzActiveEagerFalseVariable_32_1_s0_ I117 (c255_r, c255_a, c247_r, c247_a0d[31:0], c247_a1d[31:0], c254_r, c254_a, c250_r, c250_a0d[31:0], c250_a1d[31:0]);
  BrzActiveEagerFalseVariable_1_1_s0_ I118 (c257_r, c257_a, c246_r, c246_a0d, c246_a1d, c256_r, c256_a, c249_r, c249_a0d, c249_a1d);
  BrzFork_2 I119 (c258_r, c258_a, c257_r, c257_a, c255_r, c255_a);
  BrzSynch_2 I120 (c256_r, c256_a, c254_r, c254_a, c259_r, c259_a);
  BrzAdapt_32_35_s5_false_s5_false I121 (c262_r, c262_a0d[31:0], c262_a1d[31:0], c261_r, c261_a0d[34:0], c261_a1d[34:0]);
  BrzFetch_32_s5_false I122 (c264_r, c264_a, c262_r, c262_a0d[31:0], c262_a1d[31:0], c263_r0d[31:0], c263_r1d[31:0], c263_a);
  BrzFetch_32_s5_false I123 (c267_r, c267_a, c265_r, c265_a0d[31:0], c265_a1d[31:0], c266_r0d[31:0], c266_r1d[31:0], c266_a);
  BrzConstant_2_0 I124 (c269_r, c269_a0d[1:0], c269_a1d[1:0]);
  BrzCombine_35_2_33 I125 (c270_r, c270_a0d[34:0], c270_a1d[34:0], c269_r, c269_a0d[1:0], c269_a1d[1:0], c268_r, c268_a0d[32:0], c268_a1d[32:0]);
  BrzFetch_35_s5_false I126 (c272_r, c272_a, c270_r, c270_a0d[34:0], c270_a1d[34:0], c271_r0d[34:0], c271_r1d[34:0], c271_a);
  BrzConstant_1_0 I127 (c274_r, c274_a0d, c274_a1d);
  BrzCombine_35_1_34 I128 (c275_r, c275_a0d[34:0], c275_a1d[34:0], c274_r, c274_a0d, c274_a1d, c273_r, c273_a0d[33:0], c273_a1d[33:0]);
  BrzFetch_35_s5_false I129 (c277_r, c277_a, c275_r, c275_a0d[34:0], c275_a1d[34:0], c276_r0d[34:0], c276_r1d[34:0], c276_a);
  BrzFetch_35_s5_false I130 (c280_r, c280_a, c278_r, c278_a0d[34:0], c278_a1d[34:0], c279_r0d[34:0], c279_r1d[34:0], c279_a);
  BrzFetch_1_s5_false I131 (c283_r, c283_a, c281_r, c281_a0d, c281_a1d, c282_r0d, c282_r1d, c282_a);
  BrzFetch_1_s5_false I132 (c286_r, c286_a, c284_r, c284_a0d, c284_a1d, c285_r0d, c285_r1d, c285_a);
  BrzConcur_14 I133 (c298_r, c298_a, c286_r, c286_a, c283_r, c283_a, c280_r, c280_a, c277_r, c277_a, c272_r, c272_a, c267_r, c267_a, c264_r, c264_a, c260_r, c260_a, c258_r, c258_a, c245_r, c245_a, c242_r, c242_a, c239_r, c239_a, c236_r, c236_a, c233_r, c233_a);
  BrzActiveEagerFalseVariable_35_7_s63__3b0__m11m I134 (c288_r, c288_a, a_0r, a_0a0d[34:0], a_0a1d[34:0], c287_r, c287_a, c278_r, c278_a0d[34:0], c278_a1d[34:0], c273_r, c273_a0d[33:0], c273_a1d[33:0], c268_r, c268_a0d[32:0], c268_a1d[32:0], c265_r, c265_a0d[31:0], c265_a1d[31:0], c261_r, c261_a0d[34:0], c261_a1d[34:0], c251_r, c251_a0d, c251_a1d, c248_r, c248_a0d, c248_a1d);
  BrzActiveEagerFalseVariable_36_2_s11__3b0__m13m I135 (c290_r, c290_a, b_0r, b_0a0d[35:0], b_0a1d[35:0], c289_r, c289_a, c243_r, c243_a0d[35:0], c243_a1d[35:0], c237_r, c237_a0d[3:0], c237_a1d[3:0]);
  BrzActiveEagerFalseVariable_35_1_s0_ I136 (c292_r, c292_a, c_0r, c_0a0d[34:0], c_0a1d[34:0], c291_r, c291_a, c240_r, c240_a0d[34:0], c240_a1d[34:0]);
  BrzActiveEagerFalseVariable_1_1_s0_ I137 (c294_r, c294_a, mlength_0r, mlength_0a0d, mlength_0a1d, c293_r, c293_a, c284_r, c284_a0d, c284_a1d);
  BrzActiveEagerFalseVariable_1_1_s0_ I138 (c296_r, c296_a, macc_0r, macc_0a0d, macc_0a1d, c295_r, c295_a, c281_r, c281_a0d, c281_a1d);
  BrzFork_5 I139 (c297_r, c297_a, c296_r, c296_a, c294_r, c294_a, c292_r, c292_a, c290_r, c290_a, c288_r, c288_a);
  BrzSynch_5 I140 (c295_r, c295_a, c293_r, c293_a, c291_r, c291_a, c289_r, c289_a, c287_r, c287_a, c298_r, c298_a);
  BrzSequenceOptimised_5_s4_SSSS I141 (c299_r, c299_a, c297_r, c297_a, c230_r, c230_a, c208_r, c208_a, c108_r, c108_a, c78_r, c78_a);
  BrzCallMux_32_3 I142 (c266_r0d[31:0], c266_r1d[31:0], c266_a, c106_r0d[31:0], c106_r1d[31:0], c106_a, c73_r0d[31:0], c73_r1d[31:0], c73_a, raA_0r0d[31:0], raA_0r1d[31:0], raA_0a);
  BrzCallMux_32_3 I143 (c263_r0d[31:0], c263_r1d[31:0], c263_a, c103_r0d[31:0], c103_r1d[31:0], c103_a, c68_r0d[31:0], c68_r1d[31:0], c68_a, raB_0r0d[31:0], raB_0r1d[31:0], raB_0a);
  BrzCallMux_1_2 I144 (c310_r0d, c310_r1d, c310_a, c65_r0d, c65_r1d, c65_a, rac0_0r0d, rac0_0r1d, rac0_0a);
  BrzCallDemux_32_3 I145 (c247_r, c247_a0d[31:0], c247_a1d[31:0], c81_r, c81_a0d[31:0], c81_a1d[31:0], c55_r, c55_a0d[31:0], c55_a1d[31:0], raS_0r, raS_0a0d[31:0], raS_0a1d[31:0]);
  BrzCallDemux_1_3 I146 (c246_r, c246_a0d, c246_a1d, c80_r, c80_a0d, c80_a1d, c54_r, c54_a0d, c54_a1d, racN_0r, racN_0a0d, racN_0a1d);
  BrzLoop I147 (activate_0r, activate_0a, c299_r, c299_a);
  BrzVariable_1_1_s0_ I148 (c87_r0d, c87_r1d, c87_a, c23_r, c23_a0d, c23_a1d);
  BrzVariable_1_3_s0_ I149 (c84_r0d, c84_r1d, c84_a, c42_r, c42_a0d, c42_a1d, c36_r, c36_a0d, c36_a1d, c26_r, c26_a0d, c26_a1d);
  BrzVariable_1_1_s0_ I150 (c282_r0d, c282_r1d, c282_a, c45_r, c45_a0d, c45_a1d);
  BrzVariable_1_1_s0_ I151 (c285_r0d, c285_r1d, c285_a, c77_r, c77_a0d, c77_a1d);
  BrzCallMux_1_2 I152 (c90_r0d, c90_r1d, c90_a, c110_r0d, c110_r1d, c110_a, c300_r0d, c300_r1d, c300_a);
  BrzVariable_1_2_s0_ I153 (c300_r0d, c300_r1d, c300_a, c207_r, c207_a0d, c207_a1d, c64_r, c64_a0d, c64_a1d);
  BrzCallMux_36_2 I154 (c192_r0d[35:0], c192_r1d[35:0], c192_a, c244_r0d[35:0], c244_r1d[35:0], c244_a, c301_r0d[35:0], c301_r1d[35:0], c301_a);
  BrzVariable_36_1_s9_3_2e_2e34 I155 (c301_r0d[35:0], c301_r1d[35:0], c301_a, c117_r, c117_a0d[31:0], c117_a1d[31:0]);
  BrzCallMux_36_2 I156 (c198_r0d[35:0], c198_r1d[35:0], c198_a, c232_r0d[35:0], c232_r1d[35:0], c232_a, c302_r0d[35:0], c302_r1d[35:0], c302_a);
  BrzVariable_36_1_s9_3_2e_2e34 I157 (c302_r0d[35:0], c302_r1d[35:0], c302_a, c128_r, c128_a0d[31:0], c128_a1d[31:0]);
  BrzCallMux_35_2 I158 (c204_r0d[34:0], c204_r1d[34:0], c204_a, c235_r0d[34:0], c235_r1d[34:0], c235_a, c303_r0d[34:0], c303_r1d[34:0], c303_a);
  BrzVariable_35_1_s0_ I159 (c303_r0d[34:0], c303_r1d[34:0], c303_a, c182_r, c182_a0d[34:0], c182_a1d[34:0]);
  BrzCallMux_35_2 I160 (c195_r0d[34:0], c195_r1d[34:0], c195_a, c241_r0d[34:0], c241_r1d[34:0], c241_a, c304_r0d[34:0], c304_r1d[34:0], c304_a);
  BrzVariable_35_1_s0_ I161 (c304_r0d[34:0], c304_r1d[34:0], c304_a, c184_r, c184_a0d[34:0], c184_a1d[34:0]);
  BrzVariable_36_4_s36__3b0_2e_2e3_3b2_2e_2e_m31m I162 (c120_r0d[35:0], c120_r1d[35:0], c120_a, c191_r, c191_a0d[35:0], c191_a1d[35:0], c188_r, c188_a0d[3:0], c188_a1d[3:0], c105_r, c105_a0d[31:0], c105_a1d[31:0], c71_r, c71_a0d, c71_a1d);
  BrzVariable_35_2_s12__3b0_2e_2e30 I163 (c124_r0d[34:0], c124_r1d[34:0], c124_a, c194_r, c194_a0d[34:0], c194_a1d[34:0], c70_r, c70_a0d[30:0], c70_a1d[30:0]);
  BrzVariable_36_2_s12__3b2_2e_2e33 I164 (c131_r0d[35:0], c131_r1d[35:0], c131_a, c197_r, c197_a0d[35:0], c197_a1d[35:0], c102_r, c102_a0d[31:0], c102_a1d[31:0]);
  BrzVariable_35_4_s47_2_2e_2e34_3b34_2e_2e3_m29m I165 (c134_r0d[34:0], c134_r1d[34:0], c134_a, c202_r, c202_a0d[32:0], c202_a1d[32:0], c201_r, c201_a0d, c201_a1d, c200_r, c200_a0d, c200_a1d, c67_r, c67_a0d[31:0], c67_a1d[31:0]);
  BrzVariable_35_1_s0_ I166 (c216_r0d[34:0], c216_r1d[34:0], c216_a, c160_r, c160_a0d[34:0], c160_a1d[34:0]);
  BrzVariable_35_1_s0_ I167 (c220_r0d[34:0], c220_r1d[34:0], c220_a, c163_r, c163_a0d[34:0], c163_a1d[34:0]);
  BrzVariable_35_1_s0_ I168 (c224_r0d[34:0], c224_r1d[34:0], c224_a, c166_r, c166_a0d[34:0], c166_a1d[34:0]);
  BrzVariable_35_1_s0_ I169 (c228_r0d[34:0], c228_r1d[34:0], c228_a, c169_r, c169_a0d[34:0], c169_a1d[34:0]);
  BrzVariable_35_2_s0_ I170 (c271_r0d[34:0], c271_r1d[34:0], c271_a, c214_r, c214_a0d[34:0], c214_a1d[34:0], c157_r, c157_a0d[34:0], c157_a1d[34:0]);
  BrzVariable_35_2_s0_ I171 (c253_r0d[34:0], c253_r1d[34:0], c253_a, c218_r, c218_a0d[34:0], c218_a1d[34:0], c154_r, c154_a0d[34:0], c154_a1d[34:0]);
  BrzVariable_35_2_s0_ I172 (c276_r0d[34:0], c276_r1d[34:0], c276_a, c222_r, c222_a0d[34:0], c222_a1d[34:0], c151_r, c151_a0d[34:0], c151_a1d[34:0]);
  BrzVariable_35_2_s0_ I173 (c279_r0d[34:0], c279_r1d[34:0], c279_a, c226_r, c226_a0d[34:0], c226_a1d[34:0], c148_r, c148_a0d[34:0], c148_a1d[34:0]);
  BrzVariable_32_2_s0_ I174 (c93_r0d[31:0], c93_r1d[31:0], c93_a, c48_r, c48_a0d[31:0], c48_a1d[31:0], c29_r, c29_a0d[31:0], c29_a1d[31:0]);
  BrzVariable_32_3_s16__3b_3b31_2e_2e31 I175 (c57_r0d[31:0], c57_r1d[31:0], c57_a, c51_r, c51_a0d[31:0], c51_a1d[31:0], c37_r, c37_a0d[31:0], c37_a1d[31:0], c33_r, c33_a0d, c33_a1d);
  BrzCallMux_4_2 I176 (c189_r0d[3:0], c189_r1d[3:0], c189_a, c238_r0d[3:0], c238_r1d[3:0], c238_a, c305_r0d[3:0], c305_r1d[3:0], c305_a);
  BrzVariable_4_3_s8_3_2e_2e3 I177 (c305_r0d[3:0], c305_r1d[3:0], c305_a, c175_r, c175_a0d, c175_a1d, c144_r, c144_a0d[3:0], c144_a1d[3:0], c172_r, c172_a0d[3:0], c172_a1d[3:0]);
endmodule

module Balsa_nanoSpaMultiplier (
  activate_0r, activate_0a,
  bypass_0r0d, bypass_0r1d, bypass_0a,
  bypassH_0r0d, bypassH_0r1d, bypassH_0a,
  mType_0r0d, mType_0r1d, mType_0a,
  a_0r0d, a_0r1d, a_0a,
  b_0r0d, b_0r1d, b_0a,
  c_0r0d, c_0r1d, c_0a,
  mpH_0r0d, mpH_0r1d, mpH_0a,
  mpL_0r0d, mpL_0r1d, mpL_0a,
  mZ_0r0d, mZ_0r1d, mZ_0a,
  mN_0r0d, mN_0r1d, mN_0a
);
  input activate_0r;
  output activate_0a;
  input bypass_0r0d;
  input bypass_0r1d;
  output bypass_0a;
  input bypassH_0r0d;
  input bypassH_0r1d;
  output bypassH_0a;
  input [2:0] mType_0r0d;
  input [2:0] mType_0r1d;
  output mType_0a;
  input [31:0] a_0r0d;
  input [31:0] a_0r1d;
  output a_0a;
  input [31:0] b_0r0d;
  input [31:0] b_0r1d;
  output b_0a;
  input [31:0] c_0r0d;
  input [31:0] c_0r1d;
  output c_0a;
  output [31:0] mpH_0r0d;
  output [31:0] mpH_0r1d;
  input mpH_0a;
  output [31:0] mpL_0r0d;
  output [31:0] mpL_0r1d;
  input mpL_0a;
  output mZ_0r0d;
  output mZ_0r1d;
  input mZ_0a;
  output mN_0r0d;
  output mN_0r1d;
  input mN_0a;
  wire c114_r;
  wire c114_a;
  wire c113_r;
  wire c113_a;
  wire c112_r;
  wire c112_a;
  wire c111_r;
  wire c111_a;
  wire c110_r0d;
  wire c110_r1d;
  wire c110_a;
  wire c109_r;
  wire c109_a0d;
  wire c109_a1d;
  wire c108_r;
  wire c108_a;
  wire c107_r;
  wire c107_a;
  wire c106_r;
  wire c106_a;
  wire c105_r;
  wire c105_a;
  wire c104_r0d;
  wire c104_r1d;
  wire c104_a;
  wire c103_r;
  wire c103_a0d;
  wire c103_a1d;
  wire c102_r;
  wire c102_a;
  wire c101_r;
  wire c101_a;
  wire c100_r;
  wire c100_a;
  wire c99_r;
  wire c99_a;
  wire [2:0] c98_r0d;
  wire [2:0] c98_r1d;
  wire c98_a;
  wire c97_r;
  wire [2:0] c97_a0d;
  wire [2:0] c97_a1d;
  wire c96_r;
  wire c96_a;
  wire c95_r;
  wire c95_a;
  wire c94_r;
  wire c94_a;
  wire c93_r;
  wire c93_a;
  wire [31:0] c92_r0d;
  wire [31:0] c92_r1d;
  wire c92_a;
  wire c91_r;
  wire [31:0] c91_a0d;
  wire [31:0] c91_a1d;
  wire c90_r;
  wire c90_a;
  wire c89_r;
  wire c89_a;
  wire c88_r;
  wire c88_a;
  wire c87_r;
  wire c87_a;
  wire [31:0] c86_r0d;
  wire [31:0] c86_r1d;
  wire c86_a;
  wire c85_r;
  wire [31:0] c85_a0d;
  wire [31:0] c85_a1d;
  wire c84_r;
  wire c84_a;
  wire c83_r;
  wire c83_a;
  wire c82_r;
  wire c82_a;
  wire c81_r;
  wire c81_a;
  wire [31:0] c80_r0d;
  wire [31:0] c80_r1d;
  wire c80_a;
  wire c79_r;
  wire [31:0] c79_a0d;
  wire [31:0] c79_a1d;
  wire c78_r;
  wire c78_a;
  wire c77_r;
  wire [34:0] c77_a0d;
  wire [34:0] c77_a1d;
  wire c76_r;
  wire [34:0] c76_a0d;
  wire [34:0] c76_a1d;
  wire c75_r;
  wire [34:0] c75_a0d;
  wire [34:0] c75_a1d;
  wire [34:0] c74_r0d;
  wire [34:0] c74_r1d;
  wire c74_a;
  wire [34:0] c73_r0d;
  wire [34:0] c73_r1d;
  wire c73_a;
  wire c72_r;
  wire c72_a;
  wire c71_r;
  wire [31:0] c71_a0d;
  wire [31:0] c71_a1d;
  wire c70_r;
  wire [31:0] c70_a0d;
  wire [31:0] c70_a1d;
  wire c69_r;
  wire c69_a0d;
  wire c69_a1d;
  wire [31:0] c68_r0d;
  wire [31:0] c68_r1d;
  wire c68_a;
  wire c67_r0d;
  wire c67_r1d;
  wire c67_a;
  wire c66_r;
  wire c66_a;
  wire c65_r;
  wire [34:0] c65_a0d;
  wire [34:0] c65_a1d;
  wire c64_r;
  wire [34:0] c64_a0d;
  wire [34:0] c64_a1d;
  wire c63_r;
  wire [34:0] c63_a0d;
  wire [34:0] c63_a1d;
  wire c62_r;
  wire [35:0] c62_a0d;
  wire [35:0] c62_a1d;
  wire c61_r;
  wire [34:0] c61_a0d;
  wire [34:0] c61_a1d;
  wire c60_r;
  wire c60_a0d;
  wire c60_a1d;
  wire c59_r;
  wire c59_a0d;
  wire c59_a1d;
  wire c58_r0d;
  wire c58_r1d;
  wire c58_a;
  wire c57_r;
  wire c57_a0d;
  wire c57_a1d;
  wire [34:0] c56_r0d;
  wire [34:0] c56_r1d;
  wire c56_a;
  wire [34:0] c55_r0d;
  wire [34:0] c55_r1d;
  wire c55_a;
  wire [34:0] c54_r0d;
  wire [34:0] c54_r1d;
  wire c54_a;
  wire [31:0] c53_r0d;
  wire [31:0] c53_r1d;
  wire c53_a;
  wire [31:0] c52_r0d;
  wire [31:0] c52_r1d;
  wire c52_a;
  wire c51_r0d;
  wire c51_r1d;
  wire c51_a;
  wire c50_r;
  wire [31:0] c50_a0d;
  wire [31:0] c50_a1d;
  wire c49_r;
  wire c49_a0d;
  wire c49_a1d;
  wire [31:0] c48_r0d;
  wire [31:0] c48_r1d;
  wire c48_a;
  wire [31:0] c47_r0d;
  wire [31:0] c47_r1d;
  wire c47_a;
  wire c46_r0d;
  wire c46_r1d;
  wire c46_a;
  wire c45_r0d;
  wire c45_r1d;
  wire c45_a;
  wire c44_r;
  wire c44_a;
  wire c43_r;
  wire c43_a0d;
  wire c43_a1d;
  wire c42_r0d;
  wire c42_r1d;
  wire c42_a;
  wire c41_r;
  wire c41_a;
  wire c40_r;
  wire [2:0] c40_a0d;
  wire [2:0] c40_a1d;
  wire c39_r;
  wire [31:0] c39_a0d;
  wire [31:0] c39_a1d;
  wire c38_r;
  wire [31:0] c38_a0d;
  wire [31:0] c38_a1d;
  wire c37_r;
  wire [31:0] c37_a0d;
  wire [31:0] c37_a1d;
  wire [34:0] c36_r0d;
  wire [34:0] c36_r1d;
  wire c36_a;
  wire [35:0] c35_r0d;
  wire [35:0] c35_r1d;
  wire c35_a;
  wire [34:0] c34_r0d;
  wire [34:0] c34_r1d;
  wire c34_a;
  wire c33_r0d;
  wire c33_r1d;
  wire c33_a;
  wire c32_r0d;
  wire c32_r1d;
  wire c32_a;
  wire c31_r;
  wire c31_a;
  wire c30_r;
  wire c30_a0d;
  wire c30_a1d;
  wire c29_r;
  wire c29_a0d;
  wire c29_a1d;
  wire c28_r;
  wire [31:0] c28_a0d;
  wire [31:0] c28_a1d;
  wire c27_r;
  wire [31:0] c27_a0d;
  wire [31:0] c27_a1d;
  wire c26_r;
  wire [31:0] c26_a0d;
  wire [31:0] c26_a1d;
  wire c25_r;
  wire [2:0] c25_a0d;
  wire [2:0] c25_a1d;
  wire [31:0] c24_r0d;
  wire [31:0] c24_r1d;
  wire c24_a;
  wire [31:0] c23_r0d;
  wire [31:0] c23_r1d;
  wire c23_a;
  wire [31:0] c22_r0d;
  wire [31:0] c22_r1d;
  wire c22_a;
  wire [2:0] c21_r0d;
  wire [2:0] c21_r1d;
  wire c21_a;
  wire c20_r0d;
  wire c20_r1d;
  wire c20_a;
  wire c19_r0d;
  wire c19_r1d;
  wire c19_a;
  wire c18_r;
  wire c18_a;
  wire c17_r;
  wire c17_a0d;
  wire c17_a1d;
  wire c16_r;
  wire c16_a0d;
  wire c16_a1d;
  wire c15_r;
  wire [31:0] c15_a0d;
  wire [31:0] c15_a1d;
  wire c14_r;
  wire [31:0] c14_a0d;
  wire [31:0] c14_a1d;
  wire c13_r;
  wire c13_a0d;
  wire c13_a1d;
  wire c12_r;
  wire c12_a0d;
  wire c12_a1d;
  Balsa_doByPass I0 (c18_r, c18_a, c17_r, c17_a0d, c17_a1d, c16_r, c16_a0d, c16_a1d, c15_r, c15_a0d[31:0], c15_a1d[31:0], c14_r, c14_a0d[31:0], c14_a1d[31:0], c13_r, c13_a0d, c13_a1d, c12_r, c12_a0d, c12_a1d, mpH_0r0d[31:0], mpH_0r1d[31:0], mpH_0a, mpL_0r0d[31:0], mpL_0r1d[31:0], mpL_0a, mZ_0r0d, mZ_0r1d, mZ_0a, mN_0r0d, mN_0r1d, mN_0a);
  Balsa_bypassMul I1 (c31_r, c31_a, c30_r, c30_a0d, c30_a1d, c29_r, c29_a0d, c29_a1d, c28_r, c28_a0d[31:0], c28_a1d[31:0], c27_r, c27_a0d[31:0], c27_a1d[31:0], c26_r, c26_a0d[31:0], c26_a1d[31:0], c25_r, c25_a0d[2:0], c25_a1d[2:0], c24_r0d[31:0], c24_r1d[31:0], c24_a, c23_r0d[31:0], c23_r1d[31:0], c23_a, c22_r0d[31:0], c22_r1d[31:0], c22_a, c21_r0d[2:0], c21_r1d[2:0], c21_a, c20_r0d, c20_r1d, c20_a, c19_r0d, c19_r1d, c19_a);
  Balsa_signAdj I2 (c41_r, c41_a, c40_r, c40_a0d[2:0], c40_a1d[2:0], c39_r, c39_a0d[31:0], c39_a1d[31:0], c38_r, c38_a0d[31:0], c38_a1d[31:0], c37_r, c37_a0d[31:0], c37_a1d[31:0], c36_r0d[34:0], c36_r1d[34:0], c36_a, c35_r0d[35:0], c35_r1d[35:0], c35_a, c34_r0d[34:0], c34_r1d[34:0], c34_a, c33_r0d, c33_r1d, c33_a, c32_r0d, c32_r1d, c32_a);
  Balsa_mControl10 I3 (c44_r, c44_a, c43_r, c43_a0d, c43_a1d, c42_r0d, c42_r1d, c42_a);
  Balsa_nanoMBoothR3rolled I4 (c66_r, c66_a, c65_r, c65_a0d[34:0], c65_a1d[34:0], c64_r, c64_a0d[34:0], c64_a1d[34:0], c63_r, c63_a0d[34:0], c63_a1d[34:0], c62_r, c62_a0d[35:0], c62_a1d[35:0], c61_r, c61_a0d[34:0], c61_a1d[34:0], c60_r, c60_a0d, c60_a1d, c59_r, c59_a0d, c59_a1d, c58_r0d, c58_r1d, c58_a, c57_r, c57_a0d, c57_a1d, c56_r0d[34:0], c56_r1d[34:0], c56_a, c55_r0d[34:0], c55_r1d[34:0], c55_a, c54_r0d[34:0], c54_r1d[34:0], c54_a, c53_r0d[31:0], c53_r1d[31:0], c53_a, c52_r0d[31:0], c52_r1d[31:0], c52_a, c51_r0d, c51_r1d, c51_a, c50_r, c50_a0d[31:0], c50_a1d[31:0],
		c49_r, c49_a0d, c49_a1d, c48_r0d[31:0], c48_r1d[31:0], c48_a, c47_r0d[31:0], c47_r1d[31:0], c47_a, c46_r0d, c46_r1d, c46_a, c45_r0d, c45_r1d, c45_a);
  Balsa_CPadder I5 (c72_r, c72_a, c71_r, c71_a0d[31:0], c71_a1d[31:0], c70_r, c70_a0d[31:0], c70_a1d[31:0], c69_r, c69_a0d, c69_a1d, c68_r0d[31:0], c68_r1d[31:0], c68_a, c67_r0d, c67_r1d, c67_a);
  Balsa_CSAdder__DP2 I6 (c78_r, c78_a, c77_r, c77_a0d[34:0], c77_a1d[34:0], c76_r, c76_a0d[34:0], c76_a1d[34:0], c75_r, c75_a0d[34:0], c75_a1d[34:0], c74_r0d[34:0], c74_r1d[34:0], c74_a, c73_r0d[34:0], c73_r1d[34:0], c73_a);
  BrzFetch_32_s5_false I7 (c81_r, c81_a, c79_r, c79_a0d[31:0], c79_a1d[31:0], c80_r0d[31:0], c80_r1d[31:0], c80_a);
  BrzFalseVariable_32_1_s0_ I8 (c_0r0d[31:0], c_0r1d[31:0], c_0a, c82_r, c82_a, c79_r, c79_a0d[31:0], c79_a1d[31:0]);
  BrzDecisionWait_1 I9 (c83_r, c83_a, c82_r, c82_a, c81_r, c81_a);
  BrzLoop I10 (c84_r, c84_a, c83_r, c83_a);
  BrzFetch_32_s5_false I11 (c87_r, c87_a, c85_r, c85_a0d[31:0], c85_a1d[31:0], c86_r0d[31:0], c86_r1d[31:0], c86_a);
  BrzFalseVariable_32_1_s0_ I12 (b_0r0d[31:0], b_0r1d[31:0], b_0a, c88_r, c88_a, c85_r, c85_a0d[31:0], c85_a1d[31:0]);
  BrzDecisionWait_1 I13 (c89_r, c89_a, c88_r, c88_a, c87_r, c87_a);
  BrzLoop I14 (c90_r, c90_a, c89_r, c89_a);
  BrzFetch_32_s5_false I15 (c93_r, c93_a, c91_r, c91_a0d[31:0], c91_a1d[31:0], c92_r0d[31:0], c92_r1d[31:0], c92_a);
  BrzFalseVariable_32_1_s0_ I16 (a_0r0d[31:0], a_0r1d[31:0], a_0a, c94_r, c94_a, c91_r, c91_a0d[31:0], c91_a1d[31:0]);
  BrzDecisionWait_1 I17 (c95_r, c95_a, c94_r, c94_a, c93_r, c93_a);
  BrzLoop I18 (c96_r, c96_a, c95_r, c95_a);
  BrzFetch_3_s5_false I19 (c99_r, c99_a, c97_r, c97_a0d[2:0], c97_a1d[2:0], c98_r0d[2:0], c98_r1d[2:0], c98_a);
  BrzFalseVariable_3_1_s0_ I20 (mType_0r0d[2:0], mType_0r1d[2:0], mType_0a, c100_r, c100_a, c97_r, c97_a0d[2:0], c97_a1d[2:0]);
  BrzDecisionWait_1 I21 (c101_r, c101_a, c100_r, c100_a, c99_r, c99_a);
  BrzLoop I22 (c102_r, c102_a, c101_r, c101_a);
  BrzFetch_1_s5_false I23 (c105_r, c105_a, c103_r, c103_a0d, c103_a1d, c104_r0d, c104_r1d, c104_a);
  BrzFalseVariable_1_1_s0_ I24 (bypassH_0r0d, bypassH_0r1d, bypassH_0a, c106_r, c106_a, c103_r, c103_a0d, c103_a1d);
  BrzDecisionWait_1 I25 (c107_r, c107_a, c106_r, c106_a, c105_r, c105_a);
  BrzLoop I26 (c108_r, c108_a, c107_r, c107_a);
  BrzFetch_1_s5_false I27 (c111_r, c111_a, c109_r, c109_a0d, c109_a1d, c110_r0d, c110_r1d, c110_a);
  BrzFalseVariable_1_1_s0_ I28 (bypass_0r0d, bypass_0r1d, bypass_0a, c112_r, c112_a, c109_r, c109_a0d, c109_a1d);
  BrzDecisionWait_1 I29 (c113_r, c113_a, c112_r, c112_a, c111_r, c111_a);
  BrzLoop I30 (c114_r, c114_a, c113_r, c113_a);
  BrzWireFork_13 I31 (activate_0r, activate_0a, c114_r, c114_a, c108_r, c108_a, c102_r, c102_a, c96_r, c96_a, c90_r, c90_a, c84_r, c84_a, c78_r, c78_a, c72_r, c72_a, c66_r, c66_a, c44_r, c44_a, c41_r, c41_a, c31_r, c31_a, c18_r, c18_a);
  BrzPassivatorPush_1_1 I32 (c49_r, c49_a0d, c49_a1d, c67_r0d, c67_r1d, c67_a);
  BrzPassivatorPush_32_1 I33 (c50_r, c50_a0d[31:0], c50_a1d[31:0], c68_r0d[31:0], c68_r1d[31:0], c68_a);
  BrzPassivatorPush_1_1 I34 (c69_r, c69_a0d, c69_a1d, c51_r0d, c51_r1d, c51_a);
  BrzPassivatorPush_32_1 I35 (c70_r, c70_a0d[31:0], c70_a1d[31:0], c52_r0d[31:0], c52_r1d[31:0], c52_a);
  BrzPassivatorPush_32_1 I36 (c71_r, c71_a0d[31:0], c71_a1d[31:0], c53_r0d[31:0], c53_r1d[31:0], c53_a);
  BrzPassivatorPush_35_1 I37 (c64_r, c64_a0d[34:0], c64_a1d[34:0], c73_r0d[34:0], c73_r1d[34:0], c73_a);
  BrzPassivatorPush_35_1 I38 (c65_r, c65_a0d[34:0], c65_a1d[34:0], c74_r0d[34:0], c74_r1d[34:0], c74_a);
  BrzPassivatorPush_35_1 I39 (c75_r, c75_a0d[34:0], c75_a1d[34:0], c54_r0d[34:0], c54_r1d[34:0], c54_a);
  BrzPassivatorPush_35_1 I40 (c76_r, c76_a0d[34:0], c76_a1d[34:0], c55_r0d[34:0], c55_r1d[34:0], c55_a);
  BrzPassivatorPush_35_1 I41 (c77_r, c77_a0d[34:0], c77_a1d[34:0], c56_r0d[34:0], c56_r1d[34:0], c56_a);
  BrzPassivatorPush_1_1 I42 (c57_r, c57_a0d, c57_a1d, c42_r0d, c42_r1d, c42_a);
  BrzPassivatorPush_1_1 I43 (c43_r, c43_a0d, c43_a1d, c58_r0d, c58_r1d, c58_a);
  BrzPassivatorPush_1_1 I44 (c59_r, c59_a0d, c59_a1d, c32_r0d, c32_r1d, c32_a);
  BrzPassivatorPush_1_1 I45 (c60_r, c60_a0d, c60_a1d, c33_r0d, c33_r1d, c33_a);
  BrzPassivatorPush_35_1 I46 (c61_r, c61_a0d[34:0], c61_a1d[34:0], c34_r0d[34:0], c34_r1d[34:0], c34_a);
  BrzPassivatorPush_36_1 I47 (c62_r, c62_a0d[35:0], c62_a1d[35:0], c35_r0d[35:0], c35_r1d[35:0], c35_a);
  BrzPassivatorPush_35_1 I48 (c63_r, c63_a0d[34:0], c63_a1d[34:0], c36_r0d[34:0], c36_r1d[34:0], c36_a);
  BrzPassivatorPush_32_1 I49 (c26_r, c26_a0d[31:0], c26_a1d[31:0], c80_r0d[31:0], c80_r1d[31:0], c80_a);
  BrzPassivatorPush_32_1 I50 (c27_r, c27_a0d[31:0], c27_a1d[31:0], c86_r0d[31:0], c86_r1d[31:0], c86_a);
  BrzPassivatorPush_32_1 I51 (c28_r, c28_a0d[31:0], c28_a1d[31:0], c92_r0d[31:0], c92_r1d[31:0], c92_a);
  BrzPassivatorPush_3_1 I52 (c25_r, c25_a0d[2:0], c25_a1d[2:0], c98_r0d[2:0], c98_r1d[2:0], c98_a);
  BrzPassivatorPush_1_1 I53 (c29_r, c29_a0d, c29_a1d, c104_r0d, c104_r1d, c104_a);
  BrzPassivatorPush_1_1 I54 (c30_r, c30_a0d, c30_a1d, c110_r0d, c110_r1d, c110_a);
  BrzPassivatorPush_3_1 I55 (c40_r, c40_a0d[2:0], c40_a1d[2:0], c21_r0d[2:0], c21_r1d[2:0], c21_a);
  BrzPassivatorPush_32_1 I56 (c37_r, c37_a0d[31:0], c37_a1d[31:0], c22_r0d[31:0], c22_r1d[31:0], c22_a);
  BrzPassivatorPush_32_1 I57 (c38_r, c38_a0d[31:0], c38_a1d[31:0], c23_r0d[31:0], c23_r1d[31:0], c23_a);
  BrzPassivatorPush_32_1 I58 (c39_r, c39_a0d[31:0], c39_a1d[31:0], c24_r0d[31:0], c24_r1d[31:0], c24_a);
  BrzPassivatorPush_1_1 I59 (c16_r, c16_a0d, c16_a1d, c19_r0d, c19_r1d, c19_a);
  BrzPassivatorPush_1_1 I60 (c17_r, c17_a0d, c17_a1d, c20_r0d, c20_r1d, c20_a);
  BrzPassivatorPush_1_1 I61 (c12_r, c12_a0d, c12_a1d, c45_r0d, c45_r1d, c45_a);
  BrzPassivatorPush_1_1 I62 (c13_r, c13_a0d, c13_a1d, c46_r0d, c46_r1d, c46_a);
  BrzPassivatorPush_32_1 I63 (c14_r, c14_a0d[31:0], c14_a1d[31:0], c47_r0d[31:0], c47_r1d[31:0], c47_a);
  BrzPassivatorPush_32_1 I64 (c15_r, c15_a0d[31:0], c15_a1d[31:0], c48_r0d[31:0], c48_r1d[31:0], c48_a);
endmodule

module Balsa_nmult (
  activate_0r, activate_0a,
  bypass_0r0d, bypass_0r1d, bypass_0a,
  bypassH_0r0d, bypassH_0r1d, bypassH_0a,
  mType_0r0d, mType_0r1d, mType_0a,
  a_0r0d, a_0r1d, a_0a,
  b_0r0d, b_0r1d, b_0a,
  c_0r0d, c_0r1d, c_0a,
  mpH_0r0d, mpH_0r1d, mpH_0a,
  mpL_0r0d, mpL_0r1d, mpL_0a,
  mZ_0r0d, mZ_0r1d, mZ_0a,
  mN_0r0d, mN_0r1d, mN_0a
);
  input activate_0r;
  output activate_0a;
  input bypass_0r0d;
  input bypass_0r1d;
  output bypass_0a;
  input bypassH_0r0d;
  input bypassH_0r1d;
  output bypassH_0a;
  input [2:0] mType_0r0d;
  input [2:0] mType_0r1d;
  output mType_0a;
  input [31:0] a_0r0d;
  input [31:0] a_0r1d;
  output a_0a;
  input [31:0] b_0r0d;
  input [31:0] b_0r1d;
  output b_0a;
  input [31:0] c_0r0d;
  input [31:0] c_0r1d;
  output c_0a;
  output [31:0] mpH_0r0d;
  output [31:0] mpH_0r1d;
  input mpH_0a;
  output [31:0] mpL_0r0d;
  output [31:0] mpL_0r1d;
  input mpL_0a;
  output mZ_0r0d;
  output mZ_0r1d;
  input mZ_0a;
  output mN_0r0d;
  output mN_0r1d;
  input mN_0a;
  Balsa_nanoSpaMultiplier I0 (activate_0r, activate_0a, bypass_0r0d, bypass_0r1d, bypass_0a, bypassH_0r0d, bypassH_0r1d, bypassH_0a, mType_0r0d[2:0], mType_0r1d[2:0], mType_0a, a_0r0d[31:0], a_0r1d[31:0], a_0a, b_0r0d[31:0], b_0r1d[31:0], b_0a, c_0r0d[31:0], c_0r1d[31:0], c_0a, mpH_0r0d[31:0], mpH_0r1d[31:0], mpH_0a, mpL_0r0d[31:0], mpL_0r1d[31:0], mpL_0a, mZ_0r0d, mZ_0r1d, mZ_0a, mN_0r0d, mN_0r1d, mN_0a);
endmodule

