//
// by teak gui
//
// Generated on: Wed Aug 15 16:03:48 BST 2012
//


`timescale 1ns/1ps

// tkj66m1_32_1_32 TeakJ [Many [1,32,1,32],One 66]
module tkj66m1_32_1_32 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  input i_2r0;
  input i_2r1;
  output i_2a;
  input [31:0] i_3r0;
  input [31:0] i_3r1;
  output i_3a;
  output [65:0] o_0r0;
  output [65:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r0);
  BUFF I1 (o_0r0[1:1], i_1r0[0:0]);
  BUFF I2 (o_0r0[2:2], i_1r0[1:1]);
  BUFF I3 (o_0r0[3:3], i_1r0[2:2]);
  BUFF I4 (o_0r0[4:4], i_1r0[3:3]);
  BUFF I5 (o_0r0[5:5], i_1r0[4:4]);
  BUFF I6 (o_0r0[6:6], i_1r0[5:5]);
  BUFF I7 (o_0r0[7:7], i_1r0[6:6]);
  BUFF I8 (o_0r0[8:8], i_1r0[7:7]);
  BUFF I9 (o_0r0[9:9], i_1r0[8:8]);
  BUFF I10 (o_0r0[10:10], i_1r0[9:9]);
  BUFF I11 (o_0r0[11:11], i_1r0[10:10]);
  BUFF I12 (o_0r0[12:12], i_1r0[11:11]);
  BUFF I13 (o_0r0[13:13], i_1r0[12:12]);
  BUFF I14 (o_0r0[14:14], i_1r0[13:13]);
  BUFF I15 (o_0r0[15:15], i_1r0[14:14]);
  BUFF I16 (o_0r0[16:16], i_1r0[15:15]);
  BUFF I17 (o_0r0[17:17], i_1r0[16:16]);
  BUFF I18 (o_0r0[18:18], i_1r0[17:17]);
  BUFF I19 (o_0r0[19:19], i_1r0[18:18]);
  BUFF I20 (o_0r0[20:20], i_1r0[19:19]);
  BUFF I21 (o_0r0[21:21], i_1r0[20:20]);
  BUFF I22 (o_0r0[22:22], i_1r0[21:21]);
  BUFF I23 (o_0r0[23:23], i_1r0[22:22]);
  BUFF I24 (o_0r0[24:24], i_1r0[23:23]);
  BUFF I25 (o_0r0[25:25], i_1r0[24:24]);
  BUFF I26 (o_0r0[26:26], i_1r0[25:25]);
  BUFF I27 (o_0r0[27:27], i_1r0[26:26]);
  BUFF I28 (o_0r0[28:28], i_1r0[27:27]);
  BUFF I29 (o_0r0[29:29], i_1r0[28:28]);
  BUFF I30 (o_0r0[30:30], i_1r0[29:29]);
  BUFF I31 (o_0r0[31:31], i_1r0[30:30]);
  BUFF I32 (o_0r0[32:32], i_1r0[31:31]);
  BUFF I33 (o_0r0[33:33], i_2r0);
  BUFF I34 (o_0r0[34:34], i_3r0[0:0]);
  BUFF I35 (o_0r0[35:35], i_3r0[1:1]);
  BUFF I36 (o_0r0[36:36], i_3r0[2:2]);
  BUFF I37 (o_0r0[37:37], i_3r0[3:3]);
  BUFF I38 (o_0r0[38:38], i_3r0[4:4]);
  BUFF I39 (o_0r0[39:39], i_3r0[5:5]);
  BUFF I40 (o_0r0[40:40], i_3r0[6:6]);
  BUFF I41 (o_0r0[41:41], i_3r0[7:7]);
  BUFF I42 (o_0r0[42:42], i_3r0[8:8]);
  BUFF I43 (o_0r0[43:43], i_3r0[9:9]);
  BUFF I44 (o_0r0[44:44], i_3r0[10:10]);
  BUFF I45 (o_0r0[45:45], i_3r0[11:11]);
  BUFF I46 (o_0r0[46:46], i_3r0[12:12]);
  BUFF I47 (o_0r0[47:47], i_3r0[13:13]);
  BUFF I48 (o_0r0[48:48], i_3r0[14:14]);
  BUFF I49 (o_0r0[49:49], i_3r0[15:15]);
  BUFF I50 (o_0r0[50:50], i_3r0[16:16]);
  BUFF I51 (o_0r0[51:51], i_3r0[17:17]);
  BUFF I52 (o_0r0[52:52], i_3r0[18:18]);
  BUFF I53 (o_0r0[53:53], i_3r0[19:19]);
  BUFF I54 (o_0r0[54:54], i_3r0[20:20]);
  BUFF I55 (o_0r0[55:55], i_3r0[21:21]);
  BUFF I56 (o_0r0[56:56], i_3r0[22:22]);
  BUFF I57 (o_0r0[57:57], i_3r0[23:23]);
  BUFF I58 (o_0r0[58:58], i_3r0[24:24]);
  BUFF I59 (o_0r0[59:59], i_3r0[25:25]);
  BUFF I60 (o_0r0[60:60], i_3r0[26:26]);
  BUFF I61 (o_0r0[61:61], i_3r0[27:27]);
  BUFF I62 (o_0r0[62:62], i_3r0[28:28]);
  BUFF I63 (o_0r0[63:63], i_3r0[29:29]);
  BUFF I64 (o_0r0[64:64], i_3r0[30:30]);
  BUFF I65 (o_0r0[65:65], i_3r0[31:31]);
  BUFF I66 (o_0r1[0:0], i_0r1);
  BUFF I67 (o_0r1[1:1], i_1r1[0:0]);
  BUFF I68 (o_0r1[2:2], i_1r1[1:1]);
  BUFF I69 (o_0r1[3:3], i_1r1[2:2]);
  BUFF I70 (o_0r1[4:4], i_1r1[3:3]);
  BUFF I71 (o_0r1[5:5], i_1r1[4:4]);
  BUFF I72 (o_0r1[6:6], i_1r1[5:5]);
  BUFF I73 (o_0r1[7:7], i_1r1[6:6]);
  BUFF I74 (o_0r1[8:8], i_1r1[7:7]);
  BUFF I75 (o_0r1[9:9], i_1r1[8:8]);
  BUFF I76 (o_0r1[10:10], i_1r1[9:9]);
  BUFF I77 (o_0r1[11:11], i_1r1[10:10]);
  BUFF I78 (o_0r1[12:12], i_1r1[11:11]);
  BUFF I79 (o_0r1[13:13], i_1r1[12:12]);
  BUFF I80 (o_0r1[14:14], i_1r1[13:13]);
  BUFF I81 (o_0r1[15:15], i_1r1[14:14]);
  BUFF I82 (o_0r1[16:16], i_1r1[15:15]);
  BUFF I83 (o_0r1[17:17], i_1r1[16:16]);
  BUFF I84 (o_0r1[18:18], i_1r1[17:17]);
  BUFF I85 (o_0r1[19:19], i_1r1[18:18]);
  BUFF I86 (o_0r1[20:20], i_1r1[19:19]);
  BUFF I87 (o_0r1[21:21], i_1r1[20:20]);
  BUFF I88 (o_0r1[22:22], i_1r1[21:21]);
  BUFF I89 (o_0r1[23:23], i_1r1[22:22]);
  BUFF I90 (o_0r1[24:24], i_1r1[23:23]);
  BUFF I91 (o_0r1[25:25], i_1r1[24:24]);
  BUFF I92 (o_0r1[26:26], i_1r1[25:25]);
  BUFF I93 (o_0r1[27:27], i_1r1[26:26]);
  BUFF I94 (o_0r1[28:28], i_1r1[27:27]);
  BUFF I95 (o_0r1[29:29], i_1r1[28:28]);
  BUFF I96 (o_0r1[30:30], i_1r1[29:29]);
  BUFF I97 (o_0r1[31:31], i_1r1[30:30]);
  BUFF I98 (o_0r1[32:32], i_1r1[31:31]);
  BUFF I99 (o_0r1[33:33], i_2r1);
  BUFF I100 (o_0r1[34:34], i_3r1[0:0]);
  BUFF I101 (o_0r1[35:35], i_3r1[1:1]);
  BUFF I102 (o_0r1[36:36], i_3r1[2:2]);
  BUFF I103 (o_0r1[37:37], i_3r1[3:3]);
  BUFF I104 (o_0r1[38:38], i_3r1[4:4]);
  BUFF I105 (o_0r1[39:39], i_3r1[5:5]);
  BUFF I106 (o_0r1[40:40], i_3r1[6:6]);
  BUFF I107 (o_0r1[41:41], i_3r1[7:7]);
  BUFF I108 (o_0r1[42:42], i_3r1[8:8]);
  BUFF I109 (o_0r1[43:43], i_3r1[9:9]);
  BUFF I110 (o_0r1[44:44], i_3r1[10:10]);
  BUFF I111 (o_0r1[45:45], i_3r1[11:11]);
  BUFF I112 (o_0r1[46:46], i_3r1[12:12]);
  BUFF I113 (o_0r1[47:47], i_3r1[13:13]);
  BUFF I114 (o_0r1[48:48], i_3r1[14:14]);
  BUFF I115 (o_0r1[49:49], i_3r1[15:15]);
  BUFF I116 (o_0r1[50:50], i_3r1[16:16]);
  BUFF I117 (o_0r1[51:51], i_3r1[17:17]);
  BUFF I118 (o_0r1[52:52], i_3r1[18:18]);
  BUFF I119 (o_0r1[53:53], i_3r1[19:19]);
  BUFF I120 (o_0r1[54:54], i_3r1[20:20]);
  BUFF I121 (o_0r1[55:55], i_3r1[21:21]);
  BUFF I122 (o_0r1[56:56], i_3r1[22:22]);
  BUFF I123 (o_0r1[57:57], i_3r1[23:23]);
  BUFF I124 (o_0r1[58:58], i_3r1[24:24]);
  BUFF I125 (o_0r1[59:59], i_3r1[25:25]);
  BUFF I126 (o_0r1[60:60], i_3r1[26:26]);
  BUFF I127 (o_0r1[61:61], i_3r1[27:27]);
  BUFF I128 (o_0r1[62:62], i_3r1[28:28]);
  BUFF I129 (o_0r1[63:63], i_3r1[29:29]);
  BUFF I130 (o_0r1[64:64], i_3r1[30:30]);
  BUFF I131 (o_0r1[65:65], i_3r1[31:31]);
  BUFF I132 (i_0a, o_0a);
  BUFF I133 (i_1a, o_0a);
  BUFF I134 (i_2a, o_0a);
  BUFF I135 (i_3a, o_0a);
endmodule

// tkf0mo0w0_o0w0_o0w0_o0w0 TeakF [0,0,0,0] [One 0,Many [0,0,0,0]]
module tkf0mo0w0_o0w0_o0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  input reset;
  wire [1:0] simp11_0;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  BUFF I2 (o_2r, i_0r);
  BUFF I3 (o_3r, i_0r);
  C3 I4 (simp11_0[0:0], o_0a, o_1a, o_2a);
  BUFF I5 (simp11_0[1:1], o_3a);
  C2 I6 (i_0a, simp11_0[0:0], simp11_0[1:1]);
endmodule

// tkj33m32_1 TeakJ [Many [32,1],One 33]
module tkj33m32_1 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input i_1r0;
  input i_1r1;
  output i_1a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r0[0:0]);
  BUFF I1 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I2 (o_0r0[2:2], i_0r0[2:2]);
  BUFF I3 (o_0r0[3:3], i_0r0[3:3]);
  BUFF I4 (o_0r0[4:4], i_0r0[4:4]);
  BUFF I5 (o_0r0[5:5], i_0r0[5:5]);
  BUFF I6 (o_0r0[6:6], i_0r0[6:6]);
  BUFF I7 (o_0r0[7:7], i_0r0[7:7]);
  BUFF I8 (o_0r0[8:8], i_0r0[8:8]);
  BUFF I9 (o_0r0[9:9], i_0r0[9:9]);
  BUFF I10 (o_0r0[10:10], i_0r0[10:10]);
  BUFF I11 (o_0r0[11:11], i_0r0[11:11]);
  BUFF I12 (o_0r0[12:12], i_0r0[12:12]);
  BUFF I13 (o_0r0[13:13], i_0r0[13:13]);
  BUFF I14 (o_0r0[14:14], i_0r0[14:14]);
  BUFF I15 (o_0r0[15:15], i_0r0[15:15]);
  BUFF I16 (o_0r0[16:16], i_0r0[16:16]);
  BUFF I17 (o_0r0[17:17], i_0r0[17:17]);
  BUFF I18 (o_0r0[18:18], i_0r0[18:18]);
  BUFF I19 (o_0r0[19:19], i_0r0[19:19]);
  BUFF I20 (o_0r0[20:20], i_0r0[20:20]);
  BUFF I21 (o_0r0[21:21], i_0r0[21:21]);
  BUFF I22 (o_0r0[22:22], i_0r0[22:22]);
  BUFF I23 (o_0r0[23:23], i_0r0[23:23]);
  BUFF I24 (o_0r0[24:24], i_0r0[24:24]);
  BUFF I25 (o_0r0[25:25], i_0r0[25:25]);
  BUFF I26 (o_0r0[26:26], i_0r0[26:26]);
  BUFF I27 (o_0r0[27:27], i_0r0[27:27]);
  BUFF I28 (o_0r0[28:28], i_0r0[28:28]);
  BUFF I29 (o_0r0[29:29], i_0r0[29:29]);
  BUFF I30 (o_0r0[30:30], i_0r0[30:30]);
  BUFF I31 (o_0r0[31:31], i_0r0[31:31]);
  BUFF I32 (o_0r0[32:32], i_1r0);
  BUFF I33 (o_0r1[0:0], i_0r1[0:0]);
  BUFF I34 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I35 (o_0r1[2:2], i_0r1[2:2]);
  BUFF I36 (o_0r1[3:3], i_0r1[3:3]);
  BUFF I37 (o_0r1[4:4], i_0r1[4:4]);
  BUFF I38 (o_0r1[5:5], i_0r1[5:5]);
  BUFF I39 (o_0r1[6:6], i_0r1[6:6]);
  BUFF I40 (o_0r1[7:7], i_0r1[7:7]);
  BUFF I41 (o_0r1[8:8], i_0r1[8:8]);
  BUFF I42 (o_0r1[9:9], i_0r1[9:9]);
  BUFF I43 (o_0r1[10:10], i_0r1[10:10]);
  BUFF I44 (o_0r1[11:11], i_0r1[11:11]);
  BUFF I45 (o_0r1[12:12], i_0r1[12:12]);
  BUFF I46 (o_0r1[13:13], i_0r1[13:13]);
  BUFF I47 (o_0r1[14:14], i_0r1[14:14]);
  BUFF I48 (o_0r1[15:15], i_0r1[15:15]);
  BUFF I49 (o_0r1[16:16], i_0r1[16:16]);
  BUFF I50 (o_0r1[17:17], i_0r1[17:17]);
  BUFF I51 (o_0r1[18:18], i_0r1[18:18]);
  BUFF I52 (o_0r1[19:19], i_0r1[19:19]);
  BUFF I53 (o_0r1[20:20], i_0r1[20:20]);
  BUFF I54 (o_0r1[21:21], i_0r1[21:21]);
  BUFF I55 (o_0r1[22:22], i_0r1[22:22]);
  BUFF I56 (o_0r1[23:23], i_0r1[23:23]);
  BUFF I57 (o_0r1[24:24], i_0r1[24:24]);
  BUFF I58 (o_0r1[25:25], i_0r1[25:25]);
  BUFF I59 (o_0r1[26:26], i_0r1[26:26]);
  BUFF I60 (o_0r1[27:27], i_0r1[27:27]);
  BUFF I61 (o_0r1[28:28], i_0r1[28:28]);
  BUFF I62 (o_0r1[29:29], i_0r1[29:29]);
  BUFF I63 (o_0r1[30:30], i_0r1[30:30]);
  BUFF I64 (o_0r1[31:31], i_0r1[31:31]);
  BUFF I65 (o_0r1[32:32], i_1r1);
  BUFF I66 (i_0a, o_0a);
  BUFF I67 (i_1a, o_0a);
endmodule

// tkf0mo0w0_o0w0 TeakF [0,0] [One 0,Many [0,0]]
module tkf0mo0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  C2 I2 (i_0a, o_0a, o_1a);
endmodule

// tko65m33_1xori0w32bi32w32b_2apt1o0w32bi64w1b TeakO [
//     (1,TeakOp TeakOpXor [(0,0,32),(0,32,32)]),
//     (2,TeakOAppend 1 [(1,0,32),(0,64,1)])] [One 65,One 33]
module tko65m33_1xori0w32bi32w32b_2apt1o0w32bi64w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [64:0] i_0r0;
  input [64:0] i_0r1;
  output i_0a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  wire [31:0] termf_1;
  wire [31:0] termt_1;
  wire [3:0] op1_0_0;
  wire [3:0] op1_1_0;
  wire [3:0] op1_2_0;
  wire [3:0] op1_3_0;
  wire [3:0] op1_4_0;
  wire [3:0] op1_5_0;
  wire [3:0] op1_6_0;
  wire [3:0] op1_7_0;
  wire [3:0] op1_8_0;
  wire [3:0] op1_9_0;
  wire [3:0] op1_10_0;
  wire [3:0] op1_11_0;
  wire [3:0] op1_12_0;
  wire [3:0] op1_13_0;
  wire [3:0] op1_14_0;
  wire [3:0] op1_15_0;
  wire [3:0] op1_16_0;
  wire [3:0] op1_17_0;
  wire [3:0] op1_18_0;
  wire [3:0] op1_19_0;
  wire [3:0] op1_20_0;
  wire [3:0] op1_21_0;
  wire [3:0] op1_22_0;
  wire [3:0] op1_23_0;
  wire [3:0] op1_24_0;
  wire [3:0] op1_25_0;
  wire [3:0] op1_26_0;
  wire [3:0] op1_27_0;
  wire [3:0] op1_28_0;
  wire [3:0] op1_29_0;
  wire [3:0] op1_30_0;
  wire [3:0] op1_31_0;
  C2 I0 (op1_0_0[0:0], i_0r0[32:32], i_0r0[0:0]);
  C2 I1 (op1_0_0[1:1], i_0r0[32:32], i_0r1[0:0]);
  C2 I2 (op1_0_0[2:2], i_0r1[32:32], i_0r0[0:0]);
  C2 I3 (op1_0_0[3:3], i_0r1[32:32], i_0r1[0:0]);
  OR2 I4 (termf_1[0:0], op1_0_0[0:0], op1_0_0[3:3]);
  OR2 I5 (termt_1[0:0], op1_0_0[1:1], op1_0_0[2:2]);
  C2 I6 (op1_1_0[0:0], i_0r0[33:33], i_0r0[1:1]);
  C2 I7 (op1_1_0[1:1], i_0r0[33:33], i_0r1[1:1]);
  C2 I8 (op1_1_0[2:2], i_0r1[33:33], i_0r0[1:1]);
  C2 I9 (op1_1_0[3:3], i_0r1[33:33], i_0r1[1:1]);
  OR2 I10 (termf_1[1:1], op1_1_0[0:0], op1_1_0[3:3]);
  OR2 I11 (termt_1[1:1], op1_1_0[1:1], op1_1_0[2:2]);
  C2 I12 (op1_2_0[0:0], i_0r0[34:34], i_0r0[2:2]);
  C2 I13 (op1_2_0[1:1], i_0r0[34:34], i_0r1[2:2]);
  C2 I14 (op1_2_0[2:2], i_0r1[34:34], i_0r0[2:2]);
  C2 I15 (op1_2_0[3:3], i_0r1[34:34], i_0r1[2:2]);
  OR2 I16 (termf_1[2:2], op1_2_0[0:0], op1_2_0[3:3]);
  OR2 I17 (termt_1[2:2], op1_2_0[1:1], op1_2_0[2:2]);
  C2 I18 (op1_3_0[0:0], i_0r0[35:35], i_0r0[3:3]);
  C2 I19 (op1_3_0[1:1], i_0r0[35:35], i_0r1[3:3]);
  C2 I20 (op1_3_0[2:2], i_0r1[35:35], i_0r0[3:3]);
  C2 I21 (op1_3_0[3:3], i_0r1[35:35], i_0r1[3:3]);
  OR2 I22 (termf_1[3:3], op1_3_0[0:0], op1_3_0[3:3]);
  OR2 I23 (termt_1[3:3], op1_3_0[1:1], op1_3_0[2:2]);
  C2 I24 (op1_4_0[0:0], i_0r0[36:36], i_0r0[4:4]);
  C2 I25 (op1_4_0[1:1], i_0r0[36:36], i_0r1[4:4]);
  C2 I26 (op1_4_0[2:2], i_0r1[36:36], i_0r0[4:4]);
  C2 I27 (op1_4_0[3:3], i_0r1[36:36], i_0r1[4:4]);
  OR2 I28 (termf_1[4:4], op1_4_0[0:0], op1_4_0[3:3]);
  OR2 I29 (termt_1[4:4], op1_4_0[1:1], op1_4_0[2:2]);
  C2 I30 (op1_5_0[0:0], i_0r0[37:37], i_0r0[5:5]);
  C2 I31 (op1_5_0[1:1], i_0r0[37:37], i_0r1[5:5]);
  C2 I32 (op1_5_0[2:2], i_0r1[37:37], i_0r0[5:5]);
  C2 I33 (op1_5_0[3:3], i_0r1[37:37], i_0r1[5:5]);
  OR2 I34 (termf_1[5:5], op1_5_0[0:0], op1_5_0[3:3]);
  OR2 I35 (termt_1[5:5], op1_5_0[1:1], op1_5_0[2:2]);
  C2 I36 (op1_6_0[0:0], i_0r0[38:38], i_0r0[6:6]);
  C2 I37 (op1_6_0[1:1], i_0r0[38:38], i_0r1[6:6]);
  C2 I38 (op1_6_0[2:2], i_0r1[38:38], i_0r0[6:6]);
  C2 I39 (op1_6_0[3:3], i_0r1[38:38], i_0r1[6:6]);
  OR2 I40 (termf_1[6:6], op1_6_0[0:0], op1_6_0[3:3]);
  OR2 I41 (termt_1[6:6], op1_6_0[1:1], op1_6_0[2:2]);
  C2 I42 (op1_7_0[0:0], i_0r0[39:39], i_0r0[7:7]);
  C2 I43 (op1_7_0[1:1], i_0r0[39:39], i_0r1[7:7]);
  C2 I44 (op1_7_0[2:2], i_0r1[39:39], i_0r0[7:7]);
  C2 I45 (op1_7_0[3:3], i_0r1[39:39], i_0r1[7:7]);
  OR2 I46 (termf_1[7:7], op1_7_0[0:0], op1_7_0[3:3]);
  OR2 I47 (termt_1[7:7], op1_7_0[1:1], op1_7_0[2:2]);
  C2 I48 (op1_8_0[0:0], i_0r0[40:40], i_0r0[8:8]);
  C2 I49 (op1_8_0[1:1], i_0r0[40:40], i_0r1[8:8]);
  C2 I50 (op1_8_0[2:2], i_0r1[40:40], i_0r0[8:8]);
  C2 I51 (op1_8_0[3:3], i_0r1[40:40], i_0r1[8:8]);
  OR2 I52 (termf_1[8:8], op1_8_0[0:0], op1_8_0[3:3]);
  OR2 I53 (termt_1[8:8], op1_8_0[1:1], op1_8_0[2:2]);
  C2 I54 (op1_9_0[0:0], i_0r0[41:41], i_0r0[9:9]);
  C2 I55 (op1_9_0[1:1], i_0r0[41:41], i_0r1[9:9]);
  C2 I56 (op1_9_0[2:2], i_0r1[41:41], i_0r0[9:9]);
  C2 I57 (op1_9_0[3:3], i_0r1[41:41], i_0r1[9:9]);
  OR2 I58 (termf_1[9:9], op1_9_0[0:0], op1_9_0[3:3]);
  OR2 I59 (termt_1[9:9], op1_9_0[1:1], op1_9_0[2:2]);
  C2 I60 (op1_10_0[0:0], i_0r0[42:42], i_0r0[10:10]);
  C2 I61 (op1_10_0[1:1], i_0r0[42:42], i_0r1[10:10]);
  C2 I62 (op1_10_0[2:2], i_0r1[42:42], i_0r0[10:10]);
  C2 I63 (op1_10_0[3:3], i_0r1[42:42], i_0r1[10:10]);
  OR2 I64 (termf_1[10:10], op1_10_0[0:0], op1_10_0[3:3]);
  OR2 I65 (termt_1[10:10], op1_10_0[1:1], op1_10_0[2:2]);
  C2 I66 (op1_11_0[0:0], i_0r0[43:43], i_0r0[11:11]);
  C2 I67 (op1_11_0[1:1], i_0r0[43:43], i_0r1[11:11]);
  C2 I68 (op1_11_0[2:2], i_0r1[43:43], i_0r0[11:11]);
  C2 I69 (op1_11_0[3:3], i_0r1[43:43], i_0r1[11:11]);
  OR2 I70 (termf_1[11:11], op1_11_0[0:0], op1_11_0[3:3]);
  OR2 I71 (termt_1[11:11], op1_11_0[1:1], op1_11_0[2:2]);
  C2 I72 (op1_12_0[0:0], i_0r0[44:44], i_0r0[12:12]);
  C2 I73 (op1_12_0[1:1], i_0r0[44:44], i_0r1[12:12]);
  C2 I74 (op1_12_0[2:2], i_0r1[44:44], i_0r0[12:12]);
  C2 I75 (op1_12_0[3:3], i_0r1[44:44], i_0r1[12:12]);
  OR2 I76 (termf_1[12:12], op1_12_0[0:0], op1_12_0[3:3]);
  OR2 I77 (termt_1[12:12], op1_12_0[1:1], op1_12_0[2:2]);
  C2 I78 (op1_13_0[0:0], i_0r0[45:45], i_0r0[13:13]);
  C2 I79 (op1_13_0[1:1], i_0r0[45:45], i_0r1[13:13]);
  C2 I80 (op1_13_0[2:2], i_0r1[45:45], i_0r0[13:13]);
  C2 I81 (op1_13_0[3:3], i_0r1[45:45], i_0r1[13:13]);
  OR2 I82 (termf_1[13:13], op1_13_0[0:0], op1_13_0[3:3]);
  OR2 I83 (termt_1[13:13], op1_13_0[1:1], op1_13_0[2:2]);
  C2 I84 (op1_14_0[0:0], i_0r0[46:46], i_0r0[14:14]);
  C2 I85 (op1_14_0[1:1], i_0r0[46:46], i_0r1[14:14]);
  C2 I86 (op1_14_0[2:2], i_0r1[46:46], i_0r0[14:14]);
  C2 I87 (op1_14_0[3:3], i_0r1[46:46], i_0r1[14:14]);
  OR2 I88 (termf_1[14:14], op1_14_0[0:0], op1_14_0[3:3]);
  OR2 I89 (termt_1[14:14], op1_14_0[1:1], op1_14_0[2:2]);
  C2 I90 (op1_15_0[0:0], i_0r0[47:47], i_0r0[15:15]);
  C2 I91 (op1_15_0[1:1], i_0r0[47:47], i_0r1[15:15]);
  C2 I92 (op1_15_0[2:2], i_0r1[47:47], i_0r0[15:15]);
  C2 I93 (op1_15_0[3:3], i_0r1[47:47], i_0r1[15:15]);
  OR2 I94 (termf_1[15:15], op1_15_0[0:0], op1_15_0[3:3]);
  OR2 I95 (termt_1[15:15], op1_15_0[1:1], op1_15_0[2:2]);
  C2 I96 (op1_16_0[0:0], i_0r0[48:48], i_0r0[16:16]);
  C2 I97 (op1_16_0[1:1], i_0r0[48:48], i_0r1[16:16]);
  C2 I98 (op1_16_0[2:2], i_0r1[48:48], i_0r0[16:16]);
  C2 I99 (op1_16_0[3:3], i_0r1[48:48], i_0r1[16:16]);
  OR2 I100 (termf_1[16:16], op1_16_0[0:0], op1_16_0[3:3]);
  OR2 I101 (termt_1[16:16], op1_16_0[1:1], op1_16_0[2:2]);
  C2 I102 (op1_17_0[0:0], i_0r0[49:49], i_0r0[17:17]);
  C2 I103 (op1_17_0[1:1], i_0r0[49:49], i_0r1[17:17]);
  C2 I104 (op1_17_0[2:2], i_0r1[49:49], i_0r0[17:17]);
  C2 I105 (op1_17_0[3:3], i_0r1[49:49], i_0r1[17:17]);
  OR2 I106 (termf_1[17:17], op1_17_0[0:0], op1_17_0[3:3]);
  OR2 I107 (termt_1[17:17], op1_17_0[1:1], op1_17_0[2:2]);
  C2 I108 (op1_18_0[0:0], i_0r0[50:50], i_0r0[18:18]);
  C2 I109 (op1_18_0[1:1], i_0r0[50:50], i_0r1[18:18]);
  C2 I110 (op1_18_0[2:2], i_0r1[50:50], i_0r0[18:18]);
  C2 I111 (op1_18_0[3:3], i_0r1[50:50], i_0r1[18:18]);
  OR2 I112 (termf_1[18:18], op1_18_0[0:0], op1_18_0[3:3]);
  OR2 I113 (termt_1[18:18], op1_18_0[1:1], op1_18_0[2:2]);
  C2 I114 (op1_19_0[0:0], i_0r0[51:51], i_0r0[19:19]);
  C2 I115 (op1_19_0[1:1], i_0r0[51:51], i_0r1[19:19]);
  C2 I116 (op1_19_0[2:2], i_0r1[51:51], i_0r0[19:19]);
  C2 I117 (op1_19_0[3:3], i_0r1[51:51], i_0r1[19:19]);
  OR2 I118 (termf_1[19:19], op1_19_0[0:0], op1_19_0[3:3]);
  OR2 I119 (termt_1[19:19], op1_19_0[1:1], op1_19_0[2:2]);
  C2 I120 (op1_20_0[0:0], i_0r0[52:52], i_0r0[20:20]);
  C2 I121 (op1_20_0[1:1], i_0r0[52:52], i_0r1[20:20]);
  C2 I122 (op1_20_0[2:2], i_0r1[52:52], i_0r0[20:20]);
  C2 I123 (op1_20_0[3:3], i_0r1[52:52], i_0r1[20:20]);
  OR2 I124 (termf_1[20:20], op1_20_0[0:0], op1_20_0[3:3]);
  OR2 I125 (termt_1[20:20], op1_20_0[1:1], op1_20_0[2:2]);
  C2 I126 (op1_21_0[0:0], i_0r0[53:53], i_0r0[21:21]);
  C2 I127 (op1_21_0[1:1], i_0r0[53:53], i_0r1[21:21]);
  C2 I128 (op1_21_0[2:2], i_0r1[53:53], i_0r0[21:21]);
  C2 I129 (op1_21_0[3:3], i_0r1[53:53], i_0r1[21:21]);
  OR2 I130 (termf_1[21:21], op1_21_0[0:0], op1_21_0[3:3]);
  OR2 I131 (termt_1[21:21], op1_21_0[1:1], op1_21_0[2:2]);
  C2 I132 (op1_22_0[0:0], i_0r0[54:54], i_0r0[22:22]);
  C2 I133 (op1_22_0[1:1], i_0r0[54:54], i_0r1[22:22]);
  C2 I134 (op1_22_0[2:2], i_0r1[54:54], i_0r0[22:22]);
  C2 I135 (op1_22_0[3:3], i_0r1[54:54], i_0r1[22:22]);
  OR2 I136 (termf_1[22:22], op1_22_0[0:0], op1_22_0[3:3]);
  OR2 I137 (termt_1[22:22], op1_22_0[1:1], op1_22_0[2:2]);
  C2 I138 (op1_23_0[0:0], i_0r0[55:55], i_0r0[23:23]);
  C2 I139 (op1_23_0[1:1], i_0r0[55:55], i_0r1[23:23]);
  C2 I140 (op1_23_0[2:2], i_0r1[55:55], i_0r0[23:23]);
  C2 I141 (op1_23_0[3:3], i_0r1[55:55], i_0r1[23:23]);
  OR2 I142 (termf_1[23:23], op1_23_0[0:0], op1_23_0[3:3]);
  OR2 I143 (termt_1[23:23], op1_23_0[1:1], op1_23_0[2:2]);
  C2 I144 (op1_24_0[0:0], i_0r0[56:56], i_0r0[24:24]);
  C2 I145 (op1_24_0[1:1], i_0r0[56:56], i_0r1[24:24]);
  C2 I146 (op1_24_0[2:2], i_0r1[56:56], i_0r0[24:24]);
  C2 I147 (op1_24_0[3:3], i_0r1[56:56], i_0r1[24:24]);
  OR2 I148 (termf_1[24:24], op1_24_0[0:0], op1_24_0[3:3]);
  OR2 I149 (termt_1[24:24], op1_24_0[1:1], op1_24_0[2:2]);
  C2 I150 (op1_25_0[0:0], i_0r0[57:57], i_0r0[25:25]);
  C2 I151 (op1_25_0[1:1], i_0r0[57:57], i_0r1[25:25]);
  C2 I152 (op1_25_0[2:2], i_0r1[57:57], i_0r0[25:25]);
  C2 I153 (op1_25_0[3:3], i_0r1[57:57], i_0r1[25:25]);
  OR2 I154 (termf_1[25:25], op1_25_0[0:0], op1_25_0[3:3]);
  OR2 I155 (termt_1[25:25], op1_25_0[1:1], op1_25_0[2:2]);
  C2 I156 (op1_26_0[0:0], i_0r0[58:58], i_0r0[26:26]);
  C2 I157 (op1_26_0[1:1], i_0r0[58:58], i_0r1[26:26]);
  C2 I158 (op1_26_0[2:2], i_0r1[58:58], i_0r0[26:26]);
  C2 I159 (op1_26_0[3:3], i_0r1[58:58], i_0r1[26:26]);
  OR2 I160 (termf_1[26:26], op1_26_0[0:0], op1_26_0[3:3]);
  OR2 I161 (termt_1[26:26], op1_26_0[1:1], op1_26_0[2:2]);
  C2 I162 (op1_27_0[0:0], i_0r0[59:59], i_0r0[27:27]);
  C2 I163 (op1_27_0[1:1], i_0r0[59:59], i_0r1[27:27]);
  C2 I164 (op1_27_0[2:2], i_0r1[59:59], i_0r0[27:27]);
  C2 I165 (op1_27_0[3:3], i_0r1[59:59], i_0r1[27:27]);
  OR2 I166 (termf_1[27:27], op1_27_0[0:0], op1_27_0[3:3]);
  OR2 I167 (termt_1[27:27], op1_27_0[1:1], op1_27_0[2:2]);
  C2 I168 (op1_28_0[0:0], i_0r0[60:60], i_0r0[28:28]);
  C2 I169 (op1_28_0[1:1], i_0r0[60:60], i_0r1[28:28]);
  C2 I170 (op1_28_0[2:2], i_0r1[60:60], i_0r0[28:28]);
  C2 I171 (op1_28_0[3:3], i_0r1[60:60], i_0r1[28:28]);
  OR2 I172 (termf_1[28:28], op1_28_0[0:0], op1_28_0[3:3]);
  OR2 I173 (termt_1[28:28], op1_28_0[1:1], op1_28_0[2:2]);
  C2 I174 (op1_29_0[0:0], i_0r0[61:61], i_0r0[29:29]);
  C2 I175 (op1_29_0[1:1], i_0r0[61:61], i_0r1[29:29]);
  C2 I176 (op1_29_0[2:2], i_0r1[61:61], i_0r0[29:29]);
  C2 I177 (op1_29_0[3:3], i_0r1[61:61], i_0r1[29:29]);
  OR2 I178 (termf_1[29:29], op1_29_0[0:0], op1_29_0[3:3]);
  OR2 I179 (termt_1[29:29], op1_29_0[1:1], op1_29_0[2:2]);
  C2 I180 (op1_30_0[0:0], i_0r0[62:62], i_0r0[30:30]);
  C2 I181 (op1_30_0[1:1], i_0r0[62:62], i_0r1[30:30]);
  C2 I182 (op1_30_0[2:2], i_0r1[62:62], i_0r0[30:30]);
  C2 I183 (op1_30_0[3:3], i_0r1[62:62], i_0r1[30:30]);
  OR2 I184 (termf_1[30:30], op1_30_0[0:0], op1_30_0[3:3]);
  OR2 I185 (termt_1[30:30], op1_30_0[1:1], op1_30_0[2:2]);
  C2 I186 (op1_31_0[0:0], i_0r0[63:63], i_0r0[31:31]);
  C2 I187 (op1_31_0[1:1], i_0r0[63:63], i_0r1[31:31]);
  C2 I188 (op1_31_0[2:2], i_0r1[63:63], i_0r0[31:31]);
  C2 I189 (op1_31_0[3:3], i_0r1[63:63], i_0r1[31:31]);
  OR2 I190 (termf_1[31:31], op1_31_0[0:0], op1_31_0[3:3]);
  OR2 I191 (termt_1[31:31], op1_31_0[1:1], op1_31_0[2:2]);
  BUFF I192 (o_0r0[0:0], termf_1[0:0]);
  BUFF I193 (o_0r0[1:1], termf_1[1:1]);
  BUFF I194 (o_0r0[2:2], termf_1[2:2]);
  BUFF I195 (o_0r0[3:3], termf_1[3:3]);
  BUFF I196 (o_0r0[4:4], termf_1[4:4]);
  BUFF I197 (o_0r0[5:5], termf_1[5:5]);
  BUFF I198 (o_0r0[6:6], termf_1[6:6]);
  BUFF I199 (o_0r0[7:7], termf_1[7:7]);
  BUFF I200 (o_0r0[8:8], termf_1[8:8]);
  BUFF I201 (o_0r0[9:9], termf_1[9:9]);
  BUFF I202 (o_0r0[10:10], termf_1[10:10]);
  BUFF I203 (o_0r0[11:11], termf_1[11:11]);
  BUFF I204 (o_0r0[12:12], termf_1[12:12]);
  BUFF I205 (o_0r0[13:13], termf_1[13:13]);
  BUFF I206 (o_0r0[14:14], termf_1[14:14]);
  BUFF I207 (o_0r0[15:15], termf_1[15:15]);
  BUFF I208 (o_0r0[16:16], termf_1[16:16]);
  BUFF I209 (o_0r0[17:17], termf_1[17:17]);
  BUFF I210 (o_0r0[18:18], termf_1[18:18]);
  BUFF I211 (o_0r0[19:19], termf_1[19:19]);
  BUFF I212 (o_0r0[20:20], termf_1[20:20]);
  BUFF I213 (o_0r0[21:21], termf_1[21:21]);
  BUFF I214 (o_0r0[22:22], termf_1[22:22]);
  BUFF I215 (o_0r0[23:23], termf_1[23:23]);
  BUFF I216 (o_0r0[24:24], termf_1[24:24]);
  BUFF I217 (o_0r0[25:25], termf_1[25:25]);
  BUFF I218 (o_0r0[26:26], termf_1[26:26]);
  BUFF I219 (o_0r0[27:27], termf_1[27:27]);
  BUFF I220 (o_0r0[28:28], termf_1[28:28]);
  BUFF I221 (o_0r0[29:29], termf_1[29:29]);
  BUFF I222 (o_0r0[30:30], termf_1[30:30]);
  BUFF I223 (o_0r0[31:31], termf_1[31:31]);
  BUFF I224 (o_0r0[32:32], i_0r0[64:64]);
  BUFF I225 (o_0r1[0:0], termt_1[0:0]);
  BUFF I226 (o_0r1[1:1], termt_1[1:1]);
  BUFF I227 (o_0r1[2:2], termt_1[2:2]);
  BUFF I228 (o_0r1[3:3], termt_1[3:3]);
  BUFF I229 (o_0r1[4:4], termt_1[4:4]);
  BUFF I230 (o_0r1[5:5], termt_1[5:5]);
  BUFF I231 (o_0r1[6:6], termt_1[6:6]);
  BUFF I232 (o_0r1[7:7], termt_1[7:7]);
  BUFF I233 (o_0r1[8:8], termt_1[8:8]);
  BUFF I234 (o_0r1[9:9], termt_1[9:9]);
  BUFF I235 (o_0r1[10:10], termt_1[10:10]);
  BUFF I236 (o_0r1[11:11], termt_1[11:11]);
  BUFF I237 (o_0r1[12:12], termt_1[12:12]);
  BUFF I238 (o_0r1[13:13], termt_1[13:13]);
  BUFF I239 (o_0r1[14:14], termt_1[14:14]);
  BUFF I240 (o_0r1[15:15], termt_1[15:15]);
  BUFF I241 (o_0r1[16:16], termt_1[16:16]);
  BUFF I242 (o_0r1[17:17], termt_1[17:17]);
  BUFF I243 (o_0r1[18:18], termt_1[18:18]);
  BUFF I244 (o_0r1[19:19], termt_1[19:19]);
  BUFF I245 (o_0r1[20:20], termt_1[20:20]);
  BUFF I246 (o_0r1[21:21], termt_1[21:21]);
  BUFF I247 (o_0r1[22:22], termt_1[22:22]);
  BUFF I248 (o_0r1[23:23], termt_1[23:23]);
  BUFF I249 (o_0r1[24:24], termt_1[24:24]);
  BUFF I250 (o_0r1[25:25], termt_1[25:25]);
  BUFF I251 (o_0r1[26:26], termt_1[26:26]);
  BUFF I252 (o_0r1[27:27], termt_1[27:27]);
  BUFF I253 (o_0r1[28:28], termt_1[28:28]);
  BUFF I254 (o_0r1[29:29], termt_1[29:29]);
  BUFF I255 (o_0r1[30:30], termt_1[30:30]);
  BUFF I256 (o_0r1[31:31], termt_1[31:31]);
  BUFF I257 (o_0r1[32:32], i_0r1[64:64]);
  BUFF I258 (i_0a, o_0a);
endmodule

// tkf0mo0w0_o0w0_o0w0 TeakF [0,0,0] [One 0,Many [0,0,0]]
module tkf0mo0w0_o0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  input reset;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  BUFF I2 (o_2r, i_0r);
  C3 I3 (i_0a, o_0a, o_1a, o_2a);
endmodule

// tko65m33_1ori0w32bi32w32b_2apt1o0w32bi64w1b TeakO [
//     (1,TeakOp TeakOpOr [(0,0,32),(0,32,32)]),
//     (2,TeakOAppend 1 [(1,0,32),(0,64,1)])] [One 65,One 33]
module tko65m33_1ori0w32bi32w32b_2apt1o0w32bi64w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [64:0] i_0r0;
  input [64:0] i_0r1;
  output i_0a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  wire [31:0] termf_1;
  wire [31:0] termt_1;
  wire [3:0] op1_0_0;
  wire [3:0] op1_1_0;
  wire [3:0] op1_2_0;
  wire [3:0] op1_3_0;
  wire [3:0] op1_4_0;
  wire [3:0] op1_5_0;
  wire [3:0] op1_6_0;
  wire [3:0] op1_7_0;
  wire [3:0] op1_8_0;
  wire [3:0] op1_9_0;
  wire [3:0] op1_10_0;
  wire [3:0] op1_11_0;
  wire [3:0] op1_12_0;
  wire [3:0] op1_13_0;
  wire [3:0] op1_14_0;
  wire [3:0] op1_15_0;
  wire [3:0] op1_16_0;
  wire [3:0] op1_17_0;
  wire [3:0] op1_18_0;
  wire [3:0] op1_19_0;
  wire [3:0] op1_20_0;
  wire [3:0] op1_21_0;
  wire [3:0] op1_22_0;
  wire [3:0] op1_23_0;
  wire [3:0] op1_24_0;
  wire [3:0] op1_25_0;
  wire [3:0] op1_26_0;
  wire [3:0] op1_27_0;
  wire [3:0] op1_28_0;
  wire [3:0] op1_29_0;
  wire [3:0] op1_30_0;
  wire [3:0] op1_31_0;
  C2 I0 (op1_0_0[0:0], i_0r0[32:32], i_0r0[0:0]);
  C2 I1 (op1_0_0[1:1], i_0r0[32:32], i_0r1[0:0]);
  C2 I2 (op1_0_0[2:2], i_0r1[32:32], i_0r0[0:0]);
  C2 I3 (op1_0_0[3:3], i_0r1[32:32], i_0r1[0:0]);
  BUFF I4 (termf_1[0:0], op1_0_0[0:0]);
  OR3 I5 (termt_1[0:0], op1_0_0[1:1], op1_0_0[2:2], op1_0_0[3:3]);
  C2 I6 (op1_1_0[0:0], i_0r0[33:33], i_0r0[1:1]);
  C2 I7 (op1_1_0[1:1], i_0r0[33:33], i_0r1[1:1]);
  C2 I8 (op1_1_0[2:2], i_0r1[33:33], i_0r0[1:1]);
  C2 I9 (op1_1_0[3:3], i_0r1[33:33], i_0r1[1:1]);
  BUFF I10 (termf_1[1:1], op1_1_0[0:0]);
  OR3 I11 (termt_1[1:1], op1_1_0[1:1], op1_1_0[2:2], op1_1_0[3:3]);
  C2 I12 (op1_2_0[0:0], i_0r0[34:34], i_0r0[2:2]);
  C2 I13 (op1_2_0[1:1], i_0r0[34:34], i_0r1[2:2]);
  C2 I14 (op1_2_0[2:2], i_0r1[34:34], i_0r0[2:2]);
  C2 I15 (op1_2_0[3:3], i_0r1[34:34], i_0r1[2:2]);
  BUFF I16 (termf_1[2:2], op1_2_0[0:0]);
  OR3 I17 (termt_1[2:2], op1_2_0[1:1], op1_2_0[2:2], op1_2_0[3:3]);
  C2 I18 (op1_3_0[0:0], i_0r0[35:35], i_0r0[3:3]);
  C2 I19 (op1_3_0[1:1], i_0r0[35:35], i_0r1[3:3]);
  C2 I20 (op1_3_0[2:2], i_0r1[35:35], i_0r0[3:3]);
  C2 I21 (op1_3_0[3:3], i_0r1[35:35], i_0r1[3:3]);
  BUFF I22 (termf_1[3:3], op1_3_0[0:0]);
  OR3 I23 (termt_1[3:3], op1_3_0[1:1], op1_3_0[2:2], op1_3_0[3:3]);
  C2 I24 (op1_4_0[0:0], i_0r0[36:36], i_0r0[4:4]);
  C2 I25 (op1_4_0[1:1], i_0r0[36:36], i_0r1[4:4]);
  C2 I26 (op1_4_0[2:2], i_0r1[36:36], i_0r0[4:4]);
  C2 I27 (op1_4_0[3:3], i_0r1[36:36], i_0r1[4:4]);
  BUFF I28 (termf_1[4:4], op1_4_0[0:0]);
  OR3 I29 (termt_1[4:4], op1_4_0[1:1], op1_4_0[2:2], op1_4_0[3:3]);
  C2 I30 (op1_5_0[0:0], i_0r0[37:37], i_0r0[5:5]);
  C2 I31 (op1_5_0[1:1], i_0r0[37:37], i_0r1[5:5]);
  C2 I32 (op1_5_0[2:2], i_0r1[37:37], i_0r0[5:5]);
  C2 I33 (op1_5_0[3:3], i_0r1[37:37], i_0r1[5:5]);
  BUFF I34 (termf_1[5:5], op1_5_0[0:0]);
  OR3 I35 (termt_1[5:5], op1_5_0[1:1], op1_5_0[2:2], op1_5_0[3:3]);
  C2 I36 (op1_6_0[0:0], i_0r0[38:38], i_0r0[6:6]);
  C2 I37 (op1_6_0[1:1], i_0r0[38:38], i_0r1[6:6]);
  C2 I38 (op1_6_0[2:2], i_0r1[38:38], i_0r0[6:6]);
  C2 I39 (op1_6_0[3:3], i_0r1[38:38], i_0r1[6:6]);
  BUFF I40 (termf_1[6:6], op1_6_0[0:0]);
  OR3 I41 (termt_1[6:6], op1_6_0[1:1], op1_6_0[2:2], op1_6_0[3:3]);
  C2 I42 (op1_7_0[0:0], i_0r0[39:39], i_0r0[7:7]);
  C2 I43 (op1_7_0[1:1], i_0r0[39:39], i_0r1[7:7]);
  C2 I44 (op1_7_0[2:2], i_0r1[39:39], i_0r0[7:7]);
  C2 I45 (op1_7_0[3:3], i_0r1[39:39], i_0r1[7:7]);
  BUFF I46 (termf_1[7:7], op1_7_0[0:0]);
  OR3 I47 (termt_1[7:7], op1_7_0[1:1], op1_7_0[2:2], op1_7_0[3:3]);
  C2 I48 (op1_8_0[0:0], i_0r0[40:40], i_0r0[8:8]);
  C2 I49 (op1_8_0[1:1], i_0r0[40:40], i_0r1[8:8]);
  C2 I50 (op1_8_0[2:2], i_0r1[40:40], i_0r0[8:8]);
  C2 I51 (op1_8_0[3:3], i_0r1[40:40], i_0r1[8:8]);
  BUFF I52 (termf_1[8:8], op1_8_0[0:0]);
  OR3 I53 (termt_1[8:8], op1_8_0[1:1], op1_8_0[2:2], op1_8_0[3:3]);
  C2 I54 (op1_9_0[0:0], i_0r0[41:41], i_0r0[9:9]);
  C2 I55 (op1_9_0[1:1], i_0r0[41:41], i_0r1[9:9]);
  C2 I56 (op1_9_0[2:2], i_0r1[41:41], i_0r0[9:9]);
  C2 I57 (op1_9_0[3:3], i_0r1[41:41], i_0r1[9:9]);
  BUFF I58 (termf_1[9:9], op1_9_0[0:0]);
  OR3 I59 (termt_1[9:9], op1_9_0[1:1], op1_9_0[2:2], op1_9_0[3:3]);
  C2 I60 (op1_10_0[0:0], i_0r0[42:42], i_0r0[10:10]);
  C2 I61 (op1_10_0[1:1], i_0r0[42:42], i_0r1[10:10]);
  C2 I62 (op1_10_0[2:2], i_0r1[42:42], i_0r0[10:10]);
  C2 I63 (op1_10_0[3:3], i_0r1[42:42], i_0r1[10:10]);
  BUFF I64 (termf_1[10:10], op1_10_0[0:0]);
  OR3 I65 (termt_1[10:10], op1_10_0[1:1], op1_10_0[2:2], op1_10_0[3:3]);
  C2 I66 (op1_11_0[0:0], i_0r0[43:43], i_0r0[11:11]);
  C2 I67 (op1_11_0[1:1], i_0r0[43:43], i_0r1[11:11]);
  C2 I68 (op1_11_0[2:2], i_0r1[43:43], i_0r0[11:11]);
  C2 I69 (op1_11_0[3:3], i_0r1[43:43], i_0r1[11:11]);
  BUFF I70 (termf_1[11:11], op1_11_0[0:0]);
  OR3 I71 (termt_1[11:11], op1_11_0[1:1], op1_11_0[2:2], op1_11_0[3:3]);
  C2 I72 (op1_12_0[0:0], i_0r0[44:44], i_0r0[12:12]);
  C2 I73 (op1_12_0[1:1], i_0r0[44:44], i_0r1[12:12]);
  C2 I74 (op1_12_0[2:2], i_0r1[44:44], i_0r0[12:12]);
  C2 I75 (op1_12_0[3:3], i_0r1[44:44], i_0r1[12:12]);
  BUFF I76 (termf_1[12:12], op1_12_0[0:0]);
  OR3 I77 (termt_1[12:12], op1_12_0[1:1], op1_12_0[2:2], op1_12_0[3:3]);
  C2 I78 (op1_13_0[0:0], i_0r0[45:45], i_0r0[13:13]);
  C2 I79 (op1_13_0[1:1], i_0r0[45:45], i_0r1[13:13]);
  C2 I80 (op1_13_0[2:2], i_0r1[45:45], i_0r0[13:13]);
  C2 I81 (op1_13_0[3:3], i_0r1[45:45], i_0r1[13:13]);
  BUFF I82 (termf_1[13:13], op1_13_0[0:0]);
  OR3 I83 (termt_1[13:13], op1_13_0[1:1], op1_13_0[2:2], op1_13_0[3:3]);
  C2 I84 (op1_14_0[0:0], i_0r0[46:46], i_0r0[14:14]);
  C2 I85 (op1_14_0[1:1], i_0r0[46:46], i_0r1[14:14]);
  C2 I86 (op1_14_0[2:2], i_0r1[46:46], i_0r0[14:14]);
  C2 I87 (op1_14_0[3:3], i_0r1[46:46], i_0r1[14:14]);
  BUFF I88 (termf_1[14:14], op1_14_0[0:0]);
  OR3 I89 (termt_1[14:14], op1_14_0[1:1], op1_14_0[2:2], op1_14_0[3:3]);
  C2 I90 (op1_15_0[0:0], i_0r0[47:47], i_0r0[15:15]);
  C2 I91 (op1_15_0[1:1], i_0r0[47:47], i_0r1[15:15]);
  C2 I92 (op1_15_0[2:2], i_0r1[47:47], i_0r0[15:15]);
  C2 I93 (op1_15_0[3:3], i_0r1[47:47], i_0r1[15:15]);
  BUFF I94 (termf_1[15:15], op1_15_0[0:0]);
  OR3 I95 (termt_1[15:15], op1_15_0[1:1], op1_15_0[2:2], op1_15_0[3:3]);
  C2 I96 (op1_16_0[0:0], i_0r0[48:48], i_0r0[16:16]);
  C2 I97 (op1_16_0[1:1], i_0r0[48:48], i_0r1[16:16]);
  C2 I98 (op1_16_0[2:2], i_0r1[48:48], i_0r0[16:16]);
  C2 I99 (op1_16_0[3:3], i_0r1[48:48], i_0r1[16:16]);
  BUFF I100 (termf_1[16:16], op1_16_0[0:0]);
  OR3 I101 (termt_1[16:16], op1_16_0[1:1], op1_16_0[2:2], op1_16_0[3:3]);
  C2 I102 (op1_17_0[0:0], i_0r0[49:49], i_0r0[17:17]);
  C2 I103 (op1_17_0[1:1], i_0r0[49:49], i_0r1[17:17]);
  C2 I104 (op1_17_0[2:2], i_0r1[49:49], i_0r0[17:17]);
  C2 I105 (op1_17_0[3:3], i_0r1[49:49], i_0r1[17:17]);
  BUFF I106 (termf_1[17:17], op1_17_0[0:0]);
  OR3 I107 (termt_1[17:17], op1_17_0[1:1], op1_17_0[2:2], op1_17_0[3:3]);
  C2 I108 (op1_18_0[0:0], i_0r0[50:50], i_0r0[18:18]);
  C2 I109 (op1_18_0[1:1], i_0r0[50:50], i_0r1[18:18]);
  C2 I110 (op1_18_0[2:2], i_0r1[50:50], i_0r0[18:18]);
  C2 I111 (op1_18_0[3:3], i_0r1[50:50], i_0r1[18:18]);
  BUFF I112 (termf_1[18:18], op1_18_0[0:0]);
  OR3 I113 (termt_1[18:18], op1_18_0[1:1], op1_18_0[2:2], op1_18_0[3:3]);
  C2 I114 (op1_19_0[0:0], i_0r0[51:51], i_0r0[19:19]);
  C2 I115 (op1_19_0[1:1], i_0r0[51:51], i_0r1[19:19]);
  C2 I116 (op1_19_0[2:2], i_0r1[51:51], i_0r0[19:19]);
  C2 I117 (op1_19_0[3:3], i_0r1[51:51], i_0r1[19:19]);
  BUFF I118 (termf_1[19:19], op1_19_0[0:0]);
  OR3 I119 (termt_1[19:19], op1_19_0[1:1], op1_19_0[2:2], op1_19_0[3:3]);
  C2 I120 (op1_20_0[0:0], i_0r0[52:52], i_0r0[20:20]);
  C2 I121 (op1_20_0[1:1], i_0r0[52:52], i_0r1[20:20]);
  C2 I122 (op1_20_0[2:2], i_0r1[52:52], i_0r0[20:20]);
  C2 I123 (op1_20_0[3:3], i_0r1[52:52], i_0r1[20:20]);
  BUFF I124 (termf_1[20:20], op1_20_0[0:0]);
  OR3 I125 (termt_1[20:20], op1_20_0[1:1], op1_20_0[2:2], op1_20_0[3:3]);
  C2 I126 (op1_21_0[0:0], i_0r0[53:53], i_0r0[21:21]);
  C2 I127 (op1_21_0[1:1], i_0r0[53:53], i_0r1[21:21]);
  C2 I128 (op1_21_0[2:2], i_0r1[53:53], i_0r0[21:21]);
  C2 I129 (op1_21_0[3:3], i_0r1[53:53], i_0r1[21:21]);
  BUFF I130 (termf_1[21:21], op1_21_0[0:0]);
  OR3 I131 (termt_1[21:21], op1_21_0[1:1], op1_21_0[2:2], op1_21_0[3:3]);
  C2 I132 (op1_22_0[0:0], i_0r0[54:54], i_0r0[22:22]);
  C2 I133 (op1_22_0[1:1], i_0r0[54:54], i_0r1[22:22]);
  C2 I134 (op1_22_0[2:2], i_0r1[54:54], i_0r0[22:22]);
  C2 I135 (op1_22_0[3:3], i_0r1[54:54], i_0r1[22:22]);
  BUFF I136 (termf_1[22:22], op1_22_0[0:0]);
  OR3 I137 (termt_1[22:22], op1_22_0[1:1], op1_22_0[2:2], op1_22_0[3:3]);
  C2 I138 (op1_23_0[0:0], i_0r0[55:55], i_0r0[23:23]);
  C2 I139 (op1_23_0[1:1], i_0r0[55:55], i_0r1[23:23]);
  C2 I140 (op1_23_0[2:2], i_0r1[55:55], i_0r0[23:23]);
  C2 I141 (op1_23_0[3:3], i_0r1[55:55], i_0r1[23:23]);
  BUFF I142 (termf_1[23:23], op1_23_0[0:0]);
  OR3 I143 (termt_1[23:23], op1_23_0[1:1], op1_23_0[2:2], op1_23_0[3:3]);
  C2 I144 (op1_24_0[0:0], i_0r0[56:56], i_0r0[24:24]);
  C2 I145 (op1_24_0[1:1], i_0r0[56:56], i_0r1[24:24]);
  C2 I146 (op1_24_0[2:2], i_0r1[56:56], i_0r0[24:24]);
  C2 I147 (op1_24_0[3:3], i_0r1[56:56], i_0r1[24:24]);
  BUFF I148 (termf_1[24:24], op1_24_0[0:0]);
  OR3 I149 (termt_1[24:24], op1_24_0[1:1], op1_24_0[2:2], op1_24_0[3:3]);
  C2 I150 (op1_25_0[0:0], i_0r0[57:57], i_0r0[25:25]);
  C2 I151 (op1_25_0[1:1], i_0r0[57:57], i_0r1[25:25]);
  C2 I152 (op1_25_0[2:2], i_0r1[57:57], i_0r0[25:25]);
  C2 I153 (op1_25_0[3:3], i_0r1[57:57], i_0r1[25:25]);
  BUFF I154 (termf_1[25:25], op1_25_0[0:0]);
  OR3 I155 (termt_1[25:25], op1_25_0[1:1], op1_25_0[2:2], op1_25_0[3:3]);
  C2 I156 (op1_26_0[0:0], i_0r0[58:58], i_0r0[26:26]);
  C2 I157 (op1_26_0[1:1], i_0r0[58:58], i_0r1[26:26]);
  C2 I158 (op1_26_0[2:2], i_0r1[58:58], i_0r0[26:26]);
  C2 I159 (op1_26_0[3:3], i_0r1[58:58], i_0r1[26:26]);
  BUFF I160 (termf_1[26:26], op1_26_0[0:0]);
  OR3 I161 (termt_1[26:26], op1_26_0[1:1], op1_26_0[2:2], op1_26_0[3:3]);
  C2 I162 (op1_27_0[0:0], i_0r0[59:59], i_0r0[27:27]);
  C2 I163 (op1_27_0[1:1], i_0r0[59:59], i_0r1[27:27]);
  C2 I164 (op1_27_0[2:2], i_0r1[59:59], i_0r0[27:27]);
  C2 I165 (op1_27_0[3:3], i_0r1[59:59], i_0r1[27:27]);
  BUFF I166 (termf_1[27:27], op1_27_0[0:0]);
  OR3 I167 (termt_1[27:27], op1_27_0[1:1], op1_27_0[2:2], op1_27_0[3:3]);
  C2 I168 (op1_28_0[0:0], i_0r0[60:60], i_0r0[28:28]);
  C2 I169 (op1_28_0[1:1], i_0r0[60:60], i_0r1[28:28]);
  C2 I170 (op1_28_0[2:2], i_0r1[60:60], i_0r0[28:28]);
  C2 I171 (op1_28_0[3:3], i_0r1[60:60], i_0r1[28:28]);
  BUFF I172 (termf_1[28:28], op1_28_0[0:0]);
  OR3 I173 (termt_1[28:28], op1_28_0[1:1], op1_28_0[2:2], op1_28_0[3:3]);
  C2 I174 (op1_29_0[0:0], i_0r0[61:61], i_0r0[29:29]);
  C2 I175 (op1_29_0[1:1], i_0r0[61:61], i_0r1[29:29]);
  C2 I176 (op1_29_0[2:2], i_0r1[61:61], i_0r0[29:29]);
  C2 I177 (op1_29_0[3:3], i_0r1[61:61], i_0r1[29:29]);
  BUFF I178 (termf_1[29:29], op1_29_0[0:0]);
  OR3 I179 (termt_1[29:29], op1_29_0[1:1], op1_29_0[2:2], op1_29_0[3:3]);
  C2 I180 (op1_30_0[0:0], i_0r0[62:62], i_0r0[30:30]);
  C2 I181 (op1_30_0[1:1], i_0r0[62:62], i_0r1[30:30]);
  C2 I182 (op1_30_0[2:2], i_0r1[62:62], i_0r0[30:30]);
  C2 I183 (op1_30_0[3:3], i_0r1[62:62], i_0r1[30:30]);
  BUFF I184 (termf_1[30:30], op1_30_0[0:0]);
  OR3 I185 (termt_1[30:30], op1_30_0[1:1], op1_30_0[2:2], op1_30_0[3:3]);
  C2 I186 (op1_31_0[0:0], i_0r0[63:63], i_0r0[31:31]);
  C2 I187 (op1_31_0[1:1], i_0r0[63:63], i_0r1[31:31]);
  C2 I188 (op1_31_0[2:2], i_0r1[63:63], i_0r0[31:31]);
  C2 I189 (op1_31_0[3:3], i_0r1[63:63], i_0r1[31:31]);
  BUFF I190 (termf_1[31:31], op1_31_0[0:0]);
  OR3 I191 (termt_1[31:31], op1_31_0[1:1], op1_31_0[2:2], op1_31_0[3:3]);
  BUFF I192 (o_0r0[0:0], termf_1[0:0]);
  BUFF I193 (o_0r0[1:1], termf_1[1:1]);
  BUFF I194 (o_0r0[2:2], termf_1[2:2]);
  BUFF I195 (o_0r0[3:3], termf_1[3:3]);
  BUFF I196 (o_0r0[4:4], termf_1[4:4]);
  BUFF I197 (o_0r0[5:5], termf_1[5:5]);
  BUFF I198 (o_0r0[6:6], termf_1[6:6]);
  BUFF I199 (o_0r0[7:7], termf_1[7:7]);
  BUFF I200 (o_0r0[8:8], termf_1[8:8]);
  BUFF I201 (o_0r0[9:9], termf_1[9:9]);
  BUFF I202 (o_0r0[10:10], termf_1[10:10]);
  BUFF I203 (o_0r0[11:11], termf_1[11:11]);
  BUFF I204 (o_0r0[12:12], termf_1[12:12]);
  BUFF I205 (o_0r0[13:13], termf_1[13:13]);
  BUFF I206 (o_0r0[14:14], termf_1[14:14]);
  BUFF I207 (o_0r0[15:15], termf_1[15:15]);
  BUFF I208 (o_0r0[16:16], termf_1[16:16]);
  BUFF I209 (o_0r0[17:17], termf_1[17:17]);
  BUFF I210 (o_0r0[18:18], termf_1[18:18]);
  BUFF I211 (o_0r0[19:19], termf_1[19:19]);
  BUFF I212 (o_0r0[20:20], termf_1[20:20]);
  BUFF I213 (o_0r0[21:21], termf_1[21:21]);
  BUFF I214 (o_0r0[22:22], termf_1[22:22]);
  BUFF I215 (o_0r0[23:23], termf_1[23:23]);
  BUFF I216 (o_0r0[24:24], termf_1[24:24]);
  BUFF I217 (o_0r0[25:25], termf_1[25:25]);
  BUFF I218 (o_0r0[26:26], termf_1[26:26]);
  BUFF I219 (o_0r0[27:27], termf_1[27:27]);
  BUFF I220 (o_0r0[28:28], termf_1[28:28]);
  BUFF I221 (o_0r0[29:29], termf_1[29:29]);
  BUFF I222 (o_0r0[30:30], termf_1[30:30]);
  BUFF I223 (o_0r0[31:31], termf_1[31:31]);
  BUFF I224 (o_0r0[32:32], i_0r0[64:64]);
  BUFF I225 (o_0r1[0:0], termt_1[0:0]);
  BUFF I226 (o_0r1[1:1], termt_1[1:1]);
  BUFF I227 (o_0r1[2:2], termt_1[2:2]);
  BUFF I228 (o_0r1[3:3], termt_1[3:3]);
  BUFF I229 (o_0r1[4:4], termt_1[4:4]);
  BUFF I230 (o_0r1[5:5], termt_1[5:5]);
  BUFF I231 (o_0r1[6:6], termt_1[6:6]);
  BUFF I232 (o_0r1[7:7], termt_1[7:7]);
  BUFF I233 (o_0r1[8:8], termt_1[8:8]);
  BUFF I234 (o_0r1[9:9], termt_1[9:9]);
  BUFF I235 (o_0r1[10:10], termt_1[10:10]);
  BUFF I236 (o_0r1[11:11], termt_1[11:11]);
  BUFF I237 (o_0r1[12:12], termt_1[12:12]);
  BUFF I238 (o_0r1[13:13], termt_1[13:13]);
  BUFF I239 (o_0r1[14:14], termt_1[14:14]);
  BUFF I240 (o_0r1[15:15], termt_1[15:15]);
  BUFF I241 (o_0r1[16:16], termt_1[16:16]);
  BUFF I242 (o_0r1[17:17], termt_1[17:17]);
  BUFF I243 (o_0r1[18:18], termt_1[18:18]);
  BUFF I244 (o_0r1[19:19], termt_1[19:19]);
  BUFF I245 (o_0r1[20:20], termt_1[20:20]);
  BUFF I246 (o_0r1[21:21], termt_1[21:21]);
  BUFF I247 (o_0r1[22:22], termt_1[22:22]);
  BUFF I248 (o_0r1[23:23], termt_1[23:23]);
  BUFF I249 (o_0r1[24:24], termt_1[24:24]);
  BUFF I250 (o_0r1[25:25], termt_1[25:25]);
  BUFF I251 (o_0r1[26:26], termt_1[26:26]);
  BUFF I252 (o_0r1[27:27], termt_1[27:27]);
  BUFF I253 (o_0r1[28:28], termt_1[28:28]);
  BUFF I254 (o_0r1[29:29], termt_1[29:29]);
  BUFF I255 (o_0r1[30:30], termt_1[30:30]);
  BUFF I256 (o_0r1[31:31], termt_1[31:31]);
  BUFF I257 (o_0r1[32:32], i_0r1[64:64]);
  BUFF I258 (i_0a, o_0a);
endmodule

// tko65m33_1andi0w32bi32w32b_2apt1o0w32bi64w1b TeakO [
//     (1,TeakOp TeakOpAnd [(0,0,32),(0,32,32)]),
//     (2,TeakOAppend 1 [(1,0,32),(0,64,1)])] [One 65,One 33]
module tko65m33_1andi0w32bi32w32b_2apt1o0w32bi64w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [64:0] i_0r0;
  input [64:0] i_0r1;
  output i_0a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  wire [31:0] termf_1;
  wire [31:0] termt_1;
  wire [3:0] op1_0_0;
  wire [3:0] op1_1_0;
  wire [3:0] op1_2_0;
  wire [3:0] op1_3_0;
  wire [3:0] op1_4_0;
  wire [3:0] op1_5_0;
  wire [3:0] op1_6_0;
  wire [3:0] op1_7_0;
  wire [3:0] op1_8_0;
  wire [3:0] op1_9_0;
  wire [3:0] op1_10_0;
  wire [3:0] op1_11_0;
  wire [3:0] op1_12_0;
  wire [3:0] op1_13_0;
  wire [3:0] op1_14_0;
  wire [3:0] op1_15_0;
  wire [3:0] op1_16_0;
  wire [3:0] op1_17_0;
  wire [3:0] op1_18_0;
  wire [3:0] op1_19_0;
  wire [3:0] op1_20_0;
  wire [3:0] op1_21_0;
  wire [3:0] op1_22_0;
  wire [3:0] op1_23_0;
  wire [3:0] op1_24_0;
  wire [3:0] op1_25_0;
  wire [3:0] op1_26_0;
  wire [3:0] op1_27_0;
  wire [3:0] op1_28_0;
  wire [3:0] op1_29_0;
  wire [3:0] op1_30_0;
  wire [3:0] op1_31_0;
  C2 I0 (op1_0_0[0:0], i_0r0[32:32], i_0r0[0:0]);
  C2 I1 (op1_0_0[1:1], i_0r0[32:32], i_0r1[0:0]);
  C2 I2 (op1_0_0[2:2], i_0r1[32:32], i_0r0[0:0]);
  C2 I3 (op1_0_0[3:3], i_0r1[32:32], i_0r1[0:0]);
  OR3 I4 (termf_1[0:0], op1_0_0[0:0], op1_0_0[1:1], op1_0_0[2:2]);
  BUFF I5 (termt_1[0:0], op1_0_0[3:3]);
  C2 I6 (op1_1_0[0:0], i_0r0[33:33], i_0r0[1:1]);
  C2 I7 (op1_1_0[1:1], i_0r0[33:33], i_0r1[1:1]);
  C2 I8 (op1_1_0[2:2], i_0r1[33:33], i_0r0[1:1]);
  C2 I9 (op1_1_0[3:3], i_0r1[33:33], i_0r1[1:1]);
  OR3 I10 (termf_1[1:1], op1_1_0[0:0], op1_1_0[1:1], op1_1_0[2:2]);
  BUFF I11 (termt_1[1:1], op1_1_0[3:3]);
  C2 I12 (op1_2_0[0:0], i_0r0[34:34], i_0r0[2:2]);
  C2 I13 (op1_2_0[1:1], i_0r0[34:34], i_0r1[2:2]);
  C2 I14 (op1_2_0[2:2], i_0r1[34:34], i_0r0[2:2]);
  C2 I15 (op1_2_0[3:3], i_0r1[34:34], i_0r1[2:2]);
  OR3 I16 (termf_1[2:2], op1_2_0[0:0], op1_2_0[1:1], op1_2_0[2:2]);
  BUFF I17 (termt_1[2:2], op1_2_0[3:3]);
  C2 I18 (op1_3_0[0:0], i_0r0[35:35], i_0r0[3:3]);
  C2 I19 (op1_3_0[1:1], i_0r0[35:35], i_0r1[3:3]);
  C2 I20 (op1_3_0[2:2], i_0r1[35:35], i_0r0[3:3]);
  C2 I21 (op1_3_0[3:3], i_0r1[35:35], i_0r1[3:3]);
  OR3 I22 (termf_1[3:3], op1_3_0[0:0], op1_3_0[1:1], op1_3_0[2:2]);
  BUFF I23 (termt_1[3:3], op1_3_0[3:3]);
  C2 I24 (op1_4_0[0:0], i_0r0[36:36], i_0r0[4:4]);
  C2 I25 (op1_4_0[1:1], i_0r0[36:36], i_0r1[4:4]);
  C2 I26 (op1_4_0[2:2], i_0r1[36:36], i_0r0[4:4]);
  C2 I27 (op1_4_0[3:3], i_0r1[36:36], i_0r1[4:4]);
  OR3 I28 (termf_1[4:4], op1_4_0[0:0], op1_4_0[1:1], op1_4_0[2:2]);
  BUFF I29 (termt_1[4:4], op1_4_0[3:3]);
  C2 I30 (op1_5_0[0:0], i_0r0[37:37], i_0r0[5:5]);
  C2 I31 (op1_5_0[1:1], i_0r0[37:37], i_0r1[5:5]);
  C2 I32 (op1_5_0[2:2], i_0r1[37:37], i_0r0[5:5]);
  C2 I33 (op1_5_0[3:3], i_0r1[37:37], i_0r1[5:5]);
  OR3 I34 (termf_1[5:5], op1_5_0[0:0], op1_5_0[1:1], op1_5_0[2:2]);
  BUFF I35 (termt_1[5:5], op1_5_0[3:3]);
  C2 I36 (op1_6_0[0:0], i_0r0[38:38], i_0r0[6:6]);
  C2 I37 (op1_6_0[1:1], i_0r0[38:38], i_0r1[6:6]);
  C2 I38 (op1_6_0[2:2], i_0r1[38:38], i_0r0[6:6]);
  C2 I39 (op1_6_0[3:3], i_0r1[38:38], i_0r1[6:6]);
  OR3 I40 (termf_1[6:6], op1_6_0[0:0], op1_6_0[1:1], op1_6_0[2:2]);
  BUFF I41 (termt_1[6:6], op1_6_0[3:3]);
  C2 I42 (op1_7_0[0:0], i_0r0[39:39], i_0r0[7:7]);
  C2 I43 (op1_7_0[1:1], i_0r0[39:39], i_0r1[7:7]);
  C2 I44 (op1_7_0[2:2], i_0r1[39:39], i_0r0[7:7]);
  C2 I45 (op1_7_0[3:3], i_0r1[39:39], i_0r1[7:7]);
  OR3 I46 (termf_1[7:7], op1_7_0[0:0], op1_7_0[1:1], op1_7_0[2:2]);
  BUFF I47 (termt_1[7:7], op1_7_0[3:3]);
  C2 I48 (op1_8_0[0:0], i_0r0[40:40], i_0r0[8:8]);
  C2 I49 (op1_8_0[1:1], i_0r0[40:40], i_0r1[8:8]);
  C2 I50 (op1_8_0[2:2], i_0r1[40:40], i_0r0[8:8]);
  C2 I51 (op1_8_0[3:3], i_0r1[40:40], i_0r1[8:8]);
  OR3 I52 (termf_1[8:8], op1_8_0[0:0], op1_8_0[1:1], op1_8_0[2:2]);
  BUFF I53 (termt_1[8:8], op1_8_0[3:3]);
  C2 I54 (op1_9_0[0:0], i_0r0[41:41], i_0r0[9:9]);
  C2 I55 (op1_9_0[1:1], i_0r0[41:41], i_0r1[9:9]);
  C2 I56 (op1_9_0[2:2], i_0r1[41:41], i_0r0[9:9]);
  C2 I57 (op1_9_0[3:3], i_0r1[41:41], i_0r1[9:9]);
  OR3 I58 (termf_1[9:9], op1_9_0[0:0], op1_9_0[1:1], op1_9_0[2:2]);
  BUFF I59 (termt_1[9:9], op1_9_0[3:3]);
  C2 I60 (op1_10_0[0:0], i_0r0[42:42], i_0r0[10:10]);
  C2 I61 (op1_10_0[1:1], i_0r0[42:42], i_0r1[10:10]);
  C2 I62 (op1_10_0[2:2], i_0r1[42:42], i_0r0[10:10]);
  C2 I63 (op1_10_0[3:3], i_0r1[42:42], i_0r1[10:10]);
  OR3 I64 (termf_1[10:10], op1_10_0[0:0], op1_10_0[1:1], op1_10_0[2:2]);
  BUFF I65 (termt_1[10:10], op1_10_0[3:3]);
  C2 I66 (op1_11_0[0:0], i_0r0[43:43], i_0r0[11:11]);
  C2 I67 (op1_11_0[1:1], i_0r0[43:43], i_0r1[11:11]);
  C2 I68 (op1_11_0[2:2], i_0r1[43:43], i_0r0[11:11]);
  C2 I69 (op1_11_0[3:3], i_0r1[43:43], i_0r1[11:11]);
  OR3 I70 (termf_1[11:11], op1_11_0[0:0], op1_11_0[1:1], op1_11_0[2:2]);
  BUFF I71 (termt_1[11:11], op1_11_0[3:3]);
  C2 I72 (op1_12_0[0:0], i_0r0[44:44], i_0r0[12:12]);
  C2 I73 (op1_12_0[1:1], i_0r0[44:44], i_0r1[12:12]);
  C2 I74 (op1_12_0[2:2], i_0r1[44:44], i_0r0[12:12]);
  C2 I75 (op1_12_0[3:3], i_0r1[44:44], i_0r1[12:12]);
  OR3 I76 (termf_1[12:12], op1_12_0[0:0], op1_12_0[1:1], op1_12_0[2:2]);
  BUFF I77 (termt_1[12:12], op1_12_0[3:3]);
  C2 I78 (op1_13_0[0:0], i_0r0[45:45], i_0r0[13:13]);
  C2 I79 (op1_13_0[1:1], i_0r0[45:45], i_0r1[13:13]);
  C2 I80 (op1_13_0[2:2], i_0r1[45:45], i_0r0[13:13]);
  C2 I81 (op1_13_0[3:3], i_0r1[45:45], i_0r1[13:13]);
  OR3 I82 (termf_1[13:13], op1_13_0[0:0], op1_13_0[1:1], op1_13_0[2:2]);
  BUFF I83 (termt_1[13:13], op1_13_0[3:3]);
  C2 I84 (op1_14_0[0:0], i_0r0[46:46], i_0r0[14:14]);
  C2 I85 (op1_14_0[1:1], i_0r0[46:46], i_0r1[14:14]);
  C2 I86 (op1_14_0[2:2], i_0r1[46:46], i_0r0[14:14]);
  C2 I87 (op1_14_0[3:3], i_0r1[46:46], i_0r1[14:14]);
  OR3 I88 (termf_1[14:14], op1_14_0[0:0], op1_14_0[1:1], op1_14_0[2:2]);
  BUFF I89 (termt_1[14:14], op1_14_0[3:3]);
  C2 I90 (op1_15_0[0:0], i_0r0[47:47], i_0r0[15:15]);
  C2 I91 (op1_15_0[1:1], i_0r0[47:47], i_0r1[15:15]);
  C2 I92 (op1_15_0[2:2], i_0r1[47:47], i_0r0[15:15]);
  C2 I93 (op1_15_0[3:3], i_0r1[47:47], i_0r1[15:15]);
  OR3 I94 (termf_1[15:15], op1_15_0[0:0], op1_15_0[1:1], op1_15_0[2:2]);
  BUFF I95 (termt_1[15:15], op1_15_0[3:3]);
  C2 I96 (op1_16_0[0:0], i_0r0[48:48], i_0r0[16:16]);
  C2 I97 (op1_16_0[1:1], i_0r0[48:48], i_0r1[16:16]);
  C2 I98 (op1_16_0[2:2], i_0r1[48:48], i_0r0[16:16]);
  C2 I99 (op1_16_0[3:3], i_0r1[48:48], i_0r1[16:16]);
  OR3 I100 (termf_1[16:16], op1_16_0[0:0], op1_16_0[1:1], op1_16_0[2:2]);
  BUFF I101 (termt_1[16:16], op1_16_0[3:3]);
  C2 I102 (op1_17_0[0:0], i_0r0[49:49], i_0r0[17:17]);
  C2 I103 (op1_17_0[1:1], i_0r0[49:49], i_0r1[17:17]);
  C2 I104 (op1_17_0[2:2], i_0r1[49:49], i_0r0[17:17]);
  C2 I105 (op1_17_0[3:3], i_0r1[49:49], i_0r1[17:17]);
  OR3 I106 (termf_1[17:17], op1_17_0[0:0], op1_17_0[1:1], op1_17_0[2:2]);
  BUFF I107 (termt_1[17:17], op1_17_0[3:3]);
  C2 I108 (op1_18_0[0:0], i_0r0[50:50], i_0r0[18:18]);
  C2 I109 (op1_18_0[1:1], i_0r0[50:50], i_0r1[18:18]);
  C2 I110 (op1_18_0[2:2], i_0r1[50:50], i_0r0[18:18]);
  C2 I111 (op1_18_0[3:3], i_0r1[50:50], i_0r1[18:18]);
  OR3 I112 (termf_1[18:18], op1_18_0[0:0], op1_18_0[1:1], op1_18_0[2:2]);
  BUFF I113 (termt_1[18:18], op1_18_0[3:3]);
  C2 I114 (op1_19_0[0:0], i_0r0[51:51], i_0r0[19:19]);
  C2 I115 (op1_19_0[1:1], i_0r0[51:51], i_0r1[19:19]);
  C2 I116 (op1_19_0[2:2], i_0r1[51:51], i_0r0[19:19]);
  C2 I117 (op1_19_0[3:3], i_0r1[51:51], i_0r1[19:19]);
  OR3 I118 (termf_1[19:19], op1_19_0[0:0], op1_19_0[1:1], op1_19_0[2:2]);
  BUFF I119 (termt_1[19:19], op1_19_0[3:3]);
  C2 I120 (op1_20_0[0:0], i_0r0[52:52], i_0r0[20:20]);
  C2 I121 (op1_20_0[1:1], i_0r0[52:52], i_0r1[20:20]);
  C2 I122 (op1_20_0[2:2], i_0r1[52:52], i_0r0[20:20]);
  C2 I123 (op1_20_0[3:3], i_0r1[52:52], i_0r1[20:20]);
  OR3 I124 (termf_1[20:20], op1_20_0[0:0], op1_20_0[1:1], op1_20_0[2:2]);
  BUFF I125 (termt_1[20:20], op1_20_0[3:3]);
  C2 I126 (op1_21_0[0:0], i_0r0[53:53], i_0r0[21:21]);
  C2 I127 (op1_21_0[1:1], i_0r0[53:53], i_0r1[21:21]);
  C2 I128 (op1_21_0[2:2], i_0r1[53:53], i_0r0[21:21]);
  C2 I129 (op1_21_0[3:3], i_0r1[53:53], i_0r1[21:21]);
  OR3 I130 (termf_1[21:21], op1_21_0[0:0], op1_21_0[1:1], op1_21_0[2:2]);
  BUFF I131 (termt_1[21:21], op1_21_0[3:3]);
  C2 I132 (op1_22_0[0:0], i_0r0[54:54], i_0r0[22:22]);
  C2 I133 (op1_22_0[1:1], i_0r0[54:54], i_0r1[22:22]);
  C2 I134 (op1_22_0[2:2], i_0r1[54:54], i_0r0[22:22]);
  C2 I135 (op1_22_0[3:3], i_0r1[54:54], i_0r1[22:22]);
  OR3 I136 (termf_1[22:22], op1_22_0[0:0], op1_22_0[1:1], op1_22_0[2:2]);
  BUFF I137 (termt_1[22:22], op1_22_0[3:3]);
  C2 I138 (op1_23_0[0:0], i_0r0[55:55], i_0r0[23:23]);
  C2 I139 (op1_23_0[1:1], i_0r0[55:55], i_0r1[23:23]);
  C2 I140 (op1_23_0[2:2], i_0r1[55:55], i_0r0[23:23]);
  C2 I141 (op1_23_0[3:3], i_0r1[55:55], i_0r1[23:23]);
  OR3 I142 (termf_1[23:23], op1_23_0[0:0], op1_23_0[1:1], op1_23_0[2:2]);
  BUFF I143 (termt_1[23:23], op1_23_0[3:3]);
  C2 I144 (op1_24_0[0:0], i_0r0[56:56], i_0r0[24:24]);
  C2 I145 (op1_24_0[1:1], i_0r0[56:56], i_0r1[24:24]);
  C2 I146 (op1_24_0[2:2], i_0r1[56:56], i_0r0[24:24]);
  C2 I147 (op1_24_0[3:3], i_0r1[56:56], i_0r1[24:24]);
  OR3 I148 (termf_1[24:24], op1_24_0[0:0], op1_24_0[1:1], op1_24_0[2:2]);
  BUFF I149 (termt_1[24:24], op1_24_0[3:3]);
  C2 I150 (op1_25_0[0:0], i_0r0[57:57], i_0r0[25:25]);
  C2 I151 (op1_25_0[1:1], i_0r0[57:57], i_0r1[25:25]);
  C2 I152 (op1_25_0[2:2], i_0r1[57:57], i_0r0[25:25]);
  C2 I153 (op1_25_0[3:3], i_0r1[57:57], i_0r1[25:25]);
  OR3 I154 (termf_1[25:25], op1_25_0[0:0], op1_25_0[1:1], op1_25_0[2:2]);
  BUFF I155 (termt_1[25:25], op1_25_0[3:3]);
  C2 I156 (op1_26_0[0:0], i_0r0[58:58], i_0r0[26:26]);
  C2 I157 (op1_26_0[1:1], i_0r0[58:58], i_0r1[26:26]);
  C2 I158 (op1_26_0[2:2], i_0r1[58:58], i_0r0[26:26]);
  C2 I159 (op1_26_0[3:3], i_0r1[58:58], i_0r1[26:26]);
  OR3 I160 (termf_1[26:26], op1_26_0[0:0], op1_26_0[1:1], op1_26_0[2:2]);
  BUFF I161 (termt_1[26:26], op1_26_0[3:3]);
  C2 I162 (op1_27_0[0:0], i_0r0[59:59], i_0r0[27:27]);
  C2 I163 (op1_27_0[1:1], i_0r0[59:59], i_0r1[27:27]);
  C2 I164 (op1_27_0[2:2], i_0r1[59:59], i_0r0[27:27]);
  C2 I165 (op1_27_0[3:3], i_0r1[59:59], i_0r1[27:27]);
  OR3 I166 (termf_1[27:27], op1_27_0[0:0], op1_27_0[1:1], op1_27_0[2:2]);
  BUFF I167 (termt_1[27:27], op1_27_0[3:3]);
  C2 I168 (op1_28_0[0:0], i_0r0[60:60], i_0r0[28:28]);
  C2 I169 (op1_28_0[1:1], i_0r0[60:60], i_0r1[28:28]);
  C2 I170 (op1_28_0[2:2], i_0r1[60:60], i_0r0[28:28]);
  C2 I171 (op1_28_0[3:3], i_0r1[60:60], i_0r1[28:28]);
  OR3 I172 (termf_1[28:28], op1_28_0[0:0], op1_28_0[1:1], op1_28_0[2:2]);
  BUFF I173 (termt_1[28:28], op1_28_0[3:3]);
  C2 I174 (op1_29_0[0:0], i_0r0[61:61], i_0r0[29:29]);
  C2 I175 (op1_29_0[1:1], i_0r0[61:61], i_0r1[29:29]);
  C2 I176 (op1_29_0[2:2], i_0r1[61:61], i_0r0[29:29]);
  C2 I177 (op1_29_0[3:3], i_0r1[61:61], i_0r1[29:29]);
  OR3 I178 (termf_1[29:29], op1_29_0[0:0], op1_29_0[1:1], op1_29_0[2:2]);
  BUFF I179 (termt_1[29:29], op1_29_0[3:3]);
  C2 I180 (op1_30_0[0:0], i_0r0[62:62], i_0r0[30:30]);
  C2 I181 (op1_30_0[1:1], i_0r0[62:62], i_0r1[30:30]);
  C2 I182 (op1_30_0[2:2], i_0r1[62:62], i_0r0[30:30]);
  C2 I183 (op1_30_0[3:3], i_0r1[62:62], i_0r1[30:30]);
  OR3 I184 (termf_1[30:30], op1_30_0[0:0], op1_30_0[1:1], op1_30_0[2:2]);
  BUFF I185 (termt_1[30:30], op1_30_0[3:3]);
  C2 I186 (op1_31_0[0:0], i_0r0[63:63], i_0r0[31:31]);
  C2 I187 (op1_31_0[1:1], i_0r0[63:63], i_0r1[31:31]);
  C2 I188 (op1_31_0[2:2], i_0r1[63:63], i_0r0[31:31]);
  C2 I189 (op1_31_0[3:3], i_0r1[63:63], i_0r1[31:31]);
  OR3 I190 (termf_1[31:31], op1_31_0[0:0], op1_31_0[1:1], op1_31_0[2:2]);
  BUFF I191 (termt_1[31:31], op1_31_0[3:3]);
  BUFF I192 (o_0r0[0:0], termf_1[0:0]);
  BUFF I193 (o_0r0[1:1], termf_1[1:1]);
  BUFF I194 (o_0r0[2:2], termf_1[2:2]);
  BUFF I195 (o_0r0[3:3], termf_1[3:3]);
  BUFF I196 (o_0r0[4:4], termf_1[4:4]);
  BUFF I197 (o_0r0[5:5], termf_1[5:5]);
  BUFF I198 (o_0r0[6:6], termf_1[6:6]);
  BUFF I199 (o_0r0[7:7], termf_1[7:7]);
  BUFF I200 (o_0r0[8:8], termf_1[8:8]);
  BUFF I201 (o_0r0[9:9], termf_1[9:9]);
  BUFF I202 (o_0r0[10:10], termf_1[10:10]);
  BUFF I203 (o_0r0[11:11], termf_1[11:11]);
  BUFF I204 (o_0r0[12:12], termf_1[12:12]);
  BUFF I205 (o_0r0[13:13], termf_1[13:13]);
  BUFF I206 (o_0r0[14:14], termf_1[14:14]);
  BUFF I207 (o_0r0[15:15], termf_1[15:15]);
  BUFF I208 (o_0r0[16:16], termf_1[16:16]);
  BUFF I209 (o_0r0[17:17], termf_1[17:17]);
  BUFF I210 (o_0r0[18:18], termf_1[18:18]);
  BUFF I211 (o_0r0[19:19], termf_1[19:19]);
  BUFF I212 (o_0r0[20:20], termf_1[20:20]);
  BUFF I213 (o_0r0[21:21], termf_1[21:21]);
  BUFF I214 (o_0r0[22:22], termf_1[22:22]);
  BUFF I215 (o_0r0[23:23], termf_1[23:23]);
  BUFF I216 (o_0r0[24:24], termf_1[24:24]);
  BUFF I217 (o_0r0[25:25], termf_1[25:25]);
  BUFF I218 (o_0r0[26:26], termf_1[26:26]);
  BUFF I219 (o_0r0[27:27], termf_1[27:27]);
  BUFF I220 (o_0r0[28:28], termf_1[28:28]);
  BUFF I221 (o_0r0[29:29], termf_1[29:29]);
  BUFF I222 (o_0r0[30:30], termf_1[30:30]);
  BUFF I223 (o_0r0[31:31], termf_1[31:31]);
  BUFF I224 (o_0r0[32:32], i_0r0[64:64]);
  BUFF I225 (o_0r1[0:0], termt_1[0:0]);
  BUFF I226 (o_0r1[1:1], termt_1[1:1]);
  BUFF I227 (o_0r1[2:2], termt_1[2:2]);
  BUFF I228 (o_0r1[3:3], termt_1[3:3]);
  BUFF I229 (o_0r1[4:4], termt_1[4:4]);
  BUFF I230 (o_0r1[5:5], termt_1[5:5]);
  BUFF I231 (o_0r1[6:6], termt_1[6:6]);
  BUFF I232 (o_0r1[7:7], termt_1[7:7]);
  BUFF I233 (o_0r1[8:8], termt_1[8:8]);
  BUFF I234 (o_0r1[9:9], termt_1[9:9]);
  BUFF I235 (o_0r1[10:10], termt_1[10:10]);
  BUFF I236 (o_0r1[11:11], termt_1[11:11]);
  BUFF I237 (o_0r1[12:12], termt_1[12:12]);
  BUFF I238 (o_0r1[13:13], termt_1[13:13]);
  BUFF I239 (o_0r1[14:14], termt_1[14:14]);
  BUFF I240 (o_0r1[15:15], termt_1[15:15]);
  BUFF I241 (o_0r1[16:16], termt_1[16:16]);
  BUFF I242 (o_0r1[17:17], termt_1[17:17]);
  BUFF I243 (o_0r1[18:18], termt_1[18:18]);
  BUFF I244 (o_0r1[19:19], termt_1[19:19]);
  BUFF I245 (o_0r1[20:20], termt_1[20:20]);
  BUFF I246 (o_0r1[21:21], termt_1[21:21]);
  BUFF I247 (o_0r1[22:22], termt_1[22:22]);
  BUFF I248 (o_0r1[23:23], termt_1[23:23]);
  BUFF I249 (o_0r1[24:24], termt_1[24:24]);
  BUFF I250 (o_0r1[25:25], termt_1[25:25]);
  BUFF I251 (o_0r1[26:26], termt_1[26:26]);
  BUFF I252 (o_0r1[27:27], termt_1[27:27]);
  BUFF I253 (o_0r1[28:28], termt_1[28:28]);
  BUFF I254 (o_0r1[29:29], termt_1[29:29]);
  BUFF I255 (o_0r1[30:30], termt_1[30:30]);
  BUFF I256 (o_0r1[31:31], termt_1[31:31]);
  BUFF I257 (o_0r1[32:32], i_0r1[64:64]);
  BUFF I258 (i_0a, o_0a);
endmodule

// tks4_o0w4_2m3m4m5m6m7mambo0w0_dmfo0w0_1m9o0w0_co0w0_0m8meo0w0 TeakS (0+:4) [([Imp 2 0,Imp 3 0,Imp 4 
//   0,Imp 5 0,Imp 6 0,Imp 7 0,Imp 10 0,Imp 11 0],0),([Imp 13 0,Imp 15 0],0),([Imp 1 0,Imp 9 0],0),([Imp 
//   12 0],0),([Imp 0 0,Imp 8 0,Imp 14 0],0)] [One 4,Many [0,0,0,0,0]]
module tks4_o0w4_2m3m4m5m6m7mambo0w0_dmfo0w0_1m9o0w0_co0w0_0m8meo0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire sel_4;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire gsel_4;
  wire oack_0;
  wire [7:0] match0_0;
  wire [2:0] simp131_0;
  wire [1:0] simp141_0;
  wire [1:0] simp151_0;
  wire [1:0] simp161_0;
  wire [1:0] simp171_0;
  wire [1:0] simp181_0;
  wire [1:0] simp191_0;
  wire [1:0] simp201_0;
  wire [1:0] simp211_0;
  wire [1:0] match1_0;
  wire [1:0] simp241_0;
  wire [1:0] simp251_0;
  wire [1:0] match2_0;
  wire [1:0] simp281_0;
  wire [1:0] simp291_0;
  wire match3_0;
  wire [1:0] simp321_0;
  wire [2:0] match4_0;
  wire [1:0] simp351_0;
  wire [1:0] simp361_0;
  wire [1:0] simp371_0;
  wire [3:0] comp_0;
  wire [1:0] simp481_0;
  wire [1:0] simp541_0;
  NOR3 I0 (simp131_0[0:0], match0_0[0:0], match0_0[1:1], match0_0[2:2]);
  NOR3 I1 (simp131_0[1:1], match0_0[3:3], match0_0[4:4], match0_0[5:5]);
  NOR2 I2 (simp131_0[2:2], match0_0[6:6], match0_0[7:7]);
  NAND3 I3 (sel_0, simp131_0[0:0], simp131_0[1:1], simp131_0[2:2]);
  C3 I4 (simp141_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I5 (simp141_0[1:1], i_0r0[3:3]);
  C2 I6 (match0_0[0:0], simp141_0[0:0], simp141_0[1:1]);
  C3 I7 (simp151_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I8 (simp151_0[1:1], i_0r0[3:3]);
  C2 I9 (match0_0[1:1], simp151_0[0:0], simp151_0[1:1]);
  C3 I10 (simp161_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I11 (simp161_0[1:1], i_0r0[3:3]);
  C2 I12 (match0_0[2:2], simp161_0[0:0], simp161_0[1:1]);
  C3 I13 (simp171_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I14 (simp171_0[1:1], i_0r0[3:3]);
  C2 I15 (match0_0[3:3], simp171_0[0:0], simp171_0[1:1]);
  C3 I16 (simp181_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I17 (simp181_0[1:1], i_0r0[3:3]);
  C2 I18 (match0_0[4:4], simp181_0[0:0], simp181_0[1:1]);
  C3 I19 (simp191_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I20 (simp191_0[1:1], i_0r0[3:3]);
  C2 I21 (match0_0[5:5], simp191_0[0:0], simp191_0[1:1]);
  C3 I22 (simp201_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I23 (simp201_0[1:1], i_0r1[3:3]);
  C2 I24 (match0_0[6:6], simp201_0[0:0], simp201_0[1:1]);
  C3 I25 (simp211_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I26 (simp211_0[1:1], i_0r1[3:3]);
  C2 I27 (match0_0[7:7], simp211_0[0:0], simp211_0[1:1]);
  OR2 I28 (sel_1, match1_0[0:0], match1_0[1:1]);
  C3 I29 (simp241_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I30 (simp241_0[1:1], i_0r1[3:3]);
  C2 I31 (match1_0[0:0], simp241_0[0:0], simp241_0[1:1]);
  C3 I32 (simp251_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I33 (simp251_0[1:1], i_0r1[3:3]);
  C2 I34 (match1_0[1:1], simp251_0[0:0], simp251_0[1:1]);
  OR2 I35 (sel_2, match2_0[0:0], match2_0[1:1]);
  C3 I36 (simp281_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I37 (simp281_0[1:1], i_0r0[3:3]);
  C2 I38 (match2_0[0:0], simp281_0[0:0], simp281_0[1:1]);
  C3 I39 (simp291_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I40 (simp291_0[1:1], i_0r1[3:3]);
  C2 I41 (match2_0[1:1], simp291_0[0:0], simp291_0[1:1]);
  BUFF I42 (sel_3, match3_0);
  C3 I43 (simp321_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I44 (simp321_0[1:1], i_0r1[3:3]);
  C2 I45 (match3_0, simp321_0[0:0], simp321_0[1:1]);
  OR3 I46 (sel_4, match4_0[0:0], match4_0[1:1], match4_0[2:2]);
  C3 I47 (simp351_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I48 (simp351_0[1:1], i_0r0[3:3]);
  C2 I49 (match4_0[0:0], simp351_0[0:0], simp351_0[1:1]);
  C3 I50 (simp361_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I51 (simp361_0[1:1], i_0r1[3:3]);
  C2 I52 (match4_0[1:1], simp361_0[0:0], simp361_0[1:1]);
  C3 I53 (simp371_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I54 (simp371_0[1:1], i_0r1[3:3]);
  C2 I55 (match4_0[2:2], simp371_0[0:0], simp371_0[1:1]);
  C2 I56 (gsel_0, sel_0, icomplete_0);
  C2 I57 (gsel_1, sel_1, icomplete_0);
  C2 I58 (gsel_2, sel_2, icomplete_0);
  C2 I59 (gsel_3, sel_3, icomplete_0);
  C2 I60 (gsel_4, sel_4, icomplete_0);
  OR2 I61 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I62 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I63 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I64 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  C3 I65 (simp481_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  BUFF I66 (simp481_0[1:1], comp_0[3:3]);
  C2 I67 (icomplete_0, simp481_0[0:0], simp481_0[1:1]);
  BUFF I68 (o_0r, gsel_0);
  BUFF I69 (o_1r, gsel_1);
  BUFF I70 (o_2r, gsel_2);
  BUFF I71 (o_3r, gsel_3);
  BUFF I72 (o_4r, gsel_4);
  NOR3 I73 (simp541_0[0:0], o_0a, o_1a, o_2a);
  NOR2 I74 (simp541_0[1:1], o_3a, o_4a);
  NAND2 I75 (oack_0, simp541_0[0:0], simp541_0[1:1]);
  C2 I76 (i_0a, oack_0, icomplete_0);
endmodule

// tks4_o0w4_0c8m1c8mcmdmemfo0w0_2m3m4m5m6m7mambo0w0 TeakS (0+:4) [([Imp 0 8,Imp 1 8,Imp 12 0,Imp 13 0,
//   Imp 14 0,Imp 15 0],0),([Imp 2 0,Imp 3 0,Imp 4 0,Imp 5 0,Imp 6 0,Imp 7 0,Imp 10 0,Imp 11 0],0)] [One 
//   4,Many [0,0]]
module tks4_o0w4_0c8m1c8mcmdmemfo0w0_2m3m4m5m6m7mambo0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire [5:0] match0_0;
  wire [1:0] simp71_0;
  wire [1:0] simp101_0;
  wire [1:0] simp111_0;
  wire [1:0] simp121_0;
  wire [1:0] simp131_0;
  wire [7:0] match1_0;
  wire [2:0] simp151_0;
  wire [1:0] simp161_0;
  wire [1:0] simp171_0;
  wire [1:0] simp181_0;
  wire [1:0] simp191_0;
  wire [1:0] simp201_0;
  wire [1:0] simp211_0;
  wire [1:0] simp221_0;
  wire [1:0] simp231_0;
  wire [3:0] comp_0;
  wire [1:0] simp311_0;
  NOR3 I0 (simp71_0[0:0], match0_0[0:0], match0_0[1:1], match0_0[2:2]);
  NOR3 I1 (simp71_0[1:1], match0_0[3:3], match0_0[4:4], match0_0[5:5]);
  NAND2 I2 (sel_0, simp71_0[0:0], simp71_0[1:1]);
  C3 I3 (match0_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I4 (match0_0[1:1], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I5 (simp101_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I6 (simp101_0[1:1], i_0r1[3:3]);
  C2 I7 (match0_0[2:2], simp101_0[0:0], simp101_0[1:1]);
  C3 I8 (simp111_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I9 (simp111_0[1:1], i_0r1[3:3]);
  C2 I10 (match0_0[3:3], simp111_0[0:0], simp111_0[1:1]);
  C3 I11 (simp121_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I12 (simp121_0[1:1], i_0r1[3:3]);
  C2 I13 (match0_0[4:4], simp121_0[0:0], simp121_0[1:1]);
  C3 I14 (simp131_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I15 (simp131_0[1:1], i_0r1[3:3]);
  C2 I16 (match0_0[5:5], simp131_0[0:0], simp131_0[1:1]);
  NOR3 I17 (simp151_0[0:0], match1_0[0:0], match1_0[1:1], match1_0[2:2]);
  NOR3 I18 (simp151_0[1:1], match1_0[3:3], match1_0[4:4], match1_0[5:5]);
  NOR2 I19 (simp151_0[2:2], match1_0[6:6], match1_0[7:7]);
  NAND3 I20 (sel_1, simp151_0[0:0], simp151_0[1:1], simp151_0[2:2]);
  C3 I21 (simp161_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I22 (simp161_0[1:1], i_0r0[3:3]);
  C2 I23 (match1_0[0:0], simp161_0[0:0], simp161_0[1:1]);
  C3 I24 (simp171_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I25 (simp171_0[1:1], i_0r0[3:3]);
  C2 I26 (match1_0[1:1], simp171_0[0:0], simp171_0[1:1]);
  C3 I27 (simp181_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I28 (simp181_0[1:1], i_0r0[3:3]);
  C2 I29 (match1_0[2:2], simp181_0[0:0], simp181_0[1:1]);
  C3 I30 (simp191_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I31 (simp191_0[1:1], i_0r0[3:3]);
  C2 I32 (match1_0[3:3], simp191_0[0:0], simp191_0[1:1]);
  C3 I33 (simp201_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I34 (simp201_0[1:1], i_0r0[3:3]);
  C2 I35 (match1_0[4:4], simp201_0[0:0], simp201_0[1:1]);
  C3 I36 (simp211_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I37 (simp211_0[1:1], i_0r0[3:3]);
  C2 I38 (match1_0[5:5], simp211_0[0:0], simp211_0[1:1]);
  C3 I39 (simp221_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I40 (simp221_0[1:1], i_0r1[3:3]);
  C2 I41 (match1_0[6:6], simp221_0[0:0], simp221_0[1:1]);
  C3 I42 (simp231_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I43 (simp231_0[1:1], i_0r1[3:3]);
  C2 I44 (match1_0[7:7], simp231_0[0:0], simp231_0[1:1]);
  C2 I45 (gsel_0, sel_0, icomplete_0);
  C2 I46 (gsel_1, sel_1, icomplete_0);
  OR2 I47 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I48 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I49 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I50 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  C3 I51 (simp311_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  BUFF I52 (simp311_0[1:1], comp_0[3:3]);
  C2 I53 (icomplete_0, simp311_0[0:0], simp311_0[1:1]);
  BUFF I54 (o_0r, gsel_0);
  BUFF I55 (o_1r, gsel_1);
  OR2 I56 (oack_0, o_0a, o_1a);
  C2 I57 (i_0a, oack_0, icomplete_0);
endmodule

// tkj0m0_0_0 TeakJ [Many [0,0,0],One 0]
module tkj0m0_0_0 (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  output o_0r;
  input o_0a;
  input reset;
  C3 I0 (o_0r, i_0r, i_1r, i_2r);
  BUFF I1 (i_0a, o_0a);
  BUFF I2 (i_1a, o_0a);
  BUFF I3 (i_2a, o_0a);
endmodule

// tkf65mo0w0_o0w65 TeakF [0,0] [One 65,Many [0,65]]
module tkf65mo0w0_o0w65 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [64:0] i_0r0;
  input [64:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [64:0] o_1r0;
  output [64:0] o_1r1;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire [64:0] comp_0;
  wire [21:0] simp671_0;
  wire [7:0] simp672_0;
  wire [2:0] simp673_0;
  OR2 I0 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (comp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (comp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (comp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (comp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (comp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (comp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (comp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (comp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (comp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (comp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (comp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (comp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (comp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (comp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (comp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (comp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (comp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (comp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (comp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (comp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (comp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (comp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (comp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (comp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I30 (comp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I31 (comp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I32 (comp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  OR2 I33 (comp_0[33:33], i_0r0[33:33], i_0r1[33:33]);
  OR2 I34 (comp_0[34:34], i_0r0[34:34], i_0r1[34:34]);
  OR2 I35 (comp_0[35:35], i_0r0[35:35], i_0r1[35:35]);
  OR2 I36 (comp_0[36:36], i_0r0[36:36], i_0r1[36:36]);
  OR2 I37 (comp_0[37:37], i_0r0[37:37], i_0r1[37:37]);
  OR2 I38 (comp_0[38:38], i_0r0[38:38], i_0r1[38:38]);
  OR2 I39 (comp_0[39:39], i_0r0[39:39], i_0r1[39:39]);
  OR2 I40 (comp_0[40:40], i_0r0[40:40], i_0r1[40:40]);
  OR2 I41 (comp_0[41:41], i_0r0[41:41], i_0r1[41:41]);
  OR2 I42 (comp_0[42:42], i_0r0[42:42], i_0r1[42:42]);
  OR2 I43 (comp_0[43:43], i_0r0[43:43], i_0r1[43:43]);
  OR2 I44 (comp_0[44:44], i_0r0[44:44], i_0r1[44:44]);
  OR2 I45 (comp_0[45:45], i_0r0[45:45], i_0r1[45:45]);
  OR2 I46 (comp_0[46:46], i_0r0[46:46], i_0r1[46:46]);
  OR2 I47 (comp_0[47:47], i_0r0[47:47], i_0r1[47:47]);
  OR2 I48 (comp_0[48:48], i_0r0[48:48], i_0r1[48:48]);
  OR2 I49 (comp_0[49:49], i_0r0[49:49], i_0r1[49:49]);
  OR2 I50 (comp_0[50:50], i_0r0[50:50], i_0r1[50:50]);
  OR2 I51 (comp_0[51:51], i_0r0[51:51], i_0r1[51:51]);
  OR2 I52 (comp_0[52:52], i_0r0[52:52], i_0r1[52:52]);
  OR2 I53 (comp_0[53:53], i_0r0[53:53], i_0r1[53:53]);
  OR2 I54 (comp_0[54:54], i_0r0[54:54], i_0r1[54:54]);
  OR2 I55 (comp_0[55:55], i_0r0[55:55], i_0r1[55:55]);
  OR2 I56 (comp_0[56:56], i_0r0[56:56], i_0r1[56:56]);
  OR2 I57 (comp_0[57:57], i_0r0[57:57], i_0r1[57:57]);
  OR2 I58 (comp_0[58:58], i_0r0[58:58], i_0r1[58:58]);
  OR2 I59 (comp_0[59:59], i_0r0[59:59], i_0r1[59:59]);
  OR2 I60 (comp_0[60:60], i_0r0[60:60], i_0r1[60:60]);
  OR2 I61 (comp_0[61:61], i_0r0[61:61], i_0r1[61:61]);
  OR2 I62 (comp_0[62:62], i_0r0[62:62], i_0r1[62:62]);
  OR2 I63 (comp_0[63:63], i_0r0[63:63], i_0r1[63:63]);
  OR2 I64 (comp_0[64:64], i_0r0[64:64], i_0r1[64:64]);
  C3 I65 (simp671_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I66 (simp671_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C3 I67 (simp671_0[2:2], comp_0[6:6], comp_0[7:7], comp_0[8:8]);
  C3 I68 (simp671_0[3:3], comp_0[9:9], comp_0[10:10], comp_0[11:11]);
  C3 I69 (simp671_0[4:4], comp_0[12:12], comp_0[13:13], comp_0[14:14]);
  C3 I70 (simp671_0[5:5], comp_0[15:15], comp_0[16:16], comp_0[17:17]);
  C3 I71 (simp671_0[6:6], comp_0[18:18], comp_0[19:19], comp_0[20:20]);
  C3 I72 (simp671_0[7:7], comp_0[21:21], comp_0[22:22], comp_0[23:23]);
  C3 I73 (simp671_0[8:8], comp_0[24:24], comp_0[25:25], comp_0[26:26]);
  C3 I74 (simp671_0[9:9], comp_0[27:27], comp_0[28:28], comp_0[29:29]);
  C3 I75 (simp671_0[10:10], comp_0[30:30], comp_0[31:31], comp_0[32:32]);
  C3 I76 (simp671_0[11:11], comp_0[33:33], comp_0[34:34], comp_0[35:35]);
  C3 I77 (simp671_0[12:12], comp_0[36:36], comp_0[37:37], comp_0[38:38]);
  C3 I78 (simp671_0[13:13], comp_0[39:39], comp_0[40:40], comp_0[41:41]);
  C3 I79 (simp671_0[14:14], comp_0[42:42], comp_0[43:43], comp_0[44:44]);
  C3 I80 (simp671_0[15:15], comp_0[45:45], comp_0[46:46], comp_0[47:47]);
  C3 I81 (simp671_0[16:16], comp_0[48:48], comp_0[49:49], comp_0[50:50]);
  C3 I82 (simp671_0[17:17], comp_0[51:51], comp_0[52:52], comp_0[53:53]);
  C3 I83 (simp671_0[18:18], comp_0[54:54], comp_0[55:55], comp_0[56:56]);
  C3 I84 (simp671_0[19:19], comp_0[57:57], comp_0[58:58], comp_0[59:59]);
  C3 I85 (simp671_0[20:20], comp_0[60:60], comp_0[61:61], comp_0[62:62]);
  C2 I86 (simp671_0[21:21], comp_0[63:63], comp_0[64:64]);
  C3 I87 (simp672_0[0:0], simp671_0[0:0], simp671_0[1:1], simp671_0[2:2]);
  C3 I88 (simp672_0[1:1], simp671_0[3:3], simp671_0[4:4], simp671_0[5:5]);
  C3 I89 (simp672_0[2:2], simp671_0[6:6], simp671_0[7:7], simp671_0[8:8]);
  C3 I90 (simp672_0[3:3], simp671_0[9:9], simp671_0[10:10], simp671_0[11:11]);
  C3 I91 (simp672_0[4:4], simp671_0[12:12], simp671_0[13:13], simp671_0[14:14]);
  C3 I92 (simp672_0[5:5], simp671_0[15:15], simp671_0[16:16], simp671_0[17:17]);
  C3 I93 (simp672_0[6:6], simp671_0[18:18], simp671_0[19:19], simp671_0[20:20]);
  BUFF I94 (simp672_0[7:7], simp671_0[21:21]);
  C3 I95 (simp673_0[0:0], simp672_0[0:0], simp672_0[1:1], simp672_0[2:2]);
  C3 I96 (simp673_0[1:1], simp672_0[3:3], simp672_0[4:4], simp672_0[5:5]);
  C2 I97 (simp673_0[2:2], simp672_0[6:6], simp672_0[7:7]);
  C3 I98 (icomplete_0, simp673_0[0:0], simp673_0[1:1], simp673_0[2:2]);
  BUFF I99 (o_1r0[0:0], i_0r0[0:0]);
  BUFF I100 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I101 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I102 (o_1r0[3:3], i_0r0[3:3]);
  BUFF I103 (o_1r0[4:4], i_0r0[4:4]);
  BUFF I104 (o_1r0[5:5], i_0r0[5:5]);
  BUFF I105 (o_1r0[6:6], i_0r0[6:6]);
  BUFF I106 (o_1r0[7:7], i_0r0[7:7]);
  BUFF I107 (o_1r0[8:8], i_0r0[8:8]);
  BUFF I108 (o_1r0[9:9], i_0r0[9:9]);
  BUFF I109 (o_1r0[10:10], i_0r0[10:10]);
  BUFF I110 (o_1r0[11:11], i_0r0[11:11]);
  BUFF I111 (o_1r0[12:12], i_0r0[12:12]);
  BUFF I112 (o_1r0[13:13], i_0r0[13:13]);
  BUFF I113 (o_1r0[14:14], i_0r0[14:14]);
  BUFF I114 (o_1r0[15:15], i_0r0[15:15]);
  BUFF I115 (o_1r0[16:16], i_0r0[16:16]);
  BUFF I116 (o_1r0[17:17], i_0r0[17:17]);
  BUFF I117 (o_1r0[18:18], i_0r0[18:18]);
  BUFF I118 (o_1r0[19:19], i_0r0[19:19]);
  BUFF I119 (o_1r0[20:20], i_0r0[20:20]);
  BUFF I120 (o_1r0[21:21], i_0r0[21:21]);
  BUFF I121 (o_1r0[22:22], i_0r0[22:22]);
  BUFF I122 (o_1r0[23:23], i_0r0[23:23]);
  BUFF I123 (o_1r0[24:24], i_0r0[24:24]);
  BUFF I124 (o_1r0[25:25], i_0r0[25:25]);
  BUFF I125 (o_1r0[26:26], i_0r0[26:26]);
  BUFF I126 (o_1r0[27:27], i_0r0[27:27]);
  BUFF I127 (o_1r0[28:28], i_0r0[28:28]);
  BUFF I128 (o_1r0[29:29], i_0r0[29:29]);
  BUFF I129 (o_1r0[30:30], i_0r0[30:30]);
  BUFF I130 (o_1r0[31:31], i_0r0[31:31]);
  BUFF I131 (o_1r0[32:32], i_0r0[32:32]);
  BUFF I132 (o_1r0[33:33], i_0r0[33:33]);
  BUFF I133 (o_1r0[34:34], i_0r0[34:34]);
  BUFF I134 (o_1r0[35:35], i_0r0[35:35]);
  BUFF I135 (o_1r0[36:36], i_0r0[36:36]);
  BUFF I136 (o_1r0[37:37], i_0r0[37:37]);
  BUFF I137 (o_1r0[38:38], i_0r0[38:38]);
  BUFF I138 (o_1r0[39:39], i_0r0[39:39]);
  BUFF I139 (o_1r0[40:40], i_0r0[40:40]);
  BUFF I140 (o_1r0[41:41], i_0r0[41:41]);
  BUFF I141 (o_1r0[42:42], i_0r0[42:42]);
  BUFF I142 (o_1r0[43:43], i_0r0[43:43]);
  BUFF I143 (o_1r0[44:44], i_0r0[44:44]);
  BUFF I144 (o_1r0[45:45], i_0r0[45:45]);
  BUFF I145 (o_1r0[46:46], i_0r0[46:46]);
  BUFF I146 (o_1r0[47:47], i_0r0[47:47]);
  BUFF I147 (o_1r0[48:48], i_0r0[48:48]);
  BUFF I148 (o_1r0[49:49], i_0r0[49:49]);
  BUFF I149 (o_1r0[50:50], i_0r0[50:50]);
  BUFF I150 (o_1r0[51:51], i_0r0[51:51]);
  BUFF I151 (o_1r0[52:52], i_0r0[52:52]);
  BUFF I152 (o_1r0[53:53], i_0r0[53:53]);
  BUFF I153 (o_1r0[54:54], i_0r0[54:54]);
  BUFF I154 (o_1r0[55:55], i_0r0[55:55]);
  BUFF I155 (o_1r0[56:56], i_0r0[56:56]);
  BUFF I156 (o_1r0[57:57], i_0r0[57:57]);
  BUFF I157 (o_1r0[58:58], i_0r0[58:58]);
  BUFF I158 (o_1r0[59:59], i_0r0[59:59]);
  BUFF I159 (o_1r0[60:60], i_0r0[60:60]);
  BUFF I160 (o_1r0[61:61], i_0r0[61:61]);
  BUFF I161 (o_1r0[62:62], i_0r0[62:62]);
  BUFF I162 (o_1r0[63:63], i_0r0[63:63]);
  BUFF I163 (o_1r0[64:64], i_0r0[64:64]);
  BUFF I164 (o_1r1[0:0], i_0r1[0:0]);
  BUFF I165 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I166 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I167 (o_1r1[3:3], i_0r1[3:3]);
  BUFF I168 (o_1r1[4:4], i_0r1[4:4]);
  BUFF I169 (o_1r1[5:5], i_0r1[5:5]);
  BUFF I170 (o_1r1[6:6], i_0r1[6:6]);
  BUFF I171 (o_1r1[7:7], i_0r1[7:7]);
  BUFF I172 (o_1r1[8:8], i_0r1[8:8]);
  BUFF I173 (o_1r1[9:9], i_0r1[9:9]);
  BUFF I174 (o_1r1[10:10], i_0r1[10:10]);
  BUFF I175 (o_1r1[11:11], i_0r1[11:11]);
  BUFF I176 (o_1r1[12:12], i_0r1[12:12]);
  BUFF I177 (o_1r1[13:13], i_0r1[13:13]);
  BUFF I178 (o_1r1[14:14], i_0r1[14:14]);
  BUFF I179 (o_1r1[15:15], i_0r1[15:15]);
  BUFF I180 (o_1r1[16:16], i_0r1[16:16]);
  BUFF I181 (o_1r1[17:17], i_0r1[17:17]);
  BUFF I182 (o_1r1[18:18], i_0r1[18:18]);
  BUFF I183 (o_1r1[19:19], i_0r1[19:19]);
  BUFF I184 (o_1r1[20:20], i_0r1[20:20]);
  BUFF I185 (o_1r1[21:21], i_0r1[21:21]);
  BUFF I186 (o_1r1[22:22], i_0r1[22:22]);
  BUFF I187 (o_1r1[23:23], i_0r1[23:23]);
  BUFF I188 (o_1r1[24:24], i_0r1[24:24]);
  BUFF I189 (o_1r1[25:25], i_0r1[25:25]);
  BUFF I190 (o_1r1[26:26], i_0r1[26:26]);
  BUFF I191 (o_1r1[27:27], i_0r1[27:27]);
  BUFF I192 (o_1r1[28:28], i_0r1[28:28]);
  BUFF I193 (o_1r1[29:29], i_0r1[29:29]);
  BUFF I194 (o_1r1[30:30], i_0r1[30:30]);
  BUFF I195 (o_1r1[31:31], i_0r1[31:31]);
  BUFF I196 (o_1r1[32:32], i_0r1[32:32]);
  BUFF I197 (o_1r1[33:33], i_0r1[33:33]);
  BUFF I198 (o_1r1[34:34], i_0r1[34:34]);
  BUFF I199 (o_1r1[35:35], i_0r1[35:35]);
  BUFF I200 (o_1r1[36:36], i_0r1[36:36]);
  BUFF I201 (o_1r1[37:37], i_0r1[37:37]);
  BUFF I202 (o_1r1[38:38], i_0r1[38:38]);
  BUFF I203 (o_1r1[39:39], i_0r1[39:39]);
  BUFF I204 (o_1r1[40:40], i_0r1[40:40]);
  BUFF I205 (o_1r1[41:41], i_0r1[41:41]);
  BUFF I206 (o_1r1[42:42], i_0r1[42:42]);
  BUFF I207 (o_1r1[43:43], i_0r1[43:43]);
  BUFF I208 (o_1r1[44:44], i_0r1[44:44]);
  BUFF I209 (o_1r1[45:45], i_0r1[45:45]);
  BUFF I210 (o_1r1[46:46], i_0r1[46:46]);
  BUFF I211 (o_1r1[47:47], i_0r1[47:47]);
  BUFF I212 (o_1r1[48:48], i_0r1[48:48]);
  BUFF I213 (o_1r1[49:49], i_0r1[49:49]);
  BUFF I214 (o_1r1[50:50], i_0r1[50:50]);
  BUFF I215 (o_1r1[51:51], i_0r1[51:51]);
  BUFF I216 (o_1r1[52:52], i_0r1[52:52]);
  BUFF I217 (o_1r1[53:53], i_0r1[53:53]);
  BUFF I218 (o_1r1[54:54], i_0r1[54:54]);
  BUFF I219 (o_1r1[55:55], i_0r1[55:55]);
  BUFF I220 (o_1r1[56:56], i_0r1[56:56]);
  BUFF I221 (o_1r1[57:57], i_0r1[57:57]);
  BUFF I222 (o_1r1[58:58], i_0r1[58:58]);
  BUFF I223 (o_1r1[59:59], i_0r1[59:59]);
  BUFF I224 (o_1r1[60:60], i_0r1[60:60]);
  BUFF I225 (o_1r1[61:61], i_0r1[61:61]);
  BUFF I226 (o_1r1[62:62], i_0r1[62:62]);
  BUFF I227 (o_1r1[63:63], i_0r1[63:63]);
  BUFF I228 (o_1r1[64:64], i_0r1[64:64]);
  BUFF I229 (o_0r, icomplete_0);
  C3 I230 (i_0a, icomplete_0, o_0a, o_1a);
endmodule

// tkm4x33b TeakM [Many [33,33,33,33],One 33]
module tkm4x33b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, o_0r0, o_0r1, o_0a, reset);
  input [32:0] i_0r0;
  input [32:0] i_0r1;
  output i_0a;
  input [32:0] i_1r0;
  input [32:0] i_1r1;
  output i_1a;
  input [32:0] i_2r0;
  input [32:0] i_2r1;
  output i_2a;
  input [32:0] i_3r0;
  input [32:0] i_3r1;
  output i_3a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  wire [32:0] gfint_0;
  wire [32:0] gfint_1;
  wire [32:0] gfint_2;
  wire [32:0] gfint_3;
  wire [32:0] gtint_0;
  wire [32:0] gtint_1;
  wire [32:0] gtint_2;
  wire [32:0] gtint_3;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire icomp_3;
  wire nchosen_0;
  wire [1:0] simp181_0;
  wire [1:0] simp191_0;
  wire [1:0] simp201_0;
  wire [1:0] simp211_0;
  wire [1:0] simp221_0;
  wire [1:0] simp231_0;
  wire [1:0] simp241_0;
  wire [1:0] simp251_0;
  wire [1:0] simp261_0;
  wire [1:0] simp271_0;
  wire [1:0] simp281_0;
  wire [1:0] simp291_0;
  wire [1:0] simp301_0;
  wire [1:0] simp311_0;
  wire [1:0] simp321_0;
  wire [1:0] simp331_0;
  wire [1:0] simp341_0;
  wire [1:0] simp351_0;
  wire [1:0] simp361_0;
  wire [1:0] simp371_0;
  wire [1:0] simp381_0;
  wire [1:0] simp391_0;
  wire [1:0] simp401_0;
  wire [1:0] simp411_0;
  wire [1:0] simp421_0;
  wire [1:0] simp431_0;
  wire [1:0] simp441_0;
  wire [1:0] simp451_0;
  wire [1:0] simp461_0;
  wire [1:0] simp471_0;
  wire [1:0] simp481_0;
  wire [1:0] simp491_0;
  wire [1:0] simp501_0;
  wire [1:0] simp511_0;
  wire [1:0] simp521_0;
  wire [1:0] simp531_0;
  wire [1:0] simp541_0;
  wire [1:0] simp551_0;
  wire [1:0] simp561_0;
  wire [1:0] simp571_0;
  wire [1:0] simp581_0;
  wire [1:0] simp591_0;
  wire [1:0] simp601_0;
  wire [1:0] simp611_0;
  wire [1:0] simp621_0;
  wire [1:0] simp631_0;
  wire [1:0] simp641_0;
  wire [1:0] simp651_0;
  wire [1:0] simp661_0;
  wire [1:0] simp671_0;
  wire [1:0] simp681_0;
  wire [1:0] simp691_0;
  wire [1:0] simp701_0;
  wire [1:0] simp711_0;
  wire [1:0] simp721_0;
  wire [1:0] simp731_0;
  wire [1:0] simp741_0;
  wire [1:0] simp751_0;
  wire [1:0] simp761_0;
  wire [1:0] simp771_0;
  wire [1:0] simp781_0;
  wire [1:0] simp791_0;
  wire [1:0] simp801_0;
  wire [1:0] simp811_0;
  wire [1:0] simp821_0;
  wire [1:0] simp831_0;
  wire [32:0] comp0_0;
  wire [10:0] simp3821_0;
  wire [3:0] simp3822_0;
  wire [1:0] simp3823_0;
  wire [32:0] comp1_0;
  wire [10:0] simp4171_0;
  wire [3:0] simp4172_0;
  wire [1:0] simp4173_0;
  wire [32:0] comp2_0;
  wire [10:0] simp4521_0;
  wire [3:0] simp4522_0;
  wire [1:0] simp4523_0;
  wire [32:0] comp3_0;
  wire [10:0] simp4871_0;
  wire [3:0] simp4872_0;
  wire [1:0] simp4873_0;
  wire [1:0] simp4921_0;
  NOR3 I0 (simp181_0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  INV I1 (simp181_0[1:1], gfint_3[0:0]);
  NAND2 I2 (o_0r0[0:0], simp181_0[0:0], simp181_0[1:1]);
  NOR3 I3 (simp191_0[0:0], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  INV I4 (simp191_0[1:1], gfint_3[1:1]);
  NAND2 I5 (o_0r0[1:1], simp191_0[0:0], simp191_0[1:1]);
  NOR3 I6 (simp201_0[0:0], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  INV I7 (simp201_0[1:1], gfint_3[2:2]);
  NAND2 I8 (o_0r0[2:2], simp201_0[0:0], simp201_0[1:1]);
  NOR3 I9 (simp211_0[0:0], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  INV I10 (simp211_0[1:1], gfint_3[3:3]);
  NAND2 I11 (o_0r0[3:3], simp211_0[0:0], simp211_0[1:1]);
  NOR3 I12 (simp221_0[0:0], gfint_0[4:4], gfint_1[4:4], gfint_2[4:4]);
  INV I13 (simp221_0[1:1], gfint_3[4:4]);
  NAND2 I14 (o_0r0[4:4], simp221_0[0:0], simp221_0[1:1]);
  NOR3 I15 (simp231_0[0:0], gfint_0[5:5], gfint_1[5:5], gfint_2[5:5]);
  INV I16 (simp231_0[1:1], gfint_3[5:5]);
  NAND2 I17 (o_0r0[5:5], simp231_0[0:0], simp231_0[1:1]);
  NOR3 I18 (simp241_0[0:0], gfint_0[6:6], gfint_1[6:6], gfint_2[6:6]);
  INV I19 (simp241_0[1:1], gfint_3[6:6]);
  NAND2 I20 (o_0r0[6:6], simp241_0[0:0], simp241_0[1:1]);
  NOR3 I21 (simp251_0[0:0], gfint_0[7:7], gfint_1[7:7], gfint_2[7:7]);
  INV I22 (simp251_0[1:1], gfint_3[7:7]);
  NAND2 I23 (o_0r0[7:7], simp251_0[0:0], simp251_0[1:1]);
  NOR3 I24 (simp261_0[0:0], gfint_0[8:8], gfint_1[8:8], gfint_2[8:8]);
  INV I25 (simp261_0[1:1], gfint_3[8:8]);
  NAND2 I26 (o_0r0[8:8], simp261_0[0:0], simp261_0[1:1]);
  NOR3 I27 (simp271_0[0:0], gfint_0[9:9], gfint_1[9:9], gfint_2[9:9]);
  INV I28 (simp271_0[1:1], gfint_3[9:9]);
  NAND2 I29 (o_0r0[9:9], simp271_0[0:0], simp271_0[1:1]);
  NOR3 I30 (simp281_0[0:0], gfint_0[10:10], gfint_1[10:10], gfint_2[10:10]);
  INV I31 (simp281_0[1:1], gfint_3[10:10]);
  NAND2 I32 (o_0r0[10:10], simp281_0[0:0], simp281_0[1:1]);
  NOR3 I33 (simp291_0[0:0], gfint_0[11:11], gfint_1[11:11], gfint_2[11:11]);
  INV I34 (simp291_0[1:1], gfint_3[11:11]);
  NAND2 I35 (o_0r0[11:11], simp291_0[0:0], simp291_0[1:1]);
  NOR3 I36 (simp301_0[0:0], gfint_0[12:12], gfint_1[12:12], gfint_2[12:12]);
  INV I37 (simp301_0[1:1], gfint_3[12:12]);
  NAND2 I38 (o_0r0[12:12], simp301_0[0:0], simp301_0[1:1]);
  NOR3 I39 (simp311_0[0:0], gfint_0[13:13], gfint_1[13:13], gfint_2[13:13]);
  INV I40 (simp311_0[1:1], gfint_3[13:13]);
  NAND2 I41 (o_0r0[13:13], simp311_0[0:0], simp311_0[1:1]);
  NOR3 I42 (simp321_0[0:0], gfint_0[14:14], gfint_1[14:14], gfint_2[14:14]);
  INV I43 (simp321_0[1:1], gfint_3[14:14]);
  NAND2 I44 (o_0r0[14:14], simp321_0[0:0], simp321_0[1:1]);
  NOR3 I45 (simp331_0[0:0], gfint_0[15:15], gfint_1[15:15], gfint_2[15:15]);
  INV I46 (simp331_0[1:1], gfint_3[15:15]);
  NAND2 I47 (o_0r0[15:15], simp331_0[0:0], simp331_0[1:1]);
  NOR3 I48 (simp341_0[0:0], gfint_0[16:16], gfint_1[16:16], gfint_2[16:16]);
  INV I49 (simp341_0[1:1], gfint_3[16:16]);
  NAND2 I50 (o_0r0[16:16], simp341_0[0:0], simp341_0[1:1]);
  NOR3 I51 (simp351_0[0:0], gfint_0[17:17], gfint_1[17:17], gfint_2[17:17]);
  INV I52 (simp351_0[1:1], gfint_3[17:17]);
  NAND2 I53 (o_0r0[17:17], simp351_0[0:0], simp351_0[1:1]);
  NOR3 I54 (simp361_0[0:0], gfint_0[18:18], gfint_1[18:18], gfint_2[18:18]);
  INV I55 (simp361_0[1:1], gfint_3[18:18]);
  NAND2 I56 (o_0r0[18:18], simp361_0[0:0], simp361_0[1:1]);
  NOR3 I57 (simp371_0[0:0], gfint_0[19:19], gfint_1[19:19], gfint_2[19:19]);
  INV I58 (simp371_0[1:1], gfint_3[19:19]);
  NAND2 I59 (o_0r0[19:19], simp371_0[0:0], simp371_0[1:1]);
  NOR3 I60 (simp381_0[0:0], gfint_0[20:20], gfint_1[20:20], gfint_2[20:20]);
  INV I61 (simp381_0[1:1], gfint_3[20:20]);
  NAND2 I62 (o_0r0[20:20], simp381_0[0:0], simp381_0[1:1]);
  NOR3 I63 (simp391_0[0:0], gfint_0[21:21], gfint_1[21:21], gfint_2[21:21]);
  INV I64 (simp391_0[1:1], gfint_3[21:21]);
  NAND2 I65 (o_0r0[21:21], simp391_0[0:0], simp391_0[1:1]);
  NOR3 I66 (simp401_0[0:0], gfint_0[22:22], gfint_1[22:22], gfint_2[22:22]);
  INV I67 (simp401_0[1:1], gfint_3[22:22]);
  NAND2 I68 (o_0r0[22:22], simp401_0[0:0], simp401_0[1:1]);
  NOR3 I69 (simp411_0[0:0], gfint_0[23:23], gfint_1[23:23], gfint_2[23:23]);
  INV I70 (simp411_0[1:1], gfint_3[23:23]);
  NAND2 I71 (o_0r0[23:23], simp411_0[0:0], simp411_0[1:1]);
  NOR3 I72 (simp421_0[0:0], gfint_0[24:24], gfint_1[24:24], gfint_2[24:24]);
  INV I73 (simp421_0[1:1], gfint_3[24:24]);
  NAND2 I74 (o_0r0[24:24], simp421_0[0:0], simp421_0[1:1]);
  NOR3 I75 (simp431_0[0:0], gfint_0[25:25], gfint_1[25:25], gfint_2[25:25]);
  INV I76 (simp431_0[1:1], gfint_3[25:25]);
  NAND2 I77 (o_0r0[25:25], simp431_0[0:0], simp431_0[1:1]);
  NOR3 I78 (simp441_0[0:0], gfint_0[26:26], gfint_1[26:26], gfint_2[26:26]);
  INV I79 (simp441_0[1:1], gfint_3[26:26]);
  NAND2 I80 (o_0r0[26:26], simp441_0[0:0], simp441_0[1:1]);
  NOR3 I81 (simp451_0[0:0], gfint_0[27:27], gfint_1[27:27], gfint_2[27:27]);
  INV I82 (simp451_0[1:1], gfint_3[27:27]);
  NAND2 I83 (o_0r0[27:27], simp451_0[0:0], simp451_0[1:1]);
  NOR3 I84 (simp461_0[0:0], gfint_0[28:28], gfint_1[28:28], gfint_2[28:28]);
  INV I85 (simp461_0[1:1], gfint_3[28:28]);
  NAND2 I86 (o_0r0[28:28], simp461_0[0:0], simp461_0[1:1]);
  NOR3 I87 (simp471_0[0:0], gfint_0[29:29], gfint_1[29:29], gfint_2[29:29]);
  INV I88 (simp471_0[1:1], gfint_3[29:29]);
  NAND2 I89 (o_0r0[29:29], simp471_0[0:0], simp471_0[1:1]);
  NOR3 I90 (simp481_0[0:0], gfint_0[30:30], gfint_1[30:30], gfint_2[30:30]);
  INV I91 (simp481_0[1:1], gfint_3[30:30]);
  NAND2 I92 (o_0r0[30:30], simp481_0[0:0], simp481_0[1:1]);
  NOR3 I93 (simp491_0[0:0], gfint_0[31:31], gfint_1[31:31], gfint_2[31:31]);
  INV I94 (simp491_0[1:1], gfint_3[31:31]);
  NAND2 I95 (o_0r0[31:31], simp491_0[0:0], simp491_0[1:1]);
  NOR3 I96 (simp501_0[0:0], gfint_0[32:32], gfint_1[32:32], gfint_2[32:32]);
  INV I97 (simp501_0[1:1], gfint_3[32:32]);
  NAND2 I98 (o_0r0[32:32], simp501_0[0:0], simp501_0[1:1]);
  NOR3 I99 (simp511_0[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  INV I100 (simp511_0[1:1], gtint_3[0:0]);
  NAND2 I101 (o_0r1[0:0], simp511_0[0:0], simp511_0[1:1]);
  NOR3 I102 (simp521_0[0:0], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  INV I103 (simp521_0[1:1], gtint_3[1:1]);
  NAND2 I104 (o_0r1[1:1], simp521_0[0:0], simp521_0[1:1]);
  NOR3 I105 (simp531_0[0:0], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  INV I106 (simp531_0[1:1], gtint_3[2:2]);
  NAND2 I107 (o_0r1[2:2], simp531_0[0:0], simp531_0[1:1]);
  NOR3 I108 (simp541_0[0:0], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  INV I109 (simp541_0[1:1], gtint_3[3:3]);
  NAND2 I110 (o_0r1[3:3], simp541_0[0:0], simp541_0[1:1]);
  NOR3 I111 (simp551_0[0:0], gtint_0[4:4], gtint_1[4:4], gtint_2[4:4]);
  INV I112 (simp551_0[1:1], gtint_3[4:4]);
  NAND2 I113 (o_0r1[4:4], simp551_0[0:0], simp551_0[1:1]);
  NOR3 I114 (simp561_0[0:0], gtint_0[5:5], gtint_1[5:5], gtint_2[5:5]);
  INV I115 (simp561_0[1:1], gtint_3[5:5]);
  NAND2 I116 (o_0r1[5:5], simp561_0[0:0], simp561_0[1:1]);
  NOR3 I117 (simp571_0[0:0], gtint_0[6:6], gtint_1[6:6], gtint_2[6:6]);
  INV I118 (simp571_0[1:1], gtint_3[6:6]);
  NAND2 I119 (o_0r1[6:6], simp571_0[0:0], simp571_0[1:1]);
  NOR3 I120 (simp581_0[0:0], gtint_0[7:7], gtint_1[7:7], gtint_2[7:7]);
  INV I121 (simp581_0[1:1], gtint_3[7:7]);
  NAND2 I122 (o_0r1[7:7], simp581_0[0:0], simp581_0[1:1]);
  NOR3 I123 (simp591_0[0:0], gtint_0[8:8], gtint_1[8:8], gtint_2[8:8]);
  INV I124 (simp591_0[1:1], gtint_3[8:8]);
  NAND2 I125 (o_0r1[8:8], simp591_0[0:0], simp591_0[1:1]);
  NOR3 I126 (simp601_0[0:0], gtint_0[9:9], gtint_1[9:9], gtint_2[9:9]);
  INV I127 (simp601_0[1:1], gtint_3[9:9]);
  NAND2 I128 (o_0r1[9:9], simp601_0[0:0], simp601_0[1:1]);
  NOR3 I129 (simp611_0[0:0], gtint_0[10:10], gtint_1[10:10], gtint_2[10:10]);
  INV I130 (simp611_0[1:1], gtint_3[10:10]);
  NAND2 I131 (o_0r1[10:10], simp611_0[0:0], simp611_0[1:1]);
  NOR3 I132 (simp621_0[0:0], gtint_0[11:11], gtint_1[11:11], gtint_2[11:11]);
  INV I133 (simp621_0[1:1], gtint_3[11:11]);
  NAND2 I134 (o_0r1[11:11], simp621_0[0:0], simp621_0[1:1]);
  NOR3 I135 (simp631_0[0:0], gtint_0[12:12], gtint_1[12:12], gtint_2[12:12]);
  INV I136 (simp631_0[1:1], gtint_3[12:12]);
  NAND2 I137 (o_0r1[12:12], simp631_0[0:0], simp631_0[1:1]);
  NOR3 I138 (simp641_0[0:0], gtint_0[13:13], gtint_1[13:13], gtint_2[13:13]);
  INV I139 (simp641_0[1:1], gtint_3[13:13]);
  NAND2 I140 (o_0r1[13:13], simp641_0[0:0], simp641_0[1:1]);
  NOR3 I141 (simp651_0[0:0], gtint_0[14:14], gtint_1[14:14], gtint_2[14:14]);
  INV I142 (simp651_0[1:1], gtint_3[14:14]);
  NAND2 I143 (o_0r1[14:14], simp651_0[0:0], simp651_0[1:1]);
  NOR3 I144 (simp661_0[0:0], gtint_0[15:15], gtint_1[15:15], gtint_2[15:15]);
  INV I145 (simp661_0[1:1], gtint_3[15:15]);
  NAND2 I146 (o_0r1[15:15], simp661_0[0:0], simp661_0[1:1]);
  NOR3 I147 (simp671_0[0:0], gtint_0[16:16], gtint_1[16:16], gtint_2[16:16]);
  INV I148 (simp671_0[1:1], gtint_3[16:16]);
  NAND2 I149 (o_0r1[16:16], simp671_0[0:0], simp671_0[1:1]);
  NOR3 I150 (simp681_0[0:0], gtint_0[17:17], gtint_1[17:17], gtint_2[17:17]);
  INV I151 (simp681_0[1:1], gtint_3[17:17]);
  NAND2 I152 (o_0r1[17:17], simp681_0[0:0], simp681_0[1:1]);
  NOR3 I153 (simp691_0[0:0], gtint_0[18:18], gtint_1[18:18], gtint_2[18:18]);
  INV I154 (simp691_0[1:1], gtint_3[18:18]);
  NAND2 I155 (o_0r1[18:18], simp691_0[0:0], simp691_0[1:1]);
  NOR3 I156 (simp701_0[0:0], gtint_0[19:19], gtint_1[19:19], gtint_2[19:19]);
  INV I157 (simp701_0[1:1], gtint_3[19:19]);
  NAND2 I158 (o_0r1[19:19], simp701_0[0:0], simp701_0[1:1]);
  NOR3 I159 (simp711_0[0:0], gtint_0[20:20], gtint_1[20:20], gtint_2[20:20]);
  INV I160 (simp711_0[1:1], gtint_3[20:20]);
  NAND2 I161 (o_0r1[20:20], simp711_0[0:0], simp711_0[1:1]);
  NOR3 I162 (simp721_0[0:0], gtint_0[21:21], gtint_1[21:21], gtint_2[21:21]);
  INV I163 (simp721_0[1:1], gtint_3[21:21]);
  NAND2 I164 (o_0r1[21:21], simp721_0[0:0], simp721_0[1:1]);
  NOR3 I165 (simp731_0[0:0], gtint_0[22:22], gtint_1[22:22], gtint_2[22:22]);
  INV I166 (simp731_0[1:1], gtint_3[22:22]);
  NAND2 I167 (o_0r1[22:22], simp731_0[0:0], simp731_0[1:1]);
  NOR3 I168 (simp741_0[0:0], gtint_0[23:23], gtint_1[23:23], gtint_2[23:23]);
  INV I169 (simp741_0[1:1], gtint_3[23:23]);
  NAND2 I170 (o_0r1[23:23], simp741_0[0:0], simp741_0[1:1]);
  NOR3 I171 (simp751_0[0:0], gtint_0[24:24], gtint_1[24:24], gtint_2[24:24]);
  INV I172 (simp751_0[1:1], gtint_3[24:24]);
  NAND2 I173 (o_0r1[24:24], simp751_0[0:0], simp751_0[1:1]);
  NOR3 I174 (simp761_0[0:0], gtint_0[25:25], gtint_1[25:25], gtint_2[25:25]);
  INV I175 (simp761_0[1:1], gtint_3[25:25]);
  NAND2 I176 (o_0r1[25:25], simp761_0[0:0], simp761_0[1:1]);
  NOR3 I177 (simp771_0[0:0], gtint_0[26:26], gtint_1[26:26], gtint_2[26:26]);
  INV I178 (simp771_0[1:1], gtint_3[26:26]);
  NAND2 I179 (o_0r1[26:26], simp771_0[0:0], simp771_0[1:1]);
  NOR3 I180 (simp781_0[0:0], gtint_0[27:27], gtint_1[27:27], gtint_2[27:27]);
  INV I181 (simp781_0[1:1], gtint_3[27:27]);
  NAND2 I182 (o_0r1[27:27], simp781_0[0:0], simp781_0[1:1]);
  NOR3 I183 (simp791_0[0:0], gtint_0[28:28], gtint_1[28:28], gtint_2[28:28]);
  INV I184 (simp791_0[1:1], gtint_3[28:28]);
  NAND2 I185 (o_0r1[28:28], simp791_0[0:0], simp791_0[1:1]);
  NOR3 I186 (simp801_0[0:0], gtint_0[29:29], gtint_1[29:29], gtint_2[29:29]);
  INV I187 (simp801_0[1:1], gtint_3[29:29]);
  NAND2 I188 (o_0r1[29:29], simp801_0[0:0], simp801_0[1:1]);
  NOR3 I189 (simp811_0[0:0], gtint_0[30:30], gtint_1[30:30], gtint_2[30:30]);
  INV I190 (simp811_0[1:1], gtint_3[30:30]);
  NAND2 I191 (o_0r1[30:30], simp811_0[0:0], simp811_0[1:1]);
  NOR3 I192 (simp821_0[0:0], gtint_0[31:31], gtint_1[31:31], gtint_2[31:31]);
  INV I193 (simp821_0[1:1], gtint_3[31:31]);
  NAND2 I194 (o_0r1[31:31], simp821_0[0:0], simp821_0[1:1]);
  NOR3 I195 (simp831_0[0:0], gtint_0[32:32], gtint_1[32:32], gtint_2[32:32]);
  INV I196 (simp831_0[1:1], gtint_3[32:32]);
  NAND2 I197 (o_0r1[32:32], simp831_0[0:0], simp831_0[1:1]);
  AND2 I198 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I199 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I200 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I201 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I202 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I203 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I204 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I205 (gtint_0[7:7], choice_0, i_0r1[7:7]);
  AND2 I206 (gtint_0[8:8], choice_0, i_0r1[8:8]);
  AND2 I207 (gtint_0[9:9], choice_0, i_0r1[9:9]);
  AND2 I208 (gtint_0[10:10], choice_0, i_0r1[10:10]);
  AND2 I209 (gtint_0[11:11], choice_0, i_0r1[11:11]);
  AND2 I210 (gtint_0[12:12], choice_0, i_0r1[12:12]);
  AND2 I211 (gtint_0[13:13], choice_0, i_0r1[13:13]);
  AND2 I212 (gtint_0[14:14], choice_0, i_0r1[14:14]);
  AND2 I213 (gtint_0[15:15], choice_0, i_0r1[15:15]);
  AND2 I214 (gtint_0[16:16], choice_0, i_0r1[16:16]);
  AND2 I215 (gtint_0[17:17], choice_0, i_0r1[17:17]);
  AND2 I216 (gtint_0[18:18], choice_0, i_0r1[18:18]);
  AND2 I217 (gtint_0[19:19], choice_0, i_0r1[19:19]);
  AND2 I218 (gtint_0[20:20], choice_0, i_0r1[20:20]);
  AND2 I219 (gtint_0[21:21], choice_0, i_0r1[21:21]);
  AND2 I220 (gtint_0[22:22], choice_0, i_0r1[22:22]);
  AND2 I221 (gtint_0[23:23], choice_0, i_0r1[23:23]);
  AND2 I222 (gtint_0[24:24], choice_0, i_0r1[24:24]);
  AND2 I223 (gtint_0[25:25], choice_0, i_0r1[25:25]);
  AND2 I224 (gtint_0[26:26], choice_0, i_0r1[26:26]);
  AND2 I225 (gtint_0[27:27], choice_0, i_0r1[27:27]);
  AND2 I226 (gtint_0[28:28], choice_0, i_0r1[28:28]);
  AND2 I227 (gtint_0[29:29], choice_0, i_0r1[29:29]);
  AND2 I228 (gtint_0[30:30], choice_0, i_0r1[30:30]);
  AND2 I229 (gtint_0[31:31], choice_0, i_0r1[31:31]);
  AND2 I230 (gtint_0[32:32], choice_0, i_0r1[32:32]);
  AND2 I231 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I232 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I233 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I234 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I235 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I236 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I237 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I238 (gtint_1[7:7], choice_1, i_1r1[7:7]);
  AND2 I239 (gtint_1[8:8], choice_1, i_1r1[8:8]);
  AND2 I240 (gtint_1[9:9], choice_1, i_1r1[9:9]);
  AND2 I241 (gtint_1[10:10], choice_1, i_1r1[10:10]);
  AND2 I242 (gtint_1[11:11], choice_1, i_1r1[11:11]);
  AND2 I243 (gtint_1[12:12], choice_1, i_1r1[12:12]);
  AND2 I244 (gtint_1[13:13], choice_1, i_1r1[13:13]);
  AND2 I245 (gtint_1[14:14], choice_1, i_1r1[14:14]);
  AND2 I246 (gtint_1[15:15], choice_1, i_1r1[15:15]);
  AND2 I247 (gtint_1[16:16], choice_1, i_1r1[16:16]);
  AND2 I248 (gtint_1[17:17], choice_1, i_1r1[17:17]);
  AND2 I249 (gtint_1[18:18], choice_1, i_1r1[18:18]);
  AND2 I250 (gtint_1[19:19], choice_1, i_1r1[19:19]);
  AND2 I251 (gtint_1[20:20], choice_1, i_1r1[20:20]);
  AND2 I252 (gtint_1[21:21], choice_1, i_1r1[21:21]);
  AND2 I253 (gtint_1[22:22], choice_1, i_1r1[22:22]);
  AND2 I254 (gtint_1[23:23], choice_1, i_1r1[23:23]);
  AND2 I255 (gtint_1[24:24], choice_1, i_1r1[24:24]);
  AND2 I256 (gtint_1[25:25], choice_1, i_1r1[25:25]);
  AND2 I257 (gtint_1[26:26], choice_1, i_1r1[26:26]);
  AND2 I258 (gtint_1[27:27], choice_1, i_1r1[27:27]);
  AND2 I259 (gtint_1[28:28], choice_1, i_1r1[28:28]);
  AND2 I260 (gtint_1[29:29], choice_1, i_1r1[29:29]);
  AND2 I261 (gtint_1[30:30], choice_1, i_1r1[30:30]);
  AND2 I262 (gtint_1[31:31], choice_1, i_1r1[31:31]);
  AND2 I263 (gtint_1[32:32], choice_1, i_1r1[32:32]);
  AND2 I264 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I265 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I266 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I267 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AND2 I268 (gtint_2[4:4], choice_2, i_2r1[4:4]);
  AND2 I269 (gtint_2[5:5], choice_2, i_2r1[5:5]);
  AND2 I270 (gtint_2[6:6], choice_2, i_2r1[6:6]);
  AND2 I271 (gtint_2[7:7], choice_2, i_2r1[7:7]);
  AND2 I272 (gtint_2[8:8], choice_2, i_2r1[8:8]);
  AND2 I273 (gtint_2[9:9], choice_2, i_2r1[9:9]);
  AND2 I274 (gtint_2[10:10], choice_2, i_2r1[10:10]);
  AND2 I275 (gtint_2[11:11], choice_2, i_2r1[11:11]);
  AND2 I276 (gtint_2[12:12], choice_2, i_2r1[12:12]);
  AND2 I277 (gtint_2[13:13], choice_2, i_2r1[13:13]);
  AND2 I278 (gtint_2[14:14], choice_2, i_2r1[14:14]);
  AND2 I279 (gtint_2[15:15], choice_2, i_2r1[15:15]);
  AND2 I280 (gtint_2[16:16], choice_2, i_2r1[16:16]);
  AND2 I281 (gtint_2[17:17], choice_2, i_2r1[17:17]);
  AND2 I282 (gtint_2[18:18], choice_2, i_2r1[18:18]);
  AND2 I283 (gtint_2[19:19], choice_2, i_2r1[19:19]);
  AND2 I284 (gtint_2[20:20], choice_2, i_2r1[20:20]);
  AND2 I285 (gtint_2[21:21], choice_2, i_2r1[21:21]);
  AND2 I286 (gtint_2[22:22], choice_2, i_2r1[22:22]);
  AND2 I287 (gtint_2[23:23], choice_2, i_2r1[23:23]);
  AND2 I288 (gtint_2[24:24], choice_2, i_2r1[24:24]);
  AND2 I289 (gtint_2[25:25], choice_2, i_2r1[25:25]);
  AND2 I290 (gtint_2[26:26], choice_2, i_2r1[26:26]);
  AND2 I291 (gtint_2[27:27], choice_2, i_2r1[27:27]);
  AND2 I292 (gtint_2[28:28], choice_2, i_2r1[28:28]);
  AND2 I293 (gtint_2[29:29], choice_2, i_2r1[29:29]);
  AND2 I294 (gtint_2[30:30], choice_2, i_2r1[30:30]);
  AND2 I295 (gtint_2[31:31], choice_2, i_2r1[31:31]);
  AND2 I296 (gtint_2[32:32], choice_2, i_2r1[32:32]);
  AND2 I297 (gtint_3[0:0], choice_3, i_3r1[0:0]);
  AND2 I298 (gtint_3[1:1], choice_3, i_3r1[1:1]);
  AND2 I299 (gtint_3[2:2], choice_3, i_3r1[2:2]);
  AND2 I300 (gtint_3[3:3], choice_3, i_3r1[3:3]);
  AND2 I301 (gtint_3[4:4], choice_3, i_3r1[4:4]);
  AND2 I302 (gtint_3[5:5], choice_3, i_3r1[5:5]);
  AND2 I303 (gtint_3[6:6], choice_3, i_3r1[6:6]);
  AND2 I304 (gtint_3[7:7], choice_3, i_3r1[7:7]);
  AND2 I305 (gtint_3[8:8], choice_3, i_3r1[8:8]);
  AND2 I306 (gtint_3[9:9], choice_3, i_3r1[9:9]);
  AND2 I307 (gtint_3[10:10], choice_3, i_3r1[10:10]);
  AND2 I308 (gtint_3[11:11], choice_3, i_3r1[11:11]);
  AND2 I309 (gtint_3[12:12], choice_3, i_3r1[12:12]);
  AND2 I310 (gtint_3[13:13], choice_3, i_3r1[13:13]);
  AND2 I311 (gtint_3[14:14], choice_3, i_3r1[14:14]);
  AND2 I312 (gtint_3[15:15], choice_3, i_3r1[15:15]);
  AND2 I313 (gtint_3[16:16], choice_3, i_3r1[16:16]);
  AND2 I314 (gtint_3[17:17], choice_3, i_3r1[17:17]);
  AND2 I315 (gtint_3[18:18], choice_3, i_3r1[18:18]);
  AND2 I316 (gtint_3[19:19], choice_3, i_3r1[19:19]);
  AND2 I317 (gtint_3[20:20], choice_3, i_3r1[20:20]);
  AND2 I318 (gtint_3[21:21], choice_3, i_3r1[21:21]);
  AND2 I319 (gtint_3[22:22], choice_3, i_3r1[22:22]);
  AND2 I320 (gtint_3[23:23], choice_3, i_3r1[23:23]);
  AND2 I321 (gtint_3[24:24], choice_3, i_3r1[24:24]);
  AND2 I322 (gtint_3[25:25], choice_3, i_3r1[25:25]);
  AND2 I323 (gtint_3[26:26], choice_3, i_3r1[26:26]);
  AND2 I324 (gtint_3[27:27], choice_3, i_3r1[27:27]);
  AND2 I325 (gtint_3[28:28], choice_3, i_3r1[28:28]);
  AND2 I326 (gtint_3[29:29], choice_3, i_3r1[29:29]);
  AND2 I327 (gtint_3[30:30], choice_3, i_3r1[30:30]);
  AND2 I328 (gtint_3[31:31], choice_3, i_3r1[31:31]);
  AND2 I329 (gtint_3[32:32], choice_3, i_3r1[32:32]);
  AND2 I330 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I331 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I332 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I333 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I334 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I335 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I336 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I337 (gfint_0[7:7], choice_0, i_0r0[7:7]);
  AND2 I338 (gfint_0[8:8], choice_0, i_0r0[8:8]);
  AND2 I339 (gfint_0[9:9], choice_0, i_0r0[9:9]);
  AND2 I340 (gfint_0[10:10], choice_0, i_0r0[10:10]);
  AND2 I341 (gfint_0[11:11], choice_0, i_0r0[11:11]);
  AND2 I342 (gfint_0[12:12], choice_0, i_0r0[12:12]);
  AND2 I343 (gfint_0[13:13], choice_0, i_0r0[13:13]);
  AND2 I344 (gfint_0[14:14], choice_0, i_0r0[14:14]);
  AND2 I345 (gfint_0[15:15], choice_0, i_0r0[15:15]);
  AND2 I346 (gfint_0[16:16], choice_0, i_0r0[16:16]);
  AND2 I347 (gfint_0[17:17], choice_0, i_0r0[17:17]);
  AND2 I348 (gfint_0[18:18], choice_0, i_0r0[18:18]);
  AND2 I349 (gfint_0[19:19], choice_0, i_0r0[19:19]);
  AND2 I350 (gfint_0[20:20], choice_0, i_0r0[20:20]);
  AND2 I351 (gfint_0[21:21], choice_0, i_0r0[21:21]);
  AND2 I352 (gfint_0[22:22], choice_0, i_0r0[22:22]);
  AND2 I353 (gfint_0[23:23], choice_0, i_0r0[23:23]);
  AND2 I354 (gfint_0[24:24], choice_0, i_0r0[24:24]);
  AND2 I355 (gfint_0[25:25], choice_0, i_0r0[25:25]);
  AND2 I356 (gfint_0[26:26], choice_0, i_0r0[26:26]);
  AND2 I357 (gfint_0[27:27], choice_0, i_0r0[27:27]);
  AND2 I358 (gfint_0[28:28], choice_0, i_0r0[28:28]);
  AND2 I359 (gfint_0[29:29], choice_0, i_0r0[29:29]);
  AND2 I360 (gfint_0[30:30], choice_0, i_0r0[30:30]);
  AND2 I361 (gfint_0[31:31], choice_0, i_0r0[31:31]);
  AND2 I362 (gfint_0[32:32], choice_0, i_0r0[32:32]);
  AND2 I363 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I364 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I365 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I366 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I367 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I368 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I369 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I370 (gfint_1[7:7], choice_1, i_1r0[7:7]);
  AND2 I371 (gfint_1[8:8], choice_1, i_1r0[8:8]);
  AND2 I372 (gfint_1[9:9], choice_1, i_1r0[9:9]);
  AND2 I373 (gfint_1[10:10], choice_1, i_1r0[10:10]);
  AND2 I374 (gfint_1[11:11], choice_1, i_1r0[11:11]);
  AND2 I375 (gfint_1[12:12], choice_1, i_1r0[12:12]);
  AND2 I376 (gfint_1[13:13], choice_1, i_1r0[13:13]);
  AND2 I377 (gfint_1[14:14], choice_1, i_1r0[14:14]);
  AND2 I378 (gfint_1[15:15], choice_1, i_1r0[15:15]);
  AND2 I379 (gfint_1[16:16], choice_1, i_1r0[16:16]);
  AND2 I380 (gfint_1[17:17], choice_1, i_1r0[17:17]);
  AND2 I381 (gfint_1[18:18], choice_1, i_1r0[18:18]);
  AND2 I382 (gfint_1[19:19], choice_1, i_1r0[19:19]);
  AND2 I383 (gfint_1[20:20], choice_1, i_1r0[20:20]);
  AND2 I384 (gfint_1[21:21], choice_1, i_1r0[21:21]);
  AND2 I385 (gfint_1[22:22], choice_1, i_1r0[22:22]);
  AND2 I386 (gfint_1[23:23], choice_1, i_1r0[23:23]);
  AND2 I387 (gfint_1[24:24], choice_1, i_1r0[24:24]);
  AND2 I388 (gfint_1[25:25], choice_1, i_1r0[25:25]);
  AND2 I389 (gfint_1[26:26], choice_1, i_1r0[26:26]);
  AND2 I390 (gfint_1[27:27], choice_1, i_1r0[27:27]);
  AND2 I391 (gfint_1[28:28], choice_1, i_1r0[28:28]);
  AND2 I392 (gfint_1[29:29], choice_1, i_1r0[29:29]);
  AND2 I393 (gfint_1[30:30], choice_1, i_1r0[30:30]);
  AND2 I394 (gfint_1[31:31], choice_1, i_1r0[31:31]);
  AND2 I395 (gfint_1[32:32], choice_1, i_1r0[32:32]);
  AND2 I396 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I397 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I398 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I399 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AND2 I400 (gfint_2[4:4], choice_2, i_2r0[4:4]);
  AND2 I401 (gfint_2[5:5], choice_2, i_2r0[5:5]);
  AND2 I402 (gfint_2[6:6], choice_2, i_2r0[6:6]);
  AND2 I403 (gfint_2[7:7], choice_2, i_2r0[7:7]);
  AND2 I404 (gfint_2[8:8], choice_2, i_2r0[8:8]);
  AND2 I405 (gfint_2[9:9], choice_2, i_2r0[9:9]);
  AND2 I406 (gfint_2[10:10], choice_2, i_2r0[10:10]);
  AND2 I407 (gfint_2[11:11], choice_2, i_2r0[11:11]);
  AND2 I408 (gfint_2[12:12], choice_2, i_2r0[12:12]);
  AND2 I409 (gfint_2[13:13], choice_2, i_2r0[13:13]);
  AND2 I410 (gfint_2[14:14], choice_2, i_2r0[14:14]);
  AND2 I411 (gfint_2[15:15], choice_2, i_2r0[15:15]);
  AND2 I412 (gfint_2[16:16], choice_2, i_2r0[16:16]);
  AND2 I413 (gfint_2[17:17], choice_2, i_2r0[17:17]);
  AND2 I414 (gfint_2[18:18], choice_2, i_2r0[18:18]);
  AND2 I415 (gfint_2[19:19], choice_2, i_2r0[19:19]);
  AND2 I416 (gfint_2[20:20], choice_2, i_2r0[20:20]);
  AND2 I417 (gfint_2[21:21], choice_2, i_2r0[21:21]);
  AND2 I418 (gfint_2[22:22], choice_2, i_2r0[22:22]);
  AND2 I419 (gfint_2[23:23], choice_2, i_2r0[23:23]);
  AND2 I420 (gfint_2[24:24], choice_2, i_2r0[24:24]);
  AND2 I421 (gfint_2[25:25], choice_2, i_2r0[25:25]);
  AND2 I422 (gfint_2[26:26], choice_2, i_2r0[26:26]);
  AND2 I423 (gfint_2[27:27], choice_2, i_2r0[27:27]);
  AND2 I424 (gfint_2[28:28], choice_2, i_2r0[28:28]);
  AND2 I425 (gfint_2[29:29], choice_2, i_2r0[29:29]);
  AND2 I426 (gfint_2[30:30], choice_2, i_2r0[30:30]);
  AND2 I427 (gfint_2[31:31], choice_2, i_2r0[31:31]);
  AND2 I428 (gfint_2[32:32], choice_2, i_2r0[32:32]);
  AND2 I429 (gfint_3[0:0], choice_3, i_3r0[0:0]);
  AND2 I430 (gfint_3[1:1], choice_3, i_3r0[1:1]);
  AND2 I431 (gfint_3[2:2], choice_3, i_3r0[2:2]);
  AND2 I432 (gfint_3[3:3], choice_3, i_3r0[3:3]);
  AND2 I433 (gfint_3[4:4], choice_3, i_3r0[4:4]);
  AND2 I434 (gfint_3[5:5], choice_3, i_3r0[5:5]);
  AND2 I435 (gfint_3[6:6], choice_3, i_3r0[6:6]);
  AND2 I436 (gfint_3[7:7], choice_3, i_3r0[7:7]);
  AND2 I437 (gfint_3[8:8], choice_3, i_3r0[8:8]);
  AND2 I438 (gfint_3[9:9], choice_3, i_3r0[9:9]);
  AND2 I439 (gfint_3[10:10], choice_3, i_3r0[10:10]);
  AND2 I440 (gfint_3[11:11], choice_3, i_3r0[11:11]);
  AND2 I441 (gfint_3[12:12], choice_3, i_3r0[12:12]);
  AND2 I442 (gfint_3[13:13], choice_3, i_3r0[13:13]);
  AND2 I443 (gfint_3[14:14], choice_3, i_3r0[14:14]);
  AND2 I444 (gfint_3[15:15], choice_3, i_3r0[15:15]);
  AND2 I445 (gfint_3[16:16], choice_3, i_3r0[16:16]);
  AND2 I446 (gfint_3[17:17], choice_3, i_3r0[17:17]);
  AND2 I447 (gfint_3[18:18], choice_3, i_3r0[18:18]);
  AND2 I448 (gfint_3[19:19], choice_3, i_3r0[19:19]);
  AND2 I449 (gfint_3[20:20], choice_3, i_3r0[20:20]);
  AND2 I450 (gfint_3[21:21], choice_3, i_3r0[21:21]);
  AND2 I451 (gfint_3[22:22], choice_3, i_3r0[22:22]);
  AND2 I452 (gfint_3[23:23], choice_3, i_3r0[23:23]);
  AND2 I453 (gfint_3[24:24], choice_3, i_3r0[24:24]);
  AND2 I454 (gfint_3[25:25], choice_3, i_3r0[25:25]);
  AND2 I455 (gfint_3[26:26], choice_3, i_3r0[26:26]);
  AND2 I456 (gfint_3[27:27], choice_3, i_3r0[27:27]);
  AND2 I457 (gfint_3[28:28], choice_3, i_3r0[28:28]);
  AND2 I458 (gfint_3[29:29], choice_3, i_3r0[29:29]);
  AND2 I459 (gfint_3[30:30], choice_3, i_3r0[30:30]);
  AND2 I460 (gfint_3[31:31], choice_3, i_3r0[31:31]);
  AND2 I461 (gfint_3[32:32], choice_3, i_3r0[32:32]);
  OR2 I462 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I463 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I464 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I465 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I466 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I467 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I468 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I469 (comp0_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I470 (comp0_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I471 (comp0_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I472 (comp0_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I473 (comp0_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I474 (comp0_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I475 (comp0_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I476 (comp0_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I477 (comp0_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I478 (comp0_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I479 (comp0_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I480 (comp0_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I481 (comp0_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I482 (comp0_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I483 (comp0_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I484 (comp0_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I485 (comp0_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I486 (comp0_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I487 (comp0_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I488 (comp0_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I489 (comp0_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I490 (comp0_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I491 (comp0_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I492 (comp0_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I493 (comp0_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I494 (comp0_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  C3 I495 (simp3821_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I496 (simp3821_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I497 (simp3821_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I498 (simp3821_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I499 (simp3821_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I500 (simp3821_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I501 (simp3821_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I502 (simp3821_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I503 (simp3821_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I504 (simp3821_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C3 I505 (simp3821_0[10:10], comp0_0[30:30], comp0_0[31:31], comp0_0[32:32]);
  C3 I506 (simp3822_0[0:0], simp3821_0[0:0], simp3821_0[1:1], simp3821_0[2:2]);
  C3 I507 (simp3822_0[1:1], simp3821_0[3:3], simp3821_0[4:4], simp3821_0[5:5]);
  C3 I508 (simp3822_0[2:2], simp3821_0[6:6], simp3821_0[7:7], simp3821_0[8:8]);
  C2 I509 (simp3822_0[3:3], simp3821_0[9:9], simp3821_0[10:10]);
  C3 I510 (simp3823_0[0:0], simp3822_0[0:0], simp3822_0[1:1], simp3822_0[2:2]);
  BUFF I511 (simp3823_0[1:1], simp3822_0[3:3]);
  C2 I512 (icomp_0, simp3823_0[0:0], simp3823_0[1:1]);
  OR2 I513 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I514 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I515 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I516 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I517 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I518 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I519 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  OR2 I520 (comp1_0[7:7], i_1r0[7:7], i_1r1[7:7]);
  OR2 I521 (comp1_0[8:8], i_1r0[8:8], i_1r1[8:8]);
  OR2 I522 (comp1_0[9:9], i_1r0[9:9], i_1r1[9:9]);
  OR2 I523 (comp1_0[10:10], i_1r0[10:10], i_1r1[10:10]);
  OR2 I524 (comp1_0[11:11], i_1r0[11:11], i_1r1[11:11]);
  OR2 I525 (comp1_0[12:12], i_1r0[12:12], i_1r1[12:12]);
  OR2 I526 (comp1_0[13:13], i_1r0[13:13], i_1r1[13:13]);
  OR2 I527 (comp1_0[14:14], i_1r0[14:14], i_1r1[14:14]);
  OR2 I528 (comp1_0[15:15], i_1r0[15:15], i_1r1[15:15]);
  OR2 I529 (comp1_0[16:16], i_1r0[16:16], i_1r1[16:16]);
  OR2 I530 (comp1_0[17:17], i_1r0[17:17], i_1r1[17:17]);
  OR2 I531 (comp1_0[18:18], i_1r0[18:18], i_1r1[18:18]);
  OR2 I532 (comp1_0[19:19], i_1r0[19:19], i_1r1[19:19]);
  OR2 I533 (comp1_0[20:20], i_1r0[20:20], i_1r1[20:20]);
  OR2 I534 (comp1_0[21:21], i_1r0[21:21], i_1r1[21:21]);
  OR2 I535 (comp1_0[22:22], i_1r0[22:22], i_1r1[22:22]);
  OR2 I536 (comp1_0[23:23], i_1r0[23:23], i_1r1[23:23]);
  OR2 I537 (comp1_0[24:24], i_1r0[24:24], i_1r1[24:24]);
  OR2 I538 (comp1_0[25:25], i_1r0[25:25], i_1r1[25:25]);
  OR2 I539 (comp1_0[26:26], i_1r0[26:26], i_1r1[26:26]);
  OR2 I540 (comp1_0[27:27], i_1r0[27:27], i_1r1[27:27]);
  OR2 I541 (comp1_0[28:28], i_1r0[28:28], i_1r1[28:28]);
  OR2 I542 (comp1_0[29:29], i_1r0[29:29], i_1r1[29:29]);
  OR2 I543 (comp1_0[30:30], i_1r0[30:30], i_1r1[30:30]);
  OR2 I544 (comp1_0[31:31], i_1r0[31:31], i_1r1[31:31]);
  OR2 I545 (comp1_0[32:32], i_1r0[32:32], i_1r1[32:32]);
  C3 I546 (simp4171_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I547 (simp4171_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  C3 I548 (simp4171_0[2:2], comp1_0[6:6], comp1_0[7:7], comp1_0[8:8]);
  C3 I549 (simp4171_0[3:3], comp1_0[9:9], comp1_0[10:10], comp1_0[11:11]);
  C3 I550 (simp4171_0[4:4], comp1_0[12:12], comp1_0[13:13], comp1_0[14:14]);
  C3 I551 (simp4171_0[5:5], comp1_0[15:15], comp1_0[16:16], comp1_0[17:17]);
  C3 I552 (simp4171_0[6:6], comp1_0[18:18], comp1_0[19:19], comp1_0[20:20]);
  C3 I553 (simp4171_0[7:7], comp1_0[21:21], comp1_0[22:22], comp1_0[23:23]);
  C3 I554 (simp4171_0[8:8], comp1_0[24:24], comp1_0[25:25], comp1_0[26:26]);
  C3 I555 (simp4171_0[9:9], comp1_0[27:27], comp1_0[28:28], comp1_0[29:29]);
  C3 I556 (simp4171_0[10:10], comp1_0[30:30], comp1_0[31:31], comp1_0[32:32]);
  C3 I557 (simp4172_0[0:0], simp4171_0[0:0], simp4171_0[1:1], simp4171_0[2:2]);
  C3 I558 (simp4172_0[1:1], simp4171_0[3:3], simp4171_0[4:4], simp4171_0[5:5]);
  C3 I559 (simp4172_0[2:2], simp4171_0[6:6], simp4171_0[7:7], simp4171_0[8:8]);
  C2 I560 (simp4172_0[3:3], simp4171_0[9:9], simp4171_0[10:10]);
  C3 I561 (simp4173_0[0:0], simp4172_0[0:0], simp4172_0[1:1], simp4172_0[2:2]);
  BUFF I562 (simp4173_0[1:1], simp4172_0[3:3]);
  C2 I563 (icomp_1, simp4173_0[0:0], simp4173_0[1:1]);
  OR2 I564 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I565 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I566 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2 I567 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  OR2 I568 (comp2_0[4:4], i_2r0[4:4], i_2r1[4:4]);
  OR2 I569 (comp2_0[5:5], i_2r0[5:5], i_2r1[5:5]);
  OR2 I570 (comp2_0[6:6], i_2r0[6:6], i_2r1[6:6]);
  OR2 I571 (comp2_0[7:7], i_2r0[7:7], i_2r1[7:7]);
  OR2 I572 (comp2_0[8:8], i_2r0[8:8], i_2r1[8:8]);
  OR2 I573 (comp2_0[9:9], i_2r0[9:9], i_2r1[9:9]);
  OR2 I574 (comp2_0[10:10], i_2r0[10:10], i_2r1[10:10]);
  OR2 I575 (comp2_0[11:11], i_2r0[11:11], i_2r1[11:11]);
  OR2 I576 (comp2_0[12:12], i_2r0[12:12], i_2r1[12:12]);
  OR2 I577 (comp2_0[13:13], i_2r0[13:13], i_2r1[13:13]);
  OR2 I578 (comp2_0[14:14], i_2r0[14:14], i_2r1[14:14]);
  OR2 I579 (comp2_0[15:15], i_2r0[15:15], i_2r1[15:15]);
  OR2 I580 (comp2_0[16:16], i_2r0[16:16], i_2r1[16:16]);
  OR2 I581 (comp2_0[17:17], i_2r0[17:17], i_2r1[17:17]);
  OR2 I582 (comp2_0[18:18], i_2r0[18:18], i_2r1[18:18]);
  OR2 I583 (comp2_0[19:19], i_2r0[19:19], i_2r1[19:19]);
  OR2 I584 (comp2_0[20:20], i_2r0[20:20], i_2r1[20:20]);
  OR2 I585 (comp2_0[21:21], i_2r0[21:21], i_2r1[21:21]);
  OR2 I586 (comp2_0[22:22], i_2r0[22:22], i_2r1[22:22]);
  OR2 I587 (comp2_0[23:23], i_2r0[23:23], i_2r1[23:23]);
  OR2 I588 (comp2_0[24:24], i_2r0[24:24], i_2r1[24:24]);
  OR2 I589 (comp2_0[25:25], i_2r0[25:25], i_2r1[25:25]);
  OR2 I590 (comp2_0[26:26], i_2r0[26:26], i_2r1[26:26]);
  OR2 I591 (comp2_0[27:27], i_2r0[27:27], i_2r1[27:27]);
  OR2 I592 (comp2_0[28:28], i_2r0[28:28], i_2r1[28:28]);
  OR2 I593 (comp2_0[29:29], i_2r0[29:29], i_2r1[29:29]);
  OR2 I594 (comp2_0[30:30], i_2r0[30:30], i_2r1[30:30]);
  OR2 I595 (comp2_0[31:31], i_2r0[31:31], i_2r1[31:31]);
  OR2 I596 (comp2_0[32:32], i_2r0[32:32], i_2r1[32:32]);
  C3 I597 (simp4521_0[0:0], comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C3 I598 (simp4521_0[1:1], comp2_0[3:3], comp2_0[4:4], comp2_0[5:5]);
  C3 I599 (simp4521_0[2:2], comp2_0[6:6], comp2_0[7:7], comp2_0[8:8]);
  C3 I600 (simp4521_0[3:3], comp2_0[9:9], comp2_0[10:10], comp2_0[11:11]);
  C3 I601 (simp4521_0[4:4], comp2_0[12:12], comp2_0[13:13], comp2_0[14:14]);
  C3 I602 (simp4521_0[5:5], comp2_0[15:15], comp2_0[16:16], comp2_0[17:17]);
  C3 I603 (simp4521_0[6:6], comp2_0[18:18], comp2_0[19:19], comp2_0[20:20]);
  C3 I604 (simp4521_0[7:7], comp2_0[21:21], comp2_0[22:22], comp2_0[23:23]);
  C3 I605 (simp4521_0[8:8], comp2_0[24:24], comp2_0[25:25], comp2_0[26:26]);
  C3 I606 (simp4521_0[9:9], comp2_0[27:27], comp2_0[28:28], comp2_0[29:29]);
  C3 I607 (simp4521_0[10:10], comp2_0[30:30], comp2_0[31:31], comp2_0[32:32]);
  C3 I608 (simp4522_0[0:0], simp4521_0[0:0], simp4521_0[1:1], simp4521_0[2:2]);
  C3 I609 (simp4522_0[1:1], simp4521_0[3:3], simp4521_0[4:4], simp4521_0[5:5]);
  C3 I610 (simp4522_0[2:2], simp4521_0[6:6], simp4521_0[7:7], simp4521_0[8:8]);
  C2 I611 (simp4522_0[3:3], simp4521_0[9:9], simp4521_0[10:10]);
  C3 I612 (simp4523_0[0:0], simp4522_0[0:0], simp4522_0[1:1], simp4522_0[2:2]);
  BUFF I613 (simp4523_0[1:1], simp4522_0[3:3]);
  C2 I614 (icomp_2, simp4523_0[0:0], simp4523_0[1:1]);
  OR2 I615 (comp3_0[0:0], i_3r0[0:0], i_3r1[0:0]);
  OR2 I616 (comp3_0[1:1], i_3r0[1:1], i_3r1[1:1]);
  OR2 I617 (comp3_0[2:2], i_3r0[2:2], i_3r1[2:2]);
  OR2 I618 (comp3_0[3:3], i_3r0[3:3], i_3r1[3:3]);
  OR2 I619 (comp3_0[4:4], i_3r0[4:4], i_3r1[4:4]);
  OR2 I620 (comp3_0[5:5], i_3r0[5:5], i_3r1[5:5]);
  OR2 I621 (comp3_0[6:6], i_3r0[6:6], i_3r1[6:6]);
  OR2 I622 (comp3_0[7:7], i_3r0[7:7], i_3r1[7:7]);
  OR2 I623 (comp3_0[8:8], i_3r0[8:8], i_3r1[8:8]);
  OR2 I624 (comp3_0[9:9], i_3r0[9:9], i_3r1[9:9]);
  OR2 I625 (comp3_0[10:10], i_3r0[10:10], i_3r1[10:10]);
  OR2 I626 (comp3_0[11:11], i_3r0[11:11], i_3r1[11:11]);
  OR2 I627 (comp3_0[12:12], i_3r0[12:12], i_3r1[12:12]);
  OR2 I628 (comp3_0[13:13], i_3r0[13:13], i_3r1[13:13]);
  OR2 I629 (comp3_0[14:14], i_3r0[14:14], i_3r1[14:14]);
  OR2 I630 (comp3_0[15:15], i_3r0[15:15], i_3r1[15:15]);
  OR2 I631 (comp3_0[16:16], i_3r0[16:16], i_3r1[16:16]);
  OR2 I632 (comp3_0[17:17], i_3r0[17:17], i_3r1[17:17]);
  OR2 I633 (comp3_0[18:18], i_3r0[18:18], i_3r1[18:18]);
  OR2 I634 (comp3_0[19:19], i_3r0[19:19], i_3r1[19:19]);
  OR2 I635 (comp3_0[20:20], i_3r0[20:20], i_3r1[20:20]);
  OR2 I636 (comp3_0[21:21], i_3r0[21:21], i_3r1[21:21]);
  OR2 I637 (comp3_0[22:22], i_3r0[22:22], i_3r1[22:22]);
  OR2 I638 (comp3_0[23:23], i_3r0[23:23], i_3r1[23:23]);
  OR2 I639 (comp3_0[24:24], i_3r0[24:24], i_3r1[24:24]);
  OR2 I640 (comp3_0[25:25], i_3r0[25:25], i_3r1[25:25]);
  OR2 I641 (comp3_0[26:26], i_3r0[26:26], i_3r1[26:26]);
  OR2 I642 (comp3_0[27:27], i_3r0[27:27], i_3r1[27:27]);
  OR2 I643 (comp3_0[28:28], i_3r0[28:28], i_3r1[28:28]);
  OR2 I644 (comp3_0[29:29], i_3r0[29:29], i_3r1[29:29]);
  OR2 I645 (comp3_0[30:30], i_3r0[30:30], i_3r1[30:30]);
  OR2 I646 (comp3_0[31:31], i_3r0[31:31], i_3r1[31:31]);
  OR2 I647 (comp3_0[32:32], i_3r0[32:32], i_3r1[32:32]);
  C3 I648 (simp4871_0[0:0], comp3_0[0:0], comp3_0[1:1], comp3_0[2:2]);
  C3 I649 (simp4871_0[1:1], comp3_0[3:3], comp3_0[4:4], comp3_0[5:5]);
  C3 I650 (simp4871_0[2:2], comp3_0[6:6], comp3_0[7:7], comp3_0[8:8]);
  C3 I651 (simp4871_0[3:3], comp3_0[9:9], comp3_0[10:10], comp3_0[11:11]);
  C3 I652 (simp4871_0[4:4], comp3_0[12:12], comp3_0[13:13], comp3_0[14:14]);
  C3 I653 (simp4871_0[5:5], comp3_0[15:15], comp3_0[16:16], comp3_0[17:17]);
  C3 I654 (simp4871_0[6:6], comp3_0[18:18], comp3_0[19:19], comp3_0[20:20]);
  C3 I655 (simp4871_0[7:7], comp3_0[21:21], comp3_0[22:22], comp3_0[23:23]);
  C3 I656 (simp4871_0[8:8], comp3_0[24:24], comp3_0[25:25], comp3_0[26:26]);
  C3 I657 (simp4871_0[9:9], comp3_0[27:27], comp3_0[28:28], comp3_0[29:29]);
  C3 I658 (simp4871_0[10:10], comp3_0[30:30], comp3_0[31:31], comp3_0[32:32]);
  C3 I659 (simp4872_0[0:0], simp4871_0[0:0], simp4871_0[1:1], simp4871_0[2:2]);
  C3 I660 (simp4872_0[1:1], simp4871_0[3:3], simp4871_0[4:4], simp4871_0[5:5]);
  C3 I661 (simp4872_0[2:2], simp4871_0[6:6], simp4871_0[7:7], simp4871_0[8:8]);
  C2 I662 (simp4872_0[3:3], simp4871_0[9:9], simp4871_0[10:10]);
  C3 I663 (simp4873_0[0:0], simp4872_0[0:0], simp4872_0[1:1], simp4872_0[2:2]);
  BUFF I664 (simp4873_0[1:1], simp4872_0[3:3]);
  C2 I665 (icomp_3, simp4873_0[0:0], simp4873_0[1:1]);
  C2R I666 (choice_0, icomp_0, nchosen_0, reset);
  C2R I667 (choice_1, icomp_1, nchosen_0, reset);
  C2R I668 (choice_2, icomp_2, nchosen_0, reset);
  C2R I669 (choice_3, icomp_3, nchosen_0, reset);
  NOR3 I670 (simp4921_0[0:0], choice_0, choice_1, choice_2);
  INV I671 (simp4921_0[1:1], choice_3);
  NAND2 I672 (anychoice_0, simp4921_0[0:0], simp4921_0[1:1]);
  NOR2 I673 (nchosen_0, anychoice_0, o_0a);
  C2R I674 (i_0a, choice_0, o_0a, reset);
  C2R I675 (i_1a, choice_1, o_0a, reset);
  C2R I676 (i_2a, choice_2, o_0a, reset);
  C2R I677 (i_3a, choice_3, o_0a, reset);
endmodule

// tkm4x0b TeakM [Many [0,0,0,0],One 0]
module tkm4x0b (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, i_3r, i_3a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  output o_0r;
  input o_0a;
  input reset;
  wire nchosen_0;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire [1:0] simp101_0;
  C2R I0 (choice_0, i_0r, nchosen_0, reset);
  C2R I1 (choice_1, i_1r, nchosen_0, reset);
  C2R I2 (choice_2, i_2r, nchosen_0, reset);
  C2R I3 (choice_3, i_3r, nchosen_0, reset);
  NOR2 I4 (nchosen_0, o_0r, o_0a);
  NOR3 I5 (simp101_0[0:0], choice_0, choice_1, choice_2);
  INV I6 (simp101_0[1:1], choice_3);
  NAND2 I7 (o_0r, simp101_0[0:0], simp101_0[1:1]);
  C2R I8 (i_0a, choice_0, o_0a, reset);
  C2R I9 (i_1a, choice_1, o_0a, reset);
  C2R I10 (i_2a, choice_2, o_0a, reset);
  C2R I11 (i_3a, choice_3, o_0a, reset);
endmodule

// tkf3mo0w0_o0w3 TeakF [0,0] [One 3,Many [0,3]]
module tkf3mo0w0_o0w3 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [2:0] o_1r0;
  output [2:0] o_1r1;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire [2:0] comp_0;
  OR2 I0 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I3 (icomplete_0, comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  BUFF I4 (o_1r0[0:0], i_0r0[0:0]);
  BUFF I5 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I6 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I7 (o_1r1[0:0], i_0r1[0:0]);
  BUFF I8 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I9 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I10 (o_0r, icomplete_0);
  C3 I11 (i_0a, icomplete_0, o_0a, o_1a);
endmodule

// tkm2x1b TeakM [Many [1,1],One 1]
module tkm2x1b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input i_1r0;
  input i_1r1;
  output i_1a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire gfint_0;
  wire gfint_1;
  wire gtint_0;
  wire gtint_1;
  wire choice_0;
  wire choice_1;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire nchosen_0;
  wire comp0_0;
  wire comp1_0;
  OR2 I0 (o_0r0, gfint_0, gfint_1);
  OR2 I1 (o_0r1, gtint_0, gtint_1);
  AND2 I2 (gtint_0, choice_0, i_0r1);
  AND2 I3 (gtint_1, choice_1, i_1r1);
  AND2 I4 (gfint_0, choice_0, i_0r0);
  AND2 I5 (gfint_1, choice_1, i_1r0);
  OR2 I6 (comp0_0, i_0r0, i_0r1);
  BUFF I7 (icomp_0, comp0_0);
  OR2 I8 (comp1_0, i_1r0, i_1r1);
  BUFF I9 (icomp_1, comp1_0);
  C2R I10 (choice_0, icomp_0, nchosen_0, reset);
  C2R I11 (choice_1, icomp_1, nchosen_0, reset);
  OR2 I12 (anychoice_0, choice_0, choice_1);
  NOR2 I13 (nchosen_0, anychoice_0, o_0a);
  C2R I14 (i_0a, choice_0, o_0a, reset);
  C2R I15 (i_1a, choice_1, o_0a, reset);
endmodule

// tkm2x0b TeakM [Many [0,0],One 0]
module tkm2x0b (i_0r, i_0a, i_1r, i_1a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  output o_0r;
  input o_0a;
  input reset;
  wire nchosen_0;
  wire choice_0;
  wire choice_1;
  C2R I0 (choice_0, i_0r, nchosen_0, reset);
  C2R I1 (choice_1, i_1r, nchosen_0, reset);
  NOR2 I2 (nchosen_0, o_0r, o_0a);
  OR2 I3 (o_0r, choice_0, choice_1);
  C2R I4 (i_0a, choice_0, o_0a, reset);
  C2R I5 (i_1a, choice_1, o_0a, reset);
endmodule

// tkm3x1b TeakM [Many [1,1,1],One 1]
module tkm3x1b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input i_1r0;
  input i_1r1;
  output i_1a;
  input i_2r0;
  input i_2r1;
  output i_2a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire gfint_0;
  wire gfint_1;
  wire gfint_2;
  wire gtint_0;
  wire gtint_1;
  wire gtint_2;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire nchosen_0;
  wire comp0_0;
  wire comp1_0;
  wire comp2_0;
  OR3 I0 (o_0r0, gfint_0, gfint_1, gfint_2);
  OR3 I1 (o_0r1, gtint_0, gtint_1, gtint_2);
  AND2 I2 (gtint_0, choice_0, i_0r1);
  AND2 I3 (gtint_1, choice_1, i_1r1);
  AND2 I4 (gtint_2, choice_2, i_2r1);
  AND2 I5 (gfint_0, choice_0, i_0r0);
  AND2 I6 (gfint_1, choice_1, i_1r0);
  AND2 I7 (gfint_2, choice_2, i_2r0);
  OR2 I8 (comp0_0, i_0r0, i_0r1);
  BUFF I9 (icomp_0, comp0_0);
  OR2 I10 (comp1_0, i_1r0, i_1r1);
  BUFF I11 (icomp_1, comp1_0);
  OR2 I12 (comp2_0, i_2r0, i_2r1);
  BUFF I13 (icomp_2, comp2_0);
  C2R I14 (choice_0, icomp_0, nchosen_0, reset);
  C2R I15 (choice_1, icomp_1, nchosen_0, reset);
  C2R I16 (choice_2, icomp_2, nchosen_0, reset);
  OR3 I17 (anychoice_0, choice_0, choice_1, choice_2);
  NOR2 I18 (nchosen_0, anychoice_0, o_0a);
  C2R I19 (i_0a, choice_0, o_0a, reset);
  C2R I20 (i_1a, choice_1, o_0a, reset);
  C2R I21 (i_2a, choice_2, o_0a, reset);
endmodule

// tkj8m1_7 TeakJ [Many [1,7],One 8]
module tkj8m1_7 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input [6:0] i_1r0;
  input [6:0] i_1r1;
  output i_1a;
  output [7:0] o_0r0;
  output [7:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r0);
  BUFF I1 (o_0r0[1:1], i_1r0[0:0]);
  BUFF I2 (o_0r0[2:2], i_1r0[1:1]);
  BUFF I3 (o_0r0[3:3], i_1r0[2:2]);
  BUFF I4 (o_0r0[4:4], i_1r0[3:3]);
  BUFF I5 (o_0r0[5:5], i_1r0[4:4]);
  BUFF I6 (o_0r0[6:6], i_1r0[5:5]);
  BUFF I7 (o_0r0[7:7], i_1r0[6:6]);
  BUFF I8 (o_0r1[0:0], i_0r1);
  BUFF I9 (o_0r1[1:1], i_1r1[0:0]);
  BUFF I10 (o_0r1[2:2], i_1r1[1:1]);
  BUFF I11 (o_0r1[3:3], i_1r1[2:2]);
  BUFF I12 (o_0r1[4:4], i_1r1[3:3]);
  BUFF I13 (o_0r1[5:5], i_1r1[4:4]);
  BUFF I14 (o_0r1[6:6], i_1r1[5:5]);
  BUFF I15 (o_0r1[7:7], i_1r1[6:6]);
  BUFF I16 (i_0a, o_0a);
  BUFF I17 (i_1a, o_0a);
endmodule

// tkf33mo0w0_o0w33 TeakF [0,0] [One 33,Many [0,33]]
module tkf33mo0w0_o0w33 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [32:0] i_0r0;
  input [32:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [32:0] o_1r0;
  output [32:0] o_1r1;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire [32:0] comp_0;
  wire [10:0] simp351_0;
  wire [3:0] simp352_0;
  wire [1:0] simp353_0;
  OR2 I0 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (comp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (comp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (comp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (comp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (comp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (comp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (comp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (comp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (comp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (comp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (comp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (comp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (comp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (comp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (comp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (comp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (comp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (comp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (comp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (comp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (comp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (comp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (comp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (comp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I30 (comp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I31 (comp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I32 (comp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  C3 I33 (simp351_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I34 (simp351_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C3 I35 (simp351_0[2:2], comp_0[6:6], comp_0[7:7], comp_0[8:8]);
  C3 I36 (simp351_0[3:3], comp_0[9:9], comp_0[10:10], comp_0[11:11]);
  C3 I37 (simp351_0[4:4], comp_0[12:12], comp_0[13:13], comp_0[14:14]);
  C3 I38 (simp351_0[5:5], comp_0[15:15], comp_0[16:16], comp_0[17:17]);
  C3 I39 (simp351_0[6:6], comp_0[18:18], comp_0[19:19], comp_0[20:20]);
  C3 I40 (simp351_0[7:7], comp_0[21:21], comp_0[22:22], comp_0[23:23]);
  C3 I41 (simp351_0[8:8], comp_0[24:24], comp_0[25:25], comp_0[26:26]);
  C3 I42 (simp351_0[9:9], comp_0[27:27], comp_0[28:28], comp_0[29:29]);
  C3 I43 (simp351_0[10:10], comp_0[30:30], comp_0[31:31], comp_0[32:32]);
  C3 I44 (simp352_0[0:0], simp351_0[0:0], simp351_0[1:1], simp351_0[2:2]);
  C3 I45 (simp352_0[1:1], simp351_0[3:3], simp351_0[4:4], simp351_0[5:5]);
  C3 I46 (simp352_0[2:2], simp351_0[6:6], simp351_0[7:7], simp351_0[8:8]);
  C2 I47 (simp352_0[3:3], simp351_0[9:9], simp351_0[10:10]);
  C3 I48 (simp353_0[0:0], simp352_0[0:0], simp352_0[1:1], simp352_0[2:2]);
  BUFF I49 (simp353_0[1:1], simp352_0[3:3]);
  C2 I50 (icomplete_0, simp353_0[0:0], simp353_0[1:1]);
  BUFF I51 (o_1r0[0:0], i_0r0[0:0]);
  BUFF I52 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I53 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I54 (o_1r0[3:3], i_0r0[3:3]);
  BUFF I55 (o_1r0[4:4], i_0r0[4:4]);
  BUFF I56 (o_1r0[5:5], i_0r0[5:5]);
  BUFF I57 (o_1r0[6:6], i_0r0[6:6]);
  BUFF I58 (o_1r0[7:7], i_0r0[7:7]);
  BUFF I59 (o_1r0[8:8], i_0r0[8:8]);
  BUFF I60 (o_1r0[9:9], i_0r0[9:9]);
  BUFF I61 (o_1r0[10:10], i_0r0[10:10]);
  BUFF I62 (o_1r0[11:11], i_0r0[11:11]);
  BUFF I63 (o_1r0[12:12], i_0r0[12:12]);
  BUFF I64 (o_1r0[13:13], i_0r0[13:13]);
  BUFF I65 (o_1r0[14:14], i_0r0[14:14]);
  BUFF I66 (o_1r0[15:15], i_0r0[15:15]);
  BUFF I67 (o_1r0[16:16], i_0r0[16:16]);
  BUFF I68 (o_1r0[17:17], i_0r0[17:17]);
  BUFF I69 (o_1r0[18:18], i_0r0[18:18]);
  BUFF I70 (o_1r0[19:19], i_0r0[19:19]);
  BUFF I71 (o_1r0[20:20], i_0r0[20:20]);
  BUFF I72 (o_1r0[21:21], i_0r0[21:21]);
  BUFF I73 (o_1r0[22:22], i_0r0[22:22]);
  BUFF I74 (o_1r0[23:23], i_0r0[23:23]);
  BUFF I75 (o_1r0[24:24], i_0r0[24:24]);
  BUFF I76 (o_1r0[25:25], i_0r0[25:25]);
  BUFF I77 (o_1r0[26:26], i_0r0[26:26]);
  BUFF I78 (o_1r0[27:27], i_0r0[27:27]);
  BUFF I79 (o_1r0[28:28], i_0r0[28:28]);
  BUFF I80 (o_1r0[29:29], i_0r0[29:29]);
  BUFF I81 (o_1r0[30:30], i_0r0[30:30]);
  BUFF I82 (o_1r0[31:31], i_0r0[31:31]);
  BUFF I83 (o_1r0[32:32], i_0r0[32:32]);
  BUFF I84 (o_1r1[0:0], i_0r1[0:0]);
  BUFF I85 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I86 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I87 (o_1r1[3:3], i_0r1[3:3]);
  BUFF I88 (o_1r1[4:4], i_0r1[4:4]);
  BUFF I89 (o_1r1[5:5], i_0r1[5:5]);
  BUFF I90 (o_1r1[6:6], i_0r1[6:6]);
  BUFF I91 (o_1r1[7:7], i_0r1[7:7]);
  BUFF I92 (o_1r1[8:8], i_0r1[8:8]);
  BUFF I93 (o_1r1[9:9], i_0r1[9:9]);
  BUFF I94 (o_1r1[10:10], i_0r1[10:10]);
  BUFF I95 (o_1r1[11:11], i_0r1[11:11]);
  BUFF I96 (o_1r1[12:12], i_0r1[12:12]);
  BUFF I97 (o_1r1[13:13], i_0r1[13:13]);
  BUFF I98 (o_1r1[14:14], i_0r1[14:14]);
  BUFF I99 (o_1r1[15:15], i_0r1[15:15]);
  BUFF I100 (o_1r1[16:16], i_0r1[16:16]);
  BUFF I101 (o_1r1[17:17], i_0r1[17:17]);
  BUFF I102 (o_1r1[18:18], i_0r1[18:18]);
  BUFF I103 (o_1r1[19:19], i_0r1[19:19]);
  BUFF I104 (o_1r1[20:20], i_0r1[20:20]);
  BUFF I105 (o_1r1[21:21], i_0r1[21:21]);
  BUFF I106 (o_1r1[22:22], i_0r1[22:22]);
  BUFF I107 (o_1r1[23:23], i_0r1[23:23]);
  BUFF I108 (o_1r1[24:24], i_0r1[24:24]);
  BUFF I109 (o_1r1[25:25], i_0r1[25:25]);
  BUFF I110 (o_1r1[26:26], i_0r1[26:26]);
  BUFF I111 (o_1r1[27:27], i_0r1[27:27]);
  BUFF I112 (o_1r1[28:28], i_0r1[28:28]);
  BUFF I113 (o_1r1[29:29], i_0r1[29:29]);
  BUFF I114 (o_1r1[30:30], i_0r1[30:30]);
  BUFF I115 (o_1r1[31:31], i_0r1[31:31]);
  BUFF I116 (o_1r1[32:32], i_0r1[32:32]);
  BUFF I117 (o_0r, icomplete_0);
  C3 I118 (i_0a, icomplete_0, o_0a, o_1a);
endmodule

// tkvavbvciv65_wo0w65_ro0w32o0w32o0w32o0w32o32w32o32w32o32w32o32w32o32w32o64w1o64w1o64w1o64w1o64w1o64w
//   1 TeakV "a_v-b_v-ci_v" 65 [] [0] [0,0,0,0,32,32,32,32,32,64,64,64,64,64,64] [Many [65],Many [0],Many
//    [0,0,0,0,0,0,0,0,0,0,0,0,0,0,0],Many [32,32,32,32,32,32,32,32,32,1,1,1,1,1,1]]
module tkvavbvciv65_wo0w65_ro0w32o0w32o0w32o0w32o32w32o32w32o32w32o32w32o32w32o64w1o64w1o64w1o64w1o64w1o64w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rg_5r, rg_5a, rg_6r, rg_6a, rg_7r, rg_7a, rg_8r, rg_8a, rg_9r, rg_9a, rg_10r, rg_10a, rg_11r, rg_11a, rg_12r, rg_12a, rg_13r, rg_13a, rg_14r, rg_14a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, rd_5r0, rd_5r1, rd_5a, rd_6r0, rd_6r1, rd_6a, rd_7r0, rd_7r1, rd_7a, rd_8r0, rd_8r1, rd_8a, rd_9r0, rd_9r1, rd_9a, rd_10r0, rd_10r1, rd_10a, rd_11r0, rd_11r1, rd_11a, rd_12r0, rd_12r1, rd_12a, rd_13r0, rd_13r1, rd_13a, rd_14r0, rd_14r1, rd_14a, reset);
  input [64:0] wg_0r0;
  input [64:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  input rg_5r;
  output rg_5a;
  input rg_6r;
  output rg_6a;
  input rg_7r;
  output rg_7a;
  input rg_8r;
  output rg_8a;
  input rg_9r;
  output rg_9a;
  input rg_10r;
  output rg_10a;
  input rg_11r;
  output rg_11a;
  input rg_12r;
  output rg_12a;
  input rg_13r;
  output rg_13a;
  input rg_14r;
  output rg_14a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  output [31:0] rd_3r0;
  output [31:0] rd_3r1;
  input rd_3a;
  output [31:0] rd_4r0;
  output [31:0] rd_4r1;
  input rd_4a;
  output [31:0] rd_5r0;
  output [31:0] rd_5r1;
  input rd_5a;
  output [31:0] rd_6r0;
  output [31:0] rd_6r1;
  input rd_6a;
  output [31:0] rd_7r0;
  output [31:0] rd_7r1;
  input rd_7a;
  output [31:0] rd_8r0;
  output [31:0] rd_8r1;
  input rd_8a;
  output rd_9r0;
  output rd_9r1;
  input rd_9a;
  output rd_10r0;
  output rd_10r1;
  input rd_10a;
  output rd_11r0;
  output rd_11r1;
  input rd_11a;
  output rd_12r0;
  output rd_12r1;
  input rd_12a;
  output rd_13r0;
  output rd_13r1;
  input rd_13a;
  output rd_14r0;
  output rd_14r1;
  input rd_14a;
  input reset;
  wire [64:0] wf_0;
  wire [64:0] wt_0;
  wire [64:0] df_0;
  wire [64:0] dt_0;
  wire wc_0;
  wire [64:0] wacks_0;
  wire [64:0] wenr_0;
  wire [64:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [64:0] drlgf_0;
  wire [64:0] drlgt_0;
  wire [64:0] comp0_0;
  wire [21:0] simp4691_0;
  wire [7:0] simp4692_0;
  wire [2:0] simp4693_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [64:0] conwgit_0;
  wire [64:0] conwgif_0;
  wire conwig_0;
  wire [21:0] simp8031_0;
  wire [7:0] simp8032_0;
  wire [2:0] simp8033_0;
  wire [9:0] simp13921_0;
  wire [3:0] simp13922_0;
  wire [1:0] simp13923_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (wen_0[32:32], wenr_0[32:32], nreset_0);
  AND2 I34 (wen_0[33:33], wenr_0[33:33], nreset_0);
  AND2 I35 (wen_0[34:34], wenr_0[34:34], nreset_0);
  AND2 I36 (wen_0[35:35], wenr_0[35:35], nreset_0);
  AND2 I37 (wen_0[36:36], wenr_0[36:36], nreset_0);
  AND2 I38 (wen_0[37:37], wenr_0[37:37], nreset_0);
  AND2 I39 (wen_0[38:38], wenr_0[38:38], nreset_0);
  AND2 I40 (wen_0[39:39], wenr_0[39:39], nreset_0);
  AND2 I41 (wen_0[40:40], wenr_0[40:40], nreset_0);
  AND2 I42 (wen_0[41:41], wenr_0[41:41], nreset_0);
  AND2 I43 (wen_0[42:42], wenr_0[42:42], nreset_0);
  AND2 I44 (wen_0[43:43], wenr_0[43:43], nreset_0);
  AND2 I45 (wen_0[44:44], wenr_0[44:44], nreset_0);
  AND2 I46 (wen_0[45:45], wenr_0[45:45], nreset_0);
  AND2 I47 (wen_0[46:46], wenr_0[46:46], nreset_0);
  AND2 I48 (wen_0[47:47], wenr_0[47:47], nreset_0);
  AND2 I49 (wen_0[48:48], wenr_0[48:48], nreset_0);
  AND2 I50 (wen_0[49:49], wenr_0[49:49], nreset_0);
  AND2 I51 (wen_0[50:50], wenr_0[50:50], nreset_0);
  AND2 I52 (wen_0[51:51], wenr_0[51:51], nreset_0);
  AND2 I53 (wen_0[52:52], wenr_0[52:52], nreset_0);
  AND2 I54 (wen_0[53:53], wenr_0[53:53], nreset_0);
  AND2 I55 (wen_0[54:54], wenr_0[54:54], nreset_0);
  AND2 I56 (wen_0[55:55], wenr_0[55:55], nreset_0);
  AND2 I57 (wen_0[56:56], wenr_0[56:56], nreset_0);
  AND2 I58 (wen_0[57:57], wenr_0[57:57], nreset_0);
  AND2 I59 (wen_0[58:58], wenr_0[58:58], nreset_0);
  AND2 I60 (wen_0[59:59], wenr_0[59:59], nreset_0);
  AND2 I61 (wen_0[60:60], wenr_0[60:60], nreset_0);
  AND2 I62 (wen_0[61:61], wenr_0[61:61], nreset_0);
  AND2 I63 (wen_0[62:62], wenr_0[62:62], nreset_0);
  AND2 I64 (wen_0[63:63], wenr_0[63:63], nreset_0);
  AND2 I65 (wen_0[64:64], wenr_0[64:64], nreset_0);
  AND2 I66 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I67 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I68 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I69 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I70 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I71 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I72 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I73 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I74 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I75 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I76 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I77 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I78 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I79 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I80 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I81 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I82 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I83 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I84 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I85 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I86 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I87 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I88 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I89 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I90 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I91 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I92 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I93 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I94 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I95 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I96 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I97 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I98 (drlgf_0[32:32], wf_0[32:32], wen_0[32:32]);
  AND2 I99 (drlgf_0[33:33], wf_0[33:33], wen_0[33:33]);
  AND2 I100 (drlgf_0[34:34], wf_0[34:34], wen_0[34:34]);
  AND2 I101 (drlgf_0[35:35], wf_0[35:35], wen_0[35:35]);
  AND2 I102 (drlgf_0[36:36], wf_0[36:36], wen_0[36:36]);
  AND2 I103 (drlgf_0[37:37], wf_0[37:37], wen_0[37:37]);
  AND2 I104 (drlgf_0[38:38], wf_0[38:38], wen_0[38:38]);
  AND2 I105 (drlgf_0[39:39], wf_0[39:39], wen_0[39:39]);
  AND2 I106 (drlgf_0[40:40], wf_0[40:40], wen_0[40:40]);
  AND2 I107 (drlgf_0[41:41], wf_0[41:41], wen_0[41:41]);
  AND2 I108 (drlgf_0[42:42], wf_0[42:42], wen_0[42:42]);
  AND2 I109 (drlgf_0[43:43], wf_0[43:43], wen_0[43:43]);
  AND2 I110 (drlgf_0[44:44], wf_0[44:44], wen_0[44:44]);
  AND2 I111 (drlgf_0[45:45], wf_0[45:45], wen_0[45:45]);
  AND2 I112 (drlgf_0[46:46], wf_0[46:46], wen_0[46:46]);
  AND2 I113 (drlgf_0[47:47], wf_0[47:47], wen_0[47:47]);
  AND2 I114 (drlgf_0[48:48], wf_0[48:48], wen_0[48:48]);
  AND2 I115 (drlgf_0[49:49], wf_0[49:49], wen_0[49:49]);
  AND2 I116 (drlgf_0[50:50], wf_0[50:50], wen_0[50:50]);
  AND2 I117 (drlgf_0[51:51], wf_0[51:51], wen_0[51:51]);
  AND2 I118 (drlgf_0[52:52], wf_0[52:52], wen_0[52:52]);
  AND2 I119 (drlgf_0[53:53], wf_0[53:53], wen_0[53:53]);
  AND2 I120 (drlgf_0[54:54], wf_0[54:54], wen_0[54:54]);
  AND2 I121 (drlgf_0[55:55], wf_0[55:55], wen_0[55:55]);
  AND2 I122 (drlgf_0[56:56], wf_0[56:56], wen_0[56:56]);
  AND2 I123 (drlgf_0[57:57], wf_0[57:57], wen_0[57:57]);
  AND2 I124 (drlgf_0[58:58], wf_0[58:58], wen_0[58:58]);
  AND2 I125 (drlgf_0[59:59], wf_0[59:59], wen_0[59:59]);
  AND2 I126 (drlgf_0[60:60], wf_0[60:60], wen_0[60:60]);
  AND2 I127 (drlgf_0[61:61], wf_0[61:61], wen_0[61:61]);
  AND2 I128 (drlgf_0[62:62], wf_0[62:62], wen_0[62:62]);
  AND2 I129 (drlgf_0[63:63], wf_0[63:63], wen_0[63:63]);
  AND2 I130 (drlgf_0[64:64], wf_0[64:64], wen_0[64:64]);
  AND2 I131 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I132 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I133 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I134 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I135 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I136 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I137 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I138 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I139 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I140 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I141 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I142 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I143 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I144 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I145 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I146 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I147 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I148 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I149 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I150 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I151 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I152 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I153 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I154 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I155 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I156 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I157 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I158 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I159 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I160 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I161 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I162 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  AND2 I163 (drlgt_0[32:32], wt_0[32:32], wen_0[32:32]);
  AND2 I164 (drlgt_0[33:33], wt_0[33:33], wen_0[33:33]);
  AND2 I165 (drlgt_0[34:34], wt_0[34:34], wen_0[34:34]);
  AND2 I166 (drlgt_0[35:35], wt_0[35:35], wen_0[35:35]);
  AND2 I167 (drlgt_0[36:36], wt_0[36:36], wen_0[36:36]);
  AND2 I168 (drlgt_0[37:37], wt_0[37:37], wen_0[37:37]);
  AND2 I169 (drlgt_0[38:38], wt_0[38:38], wen_0[38:38]);
  AND2 I170 (drlgt_0[39:39], wt_0[39:39], wen_0[39:39]);
  AND2 I171 (drlgt_0[40:40], wt_0[40:40], wen_0[40:40]);
  AND2 I172 (drlgt_0[41:41], wt_0[41:41], wen_0[41:41]);
  AND2 I173 (drlgt_0[42:42], wt_0[42:42], wen_0[42:42]);
  AND2 I174 (drlgt_0[43:43], wt_0[43:43], wen_0[43:43]);
  AND2 I175 (drlgt_0[44:44], wt_0[44:44], wen_0[44:44]);
  AND2 I176 (drlgt_0[45:45], wt_0[45:45], wen_0[45:45]);
  AND2 I177 (drlgt_0[46:46], wt_0[46:46], wen_0[46:46]);
  AND2 I178 (drlgt_0[47:47], wt_0[47:47], wen_0[47:47]);
  AND2 I179 (drlgt_0[48:48], wt_0[48:48], wen_0[48:48]);
  AND2 I180 (drlgt_0[49:49], wt_0[49:49], wen_0[49:49]);
  AND2 I181 (drlgt_0[50:50], wt_0[50:50], wen_0[50:50]);
  AND2 I182 (drlgt_0[51:51], wt_0[51:51], wen_0[51:51]);
  AND2 I183 (drlgt_0[52:52], wt_0[52:52], wen_0[52:52]);
  AND2 I184 (drlgt_0[53:53], wt_0[53:53], wen_0[53:53]);
  AND2 I185 (drlgt_0[54:54], wt_0[54:54], wen_0[54:54]);
  AND2 I186 (drlgt_0[55:55], wt_0[55:55], wen_0[55:55]);
  AND2 I187 (drlgt_0[56:56], wt_0[56:56], wen_0[56:56]);
  AND2 I188 (drlgt_0[57:57], wt_0[57:57], wen_0[57:57]);
  AND2 I189 (drlgt_0[58:58], wt_0[58:58], wen_0[58:58]);
  AND2 I190 (drlgt_0[59:59], wt_0[59:59], wen_0[59:59]);
  AND2 I191 (drlgt_0[60:60], wt_0[60:60], wen_0[60:60]);
  AND2 I192 (drlgt_0[61:61], wt_0[61:61], wen_0[61:61]);
  AND2 I193 (drlgt_0[62:62], wt_0[62:62], wen_0[62:62]);
  AND2 I194 (drlgt_0[63:63], wt_0[63:63], wen_0[63:63]);
  AND2 I195 (drlgt_0[64:64], wt_0[64:64], wen_0[64:64]);
  NOR2 I196 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I197 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I198 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I199 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I200 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I201 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I202 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I203 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I204 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I205 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I206 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I207 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I208 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I209 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I210 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I211 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I212 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I213 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I214 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I215 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I216 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I217 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I218 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I219 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I220 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I221 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I222 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I223 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I224 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I225 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I226 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I227 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR2 I228 (df_0[32:32], dt_0[32:32], drlgt_0[32:32]);
  NOR2 I229 (df_0[33:33], dt_0[33:33], drlgt_0[33:33]);
  NOR2 I230 (df_0[34:34], dt_0[34:34], drlgt_0[34:34]);
  NOR2 I231 (df_0[35:35], dt_0[35:35], drlgt_0[35:35]);
  NOR2 I232 (df_0[36:36], dt_0[36:36], drlgt_0[36:36]);
  NOR2 I233 (df_0[37:37], dt_0[37:37], drlgt_0[37:37]);
  NOR2 I234 (df_0[38:38], dt_0[38:38], drlgt_0[38:38]);
  NOR2 I235 (df_0[39:39], dt_0[39:39], drlgt_0[39:39]);
  NOR2 I236 (df_0[40:40], dt_0[40:40], drlgt_0[40:40]);
  NOR2 I237 (df_0[41:41], dt_0[41:41], drlgt_0[41:41]);
  NOR2 I238 (df_0[42:42], dt_0[42:42], drlgt_0[42:42]);
  NOR2 I239 (df_0[43:43], dt_0[43:43], drlgt_0[43:43]);
  NOR2 I240 (df_0[44:44], dt_0[44:44], drlgt_0[44:44]);
  NOR2 I241 (df_0[45:45], dt_0[45:45], drlgt_0[45:45]);
  NOR2 I242 (df_0[46:46], dt_0[46:46], drlgt_0[46:46]);
  NOR2 I243 (df_0[47:47], dt_0[47:47], drlgt_0[47:47]);
  NOR2 I244 (df_0[48:48], dt_0[48:48], drlgt_0[48:48]);
  NOR2 I245 (df_0[49:49], dt_0[49:49], drlgt_0[49:49]);
  NOR2 I246 (df_0[50:50], dt_0[50:50], drlgt_0[50:50]);
  NOR2 I247 (df_0[51:51], dt_0[51:51], drlgt_0[51:51]);
  NOR2 I248 (df_0[52:52], dt_0[52:52], drlgt_0[52:52]);
  NOR2 I249 (df_0[53:53], dt_0[53:53], drlgt_0[53:53]);
  NOR2 I250 (df_0[54:54], dt_0[54:54], drlgt_0[54:54]);
  NOR2 I251 (df_0[55:55], dt_0[55:55], drlgt_0[55:55]);
  NOR2 I252 (df_0[56:56], dt_0[56:56], drlgt_0[56:56]);
  NOR2 I253 (df_0[57:57], dt_0[57:57], drlgt_0[57:57]);
  NOR2 I254 (df_0[58:58], dt_0[58:58], drlgt_0[58:58]);
  NOR2 I255 (df_0[59:59], dt_0[59:59], drlgt_0[59:59]);
  NOR2 I256 (df_0[60:60], dt_0[60:60], drlgt_0[60:60]);
  NOR2 I257 (df_0[61:61], dt_0[61:61], drlgt_0[61:61]);
  NOR2 I258 (df_0[62:62], dt_0[62:62], drlgt_0[62:62]);
  NOR2 I259 (df_0[63:63], dt_0[63:63], drlgt_0[63:63]);
  NOR2 I260 (df_0[64:64], dt_0[64:64], drlgt_0[64:64]);
  NOR3 I261 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I262 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I263 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I264 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I265 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I266 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I267 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I268 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I269 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I270 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I271 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I272 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I273 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I274 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I275 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I276 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I277 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I278 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I279 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I280 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I281 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I282 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I283 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I284 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I285 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I286 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I287 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I288 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I289 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I290 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I291 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I292 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  NOR3 I293 (dt_0[32:32], df_0[32:32], drlgf_0[32:32], reset);
  NOR3 I294 (dt_0[33:33], df_0[33:33], drlgf_0[33:33], reset);
  NOR3 I295 (dt_0[34:34], df_0[34:34], drlgf_0[34:34], reset);
  NOR3 I296 (dt_0[35:35], df_0[35:35], drlgf_0[35:35], reset);
  NOR3 I297 (dt_0[36:36], df_0[36:36], drlgf_0[36:36], reset);
  NOR3 I298 (dt_0[37:37], df_0[37:37], drlgf_0[37:37], reset);
  NOR3 I299 (dt_0[38:38], df_0[38:38], drlgf_0[38:38], reset);
  NOR3 I300 (dt_0[39:39], df_0[39:39], drlgf_0[39:39], reset);
  NOR3 I301 (dt_0[40:40], df_0[40:40], drlgf_0[40:40], reset);
  NOR3 I302 (dt_0[41:41], df_0[41:41], drlgf_0[41:41], reset);
  NOR3 I303 (dt_0[42:42], df_0[42:42], drlgf_0[42:42], reset);
  NOR3 I304 (dt_0[43:43], df_0[43:43], drlgf_0[43:43], reset);
  NOR3 I305 (dt_0[44:44], df_0[44:44], drlgf_0[44:44], reset);
  NOR3 I306 (dt_0[45:45], df_0[45:45], drlgf_0[45:45], reset);
  NOR3 I307 (dt_0[46:46], df_0[46:46], drlgf_0[46:46], reset);
  NOR3 I308 (dt_0[47:47], df_0[47:47], drlgf_0[47:47], reset);
  NOR3 I309 (dt_0[48:48], df_0[48:48], drlgf_0[48:48], reset);
  NOR3 I310 (dt_0[49:49], df_0[49:49], drlgf_0[49:49], reset);
  NOR3 I311 (dt_0[50:50], df_0[50:50], drlgf_0[50:50], reset);
  NOR3 I312 (dt_0[51:51], df_0[51:51], drlgf_0[51:51], reset);
  NOR3 I313 (dt_0[52:52], df_0[52:52], drlgf_0[52:52], reset);
  NOR3 I314 (dt_0[53:53], df_0[53:53], drlgf_0[53:53], reset);
  NOR3 I315 (dt_0[54:54], df_0[54:54], drlgf_0[54:54], reset);
  NOR3 I316 (dt_0[55:55], df_0[55:55], drlgf_0[55:55], reset);
  NOR3 I317 (dt_0[56:56], df_0[56:56], drlgf_0[56:56], reset);
  NOR3 I318 (dt_0[57:57], df_0[57:57], drlgf_0[57:57], reset);
  NOR3 I319 (dt_0[58:58], df_0[58:58], drlgf_0[58:58], reset);
  NOR3 I320 (dt_0[59:59], df_0[59:59], drlgf_0[59:59], reset);
  NOR3 I321 (dt_0[60:60], df_0[60:60], drlgf_0[60:60], reset);
  NOR3 I322 (dt_0[61:61], df_0[61:61], drlgf_0[61:61], reset);
  NOR3 I323 (dt_0[62:62], df_0[62:62], drlgf_0[62:62], reset);
  NOR3 I324 (dt_0[63:63], df_0[63:63], drlgf_0[63:63], reset);
  NOR3 I325 (dt_0[64:64], df_0[64:64], drlgf_0[64:64], reset);
  AO22 I326 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I327 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I328 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I329 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I330 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I331 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I332 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I333 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I334 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I335 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I336 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I337 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I338 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I339 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I340 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I341 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I342 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I343 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I344 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I345 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I346 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I347 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I348 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I349 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I350 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I351 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I352 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I353 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I354 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I355 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I356 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I357 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  AO22 I358 (wacks_0[32:32], drlgf_0[32:32], df_0[32:32], drlgt_0[32:32], dt_0[32:32]);
  AO22 I359 (wacks_0[33:33], drlgf_0[33:33], df_0[33:33], drlgt_0[33:33], dt_0[33:33]);
  AO22 I360 (wacks_0[34:34], drlgf_0[34:34], df_0[34:34], drlgt_0[34:34], dt_0[34:34]);
  AO22 I361 (wacks_0[35:35], drlgf_0[35:35], df_0[35:35], drlgt_0[35:35], dt_0[35:35]);
  AO22 I362 (wacks_0[36:36], drlgf_0[36:36], df_0[36:36], drlgt_0[36:36], dt_0[36:36]);
  AO22 I363 (wacks_0[37:37], drlgf_0[37:37], df_0[37:37], drlgt_0[37:37], dt_0[37:37]);
  AO22 I364 (wacks_0[38:38], drlgf_0[38:38], df_0[38:38], drlgt_0[38:38], dt_0[38:38]);
  AO22 I365 (wacks_0[39:39], drlgf_0[39:39], df_0[39:39], drlgt_0[39:39], dt_0[39:39]);
  AO22 I366 (wacks_0[40:40], drlgf_0[40:40], df_0[40:40], drlgt_0[40:40], dt_0[40:40]);
  AO22 I367 (wacks_0[41:41], drlgf_0[41:41], df_0[41:41], drlgt_0[41:41], dt_0[41:41]);
  AO22 I368 (wacks_0[42:42], drlgf_0[42:42], df_0[42:42], drlgt_0[42:42], dt_0[42:42]);
  AO22 I369 (wacks_0[43:43], drlgf_0[43:43], df_0[43:43], drlgt_0[43:43], dt_0[43:43]);
  AO22 I370 (wacks_0[44:44], drlgf_0[44:44], df_0[44:44], drlgt_0[44:44], dt_0[44:44]);
  AO22 I371 (wacks_0[45:45], drlgf_0[45:45], df_0[45:45], drlgt_0[45:45], dt_0[45:45]);
  AO22 I372 (wacks_0[46:46], drlgf_0[46:46], df_0[46:46], drlgt_0[46:46], dt_0[46:46]);
  AO22 I373 (wacks_0[47:47], drlgf_0[47:47], df_0[47:47], drlgt_0[47:47], dt_0[47:47]);
  AO22 I374 (wacks_0[48:48], drlgf_0[48:48], df_0[48:48], drlgt_0[48:48], dt_0[48:48]);
  AO22 I375 (wacks_0[49:49], drlgf_0[49:49], df_0[49:49], drlgt_0[49:49], dt_0[49:49]);
  AO22 I376 (wacks_0[50:50], drlgf_0[50:50], df_0[50:50], drlgt_0[50:50], dt_0[50:50]);
  AO22 I377 (wacks_0[51:51], drlgf_0[51:51], df_0[51:51], drlgt_0[51:51], dt_0[51:51]);
  AO22 I378 (wacks_0[52:52], drlgf_0[52:52], df_0[52:52], drlgt_0[52:52], dt_0[52:52]);
  AO22 I379 (wacks_0[53:53], drlgf_0[53:53], df_0[53:53], drlgt_0[53:53], dt_0[53:53]);
  AO22 I380 (wacks_0[54:54], drlgf_0[54:54], df_0[54:54], drlgt_0[54:54], dt_0[54:54]);
  AO22 I381 (wacks_0[55:55], drlgf_0[55:55], df_0[55:55], drlgt_0[55:55], dt_0[55:55]);
  AO22 I382 (wacks_0[56:56], drlgf_0[56:56], df_0[56:56], drlgt_0[56:56], dt_0[56:56]);
  AO22 I383 (wacks_0[57:57], drlgf_0[57:57], df_0[57:57], drlgt_0[57:57], dt_0[57:57]);
  AO22 I384 (wacks_0[58:58], drlgf_0[58:58], df_0[58:58], drlgt_0[58:58], dt_0[58:58]);
  AO22 I385 (wacks_0[59:59], drlgf_0[59:59], df_0[59:59], drlgt_0[59:59], dt_0[59:59]);
  AO22 I386 (wacks_0[60:60], drlgf_0[60:60], df_0[60:60], drlgt_0[60:60], dt_0[60:60]);
  AO22 I387 (wacks_0[61:61], drlgf_0[61:61], df_0[61:61], drlgt_0[61:61], dt_0[61:61]);
  AO22 I388 (wacks_0[62:62], drlgf_0[62:62], df_0[62:62], drlgt_0[62:62], dt_0[62:62]);
  AO22 I389 (wacks_0[63:63], drlgf_0[63:63], df_0[63:63], drlgt_0[63:63], dt_0[63:63]);
  AO22 I390 (wacks_0[64:64], drlgf_0[64:64], df_0[64:64], drlgt_0[64:64], dt_0[64:64]);
  OR2 I391 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I392 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I393 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I394 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I395 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I396 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I397 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I398 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I399 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I400 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I401 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I402 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I403 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I404 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I405 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I406 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I407 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I408 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I409 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I410 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I411 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I412 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I413 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I414 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I415 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I416 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I417 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I418 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I419 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I420 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I421 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I422 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  OR2 I423 (comp0_0[32:32], wg_0r0[32:32], wg_0r1[32:32]);
  OR2 I424 (comp0_0[33:33], wg_0r0[33:33], wg_0r1[33:33]);
  OR2 I425 (comp0_0[34:34], wg_0r0[34:34], wg_0r1[34:34]);
  OR2 I426 (comp0_0[35:35], wg_0r0[35:35], wg_0r1[35:35]);
  OR2 I427 (comp0_0[36:36], wg_0r0[36:36], wg_0r1[36:36]);
  OR2 I428 (comp0_0[37:37], wg_0r0[37:37], wg_0r1[37:37]);
  OR2 I429 (comp0_0[38:38], wg_0r0[38:38], wg_0r1[38:38]);
  OR2 I430 (comp0_0[39:39], wg_0r0[39:39], wg_0r1[39:39]);
  OR2 I431 (comp0_0[40:40], wg_0r0[40:40], wg_0r1[40:40]);
  OR2 I432 (comp0_0[41:41], wg_0r0[41:41], wg_0r1[41:41]);
  OR2 I433 (comp0_0[42:42], wg_0r0[42:42], wg_0r1[42:42]);
  OR2 I434 (comp0_0[43:43], wg_0r0[43:43], wg_0r1[43:43]);
  OR2 I435 (comp0_0[44:44], wg_0r0[44:44], wg_0r1[44:44]);
  OR2 I436 (comp0_0[45:45], wg_0r0[45:45], wg_0r1[45:45]);
  OR2 I437 (comp0_0[46:46], wg_0r0[46:46], wg_0r1[46:46]);
  OR2 I438 (comp0_0[47:47], wg_0r0[47:47], wg_0r1[47:47]);
  OR2 I439 (comp0_0[48:48], wg_0r0[48:48], wg_0r1[48:48]);
  OR2 I440 (comp0_0[49:49], wg_0r0[49:49], wg_0r1[49:49]);
  OR2 I441 (comp0_0[50:50], wg_0r0[50:50], wg_0r1[50:50]);
  OR2 I442 (comp0_0[51:51], wg_0r0[51:51], wg_0r1[51:51]);
  OR2 I443 (comp0_0[52:52], wg_0r0[52:52], wg_0r1[52:52]);
  OR2 I444 (comp0_0[53:53], wg_0r0[53:53], wg_0r1[53:53]);
  OR2 I445 (comp0_0[54:54], wg_0r0[54:54], wg_0r1[54:54]);
  OR2 I446 (comp0_0[55:55], wg_0r0[55:55], wg_0r1[55:55]);
  OR2 I447 (comp0_0[56:56], wg_0r0[56:56], wg_0r1[56:56]);
  OR2 I448 (comp0_0[57:57], wg_0r0[57:57], wg_0r1[57:57]);
  OR2 I449 (comp0_0[58:58], wg_0r0[58:58], wg_0r1[58:58]);
  OR2 I450 (comp0_0[59:59], wg_0r0[59:59], wg_0r1[59:59]);
  OR2 I451 (comp0_0[60:60], wg_0r0[60:60], wg_0r1[60:60]);
  OR2 I452 (comp0_0[61:61], wg_0r0[61:61], wg_0r1[61:61]);
  OR2 I453 (comp0_0[62:62], wg_0r0[62:62], wg_0r1[62:62]);
  OR2 I454 (comp0_0[63:63], wg_0r0[63:63], wg_0r1[63:63]);
  OR2 I455 (comp0_0[64:64], wg_0r0[64:64], wg_0r1[64:64]);
  C3 I456 (simp4691_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I457 (simp4691_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I458 (simp4691_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I459 (simp4691_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I460 (simp4691_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I461 (simp4691_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I462 (simp4691_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I463 (simp4691_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I464 (simp4691_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I465 (simp4691_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C3 I466 (simp4691_0[10:10], comp0_0[30:30], comp0_0[31:31], comp0_0[32:32]);
  C3 I467 (simp4691_0[11:11], comp0_0[33:33], comp0_0[34:34], comp0_0[35:35]);
  C3 I468 (simp4691_0[12:12], comp0_0[36:36], comp0_0[37:37], comp0_0[38:38]);
  C3 I469 (simp4691_0[13:13], comp0_0[39:39], comp0_0[40:40], comp0_0[41:41]);
  C3 I470 (simp4691_0[14:14], comp0_0[42:42], comp0_0[43:43], comp0_0[44:44]);
  C3 I471 (simp4691_0[15:15], comp0_0[45:45], comp0_0[46:46], comp0_0[47:47]);
  C3 I472 (simp4691_0[16:16], comp0_0[48:48], comp0_0[49:49], comp0_0[50:50]);
  C3 I473 (simp4691_0[17:17], comp0_0[51:51], comp0_0[52:52], comp0_0[53:53]);
  C3 I474 (simp4691_0[18:18], comp0_0[54:54], comp0_0[55:55], comp0_0[56:56]);
  C3 I475 (simp4691_0[19:19], comp0_0[57:57], comp0_0[58:58], comp0_0[59:59]);
  C3 I476 (simp4691_0[20:20], comp0_0[60:60], comp0_0[61:61], comp0_0[62:62]);
  C2 I477 (simp4691_0[21:21], comp0_0[63:63], comp0_0[64:64]);
  C3 I478 (simp4692_0[0:0], simp4691_0[0:0], simp4691_0[1:1], simp4691_0[2:2]);
  C3 I479 (simp4692_0[1:1], simp4691_0[3:3], simp4691_0[4:4], simp4691_0[5:5]);
  C3 I480 (simp4692_0[2:2], simp4691_0[6:6], simp4691_0[7:7], simp4691_0[8:8]);
  C3 I481 (simp4692_0[3:3], simp4691_0[9:9], simp4691_0[10:10], simp4691_0[11:11]);
  C3 I482 (simp4692_0[4:4], simp4691_0[12:12], simp4691_0[13:13], simp4691_0[14:14]);
  C3 I483 (simp4692_0[5:5], simp4691_0[15:15], simp4691_0[16:16], simp4691_0[17:17]);
  C3 I484 (simp4692_0[6:6], simp4691_0[18:18], simp4691_0[19:19], simp4691_0[20:20]);
  BUFF I485 (simp4692_0[7:7], simp4691_0[21:21]);
  C3 I486 (simp4693_0[0:0], simp4692_0[0:0], simp4692_0[1:1], simp4692_0[2:2]);
  C3 I487 (simp4693_0[1:1], simp4692_0[3:3], simp4692_0[4:4], simp4692_0[5:5]);
  C2 I488 (simp4693_0[2:2], simp4692_0[6:6], simp4692_0[7:7]);
  C3 I489 (wc_0, simp4693_0[0:0], simp4693_0[1:1], simp4693_0[2:2]);
  AND2 I490 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I491 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I492 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I493 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I494 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I495 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I496 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I497 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I498 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I499 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I500 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I501 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I502 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I503 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I504 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I505 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I506 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I507 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I508 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I509 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I510 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I511 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I512 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I513 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I514 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I515 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I516 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I517 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I518 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I519 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I520 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I521 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I522 (conwgif_0[32:32], wg_0r0[32:32], conwig_0);
  AND2 I523 (conwgif_0[33:33], wg_0r0[33:33], conwig_0);
  AND2 I524 (conwgif_0[34:34], wg_0r0[34:34], conwig_0);
  AND2 I525 (conwgif_0[35:35], wg_0r0[35:35], conwig_0);
  AND2 I526 (conwgif_0[36:36], wg_0r0[36:36], conwig_0);
  AND2 I527 (conwgif_0[37:37], wg_0r0[37:37], conwig_0);
  AND2 I528 (conwgif_0[38:38], wg_0r0[38:38], conwig_0);
  AND2 I529 (conwgif_0[39:39], wg_0r0[39:39], conwig_0);
  AND2 I530 (conwgif_0[40:40], wg_0r0[40:40], conwig_0);
  AND2 I531 (conwgif_0[41:41], wg_0r0[41:41], conwig_0);
  AND2 I532 (conwgif_0[42:42], wg_0r0[42:42], conwig_0);
  AND2 I533 (conwgif_0[43:43], wg_0r0[43:43], conwig_0);
  AND2 I534 (conwgif_0[44:44], wg_0r0[44:44], conwig_0);
  AND2 I535 (conwgif_0[45:45], wg_0r0[45:45], conwig_0);
  AND2 I536 (conwgif_0[46:46], wg_0r0[46:46], conwig_0);
  AND2 I537 (conwgif_0[47:47], wg_0r0[47:47], conwig_0);
  AND2 I538 (conwgif_0[48:48], wg_0r0[48:48], conwig_0);
  AND2 I539 (conwgif_0[49:49], wg_0r0[49:49], conwig_0);
  AND2 I540 (conwgif_0[50:50], wg_0r0[50:50], conwig_0);
  AND2 I541 (conwgif_0[51:51], wg_0r0[51:51], conwig_0);
  AND2 I542 (conwgif_0[52:52], wg_0r0[52:52], conwig_0);
  AND2 I543 (conwgif_0[53:53], wg_0r0[53:53], conwig_0);
  AND2 I544 (conwgif_0[54:54], wg_0r0[54:54], conwig_0);
  AND2 I545 (conwgif_0[55:55], wg_0r0[55:55], conwig_0);
  AND2 I546 (conwgif_0[56:56], wg_0r0[56:56], conwig_0);
  AND2 I547 (conwgif_0[57:57], wg_0r0[57:57], conwig_0);
  AND2 I548 (conwgif_0[58:58], wg_0r0[58:58], conwig_0);
  AND2 I549 (conwgif_0[59:59], wg_0r0[59:59], conwig_0);
  AND2 I550 (conwgif_0[60:60], wg_0r0[60:60], conwig_0);
  AND2 I551 (conwgif_0[61:61], wg_0r0[61:61], conwig_0);
  AND2 I552 (conwgif_0[62:62], wg_0r0[62:62], conwig_0);
  AND2 I553 (conwgif_0[63:63], wg_0r0[63:63], conwig_0);
  AND2 I554 (conwgif_0[64:64], wg_0r0[64:64], conwig_0);
  AND2 I555 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I556 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I557 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I558 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I559 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I560 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I561 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I562 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I563 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I564 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I565 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I566 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I567 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I568 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I569 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I570 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I571 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I572 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I573 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I574 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I575 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I576 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I577 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I578 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I579 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I580 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I581 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I582 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I583 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I584 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I585 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I586 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  AND2 I587 (conwgit_0[32:32], wg_0r1[32:32], conwig_0);
  AND2 I588 (conwgit_0[33:33], wg_0r1[33:33], conwig_0);
  AND2 I589 (conwgit_0[34:34], wg_0r1[34:34], conwig_0);
  AND2 I590 (conwgit_0[35:35], wg_0r1[35:35], conwig_0);
  AND2 I591 (conwgit_0[36:36], wg_0r1[36:36], conwig_0);
  AND2 I592 (conwgit_0[37:37], wg_0r1[37:37], conwig_0);
  AND2 I593 (conwgit_0[38:38], wg_0r1[38:38], conwig_0);
  AND2 I594 (conwgit_0[39:39], wg_0r1[39:39], conwig_0);
  AND2 I595 (conwgit_0[40:40], wg_0r1[40:40], conwig_0);
  AND2 I596 (conwgit_0[41:41], wg_0r1[41:41], conwig_0);
  AND2 I597 (conwgit_0[42:42], wg_0r1[42:42], conwig_0);
  AND2 I598 (conwgit_0[43:43], wg_0r1[43:43], conwig_0);
  AND2 I599 (conwgit_0[44:44], wg_0r1[44:44], conwig_0);
  AND2 I600 (conwgit_0[45:45], wg_0r1[45:45], conwig_0);
  AND2 I601 (conwgit_0[46:46], wg_0r1[46:46], conwig_0);
  AND2 I602 (conwgit_0[47:47], wg_0r1[47:47], conwig_0);
  AND2 I603 (conwgit_0[48:48], wg_0r1[48:48], conwig_0);
  AND2 I604 (conwgit_0[49:49], wg_0r1[49:49], conwig_0);
  AND2 I605 (conwgit_0[50:50], wg_0r1[50:50], conwig_0);
  AND2 I606 (conwgit_0[51:51], wg_0r1[51:51], conwig_0);
  AND2 I607 (conwgit_0[52:52], wg_0r1[52:52], conwig_0);
  AND2 I608 (conwgit_0[53:53], wg_0r1[53:53], conwig_0);
  AND2 I609 (conwgit_0[54:54], wg_0r1[54:54], conwig_0);
  AND2 I610 (conwgit_0[55:55], wg_0r1[55:55], conwig_0);
  AND2 I611 (conwgit_0[56:56], wg_0r1[56:56], conwig_0);
  AND2 I612 (conwgit_0[57:57], wg_0r1[57:57], conwig_0);
  AND2 I613 (conwgit_0[58:58], wg_0r1[58:58], conwig_0);
  AND2 I614 (conwgit_0[59:59], wg_0r1[59:59], conwig_0);
  AND2 I615 (conwgit_0[60:60], wg_0r1[60:60], conwig_0);
  AND2 I616 (conwgit_0[61:61], wg_0r1[61:61], conwig_0);
  AND2 I617 (conwgit_0[62:62], wg_0r1[62:62], conwig_0);
  AND2 I618 (conwgit_0[63:63], wg_0r1[63:63], conwig_0);
  AND2 I619 (conwgit_0[64:64], wg_0r1[64:64], conwig_0);
  BUFF I620 (conwigc_0, wc_0);
  AO22 I621 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I622 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I623 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I624 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I625 (wenr_0[0:0], wc_0);
  BUFF I626 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I627 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I628 (wenr_0[1:1], wc_0);
  BUFF I629 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I630 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I631 (wenr_0[2:2], wc_0);
  BUFF I632 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I633 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I634 (wenr_0[3:3], wc_0);
  BUFF I635 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I636 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I637 (wenr_0[4:4], wc_0);
  BUFF I638 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I639 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I640 (wenr_0[5:5], wc_0);
  BUFF I641 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I642 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I643 (wenr_0[6:6], wc_0);
  BUFF I644 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I645 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I646 (wenr_0[7:7], wc_0);
  BUFF I647 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I648 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I649 (wenr_0[8:8], wc_0);
  BUFF I650 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I651 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I652 (wenr_0[9:9], wc_0);
  BUFF I653 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I654 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I655 (wenr_0[10:10], wc_0);
  BUFF I656 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I657 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I658 (wenr_0[11:11], wc_0);
  BUFF I659 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I660 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I661 (wenr_0[12:12], wc_0);
  BUFF I662 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I663 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I664 (wenr_0[13:13], wc_0);
  BUFF I665 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I666 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I667 (wenr_0[14:14], wc_0);
  BUFF I668 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I669 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I670 (wenr_0[15:15], wc_0);
  BUFF I671 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I672 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I673 (wenr_0[16:16], wc_0);
  BUFF I674 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I675 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I676 (wenr_0[17:17], wc_0);
  BUFF I677 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I678 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I679 (wenr_0[18:18], wc_0);
  BUFF I680 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I681 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I682 (wenr_0[19:19], wc_0);
  BUFF I683 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I684 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I685 (wenr_0[20:20], wc_0);
  BUFF I686 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I687 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I688 (wenr_0[21:21], wc_0);
  BUFF I689 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I690 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I691 (wenr_0[22:22], wc_0);
  BUFF I692 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I693 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I694 (wenr_0[23:23], wc_0);
  BUFF I695 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I696 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I697 (wenr_0[24:24], wc_0);
  BUFF I698 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I699 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I700 (wenr_0[25:25], wc_0);
  BUFF I701 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I702 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I703 (wenr_0[26:26], wc_0);
  BUFF I704 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I705 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I706 (wenr_0[27:27], wc_0);
  BUFF I707 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I708 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I709 (wenr_0[28:28], wc_0);
  BUFF I710 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I711 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I712 (wenr_0[29:29], wc_0);
  BUFF I713 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I714 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I715 (wenr_0[30:30], wc_0);
  BUFF I716 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I717 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I718 (wenr_0[31:31], wc_0);
  BUFF I719 (wf_0[32:32], conwgif_0[32:32]);
  BUFF I720 (wt_0[32:32], conwgit_0[32:32]);
  BUFF I721 (wenr_0[32:32], wc_0);
  BUFF I722 (wf_0[33:33], conwgif_0[33:33]);
  BUFF I723 (wt_0[33:33], conwgit_0[33:33]);
  BUFF I724 (wenr_0[33:33], wc_0);
  BUFF I725 (wf_0[34:34], conwgif_0[34:34]);
  BUFF I726 (wt_0[34:34], conwgit_0[34:34]);
  BUFF I727 (wenr_0[34:34], wc_0);
  BUFF I728 (wf_0[35:35], conwgif_0[35:35]);
  BUFF I729 (wt_0[35:35], conwgit_0[35:35]);
  BUFF I730 (wenr_0[35:35], wc_0);
  BUFF I731 (wf_0[36:36], conwgif_0[36:36]);
  BUFF I732 (wt_0[36:36], conwgit_0[36:36]);
  BUFF I733 (wenr_0[36:36], wc_0);
  BUFF I734 (wf_0[37:37], conwgif_0[37:37]);
  BUFF I735 (wt_0[37:37], conwgit_0[37:37]);
  BUFF I736 (wenr_0[37:37], wc_0);
  BUFF I737 (wf_0[38:38], conwgif_0[38:38]);
  BUFF I738 (wt_0[38:38], conwgit_0[38:38]);
  BUFF I739 (wenr_0[38:38], wc_0);
  BUFF I740 (wf_0[39:39], conwgif_0[39:39]);
  BUFF I741 (wt_0[39:39], conwgit_0[39:39]);
  BUFF I742 (wenr_0[39:39], wc_0);
  BUFF I743 (wf_0[40:40], conwgif_0[40:40]);
  BUFF I744 (wt_0[40:40], conwgit_0[40:40]);
  BUFF I745 (wenr_0[40:40], wc_0);
  BUFF I746 (wf_0[41:41], conwgif_0[41:41]);
  BUFF I747 (wt_0[41:41], conwgit_0[41:41]);
  BUFF I748 (wenr_0[41:41], wc_0);
  BUFF I749 (wf_0[42:42], conwgif_0[42:42]);
  BUFF I750 (wt_0[42:42], conwgit_0[42:42]);
  BUFF I751 (wenr_0[42:42], wc_0);
  BUFF I752 (wf_0[43:43], conwgif_0[43:43]);
  BUFF I753 (wt_0[43:43], conwgit_0[43:43]);
  BUFF I754 (wenr_0[43:43], wc_0);
  BUFF I755 (wf_0[44:44], conwgif_0[44:44]);
  BUFF I756 (wt_0[44:44], conwgit_0[44:44]);
  BUFF I757 (wenr_0[44:44], wc_0);
  BUFF I758 (wf_0[45:45], conwgif_0[45:45]);
  BUFF I759 (wt_0[45:45], conwgit_0[45:45]);
  BUFF I760 (wenr_0[45:45], wc_0);
  BUFF I761 (wf_0[46:46], conwgif_0[46:46]);
  BUFF I762 (wt_0[46:46], conwgit_0[46:46]);
  BUFF I763 (wenr_0[46:46], wc_0);
  BUFF I764 (wf_0[47:47], conwgif_0[47:47]);
  BUFF I765 (wt_0[47:47], conwgit_0[47:47]);
  BUFF I766 (wenr_0[47:47], wc_0);
  BUFF I767 (wf_0[48:48], conwgif_0[48:48]);
  BUFF I768 (wt_0[48:48], conwgit_0[48:48]);
  BUFF I769 (wenr_0[48:48], wc_0);
  BUFF I770 (wf_0[49:49], conwgif_0[49:49]);
  BUFF I771 (wt_0[49:49], conwgit_0[49:49]);
  BUFF I772 (wenr_0[49:49], wc_0);
  BUFF I773 (wf_0[50:50], conwgif_0[50:50]);
  BUFF I774 (wt_0[50:50], conwgit_0[50:50]);
  BUFF I775 (wenr_0[50:50], wc_0);
  BUFF I776 (wf_0[51:51], conwgif_0[51:51]);
  BUFF I777 (wt_0[51:51], conwgit_0[51:51]);
  BUFF I778 (wenr_0[51:51], wc_0);
  BUFF I779 (wf_0[52:52], conwgif_0[52:52]);
  BUFF I780 (wt_0[52:52], conwgit_0[52:52]);
  BUFF I781 (wenr_0[52:52], wc_0);
  BUFF I782 (wf_0[53:53], conwgif_0[53:53]);
  BUFF I783 (wt_0[53:53], conwgit_0[53:53]);
  BUFF I784 (wenr_0[53:53], wc_0);
  BUFF I785 (wf_0[54:54], conwgif_0[54:54]);
  BUFF I786 (wt_0[54:54], conwgit_0[54:54]);
  BUFF I787 (wenr_0[54:54], wc_0);
  BUFF I788 (wf_0[55:55], conwgif_0[55:55]);
  BUFF I789 (wt_0[55:55], conwgit_0[55:55]);
  BUFF I790 (wenr_0[55:55], wc_0);
  BUFF I791 (wf_0[56:56], conwgif_0[56:56]);
  BUFF I792 (wt_0[56:56], conwgit_0[56:56]);
  BUFF I793 (wenr_0[56:56], wc_0);
  BUFF I794 (wf_0[57:57], conwgif_0[57:57]);
  BUFF I795 (wt_0[57:57], conwgit_0[57:57]);
  BUFF I796 (wenr_0[57:57], wc_0);
  BUFF I797 (wf_0[58:58], conwgif_0[58:58]);
  BUFF I798 (wt_0[58:58], conwgit_0[58:58]);
  BUFF I799 (wenr_0[58:58], wc_0);
  BUFF I800 (wf_0[59:59], conwgif_0[59:59]);
  BUFF I801 (wt_0[59:59], conwgit_0[59:59]);
  BUFF I802 (wenr_0[59:59], wc_0);
  BUFF I803 (wf_0[60:60], conwgif_0[60:60]);
  BUFF I804 (wt_0[60:60], conwgit_0[60:60]);
  BUFF I805 (wenr_0[60:60], wc_0);
  BUFF I806 (wf_0[61:61], conwgif_0[61:61]);
  BUFF I807 (wt_0[61:61], conwgit_0[61:61]);
  BUFF I808 (wenr_0[61:61], wc_0);
  BUFF I809 (wf_0[62:62], conwgif_0[62:62]);
  BUFF I810 (wt_0[62:62], conwgit_0[62:62]);
  BUFF I811 (wenr_0[62:62], wc_0);
  BUFF I812 (wf_0[63:63], conwgif_0[63:63]);
  BUFF I813 (wt_0[63:63], conwgit_0[63:63]);
  BUFF I814 (wenr_0[63:63], wc_0);
  BUFF I815 (wf_0[64:64], conwgif_0[64:64]);
  BUFF I816 (wt_0[64:64], conwgit_0[64:64]);
  BUFF I817 (wenr_0[64:64], wc_0);
  C3 I818 (simp8031_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I819 (simp8031_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I820 (simp8031_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I821 (simp8031_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I822 (simp8031_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I823 (simp8031_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I824 (simp8031_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I825 (simp8031_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I826 (simp8031_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I827 (simp8031_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I828 (simp8031_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I829 (simp8031_0[11:11], wacks_0[32:32], wacks_0[33:33], wacks_0[34:34]);
  C3 I830 (simp8031_0[12:12], wacks_0[35:35], wacks_0[36:36], wacks_0[37:37]);
  C3 I831 (simp8031_0[13:13], wacks_0[38:38], wacks_0[39:39], wacks_0[40:40]);
  C3 I832 (simp8031_0[14:14], wacks_0[41:41], wacks_0[42:42], wacks_0[43:43]);
  C3 I833 (simp8031_0[15:15], wacks_0[44:44], wacks_0[45:45], wacks_0[46:46]);
  C3 I834 (simp8031_0[16:16], wacks_0[47:47], wacks_0[48:48], wacks_0[49:49]);
  C3 I835 (simp8031_0[17:17], wacks_0[50:50], wacks_0[51:51], wacks_0[52:52]);
  C3 I836 (simp8031_0[18:18], wacks_0[53:53], wacks_0[54:54], wacks_0[55:55]);
  C3 I837 (simp8031_0[19:19], wacks_0[56:56], wacks_0[57:57], wacks_0[58:58]);
  C3 I838 (simp8031_0[20:20], wacks_0[59:59], wacks_0[60:60], wacks_0[61:61]);
  C3 I839 (simp8031_0[21:21], wacks_0[62:62], wacks_0[63:63], wacks_0[64:64]);
  C3 I840 (simp8032_0[0:0], simp8031_0[0:0], simp8031_0[1:1], simp8031_0[2:2]);
  C3 I841 (simp8032_0[1:1], simp8031_0[3:3], simp8031_0[4:4], simp8031_0[5:5]);
  C3 I842 (simp8032_0[2:2], simp8031_0[6:6], simp8031_0[7:7], simp8031_0[8:8]);
  C3 I843 (simp8032_0[3:3], simp8031_0[9:9], simp8031_0[10:10], simp8031_0[11:11]);
  C3 I844 (simp8032_0[4:4], simp8031_0[12:12], simp8031_0[13:13], simp8031_0[14:14]);
  C3 I845 (simp8032_0[5:5], simp8031_0[15:15], simp8031_0[16:16], simp8031_0[17:17]);
  C3 I846 (simp8032_0[6:6], simp8031_0[18:18], simp8031_0[19:19], simp8031_0[20:20]);
  BUFF I847 (simp8032_0[7:7], simp8031_0[21:21]);
  C3 I848 (simp8033_0[0:0], simp8032_0[0:0], simp8032_0[1:1], simp8032_0[2:2]);
  C3 I849 (simp8033_0[1:1], simp8032_0[3:3], simp8032_0[4:4], simp8032_0[5:5]);
  C2 I850 (simp8033_0[2:2], simp8032_0[6:6], simp8032_0[7:7]);
  C3 I851 (wd_0r, simp8033_0[0:0], simp8033_0[1:1], simp8033_0[2:2]);
  AND2 I852 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I853 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I854 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I855 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I856 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I857 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I858 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I859 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I860 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I861 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I862 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I863 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I864 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I865 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I866 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I867 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I868 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I869 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I870 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I871 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I872 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I873 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I874 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I875 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I876 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I877 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I878 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I879 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I880 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I881 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I882 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I883 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I884 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I885 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I886 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I887 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I888 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I889 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I890 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I891 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I892 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I893 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I894 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I895 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I896 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I897 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I898 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I899 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I900 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I901 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I902 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I903 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I904 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I905 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I906 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I907 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I908 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I909 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I910 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I911 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I912 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I913 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I914 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I915 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I916 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I917 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I918 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I919 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I920 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I921 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I922 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I923 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I924 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I925 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I926 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I927 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I928 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I929 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I930 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I931 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I932 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I933 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I934 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I935 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I936 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I937 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I938 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I939 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I940 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I941 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I942 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I943 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I944 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I945 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I946 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I947 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I948 (rd_3r0[0:0], df_0[0:0], rg_3r);
  AND2 I949 (rd_3r0[1:1], df_0[1:1], rg_3r);
  AND2 I950 (rd_3r0[2:2], df_0[2:2], rg_3r);
  AND2 I951 (rd_3r0[3:3], df_0[3:3], rg_3r);
  AND2 I952 (rd_3r0[4:4], df_0[4:4], rg_3r);
  AND2 I953 (rd_3r0[5:5], df_0[5:5], rg_3r);
  AND2 I954 (rd_3r0[6:6], df_0[6:6], rg_3r);
  AND2 I955 (rd_3r0[7:7], df_0[7:7], rg_3r);
  AND2 I956 (rd_3r0[8:8], df_0[8:8], rg_3r);
  AND2 I957 (rd_3r0[9:9], df_0[9:9], rg_3r);
  AND2 I958 (rd_3r0[10:10], df_0[10:10], rg_3r);
  AND2 I959 (rd_3r0[11:11], df_0[11:11], rg_3r);
  AND2 I960 (rd_3r0[12:12], df_0[12:12], rg_3r);
  AND2 I961 (rd_3r0[13:13], df_0[13:13], rg_3r);
  AND2 I962 (rd_3r0[14:14], df_0[14:14], rg_3r);
  AND2 I963 (rd_3r0[15:15], df_0[15:15], rg_3r);
  AND2 I964 (rd_3r0[16:16], df_0[16:16], rg_3r);
  AND2 I965 (rd_3r0[17:17], df_0[17:17], rg_3r);
  AND2 I966 (rd_3r0[18:18], df_0[18:18], rg_3r);
  AND2 I967 (rd_3r0[19:19], df_0[19:19], rg_3r);
  AND2 I968 (rd_3r0[20:20], df_0[20:20], rg_3r);
  AND2 I969 (rd_3r0[21:21], df_0[21:21], rg_3r);
  AND2 I970 (rd_3r0[22:22], df_0[22:22], rg_3r);
  AND2 I971 (rd_3r0[23:23], df_0[23:23], rg_3r);
  AND2 I972 (rd_3r0[24:24], df_0[24:24], rg_3r);
  AND2 I973 (rd_3r0[25:25], df_0[25:25], rg_3r);
  AND2 I974 (rd_3r0[26:26], df_0[26:26], rg_3r);
  AND2 I975 (rd_3r0[27:27], df_0[27:27], rg_3r);
  AND2 I976 (rd_3r0[28:28], df_0[28:28], rg_3r);
  AND2 I977 (rd_3r0[29:29], df_0[29:29], rg_3r);
  AND2 I978 (rd_3r0[30:30], df_0[30:30], rg_3r);
  AND2 I979 (rd_3r0[31:31], df_0[31:31], rg_3r);
  AND2 I980 (rd_4r0[0:0], df_0[32:32], rg_4r);
  AND2 I981 (rd_4r0[1:1], df_0[33:33], rg_4r);
  AND2 I982 (rd_4r0[2:2], df_0[34:34], rg_4r);
  AND2 I983 (rd_4r0[3:3], df_0[35:35], rg_4r);
  AND2 I984 (rd_4r0[4:4], df_0[36:36], rg_4r);
  AND2 I985 (rd_4r0[5:5], df_0[37:37], rg_4r);
  AND2 I986 (rd_4r0[6:6], df_0[38:38], rg_4r);
  AND2 I987 (rd_4r0[7:7], df_0[39:39], rg_4r);
  AND2 I988 (rd_4r0[8:8], df_0[40:40], rg_4r);
  AND2 I989 (rd_4r0[9:9], df_0[41:41], rg_4r);
  AND2 I990 (rd_4r0[10:10], df_0[42:42], rg_4r);
  AND2 I991 (rd_4r0[11:11], df_0[43:43], rg_4r);
  AND2 I992 (rd_4r0[12:12], df_0[44:44], rg_4r);
  AND2 I993 (rd_4r0[13:13], df_0[45:45], rg_4r);
  AND2 I994 (rd_4r0[14:14], df_0[46:46], rg_4r);
  AND2 I995 (rd_4r0[15:15], df_0[47:47], rg_4r);
  AND2 I996 (rd_4r0[16:16], df_0[48:48], rg_4r);
  AND2 I997 (rd_4r0[17:17], df_0[49:49], rg_4r);
  AND2 I998 (rd_4r0[18:18], df_0[50:50], rg_4r);
  AND2 I999 (rd_4r0[19:19], df_0[51:51], rg_4r);
  AND2 I1000 (rd_4r0[20:20], df_0[52:52], rg_4r);
  AND2 I1001 (rd_4r0[21:21], df_0[53:53], rg_4r);
  AND2 I1002 (rd_4r0[22:22], df_0[54:54], rg_4r);
  AND2 I1003 (rd_4r0[23:23], df_0[55:55], rg_4r);
  AND2 I1004 (rd_4r0[24:24], df_0[56:56], rg_4r);
  AND2 I1005 (rd_4r0[25:25], df_0[57:57], rg_4r);
  AND2 I1006 (rd_4r0[26:26], df_0[58:58], rg_4r);
  AND2 I1007 (rd_4r0[27:27], df_0[59:59], rg_4r);
  AND2 I1008 (rd_4r0[28:28], df_0[60:60], rg_4r);
  AND2 I1009 (rd_4r0[29:29], df_0[61:61], rg_4r);
  AND2 I1010 (rd_4r0[30:30], df_0[62:62], rg_4r);
  AND2 I1011 (rd_4r0[31:31], df_0[63:63], rg_4r);
  AND2 I1012 (rd_5r0[0:0], df_0[32:32], rg_5r);
  AND2 I1013 (rd_5r0[1:1], df_0[33:33], rg_5r);
  AND2 I1014 (rd_5r0[2:2], df_0[34:34], rg_5r);
  AND2 I1015 (rd_5r0[3:3], df_0[35:35], rg_5r);
  AND2 I1016 (rd_5r0[4:4], df_0[36:36], rg_5r);
  AND2 I1017 (rd_5r0[5:5], df_0[37:37], rg_5r);
  AND2 I1018 (rd_5r0[6:6], df_0[38:38], rg_5r);
  AND2 I1019 (rd_5r0[7:7], df_0[39:39], rg_5r);
  AND2 I1020 (rd_5r0[8:8], df_0[40:40], rg_5r);
  AND2 I1021 (rd_5r0[9:9], df_0[41:41], rg_5r);
  AND2 I1022 (rd_5r0[10:10], df_0[42:42], rg_5r);
  AND2 I1023 (rd_5r0[11:11], df_0[43:43], rg_5r);
  AND2 I1024 (rd_5r0[12:12], df_0[44:44], rg_5r);
  AND2 I1025 (rd_5r0[13:13], df_0[45:45], rg_5r);
  AND2 I1026 (rd_5r0[14:14], df_0[46:46], rg_5r);
  AND2 I1027 (rd_5r0[15:15], df_0[47:47], rg_5r);
  AND2 I1028 (rd_5r0[16:16], df_0[48:48], rg_5r);
  AND2 I1029 (rd_5r0[17:17], df_0[49:49], rg_5r);
  AND2 I1030 (rd_5r0[18:18], df_0[50:50], rg_5r);
  AND2 I1031 (rd_5r0[19:19], df_0[51:51], rg_5r);
  AND2 I1032 (rd_5r0[20:20], df_0[52:52], rg_5r);
  AND2 I1033 (rd_5r0[21:21], df_0[53:53], rg_5r);
  AND2 I1034 (rd_5r0[22:22], df_0[54:54], rg_5r);
  AND2 I1035 (rd_5r0[23:23], df_0[55:55], rg_5r);
  AND2 I1036 (rd_5r0[24:24], df_0[56:56], rg_5r);
  AND2 I1037 (rd_5r0[25:25], df_0[57:57], rg_5r);
  AND2 I1038 (rd_5r0[26:26], df_0[58:58], rg_5r);
  AND2 I1039 (rd_5r0[27:27], df_0[59:59], rg_5r);
  AND2 I1040 (rd_5r0[28:28], df_0[60:60], rg_5r);
  AND2 I1041 (rd_5r0[29:29], df_0[61:61], rg_5r);
  AND2 I1042 (rd_5r0[30:30], df_0[62:62], rg_5r);
  AND2 I1043 (rd_5r0[31:31], df_0[63:63], rg_5r);
  AND2 I1044 (rd_6r0[0:0], df_0[32:32], rg_6r);
  AND2 I1045 (rd_6r0[1:1], df_0[33:33], rg_6r);
  AND2 I1046 (rd_6r0[2:2], df_0[34:34], rg_6r);
  AND2 I1047 (rd_6r0[3:3], df_0[35:35], rg_6r);
  AND2 I1048 (rd_6r0[4:4], df_0[36:36], rg_6r);
  AND2 I1049 (rd_6r0[5:5], df_0[37:37], rg_6r);
  AND2 I1050 (rd_6r0[6:6], df_0[38:38], rg_6r);
  AND2 I1051 (rd_6r0[7:7], df_0[39:39], rg_6r);
  AND2 I1052 (rd_6r0[8:8], df_0[40:40], rg_6r);
  AND2 I1053 (rd_6r0[9:9], df_0[41:41], rg_6r);
  AND2 I1054 (rd_6r0[10:10], df_0[42:42], rg_6r);
  AND2 I1055 (rd_6r0[11:11], df_0[43:43], rg_6r);
  AND2 I1056 (rd_6r0[12:12], df_0[44:44], rg_6r);
  AND2 I1057 (rd_6r0[13:13], df_0[45:45], rg_6r);
  AND2 I1058 (rd_6r0[14:14], df_0[46:46], rg_6r);
  AND2 I1059 (rd_6r0[15:15], df_0[47:47], rg_6r);
  AND2 I1060 (rd_6r0[16:16], df_0[48:48], rg_6r);
  AND2 I1061 (rd_6r0[17:17], df_0[49:49], rg_6r);
  AND2 I1062 (rd_6r0[18:18], df_0[50:50], rg_6r);
  AND2 I1063 (rd_6r0[19:19], df_0[51:51], rg_6r);
  AND2 I1064 (rd_6r0[20:20], df_0[52:52], rg_6r);
  AND2 I1065 (rd_6r0[21:21], df_0[53:53], rg_6r);
  AND2 I1066 (rd_6r0[22:22], df_0[54:54], rg_6r);
  AND2 I1067 (rd_6r0[23:23], df_0[55:55], rg_6r);
  AND2 I1068 (rd_6r0[24:24], df_0[56:56], rg_6r);
  AND2 I1069 (rd_6r0[25:25], df_0[57:57], rg_6r);
  AND2 I1070 (rd_6r0[26:26], df_0[58:58], rg_6r);
  AND2 I1071 (rd_6r0[27:27], df_0[59:59], rg_6r);
  AND2 I1072 (rd_6r0[28:28], df_0[60:60], rg_6r);
  AND2 I1073 (rd_6r0[29:29], df_0[61:61], rg_6r);
  AND2 I1074 (rd_6r0[30:30], df_0[62:62], rg_6r);
  AND2 I1075 (rd_6r0[31:31], df_0[63:63], rg_6r);
  AND2 I1076 (rd_7r0[0:0], df_0[32:32], rg_7r);
  AND2 I1077 (rd_7r0[1:1], df_0[33:33], rg_7r);
  AND2 I1078 (rd_7r0[2:2], df_0[34:34], rg_7r);
  AND2 I1079 (rd_7r0[3:3], df_0[35:35], rg_7r);
  AND2 I1080 (rd_7r0[4:4], df_0[36:36], rg_7r);
  AND2 I1081 (rd_7r0[5:5], df_0[37:37], rg_7r);
  AND2 I1082 (rd_7r0[6:6], df_0[38:38], rg_7r);
  AND2 I1083 (rd_7r0[7:7], df_0[39:39], rg_7r);
  AND2 I1084 (rd_7r0[8:8], df_0[40:40], rg_7r);
  AND2 I1085 (rd_7r0[9:9], df_0[41:41], rg_7r);
  AND2 I1086 (rd_7r0[10:10], df_0[42:42], rg_7r);
  AND2 I1087 (rd_7r0[11:11], df_0[43:43], rg_7r);
  AND2 I1088 (rd_7r0[12:12], df_0[44:44], rg_7r);
  AND2 I1089 (rd_7r0[13:13], df_0[45:45], rg_7r);
  AND2 I1090 (rd_7r0[14:14], df_0[46:46], rg_7r);
  AND2 I1091 (rd_7r0[15:15], df_0[47:47], rg_7r);
  AND2 I1092 (rd_7r0[16:16], df_0[48:48], rg_7r);
  AND2 I1093 (rd_7r0[17:17], df_0[49:49], rg_7r);
  AND2 I1094 (rd_7r0[18:18], df_0[50:50], rg_7r);
  AND2 I1095 (rd_7r0[19:19], df_0[51:51], rg_7r);
  AND2 I1096 (rd_7r0[20:20], df_0[52:52], rg_7r);
  AND2 I1097 (rd_7r0[21:21], df_0[53:53], rg_7r);
  AND2 I1098 (rd_7r0[22:22], df_0[54:54], rg_7r);
  AND2 I1099 (rd_7r0[23:23], df_0[55:55], rg_7r);
  AND2 I1100 (rd_7r0[24:24], df_0[56:56], rg_7r);
  AND2 I1101 (rd_7r0[25:25], df_0[57:57], rg_7r);
  AND2 I1102 (rd_7r0[26:26], df_0[58:58], rg_7r);
  AND2 I1103 (rd_7r0[27:27], df_0[59:59], rg_7r);
  AND2 I1104 (rd_7r0[28:28], df_0[60:60], rg_7r);
  AND2 I1105 (rd_7r0[29:29], df_0[61:61], rg_7r);
  AND2 I1106 (rd_7r0[30:30], df_0[62:62], rg_7r);
  AND2 I1107 (rd_7r0[31:31], df_0[63:63], rg_7r);
  AND2 I1108 (rd_8r0[0:0], df_0[32:32], rg_8r);
  AND2 I1109 (rd_8r0[1:1], df_0[33:33], rg_8r);
  AND2 I1110 (rd_8r0[2:2], df_0[34:34], rg_8r);
  AND2 I1111 (rd_8r0[3:3], df_0[35:35], rg_8r);
  AND2 I1112 (rd_8r0[4:4], df_0[36:36], rg_8r);
  AND2 I1113 (rd_8r0[5:5], df_0[37:37], rg_8r);
  AND2 I1114 (rd_8r0[6:6], df_0[38:38], rg_8r);
  AND2 I1115 (rd_8r0[7:7], df_0[39:39], rg_8r);
  AND2 I1116 (rd_8r0[8:8], df_0[40:40], rg_8r);
  AND2 I1117 (rd_8r0[9:9], df_0[41:41], rg_8r);
  AND2 I1118 (rd_8r0[10:10], df_0[42:42], rg_8r);
  AND2 I1119 (rd_8r0[11:11], df_0[43:43], rg_8r);
  AND2 I1120 (rd_8r0[12:12], df_0[44:44], rg_8r);
  AND2 I1121 (rd_8r0[13:13], df_0[45:45], rg_8r);
  AND2 I1122 (rd_8r0[14:14], df_0[46:46], rg_8r);
  AND2 I1123 (rd_8r0[15:15], df_0[47:47], rg_8r);
  AND2 I1124 (rd_8r0[16:16], df_0[48:48], rg_8r);
  AND2 I1125 (rd_8r0[17:17], df_0[49:49], rg_8r);
  AND2 I1126 (rd_8r0[18:18], df_0[50:50], rg_8r);
  AND2 I1127 (rd_8r0[19:19], df_0[51:51], rg_8r);
  AND2 I1128 (rd_8r0[20:20], df_0[52:52], rg_8r);
  AND2 I1129 (rd_8r0[21:21], df_0[53:53], rg_8r);
  AND2 I1130 (rd_8r0[22:22], df_0[54:54], rg_8r);
  AND2 I1131 (rd_8r0[23:23], df_0[55:55], rg_8r);
  AND2 I1132 (rd_8r0[24:24], df_0[56:56], rg_8r);
  AND2 I1133 (rd_8r0[25:25], df_0[57:57], rg_8r);
  AND2 I1134 (rd_8r0[26:26], df_0[58:58], rg_8r);
  AND2 I1135 (rd_8r0[27:27], df_0[59:59], rg_8r);
  AND2 I1136 (rd_8r0[28:28], df_0[60:60], rg_8r);
  AND2 I1137 (rd_8r0[29:29], df_0[61:61], rg_8r);
  AND2 I1138 (rd_8r0[30:30], df_0[62:62], rg_8r);
  AND2 I1139 (rd_8r0[31:31], df_0[63:63], rg_8r);
  AND2 I1140 (rd_9r0, df_0[64:64], rg_9r);
  AND2 I1141 (rd_10r0, df_0[64:64], rg_10r);
  AND2 I1142 (rd_11r0, df_0[64:64], rg_11r);
  AND2 I1143 (rd_12r0, df_0[64:64], rg_12r);
  AND2 I1144 (rd_13r0, df_0[64:64], rg_13r);
  AND2 I1145 (rd_14r0, df_0[64:64], rg_14r);
  AND2 I1146 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I1147 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I1148 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I1149 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I1150 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I1151 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I1152 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I1153 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I1154 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I1155 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I1156 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I1157 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I1158 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I1159 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I1160 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I1161 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I1162 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I1163 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I1164 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I1165 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I1166 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I1167 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I1168 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I1169 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I1170 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I1171 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I1172 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I1173 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I1174 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I1175 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I1176 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I1177 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I1178 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I1179 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I1180 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I1181 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I1182 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I1183 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I1184 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I1185 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I1186 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I1187 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I1188 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I1189 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I1190 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I1191 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I1192 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I1193 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I1194 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I1195 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I1196 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I1197 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I1198 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I1199 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I1200 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I1201 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I1202 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I1203 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I1204 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I1205 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I1206 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I1207 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I1208 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I1209 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I1210 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I1211 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I1212 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I1213 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I1214 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I1215 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I1216 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I1217 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I1218 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I1219 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I1220 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I1221 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I1222 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I1223 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I1224 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I1225 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I1226 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I1227 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I1228 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I1229 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I1230 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I1231 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I1232 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I1233 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I1234 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I1235 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I1236 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I1237 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I1238 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I1239 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I1240 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I1241 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  AND2 I1242 (rd_3r1[0:0], dt_0[0:0], rg_3r);
  AND2 I1243 (rd_3r1[1:1], dt_0[1:1], rg_3r);
  AND2 I1244 (rd_3r1[2:2], dt_0[2:2], rg_3r);
  AND2 I1245 (rd_3r1[3:3], dt_0[3:3], rg_3r);
  AND2 I1246 (rd_3r1[4:4], dt_0[4:4], rg_3r);
  AND2 I1247 (rd_3r1[5:5], dt_0[5:5], rg_3r);
  AND2 I1248 (rd_3r1[6:6], dt_0[6:6], rg_3r);
  AND2 I1249 (rd_3r1[7:7], dt_0[7:7], rg_3r);
  AND2 I1250 (rd_3r1[8:8], dt_0[8:8], rg_3r);
  AND2 I1251 (rd_3r1[9:9], dt_0[9:9], rg_3r);
  AND2 I1252 (rd_3r1[10:10], dt_0[10:10], rg_3r);
  AND2 I1253 (rd_3r1[11:11], dt_0[11:11], rg_3r);
  AND2 I1254 (rd_3r1[12:12], dt_0[12:12], rg_3r);
  AND2 I1255 (rd_3r1[13:13], dt_0[13:13], rg_3r);
  AND2 I1256 (rd_3r1[14:14], dt_0[14:14], rg_3r);
  AND2 I1257 (rd_3r1[15:15], dt_0[15:15], rg_3r);
  AND2 I1258 (rd_3r1[16:16], dt_0[16:16], rg_3r);
  AND2 I1259 (rd_3r1[17:17], dt_0[17:17], rg_3r);
  AND2 I1260 (rd_3r1[18:18], dt_0[18:18], rg_3r);
  AND2 I1261 (rd_3r1[19:19], dt_0[19:19], rg_3r);
  AND2 I1262 (rd_3r1[20:20], dt_0[20:20], rg_3r);
  AND2 I1263 (rd_3r1[21:21], dt_0[21:21], rg_3r);
  AND2 I1264 (rd_3r1[22:22], dt_0[22:22], rg_3r);
  AND2 I1265 (rd_3r1[23:23], dt_0[23:23], rg_3r);
  AND2 I1266 (rd_3r1[24:24], dt_0[24:24], rg_3r);
  AND2 I1267 (rd_3r1[25:25], dt_0[25:25], rg_3r);
  AND2 I1268 (rd_3r1[26:26], dt_0[26:26], rg_3r);
  AND2 I1269 (rd_3r1[27:27], dt_0[27:27], rg_3r);
  AND2 I1270 (rd_3r1[28:28], dt_0[28:28], rg_3r);
  AND2 I1271 (rd_3r1[29:29], dt_0[29:29], rg_3r);
  AND2 I1272 (rd_3r1[30:30], dt_0[30:30], rg_3r);
  AND2 I1273 (rd_3r1[31:31], dt_0[31:31], rg_3r);
  AND2 I1274 (rd_4r1[0:0], dt_0[32:32], rg_4r);
  AND2 I1275 (rd_4r1[1:1], dt_0[33:33], rg_4r);
  AND2 I1276 (rd_4r1[2:2], dt_0[34:34], rg_4r);
  AND2 I1277 (rd_4r1[3:3], dt_0[35:35], rg_4r);
  AND2 I1278 (rd_4r1[4:4], dt_0[36:36], rg_4r);
  AND2 I1279 (rd_4r1[5:5], dt_0[37:37], rg_4r);
  AND2 I1280 (rd_4r1[6:6], dt_0[38:38], rg_4r);
  AND2 I1281 (rd_4r1[7:7], dt_0[39:39], rg_4r);
  AND2 I1282 (rd_4r1[8:8], dt_0[40:40], rg_4r);
  AND2 I1283 (rd_4r1[9:9], dt_0[41:41], rg_4r);
  AND2 I1284 (rd_4r1[10:10], dt_0[42:42], rg_4r);
  AND2 I1285 (rd_4r1[11:11], dt_0[43:43], rg_4r);
  AND2 I1286 (rd_4r1[12:12], dt_0[44:44], rg_4r);
  AND2 I1287 (rd_4r1[13:13], dt_0[45:45], rg_4r);
  AND2 I1288 (rd_4r1[14:14], dt_0[46:46], rg_4r);
  AND2 I1289 (rd_4r1[15:15], dt_0[47:47], rg_4r);
  AND2 I1290 (rd_4r1[16:16], dt_0[48:48], rg_4r);
  AND2 I1291 (rd_4r1[17:17], dt_0[49:49], rg_4r);
  AND2 I1292 (rd_4r1[18:18], dt_0[50:50], rg_4r);
  AND2 I1293 (rd_4r1[19:19], dt_0[51:51], rg_4r);
  AND2 I1294 (rd_4r1[20:20], dt_0[52:52], rg_4r);
  AND2 I1295 (rd_4r1[21:21], dt_0[53:53], rg_4r);
  AND2 I1296 (rd_4r1[22:22], dt_0[54:54], rg_4r);
  AND2 I1297 (rd_4r1[23:23], dt_0[55:55], rg_4r);
  AND2 I1298 (rd_4r1[24:24], dt_0[56:56], rg_4r);
  AND2 I1299 (rd_4r1[25:25], dt_0[57:57], rg_4r);
  AND2 I1300 (rd_4r1[26:26], dt_0[58:58], rg_4r);
  AND2 I1301 (rd_4r1[27:27], dt_0[59:59], rg_4r);
  AND2 I1302 (rd_4r1[28:28], dt_0[60:60], rg_4r);
  AND2 I1303 (rd_4r1[29:29], dt_0[61:61], rg_4r);
  AND2 I1304 (rd_4r1[30:30], dt_0[62:62], rg_4r);
  AND2 I1305 (rd_4r1[31:31], dt_0[63:63], rg_4r);
  AND2 I1306 (rd_5r1[0:0], dt_0[32:32], rg_5r);
  AND2 I1307 (rd_5r1[1:1], dt_0[33:33], rg_5r);
  AND2 I1308 (rd_5r1[2:2], dt_0[34:34], rg_5r);
  AND2 I1309 (rd_5r1[3:3], dt_0[35:35], rg_5r);
  AND2 I1310 (rd_5r1[4:4], dt_0[36:36], rg_5r);
  AND2 I1311 (rd_5r1[5:5], dt_0[37:37], rg_5r);
  AND2 I1312 (rd_5r1[6:6], dt_0[38:38], rg_5r);
  AND2 I1313 (rd_5r1[7:7], dt_0[39:39], rg_5r);
  AND2 I1314 (rd_5r1[8:8], dt_0[40:40], rg_5r);
  AND2 I1315 (rd_5r1[9:9], dt_0[41:41], rg_5r);
  AND2 I1316 (rd_5r1[10:10], dt_0[42:42], rg_5r);
  AND2 I1317 (rd_5r1[11:11], dt_0[43:43], rg_5r);
  AND2 I1318 (rd_5r1[12:12], dt_0[44:44], rg_5r);
  AND2 I1319 (rd_5r1[13:13], dt_0[45:45], rg_5r);
  AND2 I1320 (rd_5r1[14:14], dt_0[46:46], rg_5r);
  AND2 I1321 (rd_5r1[15:15], dt_0[47:47], rg_5r);
  AND2 I1322 (rd_5r1[16:16], dt_0[48:48], rg_5r);
  AND2 I1323 (rd_5r1[17:17], dt_0[49:49], rg_5r);
  AND2 I1324 (rd_5r1[18:18], dt_0[50:50], rg_5r);
  AND2 I1325 (rd_5r1[19:19], dt_0[51:51], rg_5r);
  AND2 I1326 (rd_5r1[20:20], dt_0[52:52], rg_5r);
  AND2 I1327 (rd_5r1[21:21], dt_0[53:53], rg_5r);
  AND2 I1328 (rd_5r1[22:22], dt_0[54:54], rg_5r);
  AND2 I1329 (rd_5r1[23:23], dt_0[55:55], rg_5r);
  AND2 I1330 (rd_5r1[24:24], dt_0[56:56], rg_5r);
  AND2 I1331 (rd_5r1[25:25], dt_0[57:57], rg_5r);
  AND2 I1332 (rd_5r1[26:26], dt_0[58:58], rg_5r);
  AND2 I1333 (rd_5r1[27:27], dt_0[59:59], rg_5r);
  AND2 I1334 (rd_5r1[28:28], dt_0[60:60], rg_5r);
  AND2 I1335 (rd_5r1[29:29], dt_0[61:61], rg_5r);
  AND2 I1336 (rd_5r1[30:30], dt_0[62:62], rg_5r);
  AND2 I1337 (rd_5r1[31:31], dt_0[63:63], rg_5r);
  AND2 I1338 (rd_6r1[0:0], dt_0[32:32], rg_6r);
  AND2 I1339 (rd_6r1[1:1], dt_0[33:33], rg_6r);
  AND2 I1340 (rd_6r1[2:2], dt_0[34:34], rg_6r);
  AND2 I1341 (rd_6r1[3:3], dt_0[35:35], rg_6r);
  AND2 I1342 (rd_6r1[4:4], dt_0[36:36], rg_6r);
  AND2 I1343 (rd_6r1[5:5], dt_0[37:37], rg_6r);
  AND2 I1344 (rd_6r1[6:6], dt_0[38:38], rg_6r);
  AND2 I1345 (rd_6r1[7:7], dt_0[39:39], rg_6r);
  AND2 I1346 (rd_6r1[8:8], dt_0[40:40], rg_6r);
  AND2 I1347 (rd_6r1[9:9], dt_0[41:41], rg_6r);
  AND2 I1348 (rd_6r1[10:10], dt_0[42:42], rg_6r);
  AND2 I1349 (rd_6r1[11:11], dt_0[43:43], rg_6r);
  AND2 I1350 (rd_6r1[12:12], dt_0[44:44], rg_6r);
  AND2 I1351 (rd_6r1[13:13], dt_0[45:45], rg_6r);
  AND2 I1352 (rd_6r1[14:14], dt_0[46:46], rg_6r);
  AND2 I1353 (rd_6r1[15:15], dt_0[47:47], rg_6r);
  AND2 I1354 (rd_6r1[16:16], dt_0[48:48], rg_6r);
  AND2 I1355 (rd_6r1[17:17], dt_0[49:49], rg_6r);
  AND2 I1356 (rd_6r1[18:18], dt_0[50:50], rg_6r);
  AND2 I1357 (rd_6r1[19:19], dt_0[51:51], rg_6r);
  AND2 I1358 (rd_6r1[20:20], dt_0[52:52], rg_6r);
  AND2 I1359 (rd_6r1[21:21], dt_0[53:53], rg_6r);
  AND2 I1360 (rd_6r1[22:22], dt_0[54:54], rg_6r);
  AND2 I1361 (rd_6r1[23:23], dt_0[55:55], rg_6r);
  AND2 I1362 (rd_6r1[24:24], dt_0[56:56], rg_6r);
  AND2 I1363 (rd_6r1[25:25], dt_0[57:57], rg_6r);
  AND2 I1364 (rd_6r1[26:26], dt_0[58:58], rg_6r);
  AND2 I1365 (rd_6r1[27:27], dt_0[59:59], rg_6r);
  AND2 I1366 (rd_6r1[28:28], dt_0[60:60], rg_6r);
  AND2 I1367 (rd_6r1[29:29], dt_0[61:61], rg_6r);
  AND2 I1368 (rd_6r1[30:30], dt_0[62:62], rg_6r);
  AND2 I1369 (rd_6r1[31:31], dt_0[63:63], rg_6r);
  AND2 I1370 (rd_7r1[0:0], dt_0[32:32], rg_7r);
  AND2 I1371 (rd_7r1[1:1], dt_0[33:33], rg_7r);
  AND2 I1372 (rd_7r1[2:2], dt_0[34:34], rg_7r);
  AND2 I1373 (rd_7r1[3:3], dt_0[35:35], rg_7r);
  AND2 I1374 (rd_7r1[4:4], dt_0[36:36], rg_7r);
  AND2 I1375 (rd_7r1[5:5], dt_0[37:37], rg_7r);
  AND2 I1376 (rd_7r1[6:6], dt_0[38:38], rg_7r);
  AND2 I1377 (rd_7r1[7:7], dt_0[39:39], rg_7r);
  AND2 I1378 (rd_7r1[8:8], dt_0[40:40], rg_7r);
  AND2 I1379 (rd_7r1[9:9], dt_0[41:41], rg_7r);
  AND2 I1380 (rd_7r1[10:10], dt_0[42:42], rg_7r);
  AND2 I1381 (rd_7r1[11:11], dt_0[43:43], rg_7r);
  AND2 I1382 (rd_7r1[12:12], dt_0[44:44], rg_7r);
  AND2 I1383 (rd_7r1[13:13], dt_0[45:45], rg_7r);
  AND2 I1384 (rd_7r1[14:14], dt_0[46:46], rg_7r);
  AND2 I1385 (rd_7r1[15:15], dt_0[47:47], rg_7r);
  AND2 I1386 (rd_7r1[16:16], dt_0[48:48], rg_7r);
  AND2 I1387 (rd_7r1[17:17], dt_0[49:49], rg_7r);
  AND2 I1388 (rd_7r1[18:18], dt_0[50:50], rg_7r);
  AND2 I1389 (rd_7r1[19:19], dt_0[51:51], rg_7r);
  AND2 I1390 (rd_7r1[20:20], dt_0[52:52], rg_7r);
  AND2 I1391 (rd_7r1[21:21], dt_0[53:53], rg_7r);
  AND2 I1392 (rd_7r1[22:22], dt_0[54:54], rg_7r);
  AND2 I1393 (rd_7r1[23:23], dt_0[55:55], rg_7r);
  AND2 I1394 (rd_7r1[24:24], dt_0[56:56], rg_7r);
  AND2 I1395 (rd_7r1[25:25], dt_0[57:57], rg_7r);
  AND2 I1396 (rd_7r1[26:26], dt_0[58:58], rg_7r);
  AND2 I1397 (rd_7r1[27:27], dt_0[59:59], rg_7r);
  AND2 I1398 (rd_7r1[28:28], dt_0[60:60], rg_7r);
  AND2 I1399 (rd_7r1[29:29], dt_0[61:61], rg_7r);
  AND2 I1400 (rd_7r1[30:30], dt_0[62:62], rg_7r);
  AND2 I1401 (rd_7r1[31:31], dt_0[63:63], rg_7r);
  AND2 I1402 (rd_8r1[0:0], dt_0[32:32], rg_8r);
  AND2 I1403 (rd_8r1[1:1], dt_0[33:33], rg_8r);
  AND2 I1404 (rd_8r1[2:2], dt_0[34:34], rg_8r);
  AND2 I1405 (rd_8r1[3:3], dt_0[35:35], rg_8r);
  AND2 I1406 (rd_8r1[4:4], dt_0[36:36], rg_8r);
  AND2 I1407 (rd_8r1[5:5], dt_0[37:37], rg_8r);
  AND2 I1408 (rd_8r1[6:6], dt_0[38:38], rg_8r);
  AND2 I1409 (rd_8r1[7:7], dt_0[39:39], rg_8r);
  AND2 I1410 (rd_8r1[8:8], dt_0[40:40], rg_8r);
  AND2 I1411 (rd_8r1[9:9], dt_0[41:41], rg_8r);
  AND2 I1412 (rd_8r1[10:10], dt_0[42:42], rg_8r);
  AND2 I1413 (rd_8r1[11:11], dt_0[43:43], rg_8r);
  AND2 I1414 (rd_8r1[12:12], dt_0[44:44], rg_8r);
  AND2 I1415 (rd_8r1[13:13], dt_0[45:45], rg_8r);
  AND2 I1416 (rd_8r1[14:14], dt_0[46:46], rg_8r);
  AND2 I1417 (rd_8r1[15:15], dt_0[47:47], rg_8r);
  AND2 I1418 (rd_8r1[16:16], dt_0[48:48], rg_8r);
  AND2 I1419 (rd_8r1[17:17], dt_0[49:49], rg_8r);
  AND2 I1420 (rd_8r1[18:18], dt_0[50:50], rg_8r);
  AND2 I1421 (rd_8r1[19:19], dt_0[51:51], rg_8r);
  AND2 I1422 (rd_8r1[20:20], dt_0[52:52], rg_8r);
  AND2 I1423 (rd_8r1[21:21], dt_0[53:53], rg_8r);
  AND2 I1424 (rd_8r1[22:22], dt_0[54:54], rg_8r);
  AND2 I1425 (rd_8r1[23:23], dt_0[55:55], rg_8r);
  AND2 I1426 (rd_8r1[24:24], dt_0[56:56], rg_8r);
  AND2 I1427 (rd_8r1[25:25], dt_0[57:57], rg_8r);
  AND2 I1428 (rd_8r1[26:26], dt_0[58:58], rg_8r);
  AND2 I1429 (rd_8r1[27:27], dt_0[59:59], rg_8r);
  AND2 I1430 (rd_8r1[28:28], dt_0[60:60], rg_8r);
  AND2 I1431 (rd_8r1[29:29], dt_0[61:61], rg_8r);
  AND2 I1432 (rd_8r1[30:30], dt_0[62:62], rg_8r);
  AND2 I1433 (rd_8r1[31:31], dt_0[63:63], rg_8r);
  AND2 I1434 (rd_9r1, dt_0[64:64], rg_9r);
  AND2 I1435 (rd_10r1, dt_0[64:64], rg_10r);
  AND2 I1436 (rd_11r1, dt_0[64:64], rg_11r);
  AND2 I1437 (rd_12r1, dt_0[64:64], rg_12r);
  AND2 I1438 (rd_13r1, dt_0[64:64], rg_13r);
  AND2 I1439 (rd_14r1, dt_0[64:64], rg_14r);
  NOR3 I1440 (simp13921_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I1441 (simp13921_0[1:1], rg_3r, rg_4r, rg_5r);
  NOR3 I1442 (simp13921_0[2:2], rg_6r, rg_7r, rg_8r);
  NOR3 I1443 (simp13921_0[3:3], rg_9r, rg_10r, rg_11r);
  NOR3 I1444 (simp13921_0[4:4], rg_12r, rg_13r, rg_14r);
  NOR3 I1445 (simp13921_0[5:5], rg_0a, rg_1a, rg_2a);
  NOR3 I1446 (simp13921_0[6:6], rg_3a, rg_4a, rg_5a);
  NOR3 I1447 (simp13921_0[7:7], rg_6a, rg_7a, rg_8a);
  NOR3 I1448 (simp13921_0[8:8], rg_9a, rg_10a, rg_11a);
  NOR3 I1449 (simp13921_0[9:9], rg_12a, rg_13a, rg_14a);
  NAND3 I1450 (simp13922_0[0:0], simp13921_0[0:0], simp13921_0[1:1], simp13921_0[2:2]);
  NAND3 I1451 (simp13922_0[1:1], simp13921_0[3:3], simp13921_0[4:4], simp13921_0[5:5]);
  NAND3 I1452 (simp13922_0[2:2], simp13921_0[6:6], simp13921_0[7:7], simp13921_0[8:8]);
  INV I1453 (simp13922_0[3:3], simp13921_0[9:9]);
  NOR3 I1454 (simp13923_0[0:0], simp13922_0[0:0], simp13922_0[1:1], simp13922_0[2:2]);
  INV I1455 (simp13923_0[1:1], simp13922_0[3:3]);
  NAND2 I1456 (anyread_0, simp13923_0[0:0], simp13923_0[1:1]);
  BUFF I1457 (wg_0a, wd_0a);
  BUFF I1458 (rg_0a, rd_0a);
  BUFF I1459 (rg_1a, rd_1a);
  BUFF I1460 (rg_2a, rd_2a);
  BUFF I1461 (rg_3a, rd_3a);
  BUFF I1462 (rg_4a, rd_4a);
  BUFF I1463 (rg_5a, rd_5a);
  BUFF I1464 (rg_6a, rd_6a);
  BUFF I1465 (rg_7a, rd_7a);
  BUFF I1466 (rg_8a, rd_8a);
  BUFF I1467 (rg_9a, rd_9a);
  BUFF I1468 (rg_10a, rd_10a);
  BUFF I1469 (rg_11a, rd_11a);
  BUFF I1470 (rg_12a, rd_12a);
  BUFF I1471 (rg_13a, rd_13a);
  BUFF I1472 (rg_14a, rd_14a);
endmodule

// tkvaXORbresult34_wo0w34_ro0w1o33w1o32w1 TeakV "aXORb-result" 34 [] [0] [0,33,32] [Many [34],Many [0]
//   ,Many [0,0,0],Many [1,1,1]]
module tkvaXORbresult34_wo0w34_ro0w1o33w1o32w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [33:0] wg_0r0;
  input [33:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  output rd_1r0;
  output rd_1r1;
  input rd_1a;
  output rd_2r0;
  output rd_2r1;
  input rd_2a;
  input reset;
  wire [33:0] wf_0;
  wire [33:0] wt_0;
  wire [33:0] df_0;
  wire [33:0] dt_0;
  wire wc_0;
  wire [33:0] wacks_0;
  wire [33:0] wenr_0;
  wire [33:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [33:0] drlgf_0;
  wire [33:0] drlgt_0;
  wire [33:0] comp0_0;
  wire [11:0] simp2521_0;
  wire [3:0] simp2522_0;
  wire [1:0] simp2523_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [33:0] conwgit_0;
  wire [33:0] conwgif_0;
  wire conwig_0;
  wire [11:0] simp4311_0;
  wire [3:0] simp4312_0;
  wire [1:0] simp4313_0;
  wire [1:0] simp4381_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (wen_0[32:32], wenr_0[32:32], nreset_0);
  AND2 I34 (wen_0[33:33], wenr_0[33:33], nreset_0);
  AND2 I35 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I36 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I37 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I38 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I39 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I40 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I41 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I42 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I43 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I44 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I45 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I46 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I47 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I48 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I49 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I50 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I51 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I52 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I53 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I54 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I55 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I56 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I57 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I58 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I59 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I60 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I61 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I62 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I63 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I64 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I65 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I66 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I67 (drlgf_0[32:32], wf_0[32:32], wen_0[32:32]);
  AND2 I68 (drlgf_0[33:33], wf_0[33:33], wen_0[33:33]);
  AND2 I69 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I70 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I71 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I72 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I73 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I74 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I75 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I76 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I77 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I78 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I79 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I80 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I81 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I82 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I83 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I84 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I85 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I86 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I87 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I88 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I89 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I90 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I91 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I92 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I93 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I94 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I95 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I96 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I97 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I98 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I99 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I100 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  AND2 I101 (drlgt_0[32:32], wt_0[32:32], wen_0[32:32]);
  AND2 I102 (drlgt_0[33:33], wt_0[33:33], wen_0[33:33]);
  NOR2 I103 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I104 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I105 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I106 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I107 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I108 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I109 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I110 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I111 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I112 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I113 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I114 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I115 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I116 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I117 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I118 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I119 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I120 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I121 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I122 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I123 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I124 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I125 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I126 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I127 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I128 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I129 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I130 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I131 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I132 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I133 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I134 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR2 I135 (df_0[32:32], dt_0[32:32], drlgt_0[32:32]);
  NOR2 I136 (df_0[33:33], dt_0[33:33], drlgt_0[33:33]);
  NOR3 I137 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I138 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I139 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I140 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I141 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I142 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I143 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I144 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I145 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I146 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I147 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I148 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I149 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I150 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I151 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I152 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I153 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I154 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I155 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I156 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I157 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I158 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I159 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I160 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I161 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I162 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I163 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I164 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I165 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I166 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I167 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I168 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  NOR3 I169 (dt_0[32:32], df_0[32:32], drlgf_0[32:32], reset);
  NOR3 I170 (dt_0[33:33], df_0[33:33], drlgf_0[33:33], reset);
  AO22 I171 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I172 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I173 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I174 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I175 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I176 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I177 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I178 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I179 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I180 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I181 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I182 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I183 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I184 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I185 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I186 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I187 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I188 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I189 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I190 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I191 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I192 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I193 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I194 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I195 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I196 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I197 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I198 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I199 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I200 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I201 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I202 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  AO22 I203 (wacks_0[32:32], drlgf_0[32:32], df_0[32:32], drlgt_0[32:32], dt_0[32:32]);
  AO22 I204 (wacks_0[33:33], drlgf_0[33:33], df_0[33:33], drlgt_0[33:33], dt_0[33:33]);
  OR2 I205 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I206 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I207 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I208 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I209 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I210 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I211 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I212 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I213 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I214 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I215 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I216 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I217 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I218 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I219 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I220 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I221 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I222 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I223 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I224 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I225 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I226 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I227 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I228 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I229 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I230 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I231 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I232 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I233 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I234 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I235 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I236 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  OR2 I237 (comp0_0[32:32], wg_0r0[32:32], wg_0r1[32:32]);
  OR2 I238 (comp0_0[33:33], wg_0r0[33:33], wg_0r1[33:33]);
  C3 I239 (simp2521_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I240 (simp2521_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I241 (simp2521_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I242 (simp2521_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I243 (simp2521_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I244 (simp2521_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I245 (simp2521_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I246 (simp2521_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I247 (simp2521_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I248 (simp2521_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C3 I249 (simp2521_0[10:10], comp0_0[30:30], comp0_0[31:31], comp0_0[32:32]);
  BUFF I250 (simp2521_0[11:11], comp0_0[33:33]);
  C3 I251 (simp2522_0[0:0], simp2521_0[0:0], simp2521_0[1:1], simp2521_0[2:2]);
  C3 I252 (simp2522_0[1:1], simp2521_0[3:3], simp2521_0[4:4], simp2521_0[5:5]);
  C3 I253 (simp2522_0[2:2], simp2521_0[6:6], simp2521_0[7:7], simp2521_0[8:8]);
  C3 I254 (simp2522_0[3:3], simp2521_0[9:9], simp2521_0[10:10], simp2521_0[11:11]);
  C3 I255 (simp2523_0[0:0], simp2522_0[0:0], simp2522_0[1:1], simp2522_0[2:2]);
  BUFF I256 (simp2523_0[1:1], simp2522_0[3:3]);
  C2 I257 (wc_0, simp2523_0[0:0], simp2523_0[1:1]);
  AND2 I258 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I259 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I260 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I261 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I262 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I263 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I264 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I265 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I266 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I267 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I268 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I269 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I270 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I271 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I272 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I273 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I274 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I275 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I276 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I277 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I278 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I279 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I280 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I281 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I282 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I283 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I284 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I285 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I286 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I287 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I288 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I289 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I290 (conwgif_0[32:32], wg_0r0[32:32], conwig_0);
  AND2 I291 (conwgif_0[33:33], wg_0r0[33:33], conwig_0);
  AND2 I292 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I293 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I294 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I295 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I296 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I297 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I298 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I299 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I300 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I301 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I302 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I303 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I304 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I305 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I306 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I307 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I308 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I309 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I310 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I311 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I312 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I313 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I314 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I315 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I316 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I317 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I318 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I319 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I320 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I321 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I322 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I323 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  AND2 I324 (conwgit_0[32:32], wg_0r1[32:32], conwig_0);
  AND2 I325 (conwgit_0[33:33], wg_0r1[33:33], conwig_0);
  BUFF I326 (conwigc_0, wc_0);
  AO22 I327 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I328 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I329 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I330 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I331 (wenr_0[0:0], wc_0);
  BUFF I332 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I333 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I334 (wenr_0[1:1], wc_0);
  BUFF I335 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I336 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I337 (wenr_0[2:2], wc_0);
  BUFF I338 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I339 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I340 (wenr_0[3:3], wc_0);
  BUFF I341 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I342 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I343 (wenr_0[4:4], wc_0);
  BUFF I344 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I345 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I346 (wenr_0[5:5], wc_0);
  BUFF I347 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I348 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I349 (wenr_0[6:6], wc_0);
  BUFF I350 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I351 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I352 (wenr_0[7:7], wc_0);
  BUFF I353 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I354 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I355 (wenr_0[8:8], wc_0);
  BUFF I356 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I357 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I358 (wenr_0[9:9], wc_0);
  BUFF I359 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I360 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I361 (wenr_0[10:10], wc_0);
  BUFF I362 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I363 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I364 (wenr_0[11:11], wc_0);
  BUFF I365 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I366 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I367 (wenr_0[12:12], wc_0);
  BUFF I368 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I369 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I370 (wenr_0[13:13], wc_0);
  BUFF I371 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I372 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I373 (wenr_0[14:14], wc_0);
  BUFF I374 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I375 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I376 (wenr_0[15:15], wc_0);
  BUFF I377 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I378 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I379 (wenr_0[16:16], wc_0);
  BUFF I380 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I381 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I382 (wenr_0[17:17], wc_0);
  BUFF I383 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I384 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I385 (wenr_0[18:18], wc_0);
  BUFF I386 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I387 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I388 (wenr_0[19:19], wc_0);
  BUFF I389 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I390 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I391 (wenr_0[20:20], wc_0);
  BUFF I392 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I393 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I394 (wenr_0[21:21], wc_0);
  BUFF I395 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I396 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I397 (wenr_0[22:22], wc_0);
  BUFF I398 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I399 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I400 (wenr_0[23:23], wc_0);
  BUFF I401 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I402 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I403 (wenr_0[24:24], wc_0);
  BUFF I404 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I405 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I406 (wenr_0[25:25], wc_0);
  BUFF I407 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I408 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I409 (wenr_0[26:26], wc_0);
  BUFF I410 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I411 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I412 (wenr_0[27:27], wc_0);
  BUFF I413 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I414 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I415 (wenr_0[28:28], wc_0);
  BUFF I416 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I417 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I418 (wenr_0[29:29], wc_0);
  BUFF I419 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I420 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I421 (wenr_0[30:30], wc_0);
  BUFF I422 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I423 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I424 (wenr_0[31:31], wc_0);
  BUFF I425 (wf_0[32:32], conwgif_0[32:32]);
  BUFF I426 (wt_0[32:32], conwgit_0[32:32]);
  BUFF I427 (wenr_0[32:32], wc_0);
  BUFF I428 (wf_0[33:33], conwgif_0[33:33]);
  BUFF I429 (wt_0[33:33], conwgit_0[33:33]);
  BUFF I430 (wenr_0[33:33], wc_0);
  C3 I431 (simp4311_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I432 (simp4311_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I433 (simp4311_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I434 (simp4311_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I435 (simp4311_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I436 (simp4311_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I437 (simp4311_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I438 (simp4311_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I439 (simp4311_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I440 (simp4311_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I441 (simp4311_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C2 I442 (simp4311_0[11:11], wacks_0[32:32], wacks_0[33:33]);
  C3 I443 (simp4312_0[0:0], simp4311_0[0:0], simp4311_0[1:1], simp4311_0[2:2]);
  C3 I444 (simp4312_0[1:1], simp4311_0[3:3], simp4311_0[4:4], simp4311_0[5:5]);
  C3 I445 (simp4312_0[2:2], simp4311_0[6:6], simp4311_0[7:7], simp4311_0[8:8]);
  C3 I446 (simp4312_0[3:3], simp4311_0[9:9], simp4311_0[10:10], simp4311_0[11:11]);
  C3 I447 (simp4313_0[0:0], simp4312_0[0:0], simp4312_0[1:1], simp4312_0[2:2]);
  BUFF I448 (simp4313_0[1:1], simp4312_0[3:3]);
  C2 I449 (wd_0r, simp4313_0[0:0], simp4313_0[1:1]);
  AND2 I450 (rd_0r0, df_0[0:0], rg_0r);
  AND2 I451 (rd_1r0, df_0[33:33], rg_1r);
  AND2 I452 (rd_2r0, df_0[32:32], rg_2r);
  AND2 I453 (rd_0r1, dt_0[0:0], rg_0r);
  AND2 I454 (rd_1r1, dt_0[33:33], rg_1r);
  AND2 I455 (rd_2r1, dt_0[32:32], rg_2r);
  NOR3 I456 (simp4381_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I457 (simp4381_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I458 (anyread_0, simp4381_0[0:0], simp4381_0[1:1]);
  BUFF I459 (wg_0a, wd_0a);
  BUFF I460 (rg_0a, rd_0a);
  BUFF I461 (rg_1a, rd_1a);
  BUFF I462 (rg_2a, rd_2a);
endmodule

// tkj8m4_4_0 TeakJ [Many [4,4,0],One 8]
module tkj8m4_4_0 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r, i_2a, o_0r0, o_0r1, o_0a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  input [3:0] i_1r0;
  input [3:0] i_1r1;
  output i_1a;
  input i_2r;
  output i_2a;
  output [7:0] o_0r0;
  output [7:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [7:0] joinf_0;
  wire [7:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_1r0[0:0]);
  BUFF I5 (joinf_0[5:5], i_1r0[1:1]);
  BUFF I6 (joinf_0[6:6], i_1r0[2:2]);
  BUFF I7 (joinf_0[7:7], i_1r0[3:3]);
  BUFF I8 (joint_0[0:0], i_0r1[0:0]);
  BUFF I9 (joint_0[1:1], i_0r1[1:1]);
  BUFF I10 (joint_0[2:2], i_0r1[2:2]);
  BUFF I11 (joint_0[3:3], i_0r1[3:3]);
  BUFF I12 (joint_0[4:4], i_1r1[0:0]);
  BUFF I13 (joint_0[5:5], i_1r1[1:1]);
  BUFF I14 (joint_0[6:6], i_1r1[2:2]);
  BUFF I15 (joint_0[7:7], i_1r1[3:3]);
  BUFF I16 (icomplete_0, i_2r);
  C2 I17 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I18 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I19 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I20 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I21 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I22 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I23 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I24 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I25 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I26 (o_0r1[1:1], joint_0[1:1]);
  BUFF I27 (o_0r1[2:2], joint_0[2:2]);
  BUFF I28 (o_0r1[3:3], joint_0[3:3]);
  BUFF I29 (o_0r1[4:4], joint_0[4:4]);
  BUFF I30 (o_0r1[5:5], joint_0[5:5]);
  BUFF I31 (o_0r1[6:6], joint_0[6:6]);
  BUFF I32 (o_0r1[7:7], joint_0[7:7]);
  BUFF I33 (i_0a, o_0a);
  BUFF I34 (i_1a, o_0a);
  BUFF I35 (i_2a, o_0a);
endmodule

// tkj65m32_32_1 TeakJ [Many [32,32,1],One 65]
module tkj65m32_32_1 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  input i_2r0;
  input i_2r1;
  output i_2a;
  output [64:0] o_0r0;
  output [64:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r0[0:0]);
  BUFF I1 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I2 (o_0r0[2:2], i_0r0[2:2]);
  BUFF I3 (o_0r0[3:3], i_0r0[3:3]);
  BUFF I4 (o_0r0[4:4], i_0r0[4:4]);
  BUFF I5 (o_0r0[5:5], i_0r0[5:5]);
  BUFF I6 (o_0r0[6:6], i_0r0[6:6]);
  BUFF I7 (o_0r0[7:7], i_0r0[7:7]);
  BUFF I8 (o_0r0[8:8], i_0r0[8:8]);
  BUFF I9 (o_0r0[9:9], i_0r0[9:9]);
  BUFF I10 (o_0r0[10:10], i_0r0[10:10]);
  BUFF I11 (o_0r0[11:11], i_0r0[11:11]);
  BUFF I12 (o_0r0[12:12], i_0r0[12:12]);
  BUFF I13 (o_0r0[13:13], i_0r0[13:13]);
  BUFF I14 (o_0r0[14:14], i_0r0[14:14]);
  BUFF I15 (o_0r0[15:15], i_0r0[15:15]);
  BUFF I16 (o_0r0[16:16], i_0r0[16:16]);
  BUFF I17 (o_0r0[17:17], i_0r0[17:17]);
  BUFF I18 (o_0r0[18:18], i_0r0[18:18]);
  BUFF I19 (o_0r0[19:19], i_0r0[19:19]);
  BUFF I20 (o_0r0[20:20], i_0r0[20:20]);
  BUFF I21 (o_0r0[21:21], i_0r0[21:21]);
  BUFF I22 (o_0r0[22:22], i_0r0[22:22]);
  BUFF I23 (o_0r0[23:23], i_0r0[23:23]);
  BUFF I24 (o_0r0[24:24], i_0r0[24:24]);
  BUFF I25 (o_0r0[25:25], i_0r0[25:25]);
  BUFF I26 (o_0r0[26:26], i_0r0[26:26]);
  BUFF I27 (o_0r0[27:27], i_0r0[27:27]);
  BUFF I28 (o_0r0[28:28], i_0r0[28:28]);
  BUFF I29 (o_0r0[29:29], i_0r0[29:29]);
  BUFF I30 (o_0r0[30:30], i_0r0[30:30]);
  BUFF I31 (o_0r0[31:31], i_0r0[31:31]);
  BUFF I32 (o_0r0[32:32], i_1r0[0:0]);
  BUFF I33 (o_0r0[33:33], i_1r0[1:1]);
  BUFF I34 (o_0r0[34:34], i_1r0[2:2]);
  BUFF I35 (o_0r0[35:35], i_1r0[3:3]);
  BUFF I36 (o_0r0[36:36], i_1r0[4:4]);
  BUFF I37 (o_0r0[37:37], i_1r0[5:5]);
  BUFF I38 (o_0r0[38:38], i_1r0[6:6]);
  BUFF I39 (o_0r0[39:39], i_1r0[7:7]);
  BUFF I40 (o_0r0[40:40], i_1r0[8:8]);
  BUFF I41 (o_0r0[41:41], i_1r0[9:9]);
  BUFF I42 (o_0r0[42:42], i_1r0[10:10]);
  BUFF I43 (o_0r0[43:43], i_1r0[11:11]);
  BUFF I44 (o_0r0[44:44], i_1r0[12:12]);
  BUFF I45 (o_0r0[45:45], i_1r0[13:13]);
  BUFF I46 (o_0r0[46:46], i_1r0[14:14]);
  BUFF I47 (o_0r0[47:47], i_1r0[15:15]);
  BUFF I48 (o_0r0[48:48], i_1r0[16:16]);
  BUFF I49 (o_0r0[49:49], i_1r0[17:17]);
  BUFF I50 (o_0r0[50:50], i_1r0[18:18]);
  BUFF I51 (o_0r0[51:51], i_1r0[19:19]);
  BUFF I52 (o_0r0[52:52], i_1r0[20:20]);
  BUFF I53 (o_0r0[53:53], i_1r0[21:21]);
  BUFF I54 (o_0r0[54:54], i_1r0[22:22]);
  BUFF I55 (o_0r0[55:55], i_1r0[23:23]);
  BUFF I56 (o_0r0[56:56], i_1r0[24:24]);
  BUFF I57 (o_0r0[57:57], i_1r0[25:25]);
  BUFF I58 (o_0r0[58:58], i_1r0[26:26]);
  BUFF I59 (o_0r0[59:59], i_1r0[27:27]);
  BUFF I60 (o_0r0[60:60], i_1r0[28:28]);
  BUFF I61 (o_0r0[61:61], i_1r0[29:29]);
  BUFF I62 (o_0r0[62:62], i_1r0[30:30]);
  BUFF I63 (o_0r0[63:63], i_1r0[31:31]);
  BUFF I64 (o_0r0[64:64], i_2r0);
  BUFF I65 (o_0r1[0:0], i_0r1[0:0]);
  BUFF I66 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I67 (o_0r1[2:2], i_0r1[2:2]);
  BUFF I68 (o_0r1[3:3], i_0r1[3:3]);
  BUFF I69 (o_0r1[4:4], i_0r1[4:4]);
  BUFF I70 (o_0r1[5:5], i_0r1[5:5]);
  BUFF I71 (o_0r1[6:6], i_0r1[6:6]);
  BUFF I72 (o_0r1[7:7], i_0r1[7:7]);
  BUFF I73 (o_0r1[8:8], i_0r1[8:8]);
  BUFF I74 (o_0r1[9:9], i_0r1[9:9]);
  BUFF I75 (o_0r1[10:10], i_0r1[10:10]);
  BUFF I76 (o_0r1[11:11], i_0r1[11:11]);
  BUFF I77 (o_0r1[12:12], i_0r1[12:12]);
  BUFF I78 (o_0r1[13:13], i_0r1[13:13]);
  BUFF I79 (o_0r1[14:14], i_0r1[14:14]);
  BUFF I80 (o_0r1[15:15], i_0r1[15:15]);
  BUFF I81 (o_0r1[16:16], i_0r1[16:16]);
  BUFF I82 (o_0r1[17:17], i_0r1[17:17]);
  BUFF I83 (o_0r1[18:18], i_0r1[18:18]);
  BUFF I84 (o_0r1[19:19], i_0r1[19:19]);
  BUFF I85 (o_0r1[20:20], i_0r1[20:20]);
  BUFF I86 (o_0r1[21:21], i_0r1[21:21]);
  BUFF I87 (o_0r1[22:22], i_0r1[22:22]);
  BUFF I88 (o_0r1[23:23], i_0r1[23:23]);
  BUFF I89 (o_0r1[24:24], i_0r1[24:24]);
  BUFF I90 (o_0r1[25:25], i_0r1[25:25]);
  BUFF I91 (o_0r1[26:26], i_0r1[26:26]);
  BUFF I92 (o_0r1[27:27], i_0r1[27:27]);
  BUFF I93 (o_0r1[28:28], i_0r1[28:28]);
  BUFF I94 (o_0r1[29:29], i_0r1[29:29]);
  BUFF I95 (o_0r1[30:30], i_0r1[30:30]);
  BUFF I96 (o_0r1[31:31], i_0r1[31:31]);
  BUFF I97 (o_0r1[32:32], i_1r1[0:0]);
  BUFF I98 (o_0r1[33:33], i_1r1[1:1]);
  BUFF I99 (o_0r1[34:34], i_1r1[2:2]);
  BUFF I100 (o_0r1[35:35], i_1r1[3:3]);
  BUFF I101 (o_0r1[36:36], i_1r1[4:4]);
  BUFF I102 (o_0r1[37:37], i_1r1[5:5]);
  BUFF I103 (o_0r1[38:38], i_1r1[6:6]);
  BUFF I104 (o_0r1[39:39], i_1r1[7:7]);
  BUFF I105 (o_0r1[40:40], i_1r1[8:8]);
  BUFF I106 (o_0r1[41:41], i_1r1[9:9]);
  BUFF I107 (o_0r1[42:42], i_1r1[10:10]);
  BUFF I108 (o_0r1[43:43], i_1r1[11:11]);
  BUFF I109 (o_0r1[44:44], i_1r1[12:12]);
  BUFF I110 (o_0r1[45:45], i_1r1[13:13]);
  BUFF I111 (o_0r1[46:46], i_1r1[14:14]);
  BUFF I112 (o_0r1[47:47], i_1r1[15:15]);
  BUFF I113 (o_0r1[48:48], i_1r1[16:16]);
  BUFF I114 (o_0r1[49:49], i_1r1[17:17]);
  BUFF I115 (o_0r1[50:50], i_1r1[18:18]);
  BUFF I116 (o_0r1[51:51], i_1r1[19:19]);
  BUFF I117 (o_0r1[52:52], i_1r1[20:20]);
  BUFF I118 (o_0r1[53:53], i_1r1[21:21]);
  BUFF I119 (o_0r1[54:54], i_1r1[22:22]);
  BUFF I120 (o_0r1[55:55], i_1r1[23:23]);
  BUFF I121 (o_0r1[56:56], i_1r1[24:24]);
  BUFF I122 (o_0r1[57:57], i_1r1[25:25]);
  BUFF I123 (o_0r1[58:58], i_1r1[26:26]);
  BUFF I124 (o_0r1[59:59], i_1r1[27:27]);
  BUFF I125 (o_0r1[60:60], i_1r1[28:28]);
  BUFF I126 (o_0r1[61:61], i_1r1[29:29]);
  BUFF I127 (o_0r1[62:62], i_1r1[30:30]);
  BUFF I128 (o_0r1[63:63], i_1r1[31:31]);
  BUFF I129 (o_0r1[64:64], i_2r1);
  BUFF I130 (i_0a, o_0a);
  BUFF I131 (i_1a, o_0a);
  BUFF I132 (i_2a, o_0a);
endmodule

// tkj34m1_0_33 TeakJ [Many [1,0,33],One 34]
module tkj34m1_0_33 (i_0r0, i_0r1, i_0a, i_1r, i_1a, i_2r0, i_2r1, i_2a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  input [32:0] i_2r0;
  input [32:0] i_2r1;
  output i_2a;
  output [33:0] o_0r0;
  output [33:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [33:0] joinf_0;
  wire [33:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_0r0);
  BUFF I1 (joinf_0[1:1], i_2r0[0:0]);
  BUFF I2 (joinf_0[2:2], i_2r0[1:1]);
  BUFF I3 (joinf_0[3:3], i_2r0[2:2]);
  BUFF I4 (joinf_0[4:4], i_2r0[3:3]);
  BUFF I5 (joinf_0[5:5], i_2r0[4:4]);
  BUFF I6 (joinf_0[6:6], i_2r0[5:5]);
  BUFF I7 (joinf_0[7:7], i_2r0[6:6]);
  BUFF I8 (joinf_0[8:8], i_2r0[7:7]);
  BUFF I9 (joinf_0[9:9], i_2r0[8:8]);
  BUFF I10 (joinf_0[10:10], i_2r0[9:9]);
  BUFF I11 (joinf_0[11:11], i_2r0[10:10]);
  BUFF I12 (joinf_0[12:12], i_2r0[11:11]);
  BUFF I13 (joinf_0[13:13], i_2r0[12:12]);
  BUFF I14 (joinf_0[14:14], i_2r0[13:13]);
  BUFF I15 (joinf_0[15:15], i_2r0[14:14]);
  BUFF I16 (joinf_0[16:16], i_2r0[15:15]);
  BUFF I17 (joinf_0[17:17], i_2r0[16:16]);
  BUFF I18 (joinf_0[18:18], i_2r0[17:17]);
  BUFF I19 (joinf_0[19:19], i_2r0[18:18]);
  BUFF I20 (joinf_0[20:20], i_2r0[19:19]);
  BUFF I21 (joinf_0[21:21], i_2r0[20:20]);
  BUFF I22 (joinf_0[22:22], i_2r0[21:21]);
  BUFF I23 (joinf_0[23:23], i_2r0[22:22]);
  BUFF I24 (joinf_0[24:24], i_2r0[23:23]);
  BUFF I25 (joinf_0[25:25], i_2r0[24:24]);
  BUFF I26 (joinf_0[26:26], i_2r0[25:25]);
  BUFF I27 (joinf_0[27:27], i_2r0[26:26]);
  BUFF I28 (joinf_0[28:28], i_2r0[27:27]);
  BUFF I29 (joinf_0[29:29], i_2r0[28:28]);
  BUFF I30 (joinf_0[30:30], i_2r0[29:29]);
  BUFF I31 (joinf_0[31:31], i_2r0[30:30]);
  BUFF I32 (joinf_0[32:32], i_2r0[31:31]);
  BUFF I33 (joinf_0[33:33], i_2r0[32:32]);
  BUFF I34 (joint_0[0:0], i_0r1);
  BUFF I35 (joint_0[1:1], i_2r1[0:0]);
  BUFF I36 (joint_0[2:2], i_2r1[1:1]);
  BUFF I37 (joint_0[3:3], i_2r1[2:2]);
  BUFF I38 (joint_0[4:4], i_2r1[3:3]);
  BUFF I39 (joint_0[5:5], i_2r1[4:4]);
  BUFF I40 (joint_0[6:6], i_2r1[5:5]);
  BUFF I41 (joint_0[7:7], i_2r1[6:6]);
  BUFF I42 (joint_0[8:8], i_2r1[7:7]);
  BUFF I43 (joint_0[9:9], i_2r1[8:8]);
  BUFF I44 (joint_0[10:10], i_2r1[9:9]);
  BUFF I45 (joint_0[11:11], i_2r1[10:10]);
  BUFF I46 (joint_0[12:12], i_2r1[11:11]);
  BUFF I47 (joint_0[13:13], i_2r1[12:12]);
  BUFF I48 (joint_0[14:14], i_2r1[13:13]);
  BUFF I49 (joint_0[15:15], i_2r1[14:14]);
  BUFF I50 (joint_0[16:16], i_2r1[15:15]);
  BUFF I51 (joint_0[17:17], i_2r1[16:16]);
  BUFF I52 (joint_0[18:18], i_2r1[17:17]);
  BUFF I53 (joint_0[19:19], i_2r1[18:18]);
  BUFF I54 (joint_0[20:20], i_2r1[19:19]);
  BUFF I55 (joint_0[21:21], i_2r1[20:20]);
  BUFF I56 (joint_0[22:22], i_2r1[21:21]);
  BUFF I57 (joint_0[23:23], i_2r1[22:22]);
  BUFF I58 (joint_0[24:24], i_2r1[23:23]);
  BUFF I59 (joint_0[25:25], i_2r1[24:24]);
  BUFF I60 (joint_0[26:26], i_2r1[25:25]);
  BUFF I61 (joint_0[27:27], i_2r1[26:26]);
  BUFF I62 (joint_0[28:28], i_2r1[27:27]);
  BUFF I63 (joint_0[29:29], i_2r1[28:28]);
  BUFF I64 (joint_0[30:30], i_2r1[29:29]);
  BUFF I65 (joint_0[31:31], i_2r1[30:30]);
  BUFF I66 (joint_0[32:32], i_2r1[31:31]);
  BUFF I67 (joint_0[33:33], i_2r1[32:32]);
  BUFF I68 (icomplete_0, i_1r);
  C2 I69 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I70 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I71 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I72 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I73 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I74 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I75 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I76 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I77 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I78 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I79 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I80 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I81 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I82 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I83 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I84 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I85 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I86 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I87 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I88 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I89 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I90 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I91 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I92 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I93 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I94 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I95 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I96 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I97 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I98 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I99 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I100 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I101 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I102 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I103 (o_0r0[33:33], joinf_0[33:33]);
  BUFF I104 (o_0r1[1:1], joint_0[1:1]);
  BUFF I105 (o_0r1[2:2], joint_0[2:2]);
  BUFF I106 (o_0r1[3:3], joint_0[3:3]);
  BUFF I107 (o_0r1[4:4], joint_0[4:4]);
  BUFF I108 (o_0r1[5:5], joint_0[5:5]);
  BUFF I109 (o_0r1[6:6], joint_0[6:6]);
  BUFF I110 (o_0r1[7:7], joint_0[7:7]);
  BUFF I111 (o_0r1[8:8], joint_0[8:8]);
  BUFF I112 (o_0r1[9:9], joint_0[9:9]);
  BUFF I113 (o_0r1[10:10], joint_0[10:10]);
  BUFF I114 (o_0r1[11:11], joint_0[11:11]);
  BUFF I115 (o_0r1[12:12], joint_0[12:12]);
  BUFF I116 (o_0r1[13:13], joint_0[13:13]);
  BUFF I117 (o_0r1[14:14], joint_0[14:14]);
  BUFF I118 (o_0r1[15:15], joint_0[15:15]);
  BUFF I119 (o_0r1[16:16], joint_0[16:16]);
  BUFF I120 (o_0r1[17:17], joint_0[17:17]);
  BUFF I121 (o_0r1[18:18], joint_0[18:18]);
  BUFF I122 (o_0r1[19:19], joint_0[19:19]);
  BUFF I123 (o_0r1[20:20], joint_0[20:20]);
  BUFF I124 (o_0r1[21:21], joint_0[21:21]);
  BUFF I125 (o_0r1[22:22], joint_0[22:22]);
  BUFF I126 (o_0r1[23:23], joint_0[23:23]);
  BUFF I127 (o_0r1[24:24], joint_0[24:24]);
  BUFF I128 (o_0r1[25:25], joint_0[25:25]);
  BUFF I129 (o_0r1[26:26], joint_0[26:26]);
  BUFF I130 (o_0r1[27:27], joint_0[27:27]);
  BUFF I131 (o_0r1[28:28], joint_0[28:28]);
  BUFF I132 (o_0r1[29:29], joint_0[29:29]);
  BUFF I133 (o_0r1[30:30], joint_0[30:30]);
  BUFF I134 (o_0r1[31:31], joint_0[31:31]);
  BUFF I135 (o_0r1[32:32], joint_0[32:32]);
  BUFF I136 (o_0r1[33:33], joint_0[33:33]);
  BUFF I137 (i_0a, o_0a);
  BUFF I138 (i_1a, o_0a);
  BUFF I139 (i_2a, o_0a);
endmodule

// tkj3m1_1_1 TeakJ [Many [1,1,1],One 3]
module tkj3m1_1_1 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input i_1r0;
  input i_1r1;
  output i_1a;
  input i_2r0;
  input i_2r1;
  output i_2a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r0);
  BUFF I1 (o_0r0[1:1], i_1r0);
  BUFF I2 (o_0r0[2:2], i_2r0);
  BUFF I3 (o_0r1[0:0], i_0r1);
  BUFF I4 (o_0r1[1:1], i_1r1);
  BUFF I5 (o_0r1[2:2], i_2r1);
  BUFF I6 (i_0a, o_0a);
  BUFF I7 (i_1a, o_0a);
  BUFF I8 (i_2a, o_0a);
endmodule

// tko3m1_1xori0w1bi1w1b_2xort1o0w1bi2w1b TeakO [
//     (1,TeakOp TeakOpXor [(0,0,1),(0,1,1)]),
//     (2,TeakOp TeakOpXor [(1,0,1),(0,2,1)])] [One 3,One 1]
module tko3m1_1xori0w1bi1w1b_2xort1o0w1bi2w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire termf_1;
  wire termt_1;
  wire [3:0] op1_0_0;
  wire [3:0] op2_0_0;
  C2 I0 (op1_0_0[0:0], i_0r0[1:1], i_0r0[0:0]);
  C2 I1 (op1_0_0[1:1], i_0r0[1:1], i_0r1[0:0]);
  C2 I2 (op1_0_0[2:2], i_0r1[1:1], i_0r0[0:0]);
  C2 I3 (op1_0_0[3:3], i_0r1[1:1], i_0r1[0:0]);
  OR2 I4 (termf_1, op1_0_0[0:0], op1_0_0[3:3]);
  OR2 I5 (termt_1, op1_0_0[1:1], op1_0_0[2:2]);
  C2 I6 (op2_0_0[0:0], i_0r0[2:2], termf_1);
  C2 I7 (op2_0_0[1:1], i_0r0[2:2], termt_1);
  C2 I8 (op2_0_0[2:2], i_0r1[2:2], termf_1);
  C2 I9 (op2_0_0[3:3], i_0r1[2:2], termt_1);
  OR2 I10 (o_0r0, op2_0_0[0:0], op2_0_0[3:3]);
  OR2 I11 (o_0r1, op2_0_0[1:1], op2_0_0[2:2]);
  BUFF I12 (i_0a, o_0a);
endmodule

// tkf65mo0w1_o0w65 TeakF [0,0] [One 65,Many [1,65]]
module tkf65mo0w1_o0w65 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [64:0] i_0r0;
  input [64:0] i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  output [64:0] o_1r0;
  output [64:0] o_1r1;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire [64:0] comp_0;
  wire [21:0] simp671_0;
  wire [7:0] simp672_0;
  wire [2:0] simp673_0;
  OR2 I0 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (comp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (comp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (comp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (comp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (comp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (comp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (comp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (comp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (comp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (comp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (comp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (comp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (comp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (comp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (comp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (comp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (comp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (comp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (comp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (comp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (comp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (comp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (comp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (comp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I30 (comp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I31 (comp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I32 (comp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  OR2 I33 (comp_0[33:33], i_0r0[33:33], i_0r1[33:33]);
  OR2 I34 (comp_0[34:34], i_0r0[34:34], i_0r1[34:34]);
  OR2 I35 (comp_0[35:35], i_0r0[35:35], i_0r1[35:35]);
  OR2 I36 (comp_0[36:36], i_0r0[36:36], i_0r1[36:36]);
  OR2 I37 (comp_0[37:37], i_0r0[37:37], i_0r1[37:37]);
  OR2 I38 (comp_0[38:38], i_0r0[38:38], i_0r1[38:38]);
  OR2 I39 (comp_0[39:39], i_0r0[39:39], i_0r1[39:39]);
  OR2 I40 (comp_0[40:40], i_0r0[40:40], i_0r1[40:40]);
  OR2 I41 (comp_0[41:41], i_0r0[41:41], i_0r1[41:41]);
  OR2 I42 (comp_0[42:42], i_0r0[42:42], i_0r1[42:42]);
  OR2 I43 (comp_0[43:43], i_0r0[43:43], i_0r1[43:43]);
  OR2 I44 (comp_0[44:44], i_0r0[44:44], i_0r1[44:44]);
  OR2 I45 (comp_0[45:45], i_0r0[45:45], i_0r1[45:45]);
  OR2 I46 (comp_0[46:46], i_0r0[46:46], i_0r1[46:46]);
  OR2 I47 (comp_0[47:47], i_0r0[47:47], i_0r1[47:47]);
  OR2 I48 (comp_0[48:48], i_0r0[48:48], i_0r1[48:48]);
  OR2 I49 (comp_0[49:49], i_0r0[49:49], i_0r1[49:49]);
  OR2 I50 (comp_0[50:50], i_0r0[50:50], i_0r1[50:50]);
  OR2 I51 (comp_0[51:51], i_0r0[51:51], i_0r1[51:51]);
  OR2 I52 (comp_0[52:52], i_0r0[52:52], i_0r1[52:52]);
  OR2 I53 (comp_0[53:53], i_0r0[53:53], i_0r1[53:53]);
  OR2 I54 (comp_0[54:54], i_0r0[54:54], i_0r1[54:54]);
  OR2 I55 (comp_0[55:55], i_0r0[55:55], i_0r1[55:55]);
  OR2 I56 (comp_0[56:56], i_0r0[56:56], i_0r1[56:56]);
  OR2 I57 (comp_0[57:57], i_0r0[57:57], i_0r1[57:57]);
  OR2 I58 (comp_0[58:58], i_0r0[58:58], i_0r1[58:58]);
  OR2 I59 (comp_0[59:59], i_0r0[59:59], i_0r1[59:59]);
  OR2 I60 (comp_0[60:60], i_0r0[60:60], i_0r1[60:60]);
  OR2 I61 (comp_0[61:61], i_0r0[61:61], i_0r1[61:61]);
  OR2 I62 (comp_0[62:62], i_0r0[62:62], i_0r1[62:62]);
  OR2 I63 (comp_0[63:63], i_0r0[63:63], i_0r1[63:63]);
  OR2 I64 (comp_0[64:64], i_0r0[64:64], i_0r1[64:64]);
  C3 I65 (simp671_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I66 (simp671_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C3 I67 (simp671_0[2:2], comp_0[6:6], comp_0[7:7], comp_0[8:8]);
  C3 I68 (simp671_0[3:3], comp_0[9:9], comp_0[10:10], comp_0[11:11]);
  C3 I69 (simp671_0[4:4], comp_0[12:12], comp_0[13:13], comp_0[14:14]);
  C3 I70 (simp671_0[5:5], comp_0[15:15], comp_0[16:16], comp_0[17:17]);
  C3 I71 (simp671_0[6:6], comp_0[18:18], comp_0[19:19], comp_0[20:20]);
  C3 I72 (simp671_0[7:7], comp_0[21:21], comp_0[22:22], comp_0[23:23]);
  C3 I73 (simp671_0[8:8], comp_0[24:24], comp_0[25:25], comp_0[26:26]);
  C3 I74 (simp671_0[9:9], comp_0[27:27], comp_0[28:28], comp_0[29:29]);
  C3 I75 (simp671_0[10:10], comp_0[30:30], comp_0[31:31], comp_0[32:32]);
  C3 I76 (simp671_0[11:11], comp_0[33:33], comp_0[34:34], comp_0[35:35]);
  C3 I77 (simp671_0[12:12], comp_0[36:36], comp_0[37:37], comp_0[38:38]);
  C3 I78 (simp671_0[13:13], comp_0[39:39], comp_0[40:40], comp_0[41:41]);
  C3 I79 (simp671_0[14:14], comp_0[42:42], comp_0[43:43], comp_0[44:44]);
  C3 I80 (simp671_0[15:15], comp_0[45:45], comp_0[46:46], comp_0[47:47]);
  C3 I81 (simp671_0[16:16], comp_0[48:48], comp_0[49:49], comp_0[50:50]);
  C3 I82 (simp671_0[17:17], comp_0[51:51], comp_0[52:52], comp_0[53:53]);
  C3 I83 (simp671_0[18:18], comp_0[54:54], comp_0[55:55], comp_0[56:56]);
  C3 I84 (simp671_0[19:19], comp_0[57:57], comp_0[58:58], comp_0[59:59]);
  C3 I85 (simp671_0[20:20], comp_0[60:60], comp_0[61:61], comp_0[62:62]);
  C2 I86 (simp671_0[21:21], comp_0[63:63], comp_0[64:64]);
  C3 I87 (simp672_0[0:0], simp671_0[0:0], simp671_0[1:1], simp671_0[2:2]);
  C3 I88 (simp672_0[1:1], simp671_0[3:3], simp671_0[4:4], simp671_0[5:5]);
  C3 I89 (simp672_0[2:2], simp671_0[6:6], simp671_0[7:7], simp671_0[8:8]);
  C3 I90 (simp672_0[3:3], simp671_0[9:9], simp671_0[10:10], simp671_0[11:11]);
  C3 I91 (simp672_0[4:4], simp671_0[12:12], simp671_0[13:13], simp671_0[14:14]);
  C3 I92 (simp672_0[5:5], simp671_0[15:15], simp671_0[16:16], simp671_0[17:17]);
  C3 I93 (simp672_0[6:6], simp671_0[18:18], simp671_0[19:19], simp671_0[20:20]);
  BUFF I94 (simp672_0[7:7], simp671_0[21:21]);
  C3 I95 (simp673_0[0:0], simp672_0[0:0], simp672_0[1:1], simp672_0[2:2]);
  C3 I96 (simp673_0[1:1], simp672_0[3:3], simp672_0[4:4], simp672_0[5:5]);
  C2 I97 (simp673_0[2:2], simp672_0[6:6], simp672_0[7:7]);
  C3 I98 (icomplete_0, simp673_0[0:0], simp673_0[1:1], simp673_0[2:2]);
  C2 I99 (o_0r0, i_0r0[0:0], icomplete_0);
  BUFF I100 (o_1r0[0:0], i_0r0[0:0]);
  BUFF I101 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I102 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I103 (o_1r0[3:3], i_0r0[3:3]);
  BUFF I104 (o_1r0[4:4], i_0r0[4:4]);
  BUFF I105 (o_1r0[5:5], i_0r0[5:5]);
  BUFF I106 (o_1r0[6:6], i_0r0[6:6]);
  BUFF I107 (o_1r0[7:7], i_0r0[7:7]);
  BUFF I108 (o_1r0[8:8], i_0r0[8:8]);
  BUFF I109 (o_1r0[9:9], i_0r0[9:9]);
  BUFF I110 (o_1r0[10:10], i_0r0[10:10]);
  BUFF I111 (o_1r0[11:11], i_0r0[11:11]);
  BUFF I112 (o_1r0[12:12], i_0r0[12:12]);
  BUFF I113 (o_1r0[13:13], i_0r0[13:13]);
  BUFF I114 (o_1r0[14:14], i_0r0[14:14]);
  BUFF I115 (o_1r0[15:15], i_0r0[15:15]);
  BUFF I116 (o_1r0[16:16], i_0r0[16:16]);
  BUFF I117 (o_1r0[17:17], i_0r0[17:17]);
  BUFF I118 (o_1r0[18:18], i_0r0[18:18]);
  BUFF I119 (o_1r0[19:19], i_0r0[19:19]);
  BUFF I120 (o_1r0[20:20], i_0r0[20:20]);
  BUFF I121 (o_1r0[21:21], i_0r0[21:21]);
  BUFF I122 (o_1r0[22:22], i_0r0[22:22]);
  BUFF I123 (o_1r0[23:23], i_0r0[23:23]);
  BUFF I124 (o_1r0[24:24], i_0r0[24:24]);
  BUFF I125 (o_1r0[25:25], i_0r0[25:25]);
  BUFF I126 (o_1r0[26:26], i_0r0[26:26]);
  BUFF I127 (o_1r0[27:27], i_0r0[27:27]);
  BUFF I128 (o_1r0[28:28], i_0r0[28:28]);
  BUFF I129 (o_1r0[29:29], i_0r0[29:29]);
  BUFF I130 (o_1r0[30:30], i_0r0[30:30]);
  BUFF I131 (o_1r0[31:31], i_0r0[31:31]);
  BUFF I132 (o_1r0[32:32], i_0r0[32:32]);
  BUFF I133 (o_1r0[33:33], i_0r0[33:33]);
  BUFF I134 (o_1r0[34:34], i_0r0[34:34]);
  BUFF I135 (o_1r0[35:35], i_0r0[35:35]);
  BUFF I136 (o_1r0[36:36], i_0r0[36:36]);
  BUFF I137 (o_1r0[37:37], i_0r0[37:37]);
  BUFF I138 (o_1r0[38:38], i_0r0[38:38]);
  BUFF I139 (o_1r0[39:39], i_0r0[39:39]);
  BUFF I140 (o_1r0[40:40], i_0r0[40:40]);
  BUFF I141 (o_1r0[41:41], i_0r0[41:41]);
  BUFF I142 (o_1r0[42:42], i_0r0[42:42]);
  BUFF I143 (o_1r0[43:43], i_0r0[43:43]);
  BUFF I144 (o_1r0[44:44], i_0r0[44:44]);
  BUFF I145 (o_1r0[45:45], i_0r0[45:45]);
  BUFF I146 (o_1r0[46:46], i_0r0[46:46]);
  BUFF I147 (o_1r0[47:47], i_0r0[47:47]);
  BUFF I148 (o_1r0[48:48], i_0r0[48:48]);
  BUFF I149 (o_1r0[49:49], i_0r0[49:49]);
  BUFF I150 (o_1r0[50:50], i_0r0[50:50]);
  BUFF I151 (o_1r0[51:51], i_0r0[51:51]);
  BUFF I152 (o_1r0[52:52], i_0r0[52:52]);
  BUFF I153 (o_1r0[53:53], i_0r0[53:53]);
  BUFF I154 (o_1r0[54:54], i_0r0[54:54]);
  BUFF I155 (o_1r0[55:55], i_0r0[55:55]);
  BUFF I156 (o_1r0[56:56], i_0r0[56:56]);
  BUFF I157 (o_1r0[57:57], i_0r0[57:57]);
  BUFF I158 (o_1r0[58:58], i_0r0[58:58]);
  BUFF I159 (o_1r0[59:59], i_0r0[59:59]);
  BUFF I160 (o_1r0[60:60], i_0r0[60:60]);
  BUFF I161 (o_1r0[61:61], i_0r0[61:61]);
  BUFF I162 (o_1r0[62:62], i_0r0[62:62]);
  BUFF I163 (o_1r0[63:63], i_0r0[63:63]);
  BUFF I164 (o_1r0[64:64], i_0r0[64:64]);
  C2 I165 (o_0r1, i_0r1[0:0], icomplete_0);
  BUFF I166 (o_1r1[0:0], i_0r1[0:0]);
  BUFF I167 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I168 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I169 (o_1r1[3:3], i_0r1[3:3]);
  BUFF I170 (o_1r1[4:4], i_0r1[4:4]);
  BUFF I171 (o_1r1[5:5], i_0r1[5:5]);
  BUFF I172 (o_1r1[6:6], i_0r1[6:6]);
  BUFF I173 (o_1r1[7:7], i_0r1[7:7]);
  BUFF I174 (o_1r1[8:8], i_0r1[8:8]);
  BUFF I175 (o_1r1[9:9], i_0r1[9:9]);
  BUFF I176 (o_1r1[10:10], i_0r1[10:10]);
  BUFF I177 (o_1r1[11:11], i_0r1[11:11]);
  BUFF I178 (o_1r1[12:12], i_0r1[12:12]);
  BUFF I179 (o_1r1[13:13], i_0r1[13:13]);
  BUFF I180 (o_1r1[14:14], i_0r1[14:14]);
  BUFF I181 (o_1r1[15:15], i_0r1[15:15]);
  BUFF I182 (o_1r1[16:16], i_0r1[16:16]);
  BUFF I183 (o_1r1[17:17], i_0r1[17:17]);
  BUFF I184 (o_1r1[18:18], i_0r1[18:18]);
  BUFF I185 (o_1r1[19:19], i_0r1[19:19]);
  BUFF I186 (o_1r1[20:20], i_0r1[20:20]);
  BUFF I187 (o_1r1[21:21], i_0r1[21:21]);
  BUFF I188 (o_1r1[22:22], i_0r1[22:22]);
  BUFF I189 (o_1r1[23:23], i_0r1[23:23]);
  BUFF I190 (o_1r1[24:24], i_0r1[24:24]);
  BUFF I191 (o_1r1[25:25], i_0r1[25:25]);
  BUFF I192 (o_1r1[26:26], i_0r1[26:26]);
  BUFF I193 (o_1r1[27:27], i_0r1[27:27]);
  BUFF I194 (o_1r1[28:28], i_0r1[28:28]);
  BUFF I195 (o_1r1[29:29], i_0r1[29:29]);
  BUFF I196 (o_1r1[30:30], i_0r1[30:30]);
  BUFF I197 (o_1r1[31:31], i_0r1[31:31]);
  BUFF I198 (o_1r1[32:32], i_0r1[32:32]);
  BUFF I199 (o_1r1[33:33], i_0r1[33:33]);
  BUFF I200 (o_1r1[34:34], i_0r1[34:34]);
  BUFF I201 (o_1r1[35:35], i_0r1[35:35]);
  BUFF I202 (o_1r1[36:36], i_0r1[36:36]);
  BUFF I203 (o_1r1[37:37], i_0r1[37:37]);
  BUFF I204 (o_1r1[38:38], i_0r1[38:38]);
  BUFF I205 (o_1r1[39:39], i_0r1[39:39]);
  BUFF I206 (o_1r1[40:40], i_0r1[40:40]);
  BUFF I207 (o_1r1[41:41], i_0r1[41:41]);
  BUFF I208 (o_1r1[42:42], i_0r1[42:42]);
  BUFF I209 (o_1r1[43:43], i_0r1[43:43]);
  BUFF I210 (o_1r1[44:44], i_0r1[44:44]);
  BUFF I211 (o_1r1[45:45], i_0r1[45:45]);
  BUFF I212 (o_1r1[46:46], i_0r1[46:46]);
  BUFF I213 (o_1r1[47:47], i_0r1[47:47]);
  BUFF I214 (o_1r1[48:48], i_0r1[48:48]);
  BUFF I215 (o_1r1[49:49], i_0r1[49:49]);
  BUFF I216 (o_1r1[50:50], i_0r1[50:50]);
  BUFF I217 (o_1r1[51:51], i_0r1[51:51]);
  BUFF I218 (o_1r1[52:52], i_0r1[52:52]);
  BUFF I219 (o_1r1[53:53], i_0r1[53:53]);
  BUFF I220 (o_1r1[54:54], i_0r1[54:54]);
  BUFF I221 (o_1r1[55:55], i_0r1[55:55]);
  BUFF I222 (o_1r1[56:56], i_0r1[56:56]);
  BUFF I223 (o_1r1[57:57], i_0r1[57:57]);
  BUFF I224 (o_1r1[58:58], i_0r1[58:58]);
  BUFF I225 (o_1r1[59:59], i_0r1[59:59]);
  BUFF I226 (o_1r1[60:60], i_0r1[60:60]);
  BUFF I227 (o_1r1[61:61], i_0r1[61:61]);
  BUFF I228 (o_1r1[62:62], i_0r1[62:62]);
  BUFF I229 (o_1r1[63:63], i_0r1[63:63]);
  BUFF I230 (o_1r1[64:64], i_0r1[64:64]);
  C3 I231 (i_0a, icomplete_0, o_0a, o_1a);
endmodule

// tkf34mo0w32_o0w34_o1w32 TeakF [0,0,1] [One 34,Many [32,34,32]]
module tkf34mo0w32_o0w34_o1w32 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r0, o_1r1, o_1a, o_2r0, o_2r1, o_2a, reset);
  input [33:0] i_0r0;
  input [33:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  output [33:0] o_1r0;
  output [33:0] o_1r1;
  input o_1a;
  output [31:0] o_2r0;
  output [31:0] o_2r1;
  input o_2a;
  input reset;
  wire icomplete_0;
  wire [33:0] comp_0;
  wire [11:0] simp361_0;
  wire [3:0] simp362_0;
  wire [1:0] simp363_0;
  wire [1:0] simp2341_0;
  OR2 I0 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (comp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (comp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (comp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (comp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (comp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (comp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (comp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (comp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (comp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (comp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (comp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (comp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (comp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (comp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (comp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (comp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (comp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (comp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (comp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (comp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (comp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (comp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (comp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (comp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I30 (comp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I31 (comp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I32 (comp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  OR2 I33 (comp_0[33:33], i_0r0[33:33], i_0r1[33:33]);
  C3 I34 (simp361_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I35 (simp361_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C3 I36 (simp361_0[2:2], comp_0[6:6], comp_0[7:7], comp_0[8:8]);
  C3 I37 (simp361_0[3:3], comp_0[9:9], comp_0[10:10], comp_0[11:11]);
  C3 I38 (simp361_0[4:4], comp_0[12:12], comp_0[13:13], comp_0[14:14]);
  C3 I39 (simp361_0[5:5], comp_0[15:15], comp_0[16:16], comp_0[17:17]);
  C3 I40 (simp361_0[6:6], comp_0[18:18], comp_0[19:19], comp_0[20:20]);
  C3 I41 (simp361_0[7:7], comp_0[21:21], comp_0[22:22], comp_0[23:23]);
  C3 I42 (simp361_0[8:8], comp_0[24:24], comp_0[25:25], comp_0[26:26]);
  C3 I43 (simp361_0[9:9], comp_0[27:27], comp_0[28:28], comp_0[29:29]);
  C3 I44 (simp361_0[10:10], comp_0[30:30], comp_0[31:31], comp_0[32:32]);
  BUFF I45 (simp361_0[11:11], comp_0[33:33]);
  C3 I46 (simp362_0[0:0], simp361_0[0:0], simp361_0[1:1], simp361_0[2:2]);
  C3 I47 (simp362_0[1:1], simp361_0[3:3], simp361_0[4:4], simp361_0[5:5]);
  C3 I48 (simp362_0[2:2], simp361_0[6:6], simp361_0[7:7], simp361_0[8:8]);
  C3 I49 (simp362_0[3:3], simp361_0[9:9], simp361_0[10:10], simp361_0[11:11]);
  C3 I50 (simp363_0[0:0], simp362_0[0:0], simp362_0[1:1], simp362_0[2:2]);
  BUFF I51 (simp363_0[1:1], simp362_0[3:3]);
  C2 I52 (icomplete_0, simp363_0[0:0], simp363_0[1:1]);
  C2 I53 (o_0r0[0:0], i_0r0[0:0], icomplete_0);
  BUFF I54 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I55 (o_0r0[2:2], i_0r0[2:2]);
  BUFF I56 (o_0r0[3:3], i_0r0[3:3]);
  BUFF I57 (o_0r0[4:4], i_0r0[4:4]);
  BUFF I58 (o_0r0[5:5], i_0r0[5:5]);
  BUFF I59 (o_0r0[6:6], i_0r0[6:6]);
  BUFF I60 (o_0r0[7:7], i_0r0[7:7]);
  BUFF I61 (o_0r0[8:8], i_0r0[8:8]);
  BUFF I62 (o_0r0[9:9], i_0r0[9:9]);
  BUFF I63 (o_0r0[10:10], i_0r0[10:10]);
  BUFF I64 (o_0r0[11:11], i_0r0[11:11]);
  BUFF I65 (o_0r0[12:12], i_0r0[12:12]);
  BUFF I66 (o_0r0[13:13], i_0r0[13:13]);
  BUFF I67 (o_0r0[14:14], i_0r0[14:14]);
  BUFF I68 (o_0r0[15:15], i_0r0[15:15]);
  BUFF I69 (o_0r0[16:16], i_0r0[16:16]);
  BUFF I70 (o_0r0[17:17], i_0r0[17:17]);
  BUFF I71 (o_0r0[18:18], i_0r0[18:18]);
  BUFF I72 (o_0r0[19:19], i_0r0[19:19]);
  BUFF I73 (o_0r0[20:20], i_0r0[20:20]);
  BUFF I74 (o_0r0[21:21], i_0r0[21:21]);
  BUFF I75 (o_0r0[22:22], i_0r0[22:22]);
  BUFF I76 (o_0r0[23:23], i_0r0[23:23]);
  BUFF I77 (o_0r0[24:24], i_0r0[24:24]);
  BUFF I78 (o_0r0[25:25], i_0r0[25:25]);
  BUFF I79 (o_0r0[26:26], i_0r0[26:26]);
  BUFF I80 (o_0r0[27:27], i_0r0[27:27]);
  BUFF I81 (o_0r0[28:28], i_0r0[28:28]);
  BUFF I82 (o_0r0[29:29], i_0r0[29:29]);
  BUFF I83 (o_0r0[30:30], i_0r0[30:30]);
  BUFF I84 (o_0r0[31:31], i_0r0[31:31]);
  BUFF I85 (o_1r0[0:0], i_0r0[0:0]);
  BUFF I86 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I87 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I88 (o_1r0[3:3], i_0r0[3:3]);
  BUFF I89 (o_1r0[4:4], i_0r0[4:4]);
  BUFF I90 (o_1r0[5:5], i_0r0[5:5]);
  BUFF I91 (o_1r0[6:6], i_0r0[6:6]);
  BUFF I92 (o_1r0[7:7], i_0r0[7:7]);
  BUFF I93 (o_1r0[8:8], i_0r0[8:8]);
  BUFF I94 (o_1r0[9:9], i_0r0[9:9]);
  BUFF I95 (o_1r0[10:10], i_0r0[10:10]);
  BUFF I96 (o_1r0[11:11], i_0r0[11:11]);
  BUFF I97 (o_1r0[12:12], i_0r0[12:12]);
  BUFF I98 (o_1r0[13:13], i_0r0[13:13]);
  BUFF I99 (o_1r0[14:14], i_0r0[14:14]);
  BUFF I100 (o_1r0[15:15], i_0r0[15:15]);
  BUFF I101 (o_1r0[16:16], i_0r0[16:16]);
  BUFF I102 (o_1r0[17:17], i_0r0[17:17]);
  BUFF I103 (o_1r0[18:18], i_0r0[18:18]);
  BUFF I104 (o_1r0[19:19], i_0r0[19:19]);
  BUFF I105 (o_1r0[20:20], i_0r0[20:20]);
  BUFF I106 (o_1r0[21:21], i_0r0[21:21]);
  BUFF I107 (o_1r0[22:22], i_0r0[22:22]);
  BUFF I108 (o_1r0[23:23], i_0r0[23:23]);
  BUFF I109 (o_1r0[24:24], i_0r0[24:24]);
  BUFF I110 (o_1r0[25:25], i_0r0[25:25]);
  BUFF I111 (o_1r0[26:26], i_0r0[26:26]);
  BUFF I112 (o_1r0[27:27], i_0r0[27:27]);
  BUFF I113 (o_1r0[28:28], i_0r0[28:28]);
  BUFF I114 (o_1r0[29:29], i_0r0[29:29]);
  BUFF I115 (o_1r0[30:30], i_0r0[30:30]);
  BUFF I116 (o_1r0[31:31], i_0r0[31:31]);
  BUFF I117 (o_1r0[32:32], i_0r0[32:32]);
  BUFF I118 (o_1r0[33:33], i_0r0[33:33]);
  C2 I119 (o_2r0[0:0], i_0r0[1:1], icomplete_0);
  BUFF I120 (o_2r0[1:1], i_0r0[2:2]);
  BUFF I121 (o_2r0[2:2], i_0r0[3:3]);
  BUFF I122 (o_2r0[3:3], i_0r0[4:4]);
  BUFF I123 (o_2r0[4:4], i_0r0[5:5]);
  BUFF I124 (o_2r0[5:5], i_0r0[6:6]);
  BUFF I125 (o_2r0[6:6], i_0r0[7:7]);
  BUFF I126 (o_2r0[7:7], i_0r0[8:8]);
  BUFF I127 (o_2r0[8:8], i_0r0[9:9]);
  BUFF I128 (o_2r0[9:9], i_0r0[10:10]);
  BUFF I129 (o_2r0[10:10], i_0r0[11:11]);
  BUFF I130 (o_2r0[11:11], i_0r0[12:12]);
  BUFF I131 (o_2r0[12:12], i_0r0[13:13]);
  BUFF I132 (o_2r0[13:13], i_0r0[14:14]);
  BUFF I133 (o_2r0[14:14], i_0r0[15:15]);
  BUFF I134 (o_2r0[15:15], i_0r0[16:16]);
  BUFF I135 (o_2r0[16:16], i_0r0[17:17]);
  BUFF I136 (o_2r0[17:17], i_0r0[18:18]);
  BUFF I137 (o_2r0[18:18], i_0r0[19:19]);
  BUFF I138 (o_2r0[19:19], i_0r0[20:20]);
  BUFF I139 (o_2r0[20:20], i_0r0[21:21]);
  BUFF I140 (o_2r0[21:21], i_0r0[22:22]);
  BUFF I141 (o_2r0[22:22], i_0r0[23:23]);
  BUFF I142 (o_2r0[23:23], i_0r0[24:24]);
  BUFF I143 (o_2r0[24:24], i_0r0[25:25]);
  BUFF I144 (o_2r0[25:25], i_0r0[26:26]);
  BUFF I145 (o_2r0[26:26], i_0r0[27:27]);
  BUFF I146 (o_2r0[27:27], i_0r0[28:28]);
  BUFF I147 (o_2r0[28:28], i_0r0[29:29]);
  BUFF I148 (o_2r0[29:29], i_0r0[30:30]);
  BUFF I149 (o_2r0[30:30], i_0r0[31:31]);
  BUFF I150 (o_2r0[31:31], i_0r0[32:32]);
  C2 I151 (o_0r1[0:0], i_0r1[0:0], icomplete_0);
  BUFF I152 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I153 (o_0r1[2:2], i_0r1[2:2]);
  BUFF I154 (o_0r1[3:3], i_0r1[3:3]);
  BUFF I155 (o_0r1[4:4], i_0r1[4:4]);
  BUFF I156 (o_0r1[5:5], i_0r1[5:5]);
  BUFF I157 (o_0r1[6:6], i_0r1[6:6]);
  BUFF I158 (o_0r1[7:7], i_0r1[7:7]);
  BUFF I159 (o_0r1[8:8], i_0r1[8:8]);
  BUFF I160 (o_0r1[9:9], i_0r1[9:9]);
  BUFF I161 (o_0r1[10:10], i_0r1[10:10]);
  BUFF I162 (o_0r1[11:11], i_0r1[11:11]);
  BUFF I163 (o_0r1[12:12], i_0r1[12:12]);
  BUFF I164 (o_0r1[13:13], i_0r1[13:13]);
  BUFF I165 (o_0r1[14:14], i_0r1[14:14]);
  BUFF I166 (o_0r1[15:15], i_0r1[15:15]);
  BUFF I167 (o_0r1[16:16], i_0r1[16:16]);
  BUFF I168 (o_0r1[17:17], i_0r1[17:17]);
  BUFF I169 (o_0r1[18:18], i_0r1[18:18]);
  BUFF I170 (o_0r1[19:19], i_0r1[19:19]);
  BUFF I171 (o_0r1[20:20], i_0r1[20:20]);
  BUFF I172 (o_0r1[21:21], i_0r1[21:21]);
  BUFF I173 (o_0r1[22:22], i_0r1[22:22]);
  BUFF I174 (o_0r1[23:23], i_0r1[23:23]);
  BUFF I175 (o_0r1[24:24], i_0r1[24:24]);
  BUFF I176 (o_0r1[25:25], i_0r1[25:25]);
  BUFF I177 (o_0r1[26:26], i_0r1[26:26]);
  BUFF I178 (o_0r1[27:27], i_0r1[27:27]);
  BUFF I179 (o_0r1[28:28], i_0r1[28:28]);
  BUFF I180 (o_0r1[29:29], i_0r1[29:29]);
  BUFF I181 (o_0r1[30:30], i_0r1[30:30]);
  BUFF I182 (o_0r1[31:31], i_0r1[31:31]);
  BUFF I183 (o_1r1[0:0], i_0r1[0:0]);
  BUFF I184 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I185 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I186 (o_1r1[3:3], i_0r1[3:3]);
  BUFF I187 (o_1r1[4:4], i_0r1[4:4]);
  BUFF I188 (o_1r1[5:5], i_0r1[5:5]);
  BUFF I189 (o_1r1[6:6], i_0r1[6:6]);
  BUFF I190 (o_1r1[7:7], i_0r1[7:7]);
  BUFF I191 (o_1r1[8:8], i_0r1[8:8]);
  BUFF I192 (o_1r1[9:9], i_0r1[9:9]);
  BUFF I193 (o_1r1[10:10], i_0r1[10:10]);
  BUFF I194 (o_1r1[11:11], i_0r1[11:11]);
  BUFF I195 (o_1r1[12:12], i_0r1[12:12]);
  BUFF I196 (o_1r1[13:13], i_0r1[13:13]);
  BUFF I197 (o_1r1[14:14], i_0r1[14:14]);
  BUFF I198 (o_1r1[15:15], i_0r1[15:15]);
  BUFF I199 (o_1r1[16:16], i_0r1[16:16]);
  BUFF I200 (o_1r1[17:17], i_0r1[17:17]);
  BUFF I201 (o_1r1[18:18], i_0r1[18:18]);
  BUFF I202 (o_1r1[19:19], i_0r1[19:19]);
  BUFF I203 (o_1r1[20:20], i_0r1[20:20]);
  BUFF I204 (o_1r1[21:21], i_0r1[21:21]);
  BUFF I205 (o_1r1[22:22], i_0r1[22:22]);
  BUFF I206 (o_1r1[23:23], i_0r1[23:23]);
  BUFF I207 (o_1r1[24:24], i_0r1[24:24]);
  BUFF I208 (o_1r1[25:25], i_0r1[25:25]);
  BUFF I209 (o_1r1[26:26], i_0r1[26:26]);
  BUFF I210 (o_1r1[27:27], i_0r1[27:27]);
  BUFF I211 (o_1r1[28:28], i_0r1[28:28]);
  BUFF I212 (o_1r1[29:29], i_0r1[29:29]);
  BUFF I213 (o_1r1[30:30], i_0r1[30:30]);
  BUFF I214 (o_1r1[31:31], i_0r1[31:31]);
  BUFF I215 (o_1r1[32:32], i_0r1[32:32]);
  BUFF I216 (o_1r1[33:33], i_0r1[33:33]);
  C2 I217 (o_2r1[0:0], i_0r1[1:1], icomplete_0);
  BUFF I218 (o_2r1[1:1], i_0r1[2:2]);
  BUFF I219 (o_2r1[2:2], i_0r1[3:3]);
  BUFF I220 (o_2r1[3:3], i_0r1[4:4]);
  BUFF I221 (o_2r1[4:4], i_0r1[5:5]);
  BUFF I222 (o_2r1[5:5], i_0r1[6:6]);
  BUFF I223 (o_2r1[6:6], i_0r1[7:7]);
  BUFF I224 (o_2r1[7:7], i_0r1[8:8]);
  BUFF I225 (o_2r1[8:8], i_0r1[9:9]);
  BUFF I226 (o_2r1[9:9], i_0r1[10:10]);
  BUFF I227 (o_2r1[10:10], i_0r1[11:11]);
  BUFF I228 (o_2r1[11:11], i_0r1[12:12]);
  BUFF I229 (o_2r1[12:12], i_0r1[13:13]);
  BUFF I230 (o_2r1[13:13], i_0r1[14:14]);
  BUFF I231 (o_2r1[14:14], i_0r1[15:15]);
  BUFF I232 (o_2r1[15:15], i_0r1[16:16]);
  BUFF I233 (o_2r1[16:16], i_0r1[17:17]);
  BUFF I234 (o_2r1[17:17], i_0r1[18:18]);
  BUFF I235 (o_2r1[18:18], i_0r1[19:19]);
  BUFF I236 (o_2r1[19:19], i_0r1[20:20]);
  BUFF I237 (o_2r1[20:20], i_0r1[21:21]);
  BUFF I238 (o_2r1[21:21], i_0r1[22:22]);
  BUFF I239 (o_2r1[22:22], i_0r1[23:23]);
  BUFF I240 (o_2r1[23:23], i_0r1[24:24]);
  BUFF I241 (o_2r1[24:24], i_0r1[25:25]);
  BUFF I242 (o_2r1[25:25], i_0r1[26:26]);
  BUFF I243 (o_2r1[26:26], i_0r1[27:27]);
  BUFF I244 (o_2r1[27:27], i_0r1[28:28]);
  BUFF I245 (o_2r1[28:28], i_0r1[29:29]);
  BUFF I246 (o_2r1[29:29], i_0r1[30:30]);
  BUFF I247 (o_2r1[30:30], i_0r1[31:31]);
  BUFF I248 (o_2r1[31:31], i_0r1[32:32]);
  C3 I249 (simp2341_0[0:0], icomplete_0, o_0a, o_1a);
  BUFF I250 (simp2341_0[1:1], o_2a);
  C2 I251 (i_0a, simp2341_0[0:0], simp2341_0[1:1]);
endmodule

// tkf8mo0w4_o0w7_o0w4_o0w4 TeakF [0,0,0,0] [One 8,Many [4,7,4,4]]
module tkf8mo0w4_o0w7_o0w4_o0w4 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r0, o_1r1, o_1a, o_2r0, o_2r1, o_2a, o_3r0, o_3r1, o_3a, reset);
  input [7:0] i_0r0;
  input [7:0] i_0r1;
  output i_0a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  output [6:0] o_1r0;
  output [6:0] o_1r1;
  input o_1a;
  output [3:0] o_2r0;
  output [3:0] o_2r1;
  input o_2a;
  output [3:0] o_3r0;
  output [3:0] o_3r1;
  input o_3a;
  input reset;
  wire icomplete_0;
  wire [7:0] comp_0;
  wire [2:0] simp101_0;
  wire [1:0] simp501_0;
  OR2 I0 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (comp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (comp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  C3 I8 (simp101_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I9 (simp101_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C2 I10 (simp101_0[2:2], comp_0[6:6], comp_0[7:7]);
  C3 I11 (icomplete_0, simp101_0[0:0], simp101_0[1:1], simp101_0[2:2]);
  C2 I12 (o_0r0[0:0], i_0r0[0:0], icomplete_0);
  BUFF I13 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I14 (o_0r0[2:2], i_0r0[2:2]);
  BUFF I15 (o_0r0[3:3], i_0r0[3:3]);
  C2 I16 (o_1r0[0:0], i_0r0[0:0], icomplete_0);
  BUFF I17 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I18 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I19 (o_1r0[3:3], i_0r0[3:3]);
  BUFF I20 (o_1r0[4:4], i_0r0[4:4]);
  BUFF I21 (o_1r0[5:5], i_0r0[5:5]);
  BUFF I22 (o_1r0[6:6], i_0r0[6:6]);
  C2 I23 (o_2r0[0:0], i_0r0[0:0], icomplete_0);
  BUFF I24 (o_2r0[1:1], i_0r0[1:1]);
  BUFF I25 (o_2r0[2:2], i_0r0[2:2]);
  BUFF I26 (o_2r0[3:3], i_0r0[3:3]);
  C2 I27 (o_3r0[0:0], i_0r0[0:0], icomplete_0);
  BUFF I28 (o_3r0[1:1], i_0r0[1:1]);
  BUFF I29 (o_3r0[2:2], i_0r0[2:2]);
  BUFF I30 (o_3r0[3:3], i_0r0[3:3]);
  C2 I31 (o_0r1[0:0], i_0r1[0:0], icomplete_0);
  BUFF I32 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I33 (o_0r1[2:2], i_0r1[2:2]);
  BUFF I34 (o_0r1[3:3], i_0r1[3:3]);
  C2 I35 (o_1r1[0:0], i_0r1[0:0], icomplete_0);
  BUFF I36 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I37 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I38 (o_1r1[3:3], i_0r1[3:3]);
  BUFF I39 (o_1r1[4:4], i_0r1[4:4]);
  BUFF I40 (o_1r1[5:5], i_0r1[5:5]);
  BUFF I41 (o_1r1[6:6], i_0r1[6:6]);
  C2 I42 (o_2r1[0:0], i_0r1[0:0], icomplete_0);
  BUFF I43 (o_2r1[1:1], i_0r1[1:1]);
  BUFF I44 (o_2r1[2:2], i_0r1[2:2]);
  BUFF I45 (o_2r1[3:3], i_0r1[3:3]);
  C2 I46 (o_3r1[0:0], i_0r1[0:0], icomplete_0);
  BUFF I47 (o_3r1[1:1], i_0r1[1:1]);
  BUFF I48 (o_3r1[2:2], i_0r1[2:2]);
  BUFF I49 (o_3r1[3:3], i_0r1[3:3]);
  C3 I50 (simp501_0[0:0], icomplete_0, o_0a, o_1a);
  C2 I51 (simp501_0[1:1], o_2a, o_3a);
  C2 I52 (i_0a, simp501_0[0:0], simp501_0[1:1]);
endmodule

// tkj4m0_4 TeakJ [Many [0,4],One 4]
module tkj4m0_4 (i_0r, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  input [3:0] i_1r0;
  input [3:0] i_1r1;
  output i_1a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [3:0] joinf_0;
  wire [3:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_1r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_1r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_1r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_1r0[3:3]);
  BUFF I4 (joint_0[0:0], i_1r1[0:0]);
  BUFF I5 (joint_0[1:1], i_1r1[1:1]);
  BUFF I6 (joint_0[2:2], i_1r1[2:2]);
  BUFF I7 (joint_0[3:3], i_1r1[3:3]);
  BUFF I8 (icomplete_0, i_0r);
  C2 I9 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I10 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I11 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I12 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I13 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I14 (o_0r1[1:1], joint_0[1:1]);
  BUFF I15 (o_0r1[2:2], joint_0[2:2]);
  BUFF I16 (o_0r1[3:3], joint_0[3:3]);
  BUFF I17 (i_0a, o_0a);
  BUFF I18 (i_1a, o_0a);
endmodule

// tkj4m4_0 TeakJ [Many [4,0],One 4]
module tkj4m4_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [3:0] joinf_0;
  wire [3:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joint_0[0:0], i_0r1[0:0]);
  BUFF I5 (joint_0[1:1], i_0r1[1:1]);
  BUFF I6 (joint_0[2:2], i_0r1[2:2]);
  BUFF I7 (joint_0[3:3], i_0r1[3:3]);
  BUFF I8 (icomplete_0, i_1r);
  C2 I9 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I10 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I11 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I12 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I13 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I14 (o_0r1[1:1], joint_0[1:1]);
  BUFF I15 (o_0r1[2:2], joint_0[2:2]);
  BUFF I16 (o_0r1[3:3], joint_0[3:3]);
  BUFF I17 (i_0a, o_0a);
  BUFF I18 (i_1a, o_0a);
endmodule

// tkvctrlfisfc9_wo0w9_ro0w4o5w1o4w1o8w1 TeakV "ctrl-fi-sfc" 9 [] [0] [0,5,4,8] [Many [9],Many [0],Many
//    [0,0,0,0],Many [4,1,1,1]]
module tkvctrlfisfc9_wo0w9_ro0w4o5w1o4w1o8w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, reset);
  input [8:0] wg_0r0;
  input [8:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  output [3:0] rd_0r0;
  output [3:0] rd_0r1;
  input rd_0a;
  output rd_1r0;
  output rd_1r1;
  input rd_1a;
  output rd_2r0;
  output rd_2r1;
  input rd_2a;
  output rd_3r0;
  output rd_3r1;
  input rd_3a;
  input reset;
  wire [8:0] wf_0;
  wire [8:0] wt_0;
  wire [8:0] df_0;
  wire [8:0] dt_0;
  wire wc_0;
  wire [8:0] wacks_0;
  wire [8:0] wenr_0;
  wire [8:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [8:0] drlgf_0;
  wire [8:0] drlgt_0;
  wire [8:0] comp0_0;
  wire [2:0] simp771_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [8:0] conwgit_0;
  wire [8:0] conwgif_0;
  wire conwig_0;
  wire [3:0] simp1311_0;
  wire [1:0] simp1312_0;
  wire [2:0] simp1461_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I11 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I12 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I13 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I14 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I15 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I16 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I17 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I18 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I19 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I20 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I21 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I22 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I23 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I24 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I25 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I26 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I27 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  NOR2 I28 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I29 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I30 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I31 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I32 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I33 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I34 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I35 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I36 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR3 I37 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I38 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I39 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I40 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I41 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I42 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I43 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I44 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I45 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  AO22 I46 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I47 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I48 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I49 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I50 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I51 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I52 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I53 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I54 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  OR2 I55 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I56 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I57 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I58 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I59 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I60 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I61 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I62 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I63 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  C3 I64 (simp771_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I65 (simp771_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I66 (simp771_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I67 (wc_0, simp771_0[0:0], simp771_0[1:1], simp771_0[2:2]);
  AND2 I68 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I69 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I70 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I71 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I72 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I73 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I74 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I75 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I76 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I77 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I78 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I79 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I80 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I81 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I82 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I83 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I84 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I85 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  BUFF I86 (conwigc_0, wc_0);
  AO22 I87 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I88 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I89 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I90 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I91 (wenr_0[0:0], wc_0);
  BUFF I92 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I93 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I94 (wenr_0[1:1], wc_0);
  BUFF I95 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I96 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I97 (wenr_0[2:2], wc_0);
  BUFF I98 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I99 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I100 (wenr_0[3:3], wc_0);
  BUFF I101 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I102 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I103 (wenr_0[4:4], wc_0);
  BUFF I104 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I105 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I106 (wenr_0[5:5], wc_0);
  BUFF I107 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I108 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I109 (wenr_0[6:6], wc_0);
  BUFF I110 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I111 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I112 (wenr_0[7:7], wc_0);
  BUFF I113 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I114 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I115 (wenr_0[8:8], wc_0);
  C3 I116 (simp1311_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I117 (simp1311_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I118 (simp1311_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  BUFF I119 (simp1311_0[3:3], wacks_0[8:8]);
  C3 I120 (simp1312_0[0:0], simp1311_0[0:0], simp1311_0[1:1], simp1311_0[2:2]);
  BUFF I121 (simp1312_0[1:1], simp1311_0[3:3]);
  C2 I122 (wd_0r, simp1312_0[0:0], simp1312_0[1:1]);
  AND2 I123 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I124 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I125 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I126 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I127 (rd_1r0, df_0[5:5], rg_1r);
  AND2 I128 (rd_2r0, df_0[4:4], rg_2r);
  AND2 I129 (rd_3r0, df_0[8:8], rg_3r);
  AND2 I130 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I131 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I132 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I133 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I134 (rd_1r1, dt_0[5:5], rg_1r);
  AND2 I135 (rd_2r1, dt_0[4:4], rg_2r);
  AND2 I136 (rd_3r1, dt_0[8:8], rg_3r);
  NOR3 I137 (simp1461_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I138 (simp1461_0[1:1], rg_3r, rg_0a, rg_1a);
  NOR2 I139 (simp1461_0[2:2], rg_2a, rg_3a);
  NAND3 I140 (anyread_0, simp1461_0[0:0], simp1461_0[1:1], simp1461_0[2:2]);
  BUFF I141 (wg_0a, wd_0a);
  BUFF I142 (rg_0a, rd_0a);
  BUFF I143 (rg_1a, rd_1a);
  BUFF I144 (rg_2a, rd_2a);
  BUFF I145 (rg_3a, rd_3a);
endmodule

// tko34m34_1xori0w1bi0w1b_2apt1o0w1bi1w33b TeakO [
//     (1,TeakOp TeakOpXor [(0,0,1),(0,0,1)]),
//     (2,TeakOAppend 1 [(1,0,1),(0,1,33)])] [One 34,One 34]
module tko34m34_1xori0w1bi0w1b_2apt1o0w1bi1w33b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [33:0] i_0r0;
  input [33:0] i_0r1;
  output i_0a;
  output [33:0] o_0r0;
  output [33:0] o_0r1;
  input o_0a;
  input reset;
  wire termf_1;
  wire termt_1;
  wire [3:0] op1_0_0;
  C2 I0 (op1_0_0[0:0], i_0r0[0:0], i_0r0[0:0]);
  C2 I1 (op1_0_0[1:1], i_0r0[0:0], i_0r1[0:0]);
  C2 I2 (op1_0_0[2:2], i_0r1[0:0], i_0r0[0:0]);
  C2 I3 (op1_0_0[3:3], i_0r1[0:0], i_0r1[0:0]);
  OR2 I4 (termf_1, op1_0_0[0:0], op1_0_0[3:3]);
  OR2 I5 (termt_1, op1_0_0[1:1], op1_0_0[2:2]);
  BUFF I6 (o_0r0[0:0], termf_1);
  BUFF I7 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I8 (o_0r0[2:2], i_0r0[2:2]);
  BUFF I9 (o_0r0[3:3], i_0r0[3:3]);
  BUFF I10 (o_0r0[4:4], i_0r0[4:4]);
  BUFF I11 (o_0r0[5:5], i_0r0[5:5]);
  BUFF I12 (o_0r0[6:6], i_0r0[6:6]);
  BUFF I13 (o_0r0[7:7], i_0r0[7:7]);
  BUFF I14 (o_0r0[8:8], i_0r0[8:8]);
  BUFF I15 (o_0r0[9:9], i_0r0[9:9]);
  BUFF I16 (o_0r0[10:10], i_0r0[10:10]);
  BUFF I17 (o_0r0[11:11], i_0r0[11:11]);
  BUFF I18 (o_0r0[12:12], i_0r0[12:12]);
  BUFF I19 (o_0r0[13:13], i_0r0[13:13]);
  BUFF I20 (o_0r0[14:14], i_0r0[14:14]);
  BUFF I21 (o_0r0[15:15], i_0r0[15:15]);
  BUFF I22 (o_0r0[16:16], i_0r0[16:16]);
  BUFF I23 (o_0r0[17:17], i_0r0[17:17]);
  BUFF I24 (o_0r0[18:18], i_0r0[18:18]);
  BUFF I25 (o_0r0[19:19], i_0r0[19:19]);
  BUFF I26 (o_0r0[20:20], i_0r0[20:20]);
  BUFF I27 (o_0r0[21:21], i_0r0[21:21]);
  BUFF I28 (o_0r0[22:22], i_0r0[22:22]);
  BUFF I29 (o_0r0[23:23], i_0r0[23:23]);
  BUFF I30 (o_0r0[24:24], i_0r0[24:24]);
  BUFF I31 (o_0r0[25:25], i_0r0[25:25]);
  BUFF I32 (o_0r0[26:26], i_0r0[26:26]);
  BUFF I33 (o_0r0[27:27], i_0r0[27:27]);
  BUFF I34 (o_0r0[28:28], i_0r0[28:28]);
  BUFF I35 (o_0r0[29:29], i_0r0[29:29]);
  BUFF I36 (o_0r0[30:30], i_0r0[30:30]);
  BUFF I37 (o_0r0[31:31], i_0r0[31:31]);
  BUFF I38 (o_0r0[32:32], i_0r0[32:32]);
  BUFF I39 (o_0r0[33:33], i_0r0[33:33]);
  BUFF I40 (o_0r1[0:0], termt_1);
  BUFF I41 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I42 (o_0r1[2:2], i_0r1[2:2]);
  BUFF I43 (o_0r1[3:3], i_0r1[3:3]);
  BUFF I44 (o_0r1[4:4], i_0r1[4:4]);
  BUFF I45 (o_0r1[5:5], i_0r1[5:5]);
  BUFF I46 (o_0r1[6:6], i_0r1[6:6]);
  BUFF I47 (o_0r1[7:7], i_0r1[7:7]);
  BUFF I48 (o_0r1[8:8], i_0r1[8:8]);
  BUFF I49 (o_0r1[9:9], i_0r1[9:9]);
  BUFF I50 (o_0r1[10:10], i_0r1[10:10]);
  BUFF I51 (o_0r1[11:11], i_0r1[11:11]);
  BUFF I52 (o_0r1[12:12], i_0r1[12:12]);
  BUFF I53 (o_0r1[13:13], i_0r1[13:13]);
  BUFF I54 (o_0r1[14:14], i_0r1[14:14]);
  BUFF I55 (o_0r1[15:15], i_0r1[15:15]);
  BUFF I56 (o_0r1[16:16], i_0r1[16:16]);
  BUFF I57 (o_0r1[17:17], i_0r1[17:17]);
  BUFF I58 (o_0r1[18:18], i_0r1[18:18]);
  BUFF I59 (o_0r1[19:19], i_0r1[19:19]);
  BUFF I60 (o_0r1[20:20], i_0r1[20:20]);
  BUFF I61 (o_0r1[21:21], i_0r1[21:21]);
  BUFF I62 (o_0r1[22:22], i_0r1[22:22]);
  BUFF I63 (o_0r1[23:23], i_0r1[23:23]);
  BUFF I64 (o_0r1[24:24], i_0r1[24:24]);
  BUFF I65 (o_0r1[25:25], i_0r1[25:25]);
  BUFF I66 (o_0r1[26:26], i_0r1[26:26]);
  BUFF I67 (o_0r1[27:27], i_0r1[27:27]);
  BUFF I68 (o_0r1[28:28], i_0r1[28:28]);
  BUFF I69 (o_0r1[29:29], i_0r1[29:29]);
  BUFF I70 (o_0r1[30:30], i_0r1[30:30]);
  BUFF I71 (o_0r1[31:31], i_0r1[31:31]);
  BUFF I72 (o_0r1[32:32], i_0r1[32:32]);
  BUFF I73 (o_0r1[33:33], i_0r1[33:33]);
  BUFF I74 (i_0a, o_0a);
endmodule

// tko8m9_1api0w8bi0w1b TeakO [
//     (1,TeakOAppend 1 [(0,0,8),(0,0,1)])] [One 8,One 9]
module tko8m9_1api0w8bi0w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [7:0] i_0r0;
  input [7:0] i_0r1;
  output i_0a;
  output [8:0] o_0r0;
  output [8:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r0[0:0]);
  BUFF I1 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I2 (o_0r0[2:2], i_0r0[2:2]);
  BUFF I3 (o_0r0[3:3], i_0r0[3:3]);
  BUFF I4 (o_0r0[4:4], i_0r0[4:4]);
  BUFF I5 (o_0r0[5:5], i_0r0[5:5]);
  BUFF I6 (o_0r0[6:6], i_0r0[6:6]);
  BUFF I7 (o_0r0[7:7], i_0r0[7:7]);
  BUFF I8 (o_0r0[8:8], i_0r0[0:0]);
  BUFF I9 (o_0r1[0:0], i_0r1[0:0]);
  BUFF I10 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I11 (o_0r1[2:2], i_0r1[2:2]);
  BUFF I12 (o_0r1[3:3], i_0r1[3:3]);
  BUFF I13 (o_0r1[4:4], i_0r1[4:4]);
  BUFF I14 (o_0r1[5:5], i_0r1[5:5]);
  BUFF I15 (o_0r1[6:6], i_0r1[6:6]);
  BUFF I16 (o_0r1[7:7], i_0r1[7:7]);
  BUFF I17 (o_0r1[8:8], i_0r1[0:0]);
  BUFF I18 (i_0a, o_0a);
endmodule

// tkj33m1_32 TeakJ [Many [1,32],One 33]
module tkj33m1_32 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r0);
  BUFF I1 (o_0r0[1:1], i_1r0[0:0]);
  BUFF I2 (o_0r0[2:2], i_1r0[1:1]);
  BUFF I3 (o_0r0[3:3], i_1r0[2:2]);
  BUFF I4 (o_0r0[4:4], i_1r0[3:3]);
  BUFF I5 (o_0r0[5:5], i_1r0[4:4]);
  BUFF I6 (o_0r0[6:6], i_1r0[5:5]);
  BUFF I7 (o_0r0[7:7], i_1r0[6:6]);
  BUFF I8 (o_0r0[8:8], i_1r0[7:7]);
  BUFF I9 (o_0r0[9:9], i_1r0[8:8]);
  BUFF I10 (o_0r0[10:10], i_1r0[9:9]);
  BUFF I11 (o_0r0[11:11], i_1r0[10:10]);
  BUFF I12 (o_0r0[12:12], i_1r0[11:11]);
  BUFF I13 (o_0r0[13:13], i_1r0[12:12]);
  BUFF I14 (o_0r0[14:14], i_1r0[13:13]);
  BUFF I15 (o_0r0[15:15], i_1r0[14:14]);
  BUFF I16 (o_0r0[16:16], i_1r0[15:15]);
  BUFF I17 (o_0r0[17:17], i_1r0[16:16]);
  BUFF I18 (o_0r0[18:18], i_1r0[17:17]);
  BUFF I19 (o_0r0[19:19], i_1r0[18:18]);
  BUFF I20 (o_0r0[20:20], i_1r0[19:19]);
  BUFF I21 (o_0r0[21:21], i_1r0[20:20]);
  BUFF I22 (o_0r0[22:22], i_1r0[21:21]);
  BUFF I23 (o_0r0[23:23], i_1r0[22:22]);
  BUFF I24 (o_0r0[24:24], i_1r0[23:23]);
  BUFF I25 (o_0r0[25:25], i_1r0[24:24]);
  BUFF I26 (o_0r0[26:26], i_1r0[25:25]);
  BUFF I27 (o_0r0[27:27], i_1r0[26:26]);
  BUFF I28 (o_0r0[28:28], i_1r0[27:27]);
  BUFF I29 (o_0r0[29:29], i_1r0[28:28]);
  BUFF I30 (o_0r0[30:30], i_1r0[29:29]);
  BUFF I31 (o_0r0[31:31], i_1r0[30:30]);
  BUFF I32 (o_0r0[32:32], i_1r0[31:31]);
  BUFF I33 (o_0r1[0:0], i_0r1);
  BUFF I34 (o_0r1[1:1], i_1r1[0:0]);
  BUFF I35 (o_0r1[2:2], i_1r1[1:1]);
  BUFF I36 (o_0r1[3:3], i_1r1[2:2]);
  BUFF I37 (o_0r1[4:4], i_1r1[3:3]);
  BUFF I38 (o_0r1[5:5], i_1r1[4:4]);
  BUFF I39 (o_0r1[6:6], i_1r1[5:5]);
  BUFF I40 (o_0r1[7:7], i_1r1[6:6]);
  BUFF I41 (o_0r1[8:8], i_1r1[7:7]);
  BUFF I42 (o_0r1[9:9], i_1r1[8:8]);
  BUFF I43 (o_0r1[10:10], i_1r1[9:9]);
  BUFF I44 (o_0r1[11:11], i_1r1[10:10]);
  BUFF I45 (o_0r1[12:12], i_1r1[11:11]);
  BUFF I46 (o_0r1[13:13], i_1r1[12:12]);
  BUFF I47 (o_0r1[14:14], i_1r1[13:13]);
  BUFF I48 (o_0r1[15:15], i_1r1[14:14]);
  BUFF I49 (o_0r1[16:16], i_1r1[15:15]);
  BUFF I50 (o_0r1[17:17], i_1r1[16:16]);
  BUFF I51 (o_0r1[18:18], i_1r1[17:17]);
  BUFF I52 (o_0r1[19:19], i_1r1[18:18]);
  BUFF I53 (o_0r1[20:20], i_1r1[19:19]);
  BUFF I54 (o_0r1[21:21], i_1r1[20:20]);
  BUFF I55 (o_0r1[22:22], i_1r1[21:21]);
  BUFF I56 (o_0r1[23:23], i_1r1[22:22]);
  BUFF I57 (o_0r1[24:24], i_1r1[23:23]);
  BUFF I58 (o_0r1[25:25], i_1r1[24:24]);
  BUFF I59 (o_0r1[26:26], i_1r1[25:25]);
  BUFF I60 (o_0r1[27:27], i_1r1[26:26]);
  BUFF I61 (o_0r1[28:28], i_1r1[27:27]);
  BUFF I62 (o_0r1[29:29], i_1r1[28:28]);
  BUFF I63 (o_0r1[30:30], i_1r1[29:29]);
  BUFF I64 (o_0r1[31:31], i_1r1[30:30]);
  BUFF I65 (o_0r1[32:32], i_1r1[31:31]);
  BUFF I66 (i_0a, o_0a);
  BUFF I67 (i_1a, o_0a);
endmodule

// tks4_o0w4_0c8m1c8mcmdmemfo0w0_5m6m7o0w0_2m3mam4mbo0w4 TeakS (0+:4) [([Imp 0 8,Imp 1 8,Imp 12 0,Imp 1
//   3 0,Imp 14 0,Imp 15 0],0),([Imp 5 0,Imp 6 0,Imp 7 0],0),([Imp 2 0,Imp 3 0,Imp 10 0,Imp 4 0,Imp 11 0]
//   ,0)] [One 4,Many [0,0,4]]
module tks4_o0w4_0c8m1c8mcmdmemfo0w0_5m6m7o0w0_2m3mam4mbo0w4 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r0, o_2r1, o_2a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output [3:0] o_2r0;
  output [3:0] o_2r1;
  input o_2a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire oack_0;
  wire [5:0] match0_0;
  wire [1:0] simp91_0;
  wire [1:0] simp121_0;
  wire [1:0] simp131_0;
  wire [1:0] simp141_0;
  wire [1:0] simp151_0;
  wire [2:0] match1_0;
  wire [1:0] simp181_0;
  wire [1:0] simp191_0;
  wire [1:0] simp201_0;
  wire [4:0] match2_0;
  wire [1:0] simp221_0;
  wire [1:0] simp231_0;
  wire [1:0] simp241_0;
  wire [1:0] simp251_0;
  wire [1:0] simp261_0;
  wire [1:0] simp271_0;
  wire [3:0] comp_0;
  wire [1:0] simp361_0;
  NOR3 I0 (simp91_0[0:0], match0_0[0:0], match0_0[1:1], match0_0[2:2]);
  NOR3 I1 (simp91_0[1:1], match0_0[3:3], match0_0[4:4], match0_0[5:5]);
  NAND2 I2 (sel_0, simp91_0[0:0], simp91_0[1:1]);
  C3 I3 (match0_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I4 (match0_0[1:1], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I5 (simp121_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I6 (simp121_0[1:1], i_0r1[3:3]);
  C2 I7 (match0_0[2:2], simp121_0[0:0], simp121_0[1:1]);
  C3 I8 (simp131_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I9 (simp131_0[1:1], i_0r1[3:3]);
  C2 I10 (match0_0[3:3], simp131_0[0:0], simp131_0[1:1]);
  C3 I11 (simp141_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I12 (simp141_0[1:1], i_0r1[3:3]);
  C2 I13 (match0_0[4:4], simp141_0[0:0], simp141_0[1:1]);
  C3 I14 (simp151_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I15 (simp151_0[1:1], i_0r1[3:3]);
  C2 I16 (match0_0[5:5], simp151_0[0:0], simp151_0[1:1]);
  OR3 I17 (sel_1, match1_0[0:0], match1_0[1:1], match1_0[2:2]);
  C3 I18 (simp181_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I19 (simp181_0[1:1], i_0r0[3:3]);
  C2 I20 (match1_0[0:0], simp181_0[0:0], simp181_0[1:1]);
  C3 I21 (simp191_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I22 (simp191_0[1:1], i_0r0[3:3]);
  C2 I23 (match1_0[1:1], simp191_0[0:0], simp191_0[1:1]);
  C3 I24 (simp201_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I25 (simp201_0[1:1], i_0r0[3:3]);
  C2 I26 (match1_0[2:2], simp201_0[0:0], simp201_0[1:1]);
  NOR3 I27 (simp221_0[0:0], match2_0[0:0], match2_0[1:1], match2_0[2:2]);
  NOR2 I28 (simp221_0[1:1], match2_0[3:3], match2_0[4:4]);
  NAND2 I29 (sel_2, simp221_0[0:0], simp221_0[1:1]);
  C3 I30 (simp231_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I31 (simp231_0[1:1], i_0r0[3:3]);
  C2 I32 (match2_0[0:0], simp231_0[0:0], simp231_0[1:1]);
  C3 I33 (simp241_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I34 (simp241_0[1:1], i_0r0[3:3]);
  C2 I35 (match2_0[1:1], simp241_0[0:0], simp241_0[1:1]);
  C3 I36 (simp251_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I37 (simp251_0[1:1], i_0r1[3:3]);
  C2 I38 (match2_0[2:2], simp251_0[0:0], simp251_0[1:1]);
  C3 I39 (simp261_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I40 (simp261_0[1:1], i_0r0[3:3]);
  C2 I41 (match2_0[3:3], simp261_0[0:0], simp261_0[1:1]);
  C3 I42 (simp271_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I43 (simp271_0[1:1], i_0r1[3:3]);
  C2 I44 (match2_0[4:4], simp271_0[0:0], simp271_0[1:1]);
  C2 I45 (gsel_0, sel_0, icomplete_0);
  C2 I46 (gsel_1, sel_1, icomplete_0);
  C2 I47 (gsel_2, sel_2, icomplete_0);
  OR2 I48 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I49 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I50 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I51 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  C3 I52 (simp361_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  BUFF I53 (simp361_0[1:1], comp_0[3:3]);
  C2 I54 (icomplete_0, simp361_0[0:0], simp361_0[1:1]);
  C2 I55 (o_2r0[0:0], i_0r0[0:0], gsel_2);
  C2 I56 (o_2r0[1:1], i_0r0[1:1], gsel_2);
  C2 I57 (o_2r0[2:2], i_0r0[2:2], gsel_2);
  C2 I58 (o_2r0[3:3], i_0r0[3:3], gsel_2);
  C2 I59 (o_2r1[0:0], i_0r1[0:0], gsel_2);
  C2 I60 (o_2r1[1:1], i_0r1[1:1], gsel_2);
  C2 I61 (o_2r1[2:2], i_0r1[2:2], gsel_2);
  C2 I62 (o_2r1[3:3], i_0r1[3:3], gsel_2);
  BUFF I63 (o_0r, gsel_0);
  BUFF I64 (o_1r, gsel_1);
  OR3 I65 (oack_0, o_0a, o_1a, o_2a);
  C2 I66 (i_0a, oack_0, icomplete_0);
endmodule

// tkm2x33b TeakM [Many [33,33],One 33]
module tkm2x33b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [32:0] i_0r0;
  input [32:0] i_0r1;
  output i_0a;
  input [32:0] i_1r0;
  input [32:0] i_1r1;
  output i_1a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  wire [32:0] gfint_0;
  wire [32:0] gfint_1;
  wire [32:0] gtint_0;
  wire [32:0] gtint_1;
  wire choice_0;
  wire choice_1;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire nchosen_0;
  wire [32:0] comp0_0;
  wire [10:0] simp2421_0;
  wire [3:0] simp2422_0;
  wire [1:0] simp2423_0;
  wire [32:0] comp1_0;
  wire [10:0] simp2771_0;
  wire [3:0] simp2772_0;
  wire [1:0] simp2773_0;
  OR2 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0]);
  OR2 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1]);
  OR2 I2 (o_0r0[2:2], gfint_0[2:2], gfint_1[2:2]);
  OR2 I3 (o_0r0[3:3], gfint_0[3:3], gfint_1[3:3]);
  OR2 I4 (o_0r0[4:4], gfint_0[4:4], gfint_1[4:4]);
  OR2 I5 (o_0r0[5:5], gfint_0[5:5], gfint_1[5:5]);
  OR2 I6 (o_0r0[6:6], gfint_0[6:6], gfint_1[6:6]);
  OR2 I7 (o_0r0[7:7], gfint_0[7:7], gfint_1[7:7]);
  OR2 I8 (o_0r0[8:8], gfint_0[8:8], gfint_1[8:8]);
  OR2 I9 (o_0r0[9:9], gfint_0[9:9], gfint_1[9:9]);
  OR2 I10 (o_0r0[10:10], gfint_0[10:10], gfint_1[10:10]);
  OR2 I11 (o_0r0[11:11], gfint_0[11:11], gfint_1[11:11]);
  OR2 I12 (o_0r0[12:12], gfint_0[12:12], gfint_1[12:12]);
  OR2 I13 (o_0r0[13:13], gfint_0[13:13], gfint_1[13:13]);
  OR2 I14 (o_0r0[14:14], gfint_0[14:14], gfint_1[14:14]);
  OR2 I15 (o_0r0[15:15], gfint_0[15:15], gfint_1[15:15]);
  OR2 I16 (o_0r0[16:16], gfint_0[16:16], gfint_1[16:16]);
  OR2 I17 (o_0r0[17:17], gfint_0[17:17], gfint_1[17:17]);
  OR2 I18 (o_0r0[18:18], gfint_0[18:18], gfint_1[18:18]);
  OR2 I19 (o_0r0[19:19], gfint_0[19:19], gfint_1[19:19]);
  OR2 I20 (o_0r0[20:20], gfint_0[20:20], gfint_1[20:20]);
  OR2 I21 (o_0r0[21:21], gfint_0[21:21], gfint_1[21:21]);
  OR2 I22 (o_0r0[22:22], gfint_0[22:22], gfint_1[22:22]);
  OR2 I23 (o_0r0[23:23], gfint_0[23:23], gfint_1[23:23]);
  OR2 I24 (o_0r0[24:24], gfint_0[24:24], gfint_1[24:24]);
  OR2 I25 (o_0r0[25:25], gfint_0[25:25], gfint_1[25:25]);
  OR2 I26 (o_0r0[26:26], gfint_0[26:26], gfint_1[26:26]);
  OR2 I27 (o_0r0[27:27], gfint_0[27:27], gfint_1[27:27]);
  OR2 I28 (o_0r0[28:28], gfint_0[28:28], gfint_1[28:28]);
  OR2 I29 (o_0r0[29:29], gfint_0[29:29], gfint_1[29:29]);
  OR2 I30 (o_0r0[30:30], gfint_0[30:30], gfint_1[30:30]);
  OR2 I31 (o_0r0[31:31], gfint_0[31:31], gfint_1[31:31]);
  OR2 I32 (o_0r0[32:32], gfint_0[32:32], gfint_1[32:32]);
  OR2 I33 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0]);
  OR2 I34 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1]);
  OR2 I35 (o_0r1[2:2], gtint_0[2:2], gtint_1[2:2]);
  OR2 I36 (o_0r1[3:3], gtint_0[3:3], gtint_1[3:3]);
  OR2 I37 (o_0r1[4:4], gtint_0[4:4], gtint_1[4:4]);
  OR2 I38 (o_0r1[5:5], gtint_0[5:5], gtint_1[5:5]);
  OR2 I39 (o_0r1[6:6], gtint_0[6:6], gtint_1[6:6]);
  OR2 I40 (o_0r1[7:7], gtint_0[7:7], gtint_1[7:7]);
  OR2 I41 (o_0r1[8:8], gtint_0[8:8], gtint_1[8:8]);
  OR2 I42 (o_0r1[9:9], gtint_0[9:9], gtint_1[9:9]);
  OR2 I43 (o_0r1[10:10], gtint_0[10:10], gtint_1[10:10]);
  OR2 I44 (o_0r1[11:11], gtint_0[11:11], gtint_1[11:11]);
  OR2 I45 (o_0r1[12:12], gtint_0[12:12], gtint_1[12:12]);
  OR2 I46 (o_0r1[13:13], gtint_0[13:13], gtint_1[13:13]);
  OR2 I47 (o_0r1[14:14], gtint_0[14:14], gtint_1[14:14]);
  OR2 I48 (o_0r1[15:15], gtint_0[15:15], gtint_1[15:15]);
  OR2 I49 (o_0r1[16:16], gtint_0[16:16], gtint_1[16:16]);
  OR2 I50 (o_0r1[17:17], gtint_0[17:17], gtint_1[17:17]);
  OR2 I51 (o_0r1[18:18], gtint_0[18:18], gtint_1[18:18]);
  OR2 I52 (o_0r1[19:19], gtint_0[19:19], gtint_1[19:19]);
  OR2 I53 (o_0r1[20:20], gtint_0[20:20], gtint_1[20:20]);
  OR2 I54 (o_0r1[21:21], gtint_0[21:21], gtint_1[21:21]);
  OR2 I55 (o_0r1[22:22], gtint_0[22:22], gtint_1[22:22]);
  OR2 I56 (o_0r1[23:23], gtint_0[23:23], gtint_1[23:23]);
  OR2 I57 (o_0r1[24:24], gtint_0[24:24], gtint_1[24:24]);
  OR2 I58 (o_0r1[25:25], gtint_0[25:25], gtint_1[25:25]);
  OR2 I59 (o_0r1[26:26], gtint_0[26:26], gtint_1[26:26]);
  OR2 I60 (o_0r1[27:27], gtint_0[27:27], gtint_1[27:27]);
  OR2 I61 (o_0r1[28:28], gtint_0[28:28], gtint_1[28:28]);
  OR2 I62 (o_0r1[29:29], gtint_0[29:29], gtint_1[29:29]);
  OR2 I63 (o_0r1[30:30], gtint_0[30:30], gtint_1[30:30]);
  OR2 I64 (o_0r1[31:31], gtint_0[31:31], gtint_1[31:31]);
  OR2 I65 (o_0r1[32:32], gtint_0[32:32], gtint_1[32:32]);
  AND2 I66 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I67 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I68 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I69 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I70 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I71 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I72 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I73 (gtint_0[7:7], choice_0, i_0r1[7:7]);
  AND2 I74 (gtint_0[8:8], choice_0, i_0r1[8:8]);
  AND2 I75 (gtint_0[9:9], choice_0, i_0r1[9:9]);
  AND2 I76 (gtint_0[10:10], choice_0, i_0r1[10:10]);
  AND2 I77 (gtint_0[11:11], choice_0, i_0r1[11:11]);
  AND2 I78 (gtint_0[12:12], choice_0, i_0r1[12:12]);
  AND2 I79 (gtint_0[13:13], choice_0, i_0r1[13:13]);
  AND2 I80 (gtint_0[14:14], choice_0, i_0r1[14:14]);
  AND2 I81 (gtint_0[15:15], choice_0, i_0r1[15:15]);
  AND2 I82 (gtint_0[16:16], choice_0, i_0r1[16:16]);
  AND2 I83 (gtint_0[17:17], choice_0, i_0r1[17:17]);
  AND2 I84 (gtint_0[18:18], choice_0, i_0r1[18:18]);
  AND2 I85 (gtint_0[19:19], choice_0, i_0r1[19:19]);
  AND2 I86 (gtint_0[20:20], choice_0, i_0r1[20:20]);
  AND2 I87 (gtint_0[21:21], choice_0, i_0r1[21:21]);
  AND2 I88 (gtint_0[22:22], choice_0, i_0r1[22:22]);
  AND2 I89 (gtint_0[23:23], choice_0, i_0r1[23:23]);
  AND2 I90 (gtint_0[24:24], choice_0, i_0r1[24:24]);
  AND2 I91 (gtint_0[25:25], choice_0, i_0r1[25:25]);
  AND2 I92 (gtint_0[26:26], choice_0, i_0r1[26:26]);
  AND2 I93 (gtint_0[27:27], choice_0, i_0r1[27:27]);
  AND2 I94 (gtint_0[28:28], choice_0, i_0r1[28:28]);
  AND2 I95 (gtint_0[29:29], choice_0, i_0r1[29:29]);
  AND2 I96 (gtint_0[30:30], choice_0, i_0r1[30:30]);
  AND2 I97 (gtint_0[31:31], choice_0, i_0r1[31:31]);
  AND2 I98 (gtint_0[32:32], choice_0, i_0r1[32:32]);
  AND2 I99 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I100 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I101 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I102 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I103 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I104 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I105 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I106 (gtint_1[7:7], choice_1, i_1r1[7:7]);
  AND2 I107 (gtint_1[8:8], choice_1, i_1r1[8:8]);
  AND2 I108 (gtint_1[9:9], choice_1, i_1r1[9:9]);
  AND2 I109 (gtint_1[10:10], choice_1, i_1r1[10:10]);
  AND2 I110 (gtint_1[11:11], choice_1, i_1r1[11:11]);
  AND2 I111 (gtint_1[12:12], choice_1, i_1r1[12:12]);
  AND2 I112 (gtint_1[13:13], choice_1, i_1r1[13:13]);
  AND2 I113 (gtint_1[14:14], choice_1, i_1r1[14:14]);
  AND2 I114 (gtint_1[15:15], choice_1, i_1r1[15:15]);
  AND2 I115 (gtint_1[16:16], choice_1, i_1r1[16:16]);
  AND2 I116 (gtint_1[17:17], choice_1, i_1r1[17:17]);
  AND2 I117 (gtint_1[18:18], choice_1, i_1r1[18:18]);
  AND2 I118 (gtint_1[19:19], choice_1, i_1r1[19:19]);
  AND2 I119 (gtint_1[20:20], choice_1, i_1r1[20:20]);
  AND2 I120 (gtint_1[21:21], choice_1, i_1r1[21:21]);
  AND2 I121 (gtint_1[22:22], choice_1, i_1r1[22:22]);
  AND2 I122 (gtint_1[23:23], choice_1, i_1r1[23:23]);
  AND2 I123 (gtint_1[24:24], choice_1, i_1r1[24:24]);
  AND2 I124 (gtint_1[25:25], choice_1, i_1r1[25:25]);
  AND2 I125 (gtint_1[26:26], choice_1, i_1r1[26:26]);
  AND2 I126 (gtint_1[27:27], choice_1, i_1r1[27:27]);
  AND2 I127 (gtint_1[28:28], choice_1, i_1r1[28:28]);
  AND2 I128 (gtint_1[29:29], choice_1, i_1r1[29:29]);
  AND2 I129 (gtint_1[30:30], choice_1, i_1r1[30:30]);
  AND2 I130 (gtint_1[31:31], choice_1, i_1r1[31:31]);
  AND2 I131 (gtint_1[32:32], choice_1, i_1r1[32:32]);
  AND2 I132 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I133 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I134 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I135 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I136 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I137 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I138 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I139 (gfint_0[7:7], choice_0, i_0r0[7:7]);
  AND2 I140 (gfint_0[8:8], choice_0, i_0r0[8:8]);
  AND2 I141 (gfint_0[9:9], choice_0, i_0r0[9:9]);
  AND2 I142 (gfint_0[10:10], choice_0, i_0r0[10:10]);
  AND2 I143 (gfint_0[11:11], choice_0, i_0r0[11:11]);
  AND2 I144 (gfint_0[12:12], choice_0, i_0r0[12:12]);
  AND2 I145 (gfint_0[13:13], choice_0, i_0r0[13:13]);
  AND2 I146 (gfint_0[14:14], choice_0, i_0r0[14:14]);
  AND2 I147 (gfint_0[15:15], choice_0, i_0r0[15:15]);
  AND2 I148 (gfint_0[16:16], choice_0, i_0r0[16:16]);
  AND2 I149 (gfint_0[17:17], choice_0, i_0r0[17:17]);
  AND2 I150 (gfint_0[18:18], choice_0, i_0r0[18:18]);
  AND2 I151 (gfint_0[19:19], choice_0, i_0r0[19:19]);
  AND2 I152 (gfint_0[20:20], choice_0, i_0r0[20:20]);
  AND2 I153 (gfint_0[21:21], choice_0, i_0r0[21:21]);
  AND2 I154 (gfint_0[22:22], choice_0, i_0r0[22:22]);
  AND2 I155 (gfint_0[23:23], choice_0, i_0r0[23:23]);
  AND2 I156 (gfint_0[24:24], choice_0, i_0r0[24:24]);
  AND2 I157 (gfint_0[25:25], choice_0, i_0r0[25:25]);
  AND2 I158 (gfint_0[26:26], choice_0, i_0r0[26:26]);
  AND2 I159 (gfint_0[27:27], choice_0, i_0r0[27:27]);
  AND2 I160 (gfint_0[28:28], choice_0, i_0r0[28:28]);
  AND2 I161 (gfint_0[29:29], choice_0, i_0r0[29:29]);
  AND2 I162 (gfint_0[30:30], choice_0, i_0r0[30:30]);
  AND2 I163 (gfint_0[31:31], choice_0, i_0r0[31:31]);
  AND2 I164 (gfint_0[32:32], choice_0, i_0r0[32:32]);
  AND2 I165 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I166 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I167 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I168 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I169 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I170 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I171 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I172 (gfint_1[7:7], choice_1, i_1r0[7:7]);
  AND2 I173 (gfint_1[8:8], choice_1, i_1r0[8:8]);
  AND2 I174 (gfint_1[9:9], choice_1, i_1r0[9:9]);
  AND2 I175 (gfint_1[10:10], choice_1, i_1r0[10:10]);
  AND2 I176 (gfint_1[11:11], choice_1, i_1r0[11:11]);
  AND2 I177 (gfint_1[12:12], choice_1, i_1r0[12:12]);
  AND2 I178 (gfint_1[13:13], choice_1, i_1r0[13:13]);
  AND2 I179 (gfint_1[14:14], choice_1, i_1r0[14:14]);
  AND2 I180 (gfint_1[15:15], choice_1, i_1r0[15:15]);
  AND2 I181 (gfint_1[16:16], choice_1, i_1r0[16:16]);
  AND2 I182 (gfint_1[17:17], choice_1, i_1r0[17:17]);
  AND2 I183 (gfint_1[18:18], choice_1, i_1r0[18:18]);
  AND2 I184 (gfint_1[19:19], choice_1, i_1r0[19:19]);
  AND2 I185 (gfint_1[20:20], choice_1, i_1r0[20:20]);
  AND2 I186 (gfint_1[21:21], choice_1, i_1r0[21:21]);
  AND2 I187 (gfint_1[22:22], choice_1, i_1r0[22:22]);
  AND2 I188 (gfint_1[23:23], choice_1, i_1r0[23:23]);
  AND2 I189 (gfint_1[24:24], choice_1, i_1r0[24:24]);
  AND2 I190 (gfint_1[25:25], choice_1, i_1r0[25:25]);
  AND2 I191 (gfint_1[26:26], choice_1, i_1r0[26:26]);
  AND2 I192 (gfint_1[27:27], choice_1, i_1r0[27:27]);
  AND2 I193 (gfint_1[28:28], choice_1, i_1r0[28:28]);
  AND2 I194 (gfint_1[29:29], choice_1, i_1r0[29:29]);
  AND2 I195 (gfint_1[30:30], choice_1, i_1r0[30:30]);
  AND2 I196 (gfint_1[31:31], choice_1, i_1r0[31:31]);
  AND2 I197 (gfint_1[32:32], choice_1, i_1r0[32:32]);
  OR2 I198 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I199 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I200 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I201 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I202 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I203 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I204 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I205 (comp0_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I206 (comp0_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I207 (comp0_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I208 (comp0_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I209 (comp0_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I210 (comp0_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I211 (comp0_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I212 (comp0_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I213 (comp0_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I214 (comp0_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I215 (comp0_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I216 (comp0_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I217 (comp0_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I218 (comp0_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I219 (comp0_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I220 (comp0_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I221 (comp0_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I222 (comp0_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I223 (comp0_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I224 (comp0_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I225 (comp0_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I226 (comp0_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I227 (comp0_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I228 (comp0_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I229 (comp0_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I230 (comp0_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  C3 I231 (simp2421_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I232 (simp2421_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I233 (simp2421_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I234 (simp2421_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I235 (simp2421_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I236 (simp2421_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I237 (simp2421_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I238 (simp2421_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I239 (simp2421_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I240 (simp2421_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C3 I241 (simp2421_0[10:10], comp0_0[30:30], comp0_0[31:31], comp0_0[32:32]);
  C3 I242 (simp2422_0[0:0], simp2421_0[0:0], simp2421_0[1:1], simp2421_0[2:2]);
  C3 I243 (simp2422_0[1:1], simp2421_0[3:3], simp2421_0[4:4], simp2421_0[5:5]);
  C3 I244 (simp2422_0[2:2], simp2421_0[6:6], simp2421_0[7:7], simp2421_0[8:8]);
  C2 I245 (simp2422_0[3:3], simp2421_0[9:9], simp2421_0[10:10]);
  C3 I246 (simp2423_0[0:0], simp2422_0[0:0], simp2422_0[1:1], simp2422_0[2:2]);
  BUFF I247 (simp2423_0[1:1], simp2422_0[3:3]);
  C2 I248 (icomp_0, simp2423_0[0:0], simp2423_0[1:1]);
  OR2 I249 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I250 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I251 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I252 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I253 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I254 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I255 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  OR2 I256 (comp1_0[7:7], i_1r0[7:7], i_1r1[7:7]);
  OR2 I257 (comp1_0[8:8], i_1r0[8:8], i_1r1[8:8]);
  OR2 I258 (comp1_0[9:9], i_1r0[9:9], i_1r1[9:9]);
  OR2 I259 (comp1_0[10:10], i_1r0[10:10], i_1r1[10:10]);
  OR2 I260 (comp1_0[11:11], i_1r0[11:11], i_1r1[11:11]);
  OR2 I261 (comp1_0[12:12], i_1r0[12:12], i_1r1[12:12]);
  OR2 I262 (comp1_0[13:13], i_1r0[13:13], i_1r1[13:13]);
  OR2 I263 (comp1_0[14:14], i_1r0[14:14], i_1r1[14:14]);
  OR2 I264 (comp1_0[15:15], i_1r0[15:15], i_1r1[15:15]);
  OR2 I265 (comp1_0[16:16], i_1r0[16:16], i_1r1[16:16]);
  OR2 I266 (comp1_0[17:17], i_1r0[17:17], i_1r1[17:17]);
  OR2 I267 (comp1_0[18:18], i_1r0[18:18], i_1r1[18:18]);
  OR2 I268 (comp1_0[19:19], i_1r0[19:19], i_1r1[19:19]);
  OR2 I269 (comp1_0[20:20], i_1r0[20:20], i_1r1[20:20]);
  OR2 I270 (comp1_0[21:21], i_1r0[21:21], i_1r1[21:21]);
  OR2 I271 (comp1_0[22:22], i_1r0[22:22], i_1r1[22:22]);
  OR2 I272 (comp1_0[23:23], i_1r0[23:23], i_1r1[23:23]);
  OR2 I273 (comp1_0[24:24], i_1r0[24:24], i_1r1[24:24]);
  OR2 I274 (comp1_0[25:25], i_1r0[25:25], i_1r1[25:25]);
  OR2 I275 (comp1_0[26:26], i_1r0[26:26], i_1r1[26:26]);
  OR2 I276 (comp1_0[27:27], i_1r0[27:27], i_1r1[27:27]);
  OR2 I277 (comp1_0[28:28], i_1r0[28:28], i_1r1[28:28]);
  OR2 I278 (comp1_0[29:29], i_1r0[29:29], i_1r1[29:29]);
  OR2 I279 (comp1_0[30:30], i_1r0[30:30], i_1r1[30:30]);
  OR2 I280 (comp1_0[31:31], i_1r0[31:31], i_1r1[31:31]);
  OR2 I281 (comp1_0[32:32], i_1r0[32:32], i_1r1[32:32]);
  C3 I282 (simp2771_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I283 (simp2771_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  C3 I284 (simp2771_0[2:2], comp1_0[6:6], comp1_0[7:7], comp1_0[8:8]);
  C3 I285 (simp2771_0[3:3], comp1_0[9:9], comp1_0[10:10], comp1_0[11:11]);
  C3 I286 (simp2771_0[4:4], comp1_0[12:12], comp1_0[13:13], comp1_0[14:14]);
  C3 I287 (simp2771_0[5:5], comp1_0[15:15], comp1_0[16:16], comp1_0[17:17]);
  C3 I288 (simp2771_0[6:6], comp1_0[18:18], comp1_0[19:19], comp1_0[20:20]);
  C3 I289 (simp2771_0[7:7], comp1_0[21:21], comp1_0[22:22], comp1_0[23:23]);
  C3 I290 (simp2771_0[8:8], comp1_0[24:24], comp1_0[25:25], comp1_0[26:26]);
  C3 I291 (simp2771_0[9:9], comp1_0[27:27], comp1_0[28:28], comp1_0[29:29]);
  C3 I292 (simp2771_0[10:10], comp1_0[30:30], comp1_0[31:31], comp1_0[32:32]);
  C3 I293 (simp2772_0[0:0], simp2771_0[0:0], simp2771_0[1:1], simp2771_0[2:2]);
  C3 I294 (simp2772_0[1:1], simp2771_0[3:3], simp2771_0[4:4], simp2771_0[5:5]);
  C3 I295 (simp2772_0[2:2], simp2771_0[6:6], simp2771_0[7:7], simp2771_0[8:8]);
  C2 I296 (simp2772_0[3:3], simp2771_0[9:9], simp2771_0[10:10]);
  C3 I297 (simp2773_0[0:0], simp2772_0[0:0], simp2772_0[1:1], simp2772_0[2:2]);
  BUFF I298 (simp2773_0[1:1], simp2772_0[3:3]);
  C2 I299 (icomp_1, simp2773_0[0:0], simp2773_0[1:1]);
  C2R I300 (choice_0, icomp_0, nchosen_0, reset);
  C2R I301 (choice_1, icomp_1, nchosen_0, reset);
  OR2 I302 (anychoice_0, choice_0, choice_1);
  NOR2 I303 (nchosen_0, anychoice_0, o_0a);
  C2R I304 (i_0a, choice_0, o_0a, reset);
  C2R I305 (i_1a, choice_1, o_0a, reset);
endmodule

// tko4m1_1nm1b1_2nm1b0_3mx2o3o10_4o11_i0w4bt1o0w1bt2o0w1b TeakO [
//     (1,TeakOConstant 1 1),
//     (2,TeakOConstant 1 0),
//     (3,TeakOMux [[Imp 2 0,Imp 3 0,Imp 10 0],[Imp 4 0,Imp 11 0]] [(0,0,4),(1,0,1),(2,0,1)])] [One 4,One
//    1]
module tko4m1_1nm1b1_2nm1b0_3mx2o3o10_4o11_i0w4bt1o0w1bt2o0w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [3:0] gocomp_0;
  wire [1:0] simp61_0;
  wire termf_1;
  wire termf_2;
  wire termt_1;
  wire termt_2;
  wire gfint3_0;
  wire gfint3_1;
  wire gtint3_0;
  wire gtint3_1;
  wire selcomp3_0;
  wire selcomp3_1;
  wire sel3_0;
  wire sel3_1;
  wire selg3_0;
  wire selg3_1;
  wire icomplete3_0;
  wire scomplete3_0;
  wire comp30_0;
  wire comp31_0;
  wire [3:0] dcomp3_0;
  wire [1:0] simp401_0;
  wire [2:0] match30_0;
  wire [1:0] simp521_0;
  wire [1:0] simp531_0;
  wire [1:0] simp541_0;
  wire [1:0] match31_0;
  wire [1:0] simp571_0;
  wire [1:0] simp581_0;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  C3 I4 (simp61_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  BUFF I5 (simp61_0[1:1], gocomp_0[3:3]);
  C2 I6 (go_0, simp61_0[0:0], simp61_0[1:1]);
  BUFF I7 (termt_1, go_0);
  GND I8 (termf_1);
  BUFF I9 (termf_2, go_0);
  GND I10 (termt_2);
  OR2 I11 (comp30_0, termf_1, termt_1);
  BUFF I12 (selcomp3_0, comp30_0);
  OR2 I13 (comp31_0, termf_2, termt_2);
  BUFF I14 (selcomp3_1, comp31_0);
  OR2 I15 (dcomp3_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I16 (dcomp3_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I17 (dcomp3_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I18 (dcomp3_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  C3 I19 (simp401_0[0:0], dcomp3_0[0:0], dcomp3_0[1:1], dcomp3_0[2:2]);
  BUFF I20 (simp401_0[1:1], dcomp3_0[3:3]);
  C2 I21 (scomplete3_0, simp401_0[0:0], simp401_0[1:1]);
  C3 I22 (icomplete3_0, scomplete3_0, selcomp3_0, selcomp3_1);
  OR2 I23 (o_0r0, gfint3_0, gfint3_1);
  OR2 I24 (o_0r1, gtint3_0, gtint3_1);
  C2R I25 (sel3_0, selg3_0, icomplete3_0, reset);
  C2R I26 (sel3_1, selg3_1, icomplete3_0, reset);
  C2R I27 (gfint3_0, sel3_0, termf_1, reset);
  C2R I28 (gfint3_1, sel3_1, termf_2, reset);
  C2R I29 (gtint3_0, sel3_0, termt_1, reset);
  C2R I30 (gtint3_1, sel3_1, termt_2, reset);
  OR3 I31 (selg3_0, match30_0[0:0], match30_0[1:1], match30_0[2:2]);
  C3 I32 (simp521_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I33 (simp521_0[1:1], i_0r0[3:3]);
  C2 I34 (match30_0[0:0], simp521_0[0:0], simp521_0[1:1]);
  C3 I35 (simp531_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I36 (simp531_0[1:1], i_0r0[3:3]);
  C2 I37 (match30_0[1:1], simp531_0[0:0], simp531_0[1:1]);
  C3 I38 (simp541_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I39 (simp541_0[1:1], i_0r1[3:3]);
  C2 I40 (match30_0[2:2], simp541_0[0:0], simp541_0[1:1]);
  OR2 I41 (selg3_1, match31_0[0:0], match31_0[1:1]);
  C3 I42 (simp571_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I43 (simp571_0[1:1], i_0r0[3:3]);
  C2 I44 (match31_0[0:0], simp571_0[0:0], simp571_0[1:1]);
  C3 I45 (simp581_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I46 (simp581_0[1:1], i_0r1[3:3]);
  C2 I47 (match31_0[1:1], simp581_0[0:0], simp581_0[1:1]);
  BUFF I48 (i_0a, o_0a);
endmodule

// tko66m33_1nm1b0_2api0w33bt1o0w1b_3nm1b0_4api33w33bt3o0w1b_5addt2o0w34bt4o0w34b_6apt5o1w33b TeakO [
//     (1,TeakOConstant 1 0),
//     (2,TeakOAppend 1 [(0,0,33),(1,0,1)]),
//     (3,TeakOConstant 1 0),
//     (4,TeakOAppend 1 [(0,33,33),(3,0,1)]),
//     (5,TeakOp TeakOpAdd [(2,0,34),(4,0,34)]),
//     (6,TeakOAppend 1 [(5,1,33)])] [One 66,One 33]
module tko66m33_1nm1b0_2api0w33bt1o0w1b_3nm1b0_4api33w33bt3o0w1b_5addt2o0w34bt4o0w34b_6apt5o1w33b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [65:0] i_0r0;
  input [65:0] i_0r1;
  output i_0a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [65:0] gocomp_0;
  wire [21:0] simp681_0;
  wire [7:0] simp682_0;
  wire [2:0] simp683_0;
  wire termf_1;
  wire [33:0] termf_2;
  wire termf_3;
  wire [33:0] termf_4;
  wire [33:0] termf_5;
  wire termt_1;
  wire [33:0] termt_2;
  wire termt_3;
  wire [33:0] termt_4;
  wire [33:0] termt_5;
  wire [33:0] cf5__0;
  wire [33:0] ct5__0;
  wire [3:0] ha5__0;
  wire [7:0] fa5_1min_0;
  wire [1:0] simp2411_0;
  wire [1:0] simp2421_0;
  wire [7:0] fa5_2min_0;
  wire [1:0] simp2541_0;
  wire [1:0] simp2551_0;
  wire [7:0] fa5_3min_0;
  wire [1:0] simp2671_0;
  wire [1:0] simp2681_0;
  wire [7:0] fa5_4min_0;
  wire [1:0] simp2801_0;
  wire [1:0] simp2811_0;
  wire [7:0] fa5_5min_0;
  wire [1:0] simp2931_0;
  wire [1:0] simp2941_0;
  wire [7:0] fa5_6min_0;
  wire [1:0] simp3061_0;
  wire [1:0] simp3071_0;
  wire [7:0] fa5_7min_0;
  wire [1:0] simp3191_0;
  wire [1:0] simp3201_0;
  wire [7:0] fa5_8min_0;
  wire [1:0] simp3321_0;
  wire [1:0] simp3331_0;
  wire [7:0] fa5_9min_0;
  wire [1:0] simp3451_0;
  wire [1:0] simp3461_0;
  wire [7:0] fa5_10min_0;
  wire [1:0] simp3581_0;
  wire [1:0] simp3591_0;
  wire [7:0] fa5_11min_0;
  wire [1:0] simp3711_0;
  wire [1:0] simp3721_0;
  wire [7:0] fa5_12min_0;
  wire [1:0] simp3841_0;
  wire [1:0] simp3851_0;
  wire [7:0] fa5_13min_0;
  wire [1:0] simp3971_0;
  wire [1:0] simp3981_0;
  wire [7:0] fa5_14min_0;
  wire [1:0] simp4101_0;
  wire [1:0] simp4111_0;
  wire [7:0] fa5_15min_0;
  wire [1:0] simp4231_0;
  wire [1:0] simp4241_0;
  wire [7:0] fa5_16min_0;
  wire [1:0] simp4361_0;
  wire [1:0] simp4371_0;
  wire [7:0] fa5_17min_0;
  wire [1:0] simp4491_0;
  wire [1:0] simp4501_0;
  wire [7:0] fa5_18min_0;
  wire [1:0] simp4621_0;
  wire [1:0] simp4631_0;
  wire [7:0] fa5_19min_0;
  wire [1:0] simp4751_0;
  wire [1:0] simp4761_0;
  wire [7:0] fa5_20min_0;
  wire [1:0] simp4881_0;
  wire [1:0] simp4891_0;
  wire [7:0] fa5_21min_0;
  wire [1:0] simp5011_0;
  wire [1:0] simp5021_0;
  wire [7:0] fa5_22min_0;
  wire [1:0] simp5141_0;
  wire [1:0] simp5151_0;
  wire [7:0] fa5_23min_0;
  wire [1:0] simp5271_0;
  wire [1:0] simp5281_0;
  wire [7:0] fa5_24min_0;
  wire [1:0] simp5401_0;
  wire [1:0] simp5411_0;
  wire [7:0] fa5_25min_0;
  wire [1:0] simp5531_0;
  wire [1:0] simp5541_0;
  wire [7:0] fa5_26min_0;
  wire [1:0] simp5661_0;
  wire [1:0] simp5671_0;
  wire [7:0] fa5_27min_0;
  wire [1:0] simp5791_0;
  wire [1:0] simp5801_0;
  wire [7:0] fa5_28min_0;
  wire [1:0] simp5921_0;
  wire [1:0] simp5931_0;
  wire [7:0] fa5_29min_0;
  wire [1:0] simp6051_0;
  wire [1:0] simp6061_0;
  wire [7:0] fa5_30min_0;
  wire [1:0] simp6181_0;
  wire [1:0] simp6191_0;
  wire [7:0] fa5_31min_0;
  wire [1:0] simp6311_0;
  wire [1:0] simp6321_0;
  wire [7:0] fa5_32min_0;
  wire [1:0] simp6441_0;
  wire [1:0] simp6451_0;
  wire [7:0] fa5_33min_0;
  wire [1:0] simp6571_0;
  wire [1:0] simp6581_0;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I30 (gocomp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I31 (gocomp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I32 (gocomp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  OR2 I33 (gocomp_0[33:33], i_0r0[33:33], i_0r1[33:33]);
  OR2 I34 (gocomp_0[34:34], i_0r0[34:34], i_0r1[34:34]);
  OR2 I35 (gocomp_0[35:35], i_0r0[35:35], i_0r1[35:35]);
  OR2 I36 (gocomp_0[36:36], i_0r0[36:36], i_0r1[36:36]);
  OR2 I37 (gocomp_0[37:37], i_0r0[37:37], i_0r1[37:37]);
  OR2 I38 (gocomp_0[38:38], i_0r0[38:38], i_0r1[38:38]);
  OR2 I39 (gocomp_0[39:39], i_0r0[39:39], i_0r1[39:39]);
  OR2 I40 (gocomp_0[40:40], i_0r0[40:40], i_0r1[40:40]);
  OR2 I41 (gocomp_0[41:41], i_0r0[41:41], i_0r1[41:41]);
  OR2 I42 (gocomp_0[42:42], i_0r0[42:42], i_0r1[42:42]);
  OR2 I43 (gocomp_0[43:43], i_0r0[43:43], i_0r1[43:43]);
  OR2 I44 (gocomp_0[44:44], i_0r0[44:44], i_0r1[44:44]);
  OR2 I45 (gocomp_0[45:45], i_0r0[45:45], i_0r1[45:45]);
  OR2 I46 (gocomp_0[46:46], i_0r0[46:46], i_0r1[46:46]);
  OR2 I47 (gocomp_0[47:47], i_0r0[47:47], i_0r1[47:47]);
  OR2 I48 (gocomp_0[48:48], i_0r0[48:48], i_0r1[48:48]);
  OR2 I49 (gocomp_0[49:49], i_0r0[49:49], i_0r1[49:49]);
  OR2 I50 (gocomp_0[50:50], i_0r0[50:50], i_0r1[50:50]);
  OR2 I51 (gocomp_0[51:51], i_0r0[51:51], i_0r1[51:51]);
  OR2 I52 (gocomp_0[52:52], i_0r0[52:52], i_0r1[52:52]);
  OR2 I53 (gocomp_0[53:53], i_0r0[53:53], i_0r1[53:53]);
  OR2 I54 (gocomp_0[54:54], i_0r0[54:54], i_0r1[54:54]);
  OR2 I55 (gocomp_0[55:55], i_0r0[55:55], i_0r1[55:55]);
  OR2 I56 (gocomp_0[56:56], i_0r0[56:56], i_0r1[56:56]);
  OR2 I57 (gocomp_0[57:57], i_0r0[57:57], i_0r1[57:57]);
  OR2 I58 (gocomp_0[58:58], i_0r0[58:58], i_0r1[58:58]);
  OR2 I59 (gocomp_0[59:59], i_0r0[59:59], i_0r1[59:59]);
  OR2 I60 (gocomp_0[60:60], i_0r0[60:60], i_0r1[60:60]);
  OR2 I61 (gocomp_0[61:61], i_0r0[61:61], i_0r1[61:61]);
  OR2 I62 (gocomp_0[62:62], i_0r0[62:62], i_0r1[62:62]);
  OR2 I63 (gocomp_0[63:63], i_0r0[63:63], i_0r1[63:63]);
  OR2 I64 (gocomp_0[64:64], i_0r0[64:64], i_0r1[64:64]);
  OR2 I65 (gocomp_0[65:65], i_0r0[65:65], i_0r1[65:65]);
  C3 I66 (simp681_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  C3 I67 (simp681_0[1:1], gocomp_0[3:3], gocomp_0[4:4], gocomp_0[5:5]);
  C3 I68 (simp681_0[2:2], gocomp_0[6:6], gocomp_0[7:7], gocomp_0[8:8]);
  C3 I69 (simp681_0[3:3], gocomp_0[9:9], gocomp_0[10:10], gocomp_0[11:11]);
  C3 I70 (simp681_0[4:4], gocomp_0[12:12], gocomp_0[13:13], gocomp_0[14:14]);
  C3 I71 (simp681_0[5:5], gocomp_0[15:15], gocomp_0[16:16], gocomp_0[17:17]);
  C3 I72 (simp681_0[6:6], gocomp_0[18:18], gocomp_0[19:19], gocomp_0[20:20]);
  C3 I73 (simp681_0[7:7], gocomp_0[21:21], gocomp_0[22:22], gocomp_0[23:23]);
  C3 I74 (simp681_0[8:8], gocomp_0[24:24], gocomp_0[25:25], gocomp_0[26:26]);
  C3 I75 (simp681_0[9:9], gocomp_0[27:27], gocomp_0[28:28], gocomp_0[29:29]);
  C3 I76 (simp681_0[10:10], gocomp_0[30:30], gocomp_0[31:31], gocomp_0[32:32]);
  C3 I77 (simp681_0[11:11], gocomp_0[33:33], gocomp_0[34:34], gocomp_0[35:35]);
  C3 I78 (simp681_0[12:12], gocomp_0[36:36], gocomp_0[37:37], gocomp_0[38:38]);
  C3 I79 (simp681_0[13:13], gocomp_0[39:39], gocomp_0[40:40], gocomp_0[41:41]);
  C3 I80 (simp681_0[14:14], gocomp_0[42:42], gocomp_0[43:43], gocomp_0[44:44]);
  C3 I81 (simp681_0[15:15], gocomp_0[45:45], gocomp_0[46:46], gocomp_0[47:47]);
  C3 I82 (simp681_0[16:16], gocomp_0[48:48], gocomp_0[49:49], gocomp_0[50:50]);
  C3 I83 (simp681_0[17:17], gocomp_0[51:51], gocomp_0[52:52], gocomp_0[53:53]);
  C3 I84 (simp681_0[18:18], gocomp_0[54:54], gocomp_0[55:55], gocomp_0[56:56]);
  C3 I85 (simp681_0[19:19], gocomp_0[57:57], gocomp_0[58:58], gocomp_0[59:59]);
  C3 I86 (simp681_0[20:20], gocomp_0[60:60], gocomp_0[61:61], gocomp_0[62:62]);
  C3 I87 (simp681_0[21:21], gocomp_0[63:63], gocomp_0[64:64], gocomp_0[65:65]);
  C3 I88 (simp682_0[0:0], simp681_0[0:0], simp681_0[1:1], simp681_0[2:2]);
  C3 I89 (simp682_0[1:1], simp681_0[3:3], simp681_0[4:4], simp681_0[5:5]);
  C3 I90 (simp682_0[2:2], simp681_0[6:6], simp681_0[7:7], simp681_0[8:8]);
  C3 I91 (simp682_0[3:3], simp681_0[9:9], simp681_0[10:10], simp681_0[11:11]);
  C3 I92 (simp682_0[4:4], simp681_0[12:12], simp681_0[13:13], simp681_0[14:14]);
  C3 I93 (simp682_0[5:5], simp681_0[15:15], simp681_0[16:16], simp681_0[17:17]);
  C3 I94 (simp682_0[6:6], simp681_0[18:18], simp681_0[19:19], simp681_0[20:20]);
  BUFF I95 (simp682_0[7:7], simp681_0[21:21]);
  C3 I96 (simp683_0[0:0], simp682_0[0:0], simp682_0[1:1], simp682_0[2:2]);
  C3 I97 (simp683_0[1:1], simp682_0[3:3], simp682_0[4:4], simp682_0[5:5]);
  C2 I98 (simp683_0[2:2], simp682_0[6:6], simp682_0[7:7]);
  C3 I99 (go_0, simp683_0[0:0], simp683_0[1:1], simp683_0[2:2]);
  BUFF I100 (termf_1, go_0);
  GND I101 (termt_1);
  BUFF I102 (termf_2[0:0], i_0r0[0:0]);
  BUFF I103 (termf_2[1:1], i_0r0[1:1]);
  BUFF I104 (termf_2[2:2], i_0r0[2:2]);
  BUFF I105 (termf_2[3:3], i_0r0[3:3]);
  BUFF I106 (termf_2[4:4], i_0r0[4:4]);
  BUFF I107 (termf_2[5:5], i_0r0[5:5]);
  BUFF I108 (termf_2[6:6], i_0r0[6:6]);
  BUFF I109 (termf_2[7:7], i_0r0[7:7]);
  BUFF I110 (termf_2[8:8], i_0r0[8:8]);
  BUFF I111 (termf_2[9:9], i_0r0[9:9]);
  BUFF I112 (termf_2[10:10], i_0r0[10:10]);
  BUFF I113 (termf_2[11:11], i_0r0[11:11]);
  BUFF I114 (termf_2[12:12], i_0r0[12:12]);
  BUFF I115 (termf_2[13:13], i_0r0[13:13]);
  BUFF I116 (termf_2[14:14], i_0r0[14:14]);
  BUFF I117 (termf_2[15:15], i_0r0[15:15]);
  BUFF I118 (termf_2[16:16], i_0r0[16:16]);
  BUFF I119 (termf_2[17:17], i_0r0[17:17]);
  BUFF I120 (termf_2[18:18], i_0r0[18:18]);
  BUFF I121 (termf_2[19:19], i_0r0[19:19]);
  BUFF I122 (termf_2[20:20], i_0r0[20:20]);
  BUFF I123 (termf_2[21:21], i_0r0[21:21]);
  BUFF I124 (termf_2[22:22], i_0r0[22:22]);
  BUFF I125 (termf_2[23:23], i_0r0[23:23]);
  BUFF I126 (termf_2[24:24], i_0r0[24:24]);
  BUFF I127 (termf_2[25:25], i_0r0[25:25]);
  BUFF I128 (termf_2[26:26], i_0r0[26:26]);
  BUFF I129 (termf_2[27:27], i_0r0[27:27]);
  BUFF I130 (termf_2[28:28], i_0r0[28:28]);
  BUFF I131 (termf_2[29:29], i_0r0[29:29]);
  BUFF I132 (termf_2[30:30], i_0r0[30:30]);
  BUFF I133 (termf_2[31:31], i_0r0[31:31]);
  BUFF I134 (termf_2[32:32], i_0r0[32:32]);
  BUFF I135 (termf_2[33:33], termf_1);
  BUFF I136 (termt_2[0:0], i_0r1[0:0]);
  BUFF I137 (termt_2[1:1], i_0r1[1:1]);
  BUFF I138 (termt_2[2:2], i_0r1[2:2]);
  BUFF I139 (termt_2[3:3], i_0r1[3:3]);
  BUFF I140 (termt_2[4:4], i_0r1[4:4]);
  BUFF I141 (termt_2[5:5], i_0r1[5:5]);
  BUFF I142 (termt_2[6:6], i_0r1[6:6]);
  BUFF I143 (termt_2[7:7], i_0r1[7:7]);
  BUFF I144 (termt_2[8:8], i_0r1[8:8]);
  BUFF I145 (termt_2[9:9], i_0r1[9:9]);
  BUFF I146 (termt_2[10:10], i_0r1[10:10]);
  BUFF I147 (termt_2[11:11], i_0r1[11:11]);
  BUFF I148 (termt_2[12:12], i_0r1[12:12]);
  BUFF I149 (termt_2[13:13], i_0r1[13:13]);
  BUFF I150 (termt_2[14:14], i_0r1[14:14]);
  BUFF I151 (termt_2[15:15], i_0r1[15:15]);
  BUFF I152 (termt_2[16:16], i_0r1[16:16]);
  BUFF I153 (termt_2[17:17], i_0r1[17:17]);
  BUFF I154 (termt_2[18:18], i_0r1[18:18]);
  BUFF I155 (termt_2[19:19], i_0r1[19:19]);
  BUFF I156 (termt_2[20:20], i_0r1[20:20]);
  BUFF I157 (termt_2[21:21], i_0r1[21:21]);
  BUFF I158 (termt_2[22:22], i_0r1[22:22]);
  BUFF I159 (termt_2[23:23], i_0r1[23:23]);
  BUFF I160 (termt_2[24:24], i_0r1[24:24]);
  BUFF I161 (termt_2[25:25], i_0r1[25:25]);
  BUFF I162 (termt_2[26:26], i_0r1[26:26]);
  BUFF I163 (termt_2[27:27], i_0r1[27:27]);
  BUFF I164 (termt_2[28:28], i_0r1[28:28]);
  BUFF I165 (termt_2[29:29], i_0r1[29:29]);
  BUFF I166 (termt_2[30:30], i_0r1[30:30]);
  BUFF I167 (termt_2[31:31], i_0r1[31:31]);
  BUFF I168 (termt_2[32:32], i_0r1[32:32]);
  BUFF I169 (termt_2[33:33], termt_1);
  BUFF I170 (termf_3, go_0);
  GND I171 (termt_3);
  BUFF I172 (termf_4[0:0], i_0r0[33:33]);
  BUFF I173 (termf_4[1:1], i_0r0[34:34]);
  BUFF I174 (termf_4[2:2], i_0r0[35:35]);
  BUFF I175 (termf_4[3:3], i_0r0[36:36]);
  BUFF I176 (termf_4[4:4], i_0r0[37:37]);
  BUFF I177 (termf_4[5:5], i_0r0[38:38]);
  BUFF I178 (termf_4[6:6], i_0r0[39:39]);
  BUFF I179 (termf_4[7:7], i_0r0[40:40]);
  BUFF I180 (termf_4[8:8], i_0r0[41:41]);
  BUFF I181 (termf_4[9:9], i_0r0[42:42]);
  BUFF I182 (termf_4[10:10], i_0r0[43:43]);
  BUFF I183 (termf_4[11:11], i_0r0[44:44]);
  BUFF I184 (termf_4[12:12], i_0r0[45:45]);
  BUFF I185 (termf_4[13:13], i_0r0[46:46]);
  BUFF I186 (termf_4[14:14], i_0r0[47:47]);
  BUFF I187 (termf_4[15:15], i_0r0[48:48]);
  BUFF I188 (termf_4[16:16], i_0r0[49:49]);
  BUFF I189 (termf_4[17:17], i_0r0[50:50]);
  BUFF I190 (termf_4[18:18], i_0r0[51:51]);
  BUFF I191 (termf_4[19:19], i_0r0[52:52]);
  BUFF I192 (termf_4[20:20], i_0r0[53:53]);
  BUFF I193 (termf_4[21:21], i_0r0[54:54]);
  BUFF I194 (termf_4[22:22], i_0r0[55:55]);
  BUFF I195 (termf_4[23:23], i_0r0[56:56]);
  BUFF I196 (termf_4[24:24], i_0r0[57:57]);
  BUFF I197 (termf_4[25:25], i_0r0[58:58]);
  BUFF I198 (termf_4[26:26], i_0r0[59:59]);
  BUFF I199 (termf_4[27:27], i_0r0[60:60]);
  BUFF I200 (termf_4[28:28], i_0r0[61:61]);
  BUFF I201 (termf_4[29:29], i_0r0[62:62]);
  BUFF I202 (termf_4[30:30], i_0r0[63:63]);
  BUFF I203 (termf_4[31:31], i_0r0[64:64]);
  BUFF I204 (termf_4[32:32], i_0r0[65:65]);
  BUFF I205 (termf_4[33:33], termf_3);
  BUFF I206 (termt_4[0:0], i_0r1[33:33]);
  BUFF I207 (termt_4[1:1], i_0r1[34:34]);
  BUFF I208 (termt_4[2:2], i_0r1[35:35]);
  BUFF I209 (termt_4[3:3], i_0r1[36:36]);
  BUFF I210 (termt_4[4:4], i_0r1[37:37]);
  BUFF I211 (termt_4[5:5], i_0r1[38:38]);
  BUFF I212 (termt_4[6:6], i_0r1[39:39]);
  BUFF I213 (termt_4[7:7], i_0r1[40:40]);
  BUFF I214 (termt_4[8:8], i_0r1[41:41]);
  BUFF I215 (termt_4[9:9], i_0r1[42:42]);
  BUFF I216 (termt_4[10:10], i_0r1[43:43]);
  BUFF I217 (termt_4[11:11], i_0r1[44:44]);
  BUFF I218 (termt_4[12:12], i_0r1[45:45]);
  BUFF I219 (termt_4[13:13], i_0r1[46:46]);
  BUFF I220 (termt_4[14:14], i_0r1[47:47]);
  BUFF I221 (termt_4[15:15], i_0r1[48:48]);
  BUFF I222 (termt_4[16:16], i_0r1[49:49]);
  BUFF I223 (termt_4[17:17], i_0r1[50:50]);
  BUFF I224 (termt_4[18:18], i_0r1[51:51]);
  BUFF I225 (termt_4[19:19], i_0r1[52:52]);
  BUFF I226 (termt_4[20:20], i_0r1[53:53]);
  BUFF I227 (termt_4[21:21], i_0r1[54:54]);
  BUFF I228 (termt_4[22:22], i_0r1[55:55]);
  BUFF I229 (termt_4[23:23], i_0r1[56:56]);
  BUFF I230 (termt_4[24:24], i_0r1[57:57]);
  BUFF I231 (termt_4[25:25], i_0r1[58:58]);
  BUFF I232 (termt_4[26:26], i_0r1[59:59]);
  BUFF I233 (termt_4[27:27], i_0r1[60:60]);
  BUFF I234 (termt_4[28:28], i_0r1[61:61]);
  BUFF I235 (termt_4[29:29], i_0r1[62:62]);
  BUFF I236 (termt_4[30:30], i_0r1[63:63]);
  BUFF I237 (termt_4[31:31], i_0r1[64:64]);
  BUFF I238 (termt_4[32:32], i_0r1[65:65]);
  BUFF I239 (termt_4[33:33], termt_3);
  C2 I240 (ha5__0[0:0], termf_4[0:0], termf_2[0:0]);
  C2 I241 (ha5__0[1:1], termf_4[0:0], termt_2[0:0]);
  C2 I242 (ha5__0[2:2], termt_4[0:0], termf_2[0:0]);
  C2 I243 (ha5__0[3:3], termt_4[0:0], termt_2[0:0]);
  OR3 I244 (cf5__0[0:0], ha5__0[0:0], ha5__0[1:1], ha5__0[2:2]);
  BUFF I245 (ct5__0[0:0], ha5__0[3:3]);
  OR2 I246 (termf_5[0:0], ha5__0[0:0], ha5__0[3:3]);
  OR2 I247 (termt_5[0:0], ha5__0[1:1], ha5__0[2:2]);
  C3 I248 (fa5_1min_0[0:0], cf5__0[0:0], termf_4[1:1], termf_2[1:1]);
  C3 I249 (fa5_1min_0[1:1], cf5__0[0:0], termf_4[1:1], termt_2[1:1]);
  C3 I250 (fa5_1min_0[2:2], cf5__0[0:0], termt_4[1:1], termf_2[1:1]);
  C3 I251 (fa5_1min_0[3:3], cf5__0[0:0], termt_4[1:1], termt_2[1:1]);
  C3 I252 (fa5_1min_0[4:4], ct5__0[0:0], termf_4[1:1], termf_2[1:1]);
  C3 I253 (fa5_1min_0[5:5], ct5__0[0:0], termf_4[1:1], termt_2[1:1]);
  C3 I254 (fa5_1min_0[6:6], ct5__0[0:0], termt_4[1:1], termf_2[1:1]);
  C3 I255 (fa5_1min_0[7:7], ct5__0[0:0], termt_4[1:1], termt_2[1:1]);
  NOR3 I256 (simp2411_0[0:0], fa5_1min_0[0:0], fa5_1min_0[3:3], fa5_1min_0[5:5]);
  INV I257 (simp2411_0[1:1], fa5_1min_0[6:6]);
  NAND2 I258 (termf_5[1:1], simp2411_0[0:0], simp2411_0[1:1]);
  NOR3 I259 (simp2421_0[0:0], fa5_1min_0[1:1], fa5_1min_0[2:2], fa5_1min_0[4:4]);
  INV I260 (simp2421_0[1:1], fa5_1min_0[7:7]);
  NAND2 I261 (termt_5[1:1], simp2421_0[0:0], simp2421_0[1:1]);
  AO222 I262 (ct5__0[1:1], termt_2[1:1], termt_4[1:1], termt_2[1:1], ct5__0[0:0], termt_4[1:1], ct5__0[0:0]);
  AO222 I263 (cf5__0[1:1], termf_2[1:1], termf_4[1:1], termf_2[1:1], cf5__0[0:0], termf_4[1:1], cf5__0[0:0]);
  C3 I264 (fa5_2min_0[0:0], cf5__0[1:1], termf_4[2:2], termf_2[2:2]);
  C3 I265 (fa5_2min_0[1:1], cf5__0[1:1], termf_4[2:2], termt_2[2:2]);
  C3 I266 (fa5_2min_0[2:2], cf5__0[1:1], termt_4[2:2], termf_2[2:2]);
  C3 I267 (fa5_2min_0[3:3], cf5__0[1:1], termt_4[2:2], termt_2[2:2]);
  C3 I268 (fa5_2min_0[4:4], ct5__0[1:1], termf_4[2:2], termf_2[2:2]);
  C3 I269 (fa5_2min_0[5:5], ct5__0[1:1], termf_4[2:2], termt_2[2:2]);
  C3 I270 (fa5_2min_0[6:6], ct5__0[1:1], termt_4[2:2], termf_2[2:2]);
  C3 I271 (fa5_2min_0[7:7], ct5__0[1:1], termt_4[2:2], termt_2[2:2]);
  NOR3 I272 (simp2541_0[0:0], fa5_2min_0[0:0], fa5_2min_0[3:3], fa5_2min_0[5:5]);
  INV I273 (simp2541_0[1:1], fa5_2min_0[6:6]);
  NAND2 I274 (termf_5[2:2], simp2541_0[0:0], simp2541_0[1:1]);
  NOR3 I275 (simp2551_0[0:0], fa5_2min_0[1:1], fa5_2min_0[2:2], fa5_2min_0[4:4]);
  INV I276 (simp2551_0[1:1], fa5_2min_0[7:7]);
  NAND2 I277 (termt_5[2:2], simp2551_0[0:0], simp2551_0[1:1]);
  AO222 I278 (ct5__0[2:2], termt_2[2:2], termt_4[2:2], termt_2[2:2], ct5__0[1:1], termt_4[2:2], ct5__0[1:1]);
  AO222 I279 (cf5__0[2:2], termf_2[2:2], termf_4[2:2], termf_2[2:2], cf5__0[1:1], termf_4[2:2], cf5__0[1:1]);
  C3 I280 (fa5_3min_0[0:0], cf5__0[2:2], termf_4[3:3], termf_2[3:3]);
  C3 I281 (fa5_3min_0[1:1], cf5__0[2:2], termf_4[3:3], termt_2[3:3]);
  C3 I282 (fa5_3min_0[2:2], cf5__0[2:2], termt_4[3:3], termf_2[3:3]);
  C3 I283 (fa5_3min_0[3:3], cf5__0[2:2], termt_4[3:3], termt_2[3:3]);
  C3 I284 (fa5_3min_0[4:4], ct5__0[2:2], termf_4[3:3], termf_2[3:3]);
  C3 I285 (fa5_3min_0[5:5], ct5__0[2:2], termf_4[3:3], termt_2[3:3]);
  C3 I286 (fa5_3min_0[6:6], ct5__0[2:2], termt_4[3:3], termf_2[3:3]);
  C3 I287 (fa5_3min_0[7:7], ct5__0[2:2], termt_4[3:3], termt_2[3:3]);
  NOR3 I288 (simp2671_0[0:0], fa5_3min_0[0:0], fa5_3min_0[3:3], fa5_3min_0[5:5]);
  INV I289 (simp2671_0[1:1], fa5_3min_0[6:6]);
  NAND2 I290 (termf_5[3:3], simp2671_0[0:0], simp2671_0[1:1]);
  NOR3 I291 (simp2681_0[0:0], fa5_3min_0[1:1], fa5_3min_0[2:2], fa5_3min_0[4:4]);
  INV I292 (simp2681_0[1:1], fa5_3min_0[7:7]);
  NAND2 I293 (termt_5[3:3], simp2681_0[0:0], simp2681_0[1:1]);
  AO222 I294 (ct5__0[3:3], termt_2[3:3], termt_4[3:3], termt_2[3:3], ct5__0[2:2], termt_4[3:3], ct5__0[2:2]);
  AO222 I295 (cf5__0[3:3], termf_2[3:3], termf_4[3:3], termf_2[3:3], cf5__0[2:2], termf_4[3:3], cf5__0[2:2]);
  C3 I296 (fa5_4min_0[0:0], cf5__0[3:3], termf_4[4:4], termf_2[4:4]);
  C3 I297 (fa5_4min_0[1:1], cf5__0[3:3], termf_4[4:4], termt_2[4:4]);
  C3 I298 (fa5_4min_0[2:2], cf5__0[3:3], termt_4[4:4], termf_2[4:4]);
  C3 I299 (fa5_4min_0[3:3], cf5__0[3:3], termt_4[4:4], termt_2[4:4]);
  C3 I300 (fa5_4min_0[4:4], ct5__0[3:3], termf_4[4:4], termf_2[4:4]);
  C3 I301 (fa5_4min_0[5:5], ct5__0[3:3], termf_4[4:4], termt_2[4:4]);
  C3 I302 (fa5_4min_0[6:6], ct5__0[3:3], termt_4[4:4], termf_2[4:4]);
  C3 I303 (fa5_4min_0[7:7], ct5__0[3:3], termt_4[4:4], termt_2[4:4]);
  NOR3 I304 (simp2801_0[0:0], fa5_4min_0[0:0], fa5_4min_0[3:3], fa5_4min_0[5:5]);
  INV I305 (simp2801_0[1:1], fa5_4min_0[6:6]);
  NAND2 I306 (termf_5[4:4], simp2801_0[0:0], simp2801_0[1:1]);
  NOR3 I307 (simp2811_0[0:0], fa5_4min_0[1:1], fa5_4min_0[2:2], fa5_4min_0[4:4]);
  INV I308 (simp2811_0[1:1], fa5_4min_0[7:7]);
  NAND2 I309 (termt_5[4:4], simp2811_0[0:0], simp2811_0[1:1]);
  AO222 I310 (ct5__0[4:4], termt_2[4:4], termt_4[4:4], termt_2[4:4], ct5__0[3:3], termt_4[4:4], ct5__0[3:3]);
  AO222 I311 (cf5__0[4:4], termf_2[4:4], termf_4[4:4], termf_2[4:4], cf5__0[3:3], termf_4[4:4], cf5__0[3:3]);
  C3 I312 (fa5_5min_0[0:0], cf5__0[4:4], termf_4[5:5], termf_2[5:5]);
  C3 I313 (fa5_5min_0[1:1], cf5__0[4:4], termf_4[5:5], termt_2[5:5]);
  C3 I314 (fa5_5min_0[2:2], cf5__0[4:4], termt_4[5:5], termf_2[5:5]);
  C3 I315 (fa5_5min_0[3:3], cf5__0[4:4], termt_4[5:5], termt_2[5:5]);
  C3 I316 (fa5_5min_0[4:4], ct5__0[4:4], termf_4[5:5], termf_2[5:5]);
  C3 I317 (fa5_5min_0[5:5], ct5__0[4:4], termf_4[5:5], termt_2[5:5]);
  C3 I318 (fa5_5min_0[6:6], ct5__0[4:4], termt_4[5:5], termf_2[5:5]);
  C3 I319 (fa5_5min_0[7:7], ct5__0[4:4], termt_4[5:5], termt_2[5:5]);
  NOR3 I320 (simp2931_0[0:0], fa5_5min_0[0:0], fa5_5min_0[3:3], fa5_5min_0[5:5]);
  INV I321 (simp2931_0[1:1], fa5_5min_0[6:6]);
  NAND2 I322 (termf_5[5:5], simp2931_0[0:0], simp2931_0[1:1]);
  NOR3 I323 (simp2941_0[0:0], fa5_5min_0[1:1], fa5_5min_0[2:2], fa5_5min_0[4:4]);
  INV I324 (simp2941_0[1:1], fa5_5min_0[7:7]);
  NAND2 I325 (termt_5[5:5], simp2941_0[0:0], simp2941_0[1:1]);
  AO222 I326 (ct5__0[5:5], termt_2[5:5], termt_4[5:5], termt_2[5:5], ct5__0[4:4], termt_4[5:5], ct5__0[4:4]);
  AO222 I327 (cf5__0[5:5], termf_2[5:5], termf_4[5:5], termf_2[5:5], cf5__0[4:4], termf_4[5:5], cf5__0[4:4]);
  C3 I328 (fa5_6min_0[0:0], cf5__0[5:5], termf_4[6:6], termf_2[6:6]);
  C3 I329 (fa5_6min_0[1:1], cf5__0[5:5], termf_4[6:6], termt_2[6:6]);
  C3 I330 (fa5_6min_0[2:2], cf5__0[5:5], termt_4[6:6], termf_2[6:6]);
  C3 I331 (fa5_6min_0[3:3], cf5__0[5:5], termt_4[6:6], termt_2[6:6]);
  C3 I332 (fa5_6min_0[4:4], ct5__0[5:5], termf_4[6:6], termf_2[6:6]);
  C3 I333 (fa5_6min_0[5:5], ct5__0[5:5], termf_4[6:6], termt_2[6:6]);
  C3 I334 (fa5_6min_0[6:6], ct5__0[5:5], termt_4[6:6], termf_2[6:6]);
  C3 I335 (fa5_6min_0[7:7], ct5__0[5:5], termt_4[6:6], termt_2[6:6]);
  NOR3 I336 (simp3061_0[0:0], fa5_6min_0[0:0], fa5_6min_0[3:3], fa5_6min_0[5:5]);
  INV I337 (simp3061_0[1:1], fa5_6min_0[6:6]);
  NAND2 I338 (termf_5[6:6], simp3061_0[0:0], simp3061_0[1:1]);
  NOR3 I339 (simp3071_0[0:0], fa5_6min_0[1:1], fa5_6min_0[2:2], fa5_6min_0[4:4]);
  INV I340 (simp3071_0[1:1], fa5_6min_0[7:7]);
  NAND2 I341 (termt_5[6:6], simp3071_0[0:0], simp3071_0[1:1]);
  AO222 I342 (ct5__0[6:6], termt_2[6:6], termt_4[6:6], termt_2[6:6], ct5__0[5:5], termt_4[6:6], ct5__0[5:5]);
  AO222 I343 (cf5__0[6:6], termf_2[6:6], termf_4[6:6], termf_2[6:6], cf5__0[5:5], termf_4[6:6], cf5__0[5:5]);
  C3 I344 (fa5_7min_0[0:0], cf5__0[6:6], termf_4[7:7], termf_2[7:7]);
  C3 I345 (fa5_7min_0[1:1], cf5__0[6:6], termf_4[7:7], termt_2[7:7]);
  C3 I346 (fa5_7min_0[2:2], cf5__0[6:6], termt_4[7:7], termf_2[7:7]);
  C3 I347 (fa5_7min_0[3:3], cf5__0[6:6], termt_4[7:7], termt_2[7:7]);
  C3 I348 (fa5_7min_0[4:4], ct5__0[6:6], termf_4[7:7], termf_2[7:7]);
  C3 I349 (fa5_7min_0[5:5], ct5__0[6:6], termf_4[7:7], termt_2[7:7]);
  C3 I350 (fa5_7min_0[6:6], ct5__0[6:6], termt_4[7:7], termf_2[7:7]);
  C3 I351 (fa5_7min_0[7:7], ct5__0[6:6], termt_4[7:7], termt_2[7:7]);
  NOR3 I352 (simp3191_0[0:0], fa5_7min_0[0:0], fa5_7min_0[3:3], fa5_7min_0[5:5]);
  INV I353 (simp3191_0[1:1], fa5_7min_0[6:6]);
  NAND2 I354 (termf_5[7:7], simp3191_0[0:0], simp3191_0[1:1]);
  NOR3 I355 (simp3201_0[0:0], fa5_7min_0[1:1], fa5_7min_0[2:2], fa5_7min_0[4:4]);
  INV I356 (simp3201_0[1:1], fa5_7min_0[7:7]);
  NAND2 I357 (termt_5[7:7], simp3201_0[0:0], simp3201_0[1:1]);
  AO222 I358 (ct5__0[7:7], termt_2[7:7], termt_4[7:7], termt_2[7:7], ct5__0[6:6], termt_4[7:7], ct5__0[6:6]);
  AO222 I359 (cf5__0[7:7], termf_2[7:7], termf_4[7:7], termf_2[7:7], cf5__0[6:6], termf_4[7:7], cf5__0[6:6]);
  C3 I360 (fa5_8min_0[0:0], cf5__0[7:7], termf_4[8:8], termf_2[8:8]);
  C3 I361 (fa5_8min_0[1:1], cf5__0[7:7], termf_4[8:8], termt_2[8:8]);
  C3 I362 (fa5_8min_0[2:2], cf5__0[7:7], termt_4[8:8], termf_2[8:8]);
  C3 I363 (fa5_8min_0[3:3], cf5__0[7:7], termt_4[8:8], termt_2[8:8]);
  C3 I364 (fa5_8min_0[4:4], ct5__0[7:7], termf_4[8:8], termf_2[8:8]);
  C3 I365 (fa5_8min_0[5:5], ct5__0[7:7], termf_4[8:8], termt_2[8:8]);
  C3 I366 (fa5_8min_0[6:6], ct5__0[7:7], termt_4[8:8], termf_2[8:8]);
  C3 I367 (fa5_8min_0[7:7], ct5__0[7:7], termt_4[8:8], termt_2[8:8]);
  NOR3 I368 (simp3321_0[0:0], fa5_8min_0[0:0], fa5_8min_0[3:3], fa5_8min_0[5:5]);
  INV I369 (simp3321_0[1:1], fa5_8min_0[6:6]);
  NAND2 I370 (termf_5[8:8], simp3321_0[0:0], simp3321_0[1:1]);
  NOR3 I371 (simp3331_0[0:0], fa5_8min_0[1:1], fa5_8min_0[2:2], fa5_8min_0[4:4]);
  INV I372 (simp3331_0[1:1], fa5_8min_0[7:7]);
  NAND2 I373 (termt_5[8:8], simp3331_0[0:0], simp3331_0[1:1]);
  AO222 I374 (ct5__0[8:8], termt_2[8:8], termt_4[8:8], termt_2[8:8], ct5__0[7:7], termt_4[8:8], ct5__0[7:7]);
  AO222 I375 (cf5__0[8:8], termf_2[8:8], termf_4[8:8], termf_2[8:8], cf5__0[7:7], termf_4[8:8], cf5__0[7:7]);
  C3 I376 (fa5_9min_0[0:0], cf5__0[8:8], termf_4[9:9], termf_2[9:9]);
  C3 I377 (fa5_9min_0[1:1], cf5__0[8:8], termf_4[9:9], termt_2[9:9]);
  C3 I378 (fa5_9min_0[2:2], cf5__0[8:8], termt_4[9:9], termf_2[9:9]);
  C3 I379 (fa5_9min_0[3:3], cf5__0[8:8], termt_4[9:9], termt_2[9:9]);
  C3 I380 (fa5_9min_0[4:4], ct5__0[8:8], termf_4[9:9], termf_2[9:9]);
  C3 I381 (fa5_9min_0[5:5], ct5__0[8:8], termf_4[9:9], termt_2[9:9]);
  C3 I382 (fa5_9min_0[6:6], ct5__0[8:8], termt_4[9:9], termf_2[9:9]);
  C3 I383 (fa5_9min_0[7:7], ct5__0[8:8], termt_4[9:9], termt_2[9:9]);
  NOR3 I384 (simp3451_0[0:0], fa5_9min_0[0:0], fa5_9min_0[3:3], fa5_9min_0[5:5]);
  INV I385 (simp3451_0[1:1], fa5_9min_0[6:6]);
  NAND2 I386 (termf_5[9:9], simp3451_0[0:0], simp3451_0[1:1]);
  NOR3 I387 (simp3461_0[0:0], fa5_9min_0[1:1], fa5_9min_0[2:2], fa5_9min_0[4:4]);
  INV I388 (simp3461_0[1:1], fa5_9min_0[7:7]);
  NAND2 I389 (termt_5[9:9], simp3461_0[0:0], simp3461_0[1:1]);
  AO222 I390 (ct5__0[9:9], termt_2[9:9], termt_4[9:9], termt_2[9:9], ct5__0[8:8], termt_4[9:9], ct5__0[8:8]);
  AO222 I391 (cf5__0[9:9], termf_2[9:9], termf_4[9:9], termf_2[9:9], cf5__0[8:8], termf_4[9:9], cf5__0[8:8]);
  C3 I392 (fa5_10min_0[0:0], cf5__0[9:9], termf_4[10:10], termf_2[10:10]);
  C3 I393 (fa5_10min_0[1:1], cf5__0[9:9], termf_4[10:10], termt_2[10:10]);
  C3 I394 (fa5_10min_0[2:2], cf5__0[9:9], termt_4[10:10], termf_2[10:10]);
  C3 I395 (fa5_10min_0[3:3], cf5__0[9:9], termt_4[10:10], termt_2[10:10]);
  C3 I396 (fa5_10min_0[4:4], ct5__0[9:9], termf_4[10:10], termf_2[10:10]);
  C3 I397 (fa5_10min_0[5:5], ct5__0[9:9], termf_4[10:10], termt_2[10:10]);
  C3 I398 (fa5_10min_0[6:6], ct5__0[9:9], termt_4[10:10], termf_2[10:10]);
  C3 I399 (fa5_10min_0[7:7], ct5__0[9:9], termt_4[10:10], termt_2[10:10]);
  NOR3 I400 (simp3581_0[0:0], fa5_10min_0[0:0], fa5_10min_0[3:3], fa5_10min_0[5:5]);
  INV I401 (simp3581_0[1:1], fa5_10min_0[6:6]);
  NAND2 I402 (termf_5[10:10], simp3581_0[0:0], simp3581_0[1:1]);
  NOR3 I403 (simp3591_0[0:0], fa5_10min_0[1:1], fa5_10min_0[2:2], fa5_10min_0[4:4]);
  INV I404 (simp3591_0[1:1], fa5_10min_0[7:7]);
  NAND2 I405 (termt_5[10:10], simp3591_0[0:0], simp3591_0[1:1]);
  AO222 I406 (ct5__0[10:10], termt_2[10:10], termt_4[10:10], termt_2[10:10], ct5__0[9:9], termt_4[10:10], ct5__0[9:9]);
  AO222 I407 (cf5__0[10:10], termf_2[10:10], termf_4[10:10], termf_2[10:10], cf5__0[9:9], termf_4[10:10], cf5__0[9:9]);
  C3 I408 (fa5_11min_0[0:0], cf5__0[10:10], termf_4[11:11], termf_2[11:11]);
  C3 I409 (fa5_11min_0[1:1], cf5__0[10:10], termf_4[11:11], termt_2[11:11]);
  C3 I410 (fa5_11min_0[2:2], cf5__0[10:10], termt_4[11:11], termf_2[11:11]);
  C3 I411 (fa5_11min_0[3:3], cf5__0[10:10], termt_4[11:11], termt_2[11:11]);
  C3 I412 (fa5_11min_0[4:4], ct5__0[10:10], termf_4[11:11], termf_2[11:11]);
  C3 I413 (fa5_11min_0[5:5], ct5__0[10:10], termf_4[11:11], termt_2[11:11]);
  C3 I414 (fa5_11min_0[6:6], ct5__0[10:10], termt_4[11:11], termf_2[11:11]);
  C3 I415 (fa5_11min_0[7:7], ct5__0[10:10], termt_4[11:11], termt_2[11:11]);
  NOR3 I416 (simp3711_0[0:0], fa5_11min_0[0:0], fa5_11min_0[3:3], fa5_11min_0[5:5]);
  INV I417 (simp3711_0[1:1], fa5_11min_0[6:6]);
  NAND2 I418 (termf_5[11:11], simp3711_0[0:0], simp3711_0[1:1]);
  NOR3 I419 (simp3721_0[0:0], fa5_11min_0[1:1], fa5_11min_0[2:2], fa5_11min_0[4:4]);
  INV I420 (simp3721_0[1:1], fa5_11min_0[7:7]);
  NAND2 I421 (termt_5[11:11], simp3721_0[0:0], simp3721_0[1:1]);
  AO222 I422 (ct5__0[11:11], termt_2[11:11], termt_4[11:11], termt_2[11:11], ct5__0[10:10], termt_4[11:11], ct5__0[10:10]);
  AO222 I423 (cf5__0[11:11], termf_2[11:11], termf_4[11:11], termf_2[11:11], cf5__0[10:10], termf_4[11:11], cf5__0[10:10]);
  C3 I424 (fa5_12min_0[0:0], cf5__0[11:11], termf_4[12:12], termf_2[12:12]);
  C3 I425 (fa5_12min_0[1:1], cf5__0[11:11], termf_4[12:12], termt_2[12:12]);
  C3 I426 (fa5_12min_0[2:2], cf5__0[11:11], termt_4[12:12], termf_2[12:12]);
  C3 I427 (fa5_12min_0[3:3], cf5__0[11:11], termt_4[12:12], termt_2[12:12]);
  C3 I428 (fa5_12min_0[4:4], ct5__0[11:11], termf_4[12:12], termf_2[12:12]);
  C3 I429 (fa5_12min_0[5:5], ct5__0[11:11], termf_4[12:12], termt_2[12:12]);
  C3 I430 (fa5_12min_0[6:6], ct5__0[11:11], termt_4[12:12], termf_2[12:12]);
  C3 I431 (fa5_12min_0[7:7], ct5__0[11:11], termt_4[12:12], termt_2[12:12]);
  NOR3 I432 (simp3841_0[0:0], fa5_12min_0[0:0], fa5_12min_0[3:3], fa5_12min_0[5:5]);
  INV I433 (simp3841_0[1:1], fa5_12min_0[6:6]);
  NAND2 I434 (termf_5[12:12], simp3841_0[0:0], simp3841_0[1:1]);
  NOR3 I435 (simp3851_0[0:0], fa5_12min_0[1:1], fa5_12min_0[2:2], fa5_12min_0[4:4]);
  INV I436 (simp3851_0[1:1], fa5_12min_0[7:7]);
  NAND2 I437 (termt_5[12:12], simp3851_0[0:0], simp3851_0[1:1]);
  AO222 I438 (ct5__0[12:12], termt_2[12:12], termt_4[12:12], termt_2[12:12], ct5__0[11:11], termt_4[12:12], ct5__0[11:11]);
  AO222 I439 (cf5__0[12:12], termf_2[12:12], termf_4[12:12], termf_2[12:12], cf5__0[11:11], termf_4[12:12], cf5__0[11:11]);
  C3 I440 (fa5_13min_0[0:0], cf5__0[12:12], termf_4[13:13], termf_2[13:13]);
  C3 I441 (fa5_13min_0[1:1], cf5__0[12:12], termf_4[13:13], termt_2[13:13]);
  C3 I442 (fa5_13min_0[2:2], cf5__0[12:12], termt_4[13:13], termf_2[13:13]);
  C3 I443 (fa5_13min_0[3:3], cf5__0[12:12], termt_4[13:13], termt_2[13:13]);
  C3 I444 (fa5_13min_0[4:4], ct5__0[12:12], termf_4[13:13], termf_2[13:13]);
  C3 I445 (fa5_13min_0[5:5], ct5__0[12:12], termf_4[13:13], termt_2[13:13]);
  C3 I446 (fa5_13min_0[6:6], ct5__0[12:12], termt_4[13:13], termf_2[13:13]);
  C3 I447 (fa5_13min_0[7:7], ct5__0[12:12], termt_4[13:13], termt_2[13:13]);
  NOR3 I448 (simp3971_0[0:0], fa5_13min_0[0:0], fa5_13min_0[3:3], fa5_13min_0[5:5]);
  INV I449 (simp3971_0[1:1], fa5_13min_0[6:6]);
  NAND2 I450 (termf_5[13:13], simp3971_0[0:0], simp3971_0[1:1]);
  NOR3 I451 (simp3981_0[0:0], fa5_13min_0[1:1], fa5_13min_0[2:2], fa5_13min_0[4:4]);
  INV I452 (simp3981_0[1:1], fa5_13min_0[7:7]);
  NAND2 I453 (termt_5[13:13], simp3981_0[0:0], simp3981_0[1:1]);
  AO222 I454 (ct5__0[13:13], termt_2[13:13], termt_4[13:13], termt_2[13:13], ct5__0[12:12], termt_4[13:13], ct5__0[12:12]);
  AO222 I455 (cf5__0[13:13], termf_2[13:13], termf_4[13:13], termf_2[13:13], cf5__0[12:12], termf_4[13:13], cf5__0[12:12]);
  C3 I456 (fa5_14min_0[0:0], cf5__0[13:13], termf_4[14:14], termf_2[14:14]);
  C3 I457 (fa5_14min_0[1:1], cf5__0[13:13], termf_4[14:14], termt_2[14:14]);
  C3 I458 (fa5_14min_0[2:2], cf5__0[13:13], termt_4[14:14], termf_2[14:14]);
  C3 I459 (fa5_14min_0[3:3], cf5__0[13:13], termt_4[14:14], termt_2[14:14]);
  C3 I460 (fa5_14min_0[4:4], ct5__0[13:13], termf_4[14:14], termf_2[14:14]);
  C3 I461 (fa5_14min_0[5:5], ct5__0[13:13], termf_4[14:14], termt_2[14:14]);
  C3 I462 (fa5_14min_0[6:6], ct5__0[13:13], termt_4[14:14], termf_2[14:14]);
  C3 I463 (fa5_14min_0[7:7], ct5__0[13:13], termt_4[14:14], termt_2[14:14]);
  NOR3 I464 (simp4101_0[0:0], fa5_14min_0[0:0], fa5_14min_0[3:3], fa5_14min_0[5:5]);
  INV I465 (simp4101_0[1:1], fa5_14min_0[6:6]);
  NAND2 I466 (termf_5[14:14], simp4101_0[0:0], simp4101_0[1:1]);
  NOR3 I467 (simp4111_0[0:0], fa5_14min_0[1:1], fa5_14min_0[2:2], fa5_14min_0[4:4]);
  INV I468 (simp4111_0[1:1], fa5_14min_0[7:7]);
  NAND2 I469 (termt_5[14:14], simp4111_0[0:0], simp4111_0[1:1]);
  AO222 I470 (ct5__0[14:14], termt_2[14:14], termt_4[14:14], termt_2[14:14], ct5__0[13:13], termt_4[14:14], ct5__0[13:13]);
  AO222 I471 (cf5__0[14:14], termf_2[14:14], termf_4[14:14], termf_2[14:14], cf5__0[13:13], termf_4[14:14], cf5__0[13:13]);
  C3 I472 (fa5_15min_0[0:0], cf5__0[14:14], termf_4[15:15], termf_2[15:15]);
  C3 I473 (fa5_15min_0[1:1], cf5__0[14:14], termf_4[15:15], termt_2[15:15]);
  C3 I474 (fa5_15min_0[2:2], cf5__0[14:14], termt_4[15:15], termf_2[15:15]);
  C3 I475 (fa5_15min_0[3:3], cf5__0[14:14], termt_4[15:15], termt_2[15:15]);
  C3 I476 (fa5_15min_0[4:4], ct5__0[14:14], termf_4[15:15], termf_2[15:15]);
  C3 I477 (fa5_15min_0[5:5], ct5__0[14:14], termf_4[15:15], termt_2[15:15]);
  C3 I478 (fa5_15min_0[6:6], ct5__0[14:14], termt_4[15:15], termf_2[15:15]);
  C3 I479 (fa5_15min_0[7:7], ct5__0[14:14], termt_4[15:15], termt_2[15:15]);
  NOR3 I480 (simp4231_0[0:0], fa5_15min_0[0:0], fa5_15min_0[3:3], fa5_15min_0[5:5]);
  INV I481 (simp4231_0[1:1], fa5_15min_0[6:6]);
  NAND2 I482 (termf_5[15:15], simp4231_0[0:0], simp4231_0[1:1]);
  NOR3 I483 (simp4241_0[0:0], fa5_15min_0[1:1], fa5_15min_0[2:2], fa5_15min_0[4:4]);
  INV I484 (simp4241_0[1:1], fa5_15min_0[7:7]);
  NAND2 I485 (termt_5[15:15], simp4241_0[0:0], simp4241_0[1:1]);
  AO222 I486 (ct5__0[15:15], termt_2[15:15], termt_4[15:15], termt_2[15:15], ct5__0[14:14], termt_4[15:15], ct5__0[14:14]);
  AO222 I487 (cf5__0[15:15], termf_2[15:15], termf_4[15:15], termf_2[15:15], cf5__0[14:14], termf_4[15:15], cf5__0[14:14]);
  C3 I488 (fa5_16min_0[0:0], cf5__0[15:15], termf_4[16:16], termf_2[16:16]);
  C3 I489 (fa5_16min_0[1:1], cf5__0[15:15], termf_4[16:16], termt_2[16:16]);
  C3 I490 (fa5_16min_0[2:2], cf5__0[15:15], termt_4[16:16], termf_2[16:16]);
  C3 I491 (fa5_16min_0[3:3], cf5__0[15:15], termt_4[16:16], termt_2[16:16]);
  C3 I492 (fa5_16min_0[4:4], ct5__0[15:15], termf_4[16:16], termf_2[16:16]);
  C3 I493 (fa5_16min_0[5:5], ct5__0[15:15], termf_4[16:16], termt_2[16:16]);
  C3 I494 (fa5_16min_0[6:6], ct5__0[15:15], termt_4[16:16], termf_2[16:16]);
  C3 I495 (fa5_16min_0[7:7], ct5__0[15:15], termt_4[16:16], termt_2[16:16]);
  NOR3 I496 (simp4361_0[0:0], fa5_16min_0[0:0], fa5_16min_0[3:3], fa5_16min_0[5:5]);
  INV I497 (simp4361_0[1:1], fa5_16min_0[6:6]);
  NAND2 I498 (termf_5[16:16], simp4361_0[0:0], simp4361_0[1:1]);
  NOR3 I499 (simp4371_0[0:0], fa5_16min_0[1:1], fa5_16min_0[2:2], fa5_16min_0[4:4]);
  INV I500 (simp4371_0[1:1], fa5_16min_0[7:7]);
  NAND2 I501 (termt_5[16:16], simp4371_0[0:0], simp4371_0[1:1]);
  AO222 I502 (ct5__0[16:16], termt_2[16:16], termt_4[16:16], termt_2[16:16], ct5__0[15:15], termt_4[16:16], ct5__0[15:15]);
  AO222 I503 (cf5__0[16:16], termf_2[16:16], termf_4[16:16], termf_2[16:16], cf5__0[15:15], termf_4[16:16], cf5__0[15:15]);
  C3 I504 (fa5_17min_0[0:0], cf5__0[16:16], termf_4[17:17], termf_2[17:17]);
  C3 I505 (fa5_17min_0[1:1], cf5__0[16:16], termf_4[17:17], termt_2[17:17]);
  C3 I506 (fa5_17min_0[2:2], cf5__0[16:16], termt_4[17:17], termf_2[17:17]);
  C3 I507 (fa5_17min_0[3:3], cf5__0[16:16], termt_4[17:17], termt_2[17:17]);
  C3 I508 (fa5_17min_0[4:4], ct5__0[16:16], termf_4[17:17], termf_2[17:17]);
  C3 I509 (fa5_17min_0[5:5], ct5__0[16:16], termf_4[17:17], termt_2[17:17]);
  C3 I510 (fa5_17min_0[6:6], ct5__0[16:16], termt_4[17:17], termf_2[17:17]);
  C3 I511 (fa5_17min_0[7:7], ct5__0[16:16], termt_4[17:17], termt_2[17:17]);
  NOR3 I512 (simp4491_0[0:0], fa5_17min_0[0:0], fa5_17min_0[3:3], fa5_17min_0[5:5]);
  INV I513 (simp4491_0[1:1], fa5_17min_0[6:6]);
  NAND2 I514 (termf_5[17:17], simp4491_0[0:0], simp4491_0[1:1]);
  NOR3 I515 (simp4501_0[0:0], fa5_17min_0[1:1], fa5_17min_0[2:2], fa5_17min_0[4:4]);
  INV I516 (simp4501_0[1:1], fa5_17min_0[7:7]);
  NAND2 I517 (termt_5[17:17], simp4501_0[0:0], simp4501_0[1:1]);
  AO222 I518 (ct5__0[17:17], termt_2[17:17], termt_4[17:17], termt_2[17:17], ct5__0[16:16], termt_4[17:17], ct5__0[16:16]);
  AO222 I519 (cf5__0[17:17], termf_2[17:17], termf_4[17:17], termf_2[17:17], cf5__0[16:16], termf_4[17:17], cf5__0[16:16]);
  C3 I520 (fa5_18min_0[0:0], cf5__0[17:17], termf_4[18:18], termf_2[18:18]);
  C3 I521 (fa5_18min_0[1:1], cf5__0[17:17], termf_4[18:18], termt_2[18:18]);
  C3 I522 (fa5_18min_0[2:2], cf5__0[17:17], termt_4[18:18], termf_2[18:18]);
  C3 I523 (fa5_18min_0[3:3], cf5__0[17:17], termt_4[18:18], termt_2[18:18]);
  C3 I524 (fa5_18min_0[4:4], ct5__0[17:17], termf_4[18:18], termf_2[18:18]);
  C3 I525 (fa5_18min_0[5:5], ct5__0[17:17], termf_4[18:18], termt_2[18:18]);
  C3 I526 (fa5_18min_0[6:6], ct5__0[17:17], termt_4[18:18], termf_2[18:18]);
  C3 I527 (fa5_18min_0[7:7], ct5__0[17:17], termt_4[18:18], termt_2[18:18]);
  NOR3 I528 (simp4621_0[0:0], fa5_18min_0[0:0], fa5_18min_0[3:3], fa5_18min_0[5:5]);
  INV I529 (simp4621_0[1:1], fa5_18min_0[6:6]);
  NAND2 I530 (termf_5[18:18], simp4621_0[0:0], simp4621_0[1:1]);
  NOR3 I531 (simp4631_0[0:0], fa5_18min_0[1:1], fa5_18min_0[2:2], fa5_18min_0[4:4]);
  INV I532 (simp4631_0[1:1], fa5_18min_0[7:7]);
  NAND2 I533 (termt_5[18:18], simp4631_0[0:0], simp4631_0[1:1]);
  AO222 I534 (ct5__0[18:18], termt_2[18:18], termt_4[18:18], termt_2[18:18], ct5__0[17:17], termt_4[18:18], ct5__0[17:17]);
  AO222 I535 (cf5__0[18:18], termf_2[18:18], termf_4[18:18], termf_2[18:18], cf5__0[17:17], termf_4[18:18], cf5__0[17:17]);
  C3 I536 (fa5_19min_0[0:0], cf5__0[18:18], termf_4[19:19], termf_2[19:19]);
  C3 I537 (fa5_19min_0[1:1], cf5__0[18:18], termf_4[19:19], termt_2[19:19]);
  C3 I538 (fa5_19min_0[2:2], cf5__0[18:18], termt_4[19:19], termf_2[19:19]);
  C3 I539 (fa5_19min_0[3:3], cf5__0[18:18], termt_4[19:19], termt_2[19:19]);
  C3 I540 (fa5_19min_0[4:4], ct5__0[18:18], termf_4[19:19], termf_2[19:19]);
  C3 I541 (fa5_19min_0[5:5], ct5__0[18:18], termf_4[19:19], termt_2[19:19]);
  C3 I542 (fa5_19min_0[6:6], ct5__0[18:18], termt_4[19:19], termf_2[19:19]);
  C3 I543 (fa5_19min_0[7:7], ct5__0[18:18], termt_4[19:19], termt_2[19:19]);
  NOR3 I544 (simp4751_0[0:0], fa5_19min_0[0:0], fa5_19min_0[3:3], fa5_19min_0[5:5]);
  INV I545 (simp4751_0[1:1], fa5_19min_0[6:6]);
  NAND2 I546 (termf_5[19:19], simp4751_0[0:0], simp4751_0[1:1]);
  NOR3 I547 (simp4761_0[0:0], fa5_19min_0[1:1], fa5_19min_0[2:2], fa5_19min_0[4:4]);
  INV I548 (simp4761_0[1:1], fa5_19min_0[7:7]);
  NAND2 I549 (termt_5[19:19], simp4761_0[0:0], simp4761_0[1:1]);
  AO222 I550 (ct5__0[19:19], termt_2[19:19], termt_4[19:19], termt_2[19:19], ct5__0[18:18], termt_4[19:19], ct5__0[18:18]);
  AO222 I551 (cf5__0[19:19], termf_2[19:19], termf_4[19:19], termf_2[19:19], cf5__0[18:18], termf_4[19:19], cf5__0[18:18]);
  C3 I552 (fa5_20min_0[0:0], cf5__0[19:19], termf_4[20:20], termf_2[20:20]);
  C3 I553 (fa5_20min_0[1:1], cf5__0[19:19], termf_4[20:20], termt_2[20:20]);
  C3 I554 (fa5_20min_0[2:2], cf5__0[19:19], termt_4[20:20], termf_2[20:20]);
  C3 I555 (fa5_20min_0[3:3], cf5__0[19:19], termt_4[20:20], termt_2[20:20]);
  C3 I556 (fa5_20min_0[4:4], ct5__0[19:19], termf_4[20:20], termf_2[20:20]);
  C3 I557 (fa5_20min_0[5:5], ct5__0[19:19], termf_4[20:20], termt_2[20:20]);
  C3 I558 (fa5_20min_0[6:6], ct5__0[19:19], termt_4[20:20], termf_2[20:20]);
  C3 I559 (fa5_20min_0[7:7], ct5__0[19:19], termt_4[20:20], termt_2[20:20]);
  NOR3 I560 (simp4881_0[0:0], fa5_20min_0[0:0], fa5_20min_0[3:3], fa5_20min_0[5:5]);
  INV I561 (simp4881_0[1:1], fa5_20min_0[6:6]);
  NAND2 I562 (termf_5[20:20], simp4881_0[0:0], simp4881_0[1:1]);
  NOR3 I563 (simp4891_0[0:0], fa5_20min_0[1:1], fa5_20min_0[2:2], fa5_20min_0[4:4]);
  INV I564 (simp4891_0[1:1], fa5_20min_0[7:7]);
  NAND2 I565 (termt_5[20:20], simp4891_0[0:0], simp4891_0[1:1]);
  AO222 I566 (ct5__0[20:20], termt_2[20:20], termt_4[20:20], termt_2[20:20], ct5__0[19:19], termt_4[20:20], ct5__0[19:19]);
  AO222 I567 (cf5__0[20:20], termf_2[20:20], termf_4[20:20], termf_2[20:20], cf5__0[19:19], termf_4[20:20], cf5__0[19:19]);
  C3 I568 (fa5_21min_0[0:0], cf5__0[20:20], termf_4[21:21], termf_2[21:21]);
  C3 I569 (fa5_21min_0[1:1], cf5__0[20:20], termf_4[21:21], termt_2[21:21]);
  C3 I570 (fa5_21min_0[2:2], cf5__0[20:20], termt_4[21:21], termf_2[21:21]);
  C3 I571 (fa5_21min_0[3:3], cf5__0[20:20], termt_4[21:21], termt_2[21:21]);
  C3 I572 (fa5_21min_0[4:4], ct5__0[20:20], termf_4[21:21], termf_2[21:21]);
  C3 I573 (fa5_21min_0[5:5], ct5__0[20:20], termf_4[21:21], termt_2[21:21]);
  C3 I574 (fa5_21min_0[6:6], ct5__0[20:20], termt_4[21:21], termf_2[21:21]);
  C3 I575 (fa5_21min_0[7:7], ct5__0[20:20], termt_4[21:21], termt_2[21:21]);
  NOR3 I576 (simp5011_0[0:0], fa5_21min_0[0:0], fa5_21min_0[3:3], fa5_21min_0[5:5]);
  INV I577 (simp5011_0[1:1], fa5_21min_0[6:6]);
  NAND2 I578 (termf_5[21:21], simp5011_0[0:0], simp5011_0[1:1]);
  NOR3 I579 (simp5021_0[0:0], fa5_21min_0[1:1], fa5_21min_0[2:2], fa5_21min_0[4:4]);
  INV I580 (simp5021_0[1:1], fa5_21min_0[7:7]);
  NAND2 I581 (termt_5[21:21], simp5021_0[0:0], simp5021_0[1:1]);
  AO222 I582 (ct5__0[21:21], termt_2[21:21], termt_4[21:21], termt_2[21:21], ct5__0[20:20], termt_4[21:21], ct5__0[20:20]);
  AO222 I583 (cf5__0[21:21], termf_2[21:21], termf_4[21:21], termf_2[21:21], cf5__0[20:20], termf_4[21:21], cf5__0[20:20]);
  C3 I584 (fa5_22min_0[0:0], cf5__0[21:21], termf_4[22:22], termf_2[22:22]);
  C3 I585 (fa5_22min_0[1:1], cf5__0[21:21], termf_4[22:22], termt_2[22:22]);
  C3 I586 (fa5_22min_0[2:2], cf5__0[21:21], termt_4[22:22], termf_2[22:22]);
  C3 I587 (fa5_22min_0[3:3], cf5__0[21:21], termt_4[22:22], termt_2[22:22]);
  C3 I588 (fa5_22min_0[4:4], ct5__0[21:21], termf_4[22:22], termf_2[22:22]);
  C3 I589 (fa5_22min_0[5:5], ct5__0[21:21], termf_4[22:22], termt_2[22:22]);
  C3 I590 (fa5_22min_0[6:6], ct5__0[21:21], termt_4[22:22], termf_2[22:22]);
  C3 I591 (fa5_22min_0[7:7], ct5__0[21:21], termt_4[22:22], termt_2[22:22]);
  NOR3 I592 (simp5141_0[0:0], fa5_22min_0[0:0], fa5_22min_0[3:3], fa5_22min_0[5:5]);
  INV I593 (simp5141_0[1:1], fa5_22min_0[6:6]);
  NAND2 I594 (termf_5[22:22], simp5141_0[0:0], simp5141_0[1:1]);
  NOR3 I595 (simp5151_0[0:0], fa5_22min_0[1:1], fa5_22min_0[2:2], fa5_22min_0[4:4]);
  INV I596 (simp5151_0[1:1], fa5_22min_0[7:7]);
  NAND2 I597 (termt_5[22:22], simp5151_0[0:0], simp5151_0[1:1]);
  AO222 I598 (ct5__0[22:22], termt_2[22:22], termt_4[22:22], termt_2[22:22], ct5__0[21:21], termt_4[22:22], ct5__0[21:21]);
  AO222 I599 (cf5__0[22:22], termf_2[22:22], termf_4[22:22], termf_2[22:22], cf5__0[21:21], termf_4[22:22], cf5__0[21:21]);
  C3 I600 (fa5_23min_0[0:0], cf5__0[22:22], termf_4[23:23], termf_2[23:23]);
  C3 I601 (fa5_23min_0[1:1], cf5__0[22:22], termf_4[23:23], termt_2[23:23]);
  C3 I602 (fa5_23min_0[2:2], cf5__0[22:22], termt_4[23:23], termf_2[23:23]);
  C3 I603 (fa5_23min_0[3:3], cf5__0[22:22], termt_4[23:23], termt_2[23:23]);
  C3 I604 (fa5_23min_0[4:4], ct5__0[22:22], termf_4[23:23], termf_2[23:23]);
  C3 I605 (fa5_23min_0[5:5], ct5__0[22:22], termf_4[23:23], termt_2[23:23]);
  C3 I606 (fa5_23min_0[6:6], ct5__0[22:22], termt_4[23:23], termf_2[23:23]);
  C3 I607 (fa5_23min_0[7:7], ct5__0[22:22], termt_4[23:23], termt_2[23:23]);
  NOR3 I608 (simp5271_0[0:0], fa5_23min_0[0:0], fa5_23min_0[3:3], fa5_23min_0[5:5]);
  INV I609 (simp5271_0[1:1], fa5_23min_0[6:6]);
  NAND2 I610 (termf_5[23:23], simp5271_0[0:0], simp5271_0[1:1]);
  NOR3 I611 (simp5281_0[0:0], fa5_23min_0[1:1], fa5_23min_0[2:2], fa5_23min_0[4:4]);
  INV I612 (simp5281_0[1:1], fa5_23min_0[7:7]);
  NAND2 I613 (termt_5[23:23], simp5281_0[0:0], simp5281_0[1:1]);
  AO222 I614 (ct5__0[23:23], termt_2[23:23], termt_4[23:23], termt_2[23:23], ct5__0[22:22], termt_4[23:23], ct5__0[22:22]);
  AO222 I615 (cf5__0[23:23], termf_2[23:23], termf_4[23:23], termf_2[23:23], cf5__0[22:22], termf_4[23:23], cf5__0[22:22]);
  C3 I616 (fa5_24min_0[0:0], cf5__0[23:23], termf_4[24:24], termf_2[24:24]);
  C3 I617 (fa5_24min_0[1:1], cf5__0[23:23], termf_4[24:24], termt_2[24:24]);
  C3 I618 (fa5_24min_0[2:2], cf5__0[23:23], termt_4[24:24], termf_2[24:24]);
  C3 I619 (fa5_24min_0[3:3], cf5__0[23:23], termt_4[24:24], termt_2[24:24]);
  C3 I620 (fa5_24min_0[4:4], ct5__0[23:23], termf_4[24:24], termf_2[24:24]);
  C3 I621 (fa5_24min_0[5:5], ct5__0[23:23], termf_4[24:24], termt_2[24:24]);
  C3 I622 (fa5_24min_0[6:6], ct5__0[23:23], termt_4[24:24], termf_2[24:24]);
  C3 I623 (fa5_24min_0[7:7], ct5__0[23:23], termt_4[24:24], termt_2[24:24]);
  NOR3 I624 (simp5401_0[0:0], fa5_24min_0[0:0], fa5_24min_0[3:3], fa5_24min_0[5:5]);
  INV I625 (simp5401_0[1:1], fa5_24min_0[6:6]);
  NAND2 I626 (termf_5[24:24], simp5401_0[0:0], simp5401_0[1:1]);
  NOR3 I627 (simp5411_0[0:0], fa5_24min_0[1:1], fa5_24min_0[2:2], fa5_24min_0[4:4]);
  INV I628 (simp5411_0[1:1], fa5_24min_0[7:7]);
  NAND2 I629 (termt_5[24:24], simp5411_0[0:0], simp5411_0[1:1]);
  AO222 I630 (ct5__0[24:24], termt_2[24:24], termt_4[24:24], termt_2[24:24], ct5__0[23:23], termt_4[24:24], ct5__0[23:23]);
  AO222 I631 (cf5__0[24:24], termf_2[24:24], termf_4[24:24], termf_2[24:24], cf5__0[23:23], termf_4[24:24], cf5__0[23:23]);
  C3 I632 (fa5_25min_0[0:0], cf5__0[24:24], termf_4[25:25], termf_2[25:25]);
  C3 I633 (fa5_25min_0[1:1], cf5__0[24:24], termf_4[25:25], termt_2[25:25]);
  C3 I634 (fa5_25min_0[2:2], cf5__0[24:24], termt_4[25:25], termf_2[25:25]);
  C3 I635 (fa5_25min_0[3:3], cf5__0[24:24], termt_4[25:25], termt_2[25:25]);
  C3 I636 (fa5_25min_0[4:4], ct5__0[24:24], termf_4[25:25], termf_2[25:25]);
  C3 I637 (fa5_25min_0[5:5], ct5__0[24:24], termf_4[25:25], termt_2[25:25]);
  C3 I638 (fa5_25min_0[6:6], ct5__0[24:24], termt_4[25:25], termf_2[25:25]);
  C3 I639 (fa5_25min_0[7:7], ct5__0[24:24], termt_4[25:25], termt_2[25:25]);
  NOR3 I640 (simp5531_0[0:0], fa5_25min_0[0:0], fa5_25min_0[3:3], fa5_25min_0[5:5]);
  INV I641 (simp5531_0[1:1], fa5_25min_0[6:6]);
  NAND2 I642 (termf_5[25:25], simp5531_0[0:0], simp5531_0[1:1]);
  NOR3 I643 (simp5541_0[0:0], fa5_25min_0[1:1], fa5_25min_0[2:2], fa5_25min_0[4:4]);
  INV I644 (simp5541_0[1:1], fa5_25min_0[7:7]);
  NAND2 I645 (termt_5[25:25], simp5541_0[0:0], simp5541_0[1:1]);
  AO222 I646 (ct5__0[25:25], termt_2[25:25], termt_4[25:25], termt_2[25:25], ct5__0[24:24], termt_4[25:25], ct5__0[24:24]);
  AO222 I647 (cf5__0[25:25], termf_2[25:25], termf_4[25:25], termf_2[25:25], cf5__0[24:24], termf_4[25:25], cf5__0[24:24]);
  C3 I648 (fa5_26min_0[0:0], cf5__0[25:25], termf_4[26:26], termf_2[26:26]);
  C3 I649 (fa5_26min_0[1:1], cf5__0[25:25], termf_4[26:26], termt_2[26:26]);
  C3 I650 (fa5_26min_0[2:2], cf5__0[25:25], termt_4[26:26], termf_2[26:26]);
  C3 I651 (fa5_26min_0[3:3], cf5__0[25:25], termt_4[26:26], termt_2[26:26]);
  C3 I652 (fa5_26min_0[4:4], ct5__0[25:25], termf_4[26:26], termf_2[26:26]);
  C3 I653 (fa5_26min_0[5:5], ct5__0[25:25], termf_4[26:26], termt_2[26:26]);
  C3 I654 (fa5_26min_0[6:6], ct5__0[25:25], termt_4[26:26], termf_2[26:26]);
  C3 I655 (fa5_26min_0[7:7], ct5__0[25:25], termt_4[26:26], termt_2[26:26]);
  NOR3 I656 (simp5661_0[0:0], fa5_26min_0[0:0], fa5_26min_0[3:3], fa5_26min_0[5:5]);
  INV I657 (simp5661_0[1:1], fa5_26min_0[6:6]);
  NAND2 I658 (termf_5[26:26], simp5661_0[0:0], simp5661_0[1:1]);
  NOR3 I659 (simp5671_0[0:0], fa5_26min_0[1:1], fa5_26min_0[2:2], fa5_26min_0[4:4]);
  INV I660 (simp5671_0[1:1], fa5_26min_0[7:7]);
  NAND2 I661 (termt_5[26:26], simp5671_0[0:0], simp5671_0[1:1]);
  AO222 I662 (ct5__0[26:26], termt_2[26:26], termt_4[26:26], termt_2[26:26], ct5__0[25:25], termt_4[26:26], ct5__0[25:25]);
  AO222 I663 (cf5__0[26:26], termf_2[26:26], termf_4[26:26], termf_2[26:26], cf5__0[25:25], termf_4[26:26], cf5__0[25:25]);
  C3 I664 (fa5_27min_0[0:0], cf5__0[26:26], termf_4[27:27], termf_2[27:27]);
  C3 I665 (fa5_27min_0[1:1], cf5__0[26:26], termf_4[27:27], termt_2[27:27]);
  C3 I666 (fa5_27min_0[2:2], cf5__0[26:26], termt_4[27:27], termf_2[27:27]);
  C3 I667 (fa5_27min_0[3:3], cf5__0[26:26], termt_4[27:27], termt_2[27:27]);
  C3 I668 (fa5_27min_0[4:4], ct5__0[26:26], termf_4[27:27], termf_2[27:27]);
  C3 I669 (fa5_27min_0[5:5], ct5__0[26:26], termf_4[27:27], termt_2[27:27]);
  C3 I670 (fa5_27min_0[6:6], ct5__0[26:26], termt_4[27:27], termf_2[27:27]);
  C3 I671 (fa5_27min_0[7:7], ct5__0[26:26], termt_4[27:27], termt_2[27:27]);
  NOR3 I672 (simp5791_0[0:0], fa5_27min_0[0:0], fa5_27min_0[3:3], fa5_27min_0[5:5]);
  INV I673 (simp5791_0[1:1], fa5_27min_0[6:6]);
  NAND2 I674 (termf_5[27:27], simp5791_0[0:0], simp5791_0[1:1]);
  NOR3 I675 (simp5801_0[0:0], fa5_27min_0[1:1], fa5_27min_0[2:2], fa5_27min_0[4:4]);
  INV I676 (simp5801_0[1:1], fa5_27min_0[7:7]);
  NAND2 I677 (termt_5[27:27], simp5801_0[0:0], simp5801_0[1:1]);
  AO222 I678 (ct5__0[27:27], termt_2[27:27], termt_4[27:27], termt_2[27:27], ct5__0[26:26], termt_4[27:27], ct5__0[26:26]);
  AO222 I679 (cf5__0[27:27], termf_2[27:27], termf_4[27:27], termf_2[27:27], cf5__0[26:26], termf_4[27:27], cf5__0[26:26]);
  C3 I680 (fa5_28min_0[0:0], cf5__0[27:27], termf_4[28:28], termf_2[28:28]);
  C3 I681 (fa5_28min_0[1:1], cf5__0[27:27], termf_4[28:28], termt_2[28:28]);
  C3 I682 (fa5_28min_0[2:2], cf5__0[27:27], termt_4[28:28], termf_2[28:28]);
  C3 I683 (fa5_28min_0[3:3], cf5__0[27:27], termt_4[28:28], termt_2[28:28]);
  C3 I684 (fa5_28min_0[4:4], ct5__0[27:27], termf_4[28:28], termf_2[28:28]);
  C3 I685 (fa5_28min_0[5:5], ct5__0[27:27], termf_4[28:28], termt_2[28:28]);
  C3 I686 (fa5_28min_0[6:6], ct5__0[27:27], termt_4[28:28], termf_2[28:28]);
  C3 I687 (fa5_28min_0[7:7], ct5__0[27:27], termt_4[28:28], termt_2[28:28]);
  NOR3 I688 (simp5921_0[0:0], fa5_28min_0[0:0], fa5_28min_0[3:3], fa5_28min_0[5:5]);
  INV I689 (simp5921_0[1:1], fa5_28min_0[6:6]);
  NAND2 I690 (termf_5[28:28], simp5921_0[0:0], simp5921_0[1:1]);
  NOR3 I691 (simp5931_0[0:0], fa5_28min_0[1:1], fa5_28min_0[2:2], fa5_28min_0[4:4]);
  INV I692 (simp5931_0[1:1], fa5_28min_0[7:7]);
  NAND2 I693 (termt_5[28:28], simp5931_0[0:0], simp5931_0[1:1]);
  AO222 I694 (ct5__0[28:28], termt_2[28:28], termt_4[28:28], termt_2[28:28], ct5__0[27:27], termt_4[28:28], ct5__0[27:27]);
  AO222 I695 (cf5__0[28:28], termf_2[28:28], termf_4[28:28], termf_2[28:28], cf5__0[27:27], termf_4[28:28], cf5__0[27:27]);
  C3 I696 (fa5_29min_0[0:0], cf5__0[28:28], termf_4[29:29], termf_2[29:29]);
  C3 I697 (fa5_29min_0[1:1], cf5__0[28:28], termf_4[29:29], termt_2[29:29]);
  C3 I698 (fa5_29min_0[2:2], cf5__0[28:28], termt_4[29:29], termf_2[29:29]);
  C3 I699 (fa5_29min_0[3:3], cf5__0[28:28], termt_4[29:29], termt_2[29:29]);
  C3 I700 (fa5_29min_0[4:4], ct5__0[28:28], termf_4[29:29], termf_2[29:29]);
  C3 I701 (fa5_29min_0[5:5], ct5__0[28:28], termf_4[29:29], termt_2[29:29]);
  C3 I702 (fa5_29min_0[6:6], ct5__0[28:28], termt_4[29:29], termf_2[29:29]);
  C3 I703 (fa5_29min_0[7:7], ct5__0[28:28], termt_4[29:29], termt_2[29:29]);
  NOR3 I704 (simp6051_0[0:0], fa5_29min_0[0:0], fa5_29min_0[3:3], fa5_29min_0[5:5]);
  INV I705 (simp6051_0[1:1], fa5_29min_0[6:6]);
  NAND2 I706 (termf_5[29:29], simp6051_0[0:0], simp6051_0[1:1]);
  NOR3 I707 (simp6061_0[0:0], fa5_29min_0[1:1], fa5_29min_0[2:2], fa5_29min_0[4:4]);
  INV I708 (simp6061_0[1:1], fa5_29min_0[7:7]);
  NAND2 I709 (termt_5[29:29], simp6061_0[0:0], simp6061_0[1:1]);
  AO222 I710 (ct5__0[29:29], termt_2[29:29], termt_4[29:29], termt_2[29:29], ct5__0[28:28], termt_4[29:29], ct5__0[28:28]);
  AO222 I711 (cf5__0[29:29], termf_2[29:29], termf_4[29:29], termf_2[29:29], cf5__0[28:28], termf_4[29:29], cf5__0[28:28]);
  C3 I712 (fa5_30min_0[0:0], cf5__0[29:29], termf_4[30:30], termf_2[30:30]);
  C3 I713 (fa5_30min_0[1:1], cf5__0[29:29], termf_4[30:30], termt_2[30:30]);
  C3 I714 (fa5_30min_0[2:2], cf5__0[29:29], termt_4[30:30], termf_2[30:30]);
  C3 I715 (fa5_30min_0[3:3], cf5__0[29:29], termt_4[30:30], termt_2[30:30]);
  C3 I716 (fa5_30min_0[4:4], ct5__0[29:29], termf_4[30:30], termf_2[30:30]);
  C3 I717 (fa5_30min_0[5:5], ct5__0[29:29], termf_4[30:30], termt_2[30:30]);
  C3 I718 (fa5_30min_0[6:6], ct5__0[29:29], termt_4[30:30], termf_2[30:30]);
  C3 I719 (fa5_30min_0[7:7], ct5__0[29:29], termt_4[30:30], termt_2[30:30]);
  NOR3 I720 (simp6181_0[0:0], fa5_30min_0[0:0], fa5_30min_0[3:3], fa5_30min_0[5:5]);
  INV I721 (simp6181_0[1:1], fa5_30min_0[6:6]);
  NAND2 I722 (termf_5[30:30], simp6181_0[0:0], simp6181_0[1:1]);
  NOR3 I723 (simp6191_0[0:0], fa5_30min_0[1:1], fa5_30min_0[2:2], fa5_30min_0[4:4]);
  INV I724 (simp6191_0[1:1], fa5_30min_0[7:7]);
  NAND2 I725 (termt_5[30:30], simp6191_0[0:0], simp6191_0[1:1]);
  AO222 I726 (ct5__0[30:30], termt_2[30:30], termt_4[30:30], termt_2[30:30], ct5__0[29:29], termt_4[30:30], ct5__0[29:29]);
  AO222 I727 (cf5__0[30:30], termf_2[30:30], termf_4[30:30], termf_2[30:30], cf5__0[29:29], termf_4[30:30], cf5__0[29:29]);
  C3 I728 (fa5_31min_0[0:0], cf5__0[30:30], termf_4[31:31], termf_2[31:31]);
  C3 I729 (fa5_31min_0[1:1], cf5__0[30:30], termf_4[31:31], termt_2[31:31]);
  C3 I730 (fa5_31min_0[2:2], cf5__0[30:30], termt_4[31:31], termf_2[31:31]);
  C3 I731 (fa5_31min_0[3:3], cf5__0[30:30], termt_4[31:31], termt_2[31:31]);
  C3 I732 (fa5_31min_0[4:4], ct5__0[30:30], termf_4[31:31], termf_2[31:31]);
  C3 I733 (fa5_31min_0[5:5], ct5__0[30:30], termf_4[31:31], termt_2[31:31]);
  C3 I734 (fa5_31min_0[6:6], ct5__0[30:30], termt_4[31:31], termf_2[31:31]);
  C3 I735 (fa5_31min_0[7:7], ct5__0[30:30], termt_4[31:31], termt_2[31:31]);
  NOR3 I736 (simp6311_0[0:0], fa5_31min_0[0:0], fa5_31min_0[3:3], fa5_31min_0[5:5]);
  INV I737 (simp6311_0[1:1], fa5_31min_0[6:6]);
  NAND2 I738 (termf_5[31:31], simp6311_0[0:0], simp6311_0[1:1]);
  NOR3 I739 (simp6321_0[0:0], fa5_31min_0[1:1], fa5_31min_0[2:2], fa5_31min_0[4:4]);
  INV I740 (simp6321_0[1:1], fa5_31min_0[7:7]);
  NAND2 I741 (termt_5[31:31], simp6321_0[0:0], simp6321_0[1:1]);
  AO222 I742 (ct5__0[31:31], termt_2[31:31], termt_4[31:31], termt_2[31:31], ct5__0[30:30], termt_4[31:31], ct5__0[30:30]);
  AO222 I743 (cf5__0[31:31], termf_2[31:31], termf_4[31:31], termf_2[31:31], cf5__0[30:30], termf_4[31:31], cf5__0[30:30]);
  C3 I744 (fa5_32min_0[0:0], cf5__0[31:31], termf_4[32:32], termf_2[32:32]);
  C3 I745 (fa5_32min_0[1:1], cf5__0[31:31], termf_4[32:32], termt_2[32:32]);
  C3 I746 (fa5_32min_0[2:2], cf5__0[31:31], termt_4[32:32], termf_2[32:32]);
  C3 I747 (fa5_32min_0[3:3], cf5__0[31:31], termt_4[32:32], termt_2[32:32]);
  C3 I748 (fa5_32min_0[4:4], ct5__0[31:31], termf_4[32:32], termf_2[32:32]);
  C3 I749 (fa5_32min_0[5:5], ct5__0[31:31], termf_4[32:32], termt_2[32:32]);
  C3 I750 (fa5_32min_0[6:6], ct5__0[31:31], termt_4[32:32], termf_2[32:32]);
  C3 I751 (fa5_32min_0[7:7], ct5__0[31:31], termt_4[32:32], termt_2[32:32]);
  NOR3 I752 (simp6441_0[0:0], fa5_32min_0[0:0], fa5_32min_0[3:3], fa5_32min_0[5:5]);
  INV I753 (simp6441_0[1:1], fa5_32min_0[6:6]);
  NAND2 I754 (termf_5[32:32], simp6441_0[0:0], simp6441_0[1:1]);
  NOR3 I755 (simp6451_0[0:0], fa5_32min_0[1:1], fa5_32min_0[2:2], fa5_32min_0[4:4]);
  INV I756 (simp6451_0[1:1], fa5_32min_0[7:7]);
  NAND2 I757 (termt_5[32:32], simp6451_0[0:0], simp6451_0[1:1]);
  AO222 I758 (ct5__0[32:32], termt_2[32:32], termt_4[32:32], termt_2[32:32], ct5__0[31:31], termt_4[32:32], ct5__0[31:31]);
  AO222 I759 (cf5__0[32:32], termf_2[32:32], termf_4[32:32], termf_2[32:32], cf5__0[31:31], termf_4[32:32], cf5__0[31:31]);
  C3 I760 (fa5_33min_0[0:0], cf5__0[32:32], termf_4[33:33], termf_2[33:33]);
  C3 I761 (fa5_33min_0[1:1], cf5__0[32:32], termf_4[33:33], termt_2[33:33]);
  C3 I762 (fa5_33min_0[2:2], cf5__0[32:32], termt_4[33:33], termf_2[33:33]);
  C3 I763 (fa5_33min_0[3:3], cf5__0[32:32], termt_4[33:33], termt_2[33:33]);
  C3 I764 (fa5_33min_0[4:4], ct5__0[32:32], termf_4[33:33], termf_2[33:33]);
  C3 I765 (fa5_33min_0[5:5], ct5__0[32:32], termf_4[33:33], termt_2[33:33]);
  C3 I766 (fa5_33min_0[6:6], ct5__0[32:32], termt_4[33:33], termf_2[33:33]);
  C3 I767 (fa5_33min_0[7:7], ct5__0[32:32], termt_4[33:33], termt_2[33:33]);
  NOR3 I768 (simp6571_0[0:0], fa5_33min_0[0:0], fa5_33min_0[3:3], fa5_33min_0[5:5]);
  INV I769 (simp6571_0[1:1], fa5_33min_0[6:6]);
  NAND2 I770 (termf_5[33:33], simp6571_0[0:0], simp6571_0[1:1]);
  NOR3 I771 (simp6581_0[0:0], fa5_33min_0[1:1], fa5_33min_0[2:2], fa5_33min_0[4:4]);
  INV I772 (simp6581_0[1:1], fa5_33min_0[7:7]);
  NAND2 I773 (termt_5[33:33], simp6581_0[0:0], simp6581_0[1:1]);
  AO222 I774 (ct5__0[33:33], termt_2[33:33], termt_4[33:33], termt_2[33:33], ct5__0[32:32], termt_4[33:33], ct5__0[32:32]);
  AO222 I775 (cf5__0[33:33], termf_2[33:33], termf_4[33:33], termf_2[33:33], cf5__0[32:32], termf_4[33:33], cf5__0[32:32]);
  BUFF I776 (o_0r0[0:0], termf_5[1:1]);
  BUFF I777 (o_0r0[1:1], termf_5[2:2]);
  BUFF I778 (o_0r0[2:2], termf_5[3:3]);
  BUFF I779 (o_0r0[3:3], termf_5[4:4]);
  BUFF I780 (o_0r0[4:4], termf_5[5:5]);
  BUFF I781 (o_0r0[5:5], termf_5[6:6]);
  BUFF I782 (o_0r0[6:6], termf_5[7:7]);
  BUFF I783 (o_0r0[7:7], termf_5[8:8]);
  BUFF I784 (o_0r0[8:8], termf_5[9:9]);
  BUFF I785 (o_0r0[9:9], termf_5[10:10]);
  BUFF I786 (o_0r0[10:10], termf_5[11:11]);
  BUFF I787 (o_0r0[11:11], termf_5[12:12]);
  BUFF I788 (o_0r0[12:12], termf_5[13:13]);
  BUFF I789 (o_0r0[13:13], termf_5[14:14]);
  BUFF I790 (o_0r0[14:14], termf_5[15:15]);
  BUFF I791 (o_0r0[15:15], termf_5[16:16]);
  BUFF I792 (o_0r0[16:16], termf_5[17:17]);
  BUFF I793 (o_0r0[17:17], termf_5[18:18]);
  BUFF I794 (o_0r0[18:18], termf_5[19:19]);
  BUFF I795 (o_0r0[19:19], termf_5[20:20]);
  BUFF I796 (o_0r0[20:20], termf_5[21:21]);
  BUFF I797 (o_0r0[21:21], termf_5[22:22]);
  BUFF I798 (o_0r0[22:22], termf_5[23:23]);
  BUFF I799 (o_0r0[23:23], termf_5[24:24]);
  BUFF I800 (o_0r0[24:24], termf_5[25:25]);
  BUFF I801 (o_0r0[25:25], termf_5[26:26]);
  BUFF I802 (o_0r0[26:26], termf_5[27:27]);
  BUFF I803 (o_0r0[27:27], termf_5[28:28]);
  BUFF I804 (o_0r0[28:28], termf_5[29:29]);
  BUFF I805 (o_0r0[29:29], termf_5[30:30]);
  BUFF I806 (o_0r0[30:30], termf_5[31:31]);
  BUFF I807 (o_0r0[31:31], termf_5[32:32]);
  BUFF I808 (o_0r0[32:32], termf_5[33:33]);
  BUFF I809 (o_0r1[0:0], termt_5[1:1]);
  BUFF I810 (o_0r1[1:1], termt_5[2:2]);
  BUFF I811 (o_0r1[2:2], termt_5[3:3]);
  BUFF I812 (o_0r1[3:3], termt_5[4:4]);
  BUFF I813 (o_0r1[4:4], termt_5[5:5]);
  BUFF I814 (o_0r1[5:5], termt_5[6:6]);
  BUFF I815 (o_0r1[6:6], termt_5[7:7]);
  BUFF I816 (o_0r1[7:7], termt_5[8:8]);
  BUFF I817 (o_0r1[8:8], termt_5[9:9]);
  BUFF I818 (o_0r1[9:9], termt_5[10:10]);
  BUFF I819 (o_0r1[10:10], termt_5[11:11]);
  BUFF I820 (o_0r1[11:11], termt_5[12:12]);
  BUFF I821 (o_0r1[12:12], termt_5[13:13]);
  BUFF I822 (o_0r1[13:13], termt_5[14:14]);
  BUFF I823 (o_0r1[14:14], termt_5[15:15]);
  BUFF I824 (o_0r1[15:15], termt_5[16:16]);
  BUFF I825 (o_0r1[16:16], termt_5[17:17]);
  BUFF I826 (o_0r1[17:17], termt_5[18:18]);
  BUFF I827 (o_0r1[18:18], termt_5[19:19]);
  BUFF I828 (o_0r1[19:19], termt_5[20:20]);
  BUFF I829 (o_0r1[20:20], termt_5[21:21]);
  BUFF I830 (o_0r1[21:21], termt_5[22:22]);
  BUFF I831 (o_0r1[22:22], termt_5[23:23]);
  BUFF I832 (o_0r1[23:23], termt_5[24:24]);
  BUFF I833 (o_0r1[24:24], termt_5[25:25]);
  BUFF I834 (o_0r1[25:25], termt_5[26:26]);
  BUFF I835 (o_0r1[26:26], termt_5[27:27]);
  BUFF I836 (o_0r1[27:27], termt_5[28:28]);
  BUFF I837 (o_0r1[28:28], termt_5[29:29]);
  BUFF I838 (o_0r1[29:29], termt_5[30:30]);
  BUFF I839 (o_0r1[30:30], termt_5[31:31]);
  BUFF I840 (o_0r1[31:31], termt_5[32:32]);
  BUFF I841 (o_0r1[32:32], termt_5[33:33]);
  BUFF I842 (i_0a, o_0a);
endmodule

// tkj69m32_4_32_1 TeakJ [Many [32,4,32,1],One 69]
module tkj69m32_4_32_1 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [3:0] i_1r0;
  input [3:0] i_1r1;
  output i_1a;
  input [31:0] i_2r0;
  input [31:0] i_2r1;
  output i_2a;
  input i_3r0;
  input i_3r1;
  output i_3a;
  output [68:0] o_0r0;
  output [68:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r0[0:0]);
  BUFF I1 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I2 (o_0r0[2:2], i_0r0[2:2]);
  BUFF I3 (o_0r0[3:3], i_0r0[3:3]);
  BUFF I4 (o_0r0[4:4], i_0r0[4:4]);
  BUFF I5 (o_0r0[5:5], i_0r0[5:5]);
  BUFF I6 (o_0r0[6:6], i_0r0[6:6]);
  BUFF I7 (o_0r0[7:7], i_0r0[7:7]);
  BUFF I8 (o_0r0[8:8], i_0r0[8:8]);
  BUFF I9 (o_0r0[9:9], i_0r0[9:9]);
  BUFF I10 (o_0r0[10:10], i_0r0[10:10]);
  BUFF I11 (o_0r0[11:11], i_0r0[11:11]);
  BUFF I12 (o_0r0[12:12], i_0r0[12:12]);
  BUFF I13 (o_0r0[13:13], i_0r0[13:13]);
  BUFF I14 (o_0r0[14:14], i_0r0[14:14]);
  BUFF I15 (o_0r0[15:15], i_0r0[15:15]);
  BUFF I16 (o_0r0[16:16], i_0r0[16:16]);
  BUFF I17 (o_0r0[17:17], i_0r0[17:17]);
  BUFF I18 (o_0r0[18:18], i_0r0[18:18]);
  BUFF I19 (o_0r0[19:19], i_0r0[19:19]);
  BUFF I20 (o_0r0[20:20], i_0r0[20:20]);
  BUFF I21 (o_0r0[21:21], i_0r0[21:21]);
  BUFF I22 (o_0r0[22:22], i_0r0[22:22]);
  BUFF I23 (o_0r0[23:23], i_0r0[23:23]);
  BUFF I24 (o_0r0[24:24], i_0r0[24:24]);
  BUFF I25 (o_0r0[25:25], i_0r0[25:25]);
  BUFF I26 (o_0r0[26:26], i_0r0[26:26]);
  BUFF I27 (o_0r0[27:27], i_0r0[27:27]);
  BUFF I28 (o_0r0[28:28], i_0r0[28:28]);
  BUFF I29 (o_0r0[29:29], i_0r0[29:29]);
  BUFF I30 (o_0r0[30:30], i_0r0[30:30]);
  BUFF I31 (o_0r0[31:31], i_0r0[31:31]);
  BUFF I32 (o_0r0[32:32], i_1r0[0:0]);
  BUFF I33 (o_0r0[33:33], i_1r0[1:1]);
  BUFF I34 (o_0r0[34:34], i_1r0[2:2]);
  BUFF I35 (o_0r0[35:35], i_1r0[3:3]);
  BUFF I36 (o_0r0[36:36], i_2r0[0:0]);
  BUFF I37 (o_0r0[37:37], i_2r0[1:1]);
  BUFF I38 (o_0r0[38:38], i_2r0[2:2]);
  BUFF I39 (o_0r0[39:39], i_2r0[3:3]);
  BUFF I40 (o_0r0[40:40], i_2r0[4:4]);
  BUFF I41 (o_0r0[41:41], i_2r0[5:5]);
  BUFF I42 (o_0r0[42:42], i_2r0[6:6]);
  BUFF I43 (o_0r0[43:43], i_2r0[7:7]);
  BUFF I44 (o_0r0[44:44], i_2r0[8:8]);
  BUFF I45 (o_0r0[45:45], i_2r0[9:9]);
  BUFF I46 (o_0r0[46:46], i_2r0[10:10]);
  BUFF I47 (o_0r0[47:47], i_2r0[11:11]);
  BUFF I48 (o_0r0[48:48], i_2r0[12:12]);
  BUFF I49 (o_0r0[49:49], i_2r0[13:13]);
  BUFF I50 (o_0r0[50:50], i_2r0[14:14]);
  BUFF I51 (o_0r0[51:51], i_2r0[15:15]);
  BUFF I52 (o_0r0[52:52], i_2r0[16:16]);
  BUFF I53 (o_0r0[53:53], i_2r0[17:17]);
  BUFF I54 (o_0r0[54:54], i_2r0[18:18]);
  BUFF I55 (o_0r0[55:55], i_2r0[19:19]);
  BUFF I56 (o_0r0[56:56], i_2r0[20:20]);
  BUFF I57 (o_0r0[57:57], i_2r0[21:21]);
  BUFF I58 (o_0r0[58:58], i_2r0[22:22]);
  BUFF I59 (o_0r0[59:59], i_2r0[23:23]);
  BUFF I60 (o_0r0[60:60], i_2r0[24:24]);
  BUFF I61 (o_0r0[61:61], i_2r0[25:25]);
  BUFF I62 (o_0r0[62:62], i_2r0[26:26]);
  BUFF I63 (o_0r0[63:63], i_2r0[27:27]);
  BUFF I64 (o_0r0[64:64], i_2r0[28:28]);
  BUFF I65 (o_0r0[65:65], i_2r0[29:29]);
  BUFF I66 (o_0r0[66:66], i_2r0[30:30]);
  BUFF I67 (o_0r0[67:67], i_2r0[31:31]);
  BUFF I68 (o_0r0[68:68], i_3r0);
  BUFF I69 (o_0r1[0:0], i_0r1[0:0]);
  BUFF I70 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I71 (o_0r1[2:2], i_0r1[2:2]);
  BUFF I72 (o_0r1[3:3], i_0r1[3:3]);
  BUFF I73 (o_0r1[4:4], i_0r1[4:4]);
  BUFF I74 (o_0r1[5:5], i_0r1[5:5]);
  BUFF I75 (o_0r1[6:6], i_0r1[6:6]);
  BUFF I76 (o_0r1[7:7], i_0r1[7:7]);
  BUFF I77 (o_0r1[8:8], i_0r1[8:8]);
  BUFF I78 (o_0r1[9:9], i_0r1[9:9]);
  BUFF I79 (o_0r1[10:10], i_0r1[10:10]);
  BUFF I80 (o_0r1[11:11], i_0r1[11:11]);
  BUFF I81 (o_0r1[12:12], i_0r1[12:12]);
  BUFF I82 (o_0r1[13:13], i_0r1[13:13]);
  BUFF I83 (o_0r1[14:14], i_0r1[14:14]);
  BUFF I84 (o_0r1[15:15], i_0r1[15:15]);
  BUFF I85 (o_0r1[16:16], i_0r1[16:16]);
  BUFF I86 (o_0r1[17:17], i_0r1[17:17]);
  BUFF I87 (o_0r1[18:18], i_0r1[18:18]);
  BUFF I88 (o_0r1[19:19], i_0r1[19:19]);
  BUFF I89 (o_0r1[20:20], i_0r1[20:20]);
  BUFF I90 (o_0r1[21:21], i_0r1[21:21]);
  BUFF I91 (o_0r1[22:22], i_0r1[22:22]);
  BUFF I92 (o_0r1[23:23], i_0r1[23:23]);
  BUFF I93 (o_0r1[24:24], i_0r1[24:24]);
  BUFF I94 (o_0r1[25:25], i_0r1[25:25]);
  BUFF I95 (o_0r1[26:26], i_0r1[26:26]);
  BUFF I96 (o_0r1[27:27], i_0r1[27:27]);
  BUFF I97 (o_0r1[28:28], i_0r1[28:28]);
  BUFF I98 (o_0r1[29:29], i_0r1[29:29]);
  BUFF I99 (o_0r1[30:30], i_0r1[30:30]);
  BUFF I100 (o_0r1[31:31], i_0r1[31:31]);
  BUFF I101 (o_0r1[32:32], i_1r1[0:0]);
  BUFF I102 (o_0r1[33:33], i_1r1[1:1]);
  BUFF I103 (o_0r1[34:34], i_1r1[2:2]);
  BUFF I104 (o_0r1[35:35], i_1r1[3:3]);
  BUFF I105 (o_0r1[36:36], i_2r1[0:0]);
  BUFF I106 (o_0r1[37:37], i_2r1[1:1]);
  BUFF I107 (o_0r1[38:38], i_2r1[2:2]);
  BUFF I108 (o_0r1[39:39], i_2r1[3:3]);
  BUFF I109 (o_0r1[40:40], i_2r1[4:4]);
  BUFF I110 (o_0r1[41:41], i_2r1[5:5]);
  BUFF I111 (o_0r1[42:42], i_2r1[6:6]);
  BUFF I112 (o_0r1[43:43], i_2r1[7:7]);
  BUFF I113 (o_0r1[44:44], i_2r1[8:8]);
  BUFF I114 (o_0r1[45:45], i_2r1[9:9]);
  BUFF I115 (o_0r1[46:46], i_2r1[10:10]);
  BUFF I116 (o_0r1[47:47], i_2r1[11:11]);
  BUFF I117 (o_0r1[48:48], i_2r1[12:12]);
  BUFF I118 (o_0r1[49:49], i_2r1[13:13]);
  BUFF I119 (o_0r1[50:50], i_2r1[14:14]);
  BUFF I120 (o_0r1[51:51], i_2r1[15:15]);
  BUFF I121 (o_0r1[52:52], i_2r1[16:16]);
  BUFF I122 (o_0r1[53:53], i_2r1[17:17]);
  BUFF I123 (o_0r1[54:54], i_2r1[18:18]);
  BUFF I124 (o_0r1[55:55], i_2r1[19:19]);
  BUFF I125 (o_0r1[56:56], i_2r1[20:20]);
  BUFF I126 (o_0r1[57:57], i_2r1[21:21]);
  BUFF I127 (o_0r1[58:58], i_2r1[22:22]);
  BUFF I128 (o_0r1[59:59], i_2r1[23:23]);
  BUFF I129 (o_0r1[60:60], i_2r1[24:24]);
  BUFF I130 (o_0r1[61:61], i_2r1[25:25]);
  BUFF I131 (o_0r1[62:62], i_2r1[26:26]);
  BUFF I132 (o_0r1[63:63], i_2r1[27:27]);
  BUFF I133 (o_0r1[64:64], i_2r1[28:28]);
  BUFF I134 (o_0r1[65:65], i_2r1[29:29]);
  BUFF I135 (o_0r1[66:66], i_2r1[30:30]);
  BUFF I136 (o_0r1[67:67], i_2r1[31:31]);
  BUFF I137 (o_0r1[68:68], i_3r1);
  BUFF I138 (i_0a, o_0a);
  BUFF I139 (i_1a, o_0a);
  BUFF I140 (i_2a, o_0a);
  BUFF I141 (i_3a, o_0a);
endmodule

// tko33m4_1api0w2bi0w2b TeakO [
//     (1,TeakOAppend 1 [(0,0,2),(0,0,2)])] [One 33,One 4]
module tko33m4_1api0w2bi0w2b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [32:0] i_0r0;
  input [32:0] i_0r1;
  output i_0a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r0[0:0]);
  BUFF I1 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I2 (o_0r0[2:2], i_0r0[0:0]);
  BUFF I3 (o_0r0[3:3], i_0r0[1:1]);
  BUFF I4 (o_0r1[0:0], i_0r1[0:0]);
  BUFF I5 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I6 (o_0r1[2:2], i_0r1[0:0]);
  BUFF I7 (o_0r1[3:3], i_0r1[1:1]);
  BUFF I8 (i_0a, o_0a);
endmodule

// tko69m65_1nm2b1_2nm2b2_3mx0m12o1m12o3m8o7_2o6o10o14o15_i32w4bt1o0w2bt2o0w2b_4nm2b1_5nm2b2_6mx0m14o1m
//   12o11o15_3o7_i32w4bt4o0w2bt5o0w2b_7noti36w32b_8mx2_1_t3o0w2bt7o0w32bi36w32b_9noti0w32b_10mx2_1_t6o0w
//   2bt9o0w32bi0w32b_11apt10o0w32bt8o0w32bi68w1b TeakO [
//     (1,TeakOConstant 2 1),
//     (2,TeakOConstant 2 2),
//     (3,TeakOMux [[Imp 0 12,Imp 1 12,Imp 3 8,Imp 7 0],[Imp 2 0,Imp 6 0,Imp 10 0,Imp 14 0,Imp 15 0]] [(0
//   ,32,4),(1,0,2),(2,0,2)]),
//     (4,TeakOConstant 2 1),
//     (5,TeakOConstant 2 2),
//     (6,TeakOMux [[Imp 0 14,Imp 1 12,Imp 11 0,Imp 15 0],[Imp 3 0,Imp 7 0]] [(0,32,4),(4,0,2),(5,0,2)]),
//     (7,TeakOp TeakOpNot [(0,36,32)]),
//     (8,TeakOMux [[Imp 2 0],[Imp 1 0]] [(3,0,2),(7,0,32),(0,36,32)]),
//     (9,TeakOp TeakOpNot [(0,0,32)]),
//     (10,TeakOMux [[Imp 2 0],[Imp 1 0]] [(6,0,2),(9,0,32),(0,0,32)]),
//     (11,TeakOAppend 1 [(10,0,32),(8,0,32),(0,68,1)])] [One 69,One 65]
module tko69m65_1nm2b1_2nm2b2_3mx0m12o1m12o3m8o7_2o6o10o14o15_i32w4bt1o0w2bt2o0w2b_4nm2b1_5nm2b2_6mx0m14o1m12o11o15_3o7_i32w4bt4o0w2bt5o0w2b_7noti36w32b_8mx2_1_t3o0w2bt7o0w32bi36w32b_9noti0w32b_10mx2_1_t6o0w2bt9o0w32bi0w32b_11apt10o0w32bt8o0w32bi68w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [68:0] i_0r0;
  input [68:0] i_0r1;
  output i_0a;
  output [64:0] o_0r0;
  output [64:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [68:0] gocomp_0;
  wire [22:0] simp711_0;
  wire [7:0] simp712_0;
  wire [2:0] simp713_0;
  wire [1:0] termf_1;
  wire [1:0] termf_2;
  wire [1:0] termf_3;
  wire [1:0] termf_4;
  wire [1:0] termf_5;
  wire [1:0] termf_6;
  wire [31:0] termf_7;
  wire [31:0] termf_8;
  wire [31:0] termf_9;
  wire [31:0] termf_10;
  wire [1:0] termt_1;
  wire [1:0] termt_2;
  wire [1:0] termt_3;
  wire [1:0] termt_4;
  wire [1:0] termt_5;
  wire [1:0] termt_6;
  wire [31:0] termt_7;
  wire [31:0] termt_8;
  wire [31:0] termt_9;
  wire [31:0] termt_10;
  wire [1:0] gfint3_0;
  wire [1:0] gfint3_1;
  wire [1:0] gtint3_0;
  wire [1:0] gtint3_1;
  wire selcomp3_0;
  wire selcomp3_1;
  wire sel3_0;
  wire sel3_1;
  wire selg3_0;
  wire selg3_1;
  wire icomplete3_0;
  wire scomplete3_0;
  wire [1:0] comp30_0;
  wire [1:0] comp31_0;
  wire [3:0] dcomp3_0;
  wire [1:0] simp1251_0;
  wire [3:0] match30_0;
  wire [1:0] simp1421_0;
  wire [1:0] simp1461_0;
  wire [4:0] match31_0;
  wire [1:0] simp1481_0;
  wire [1:0] simp1491_0;
  wire [1:0] simp1501_0;
  wire [1:0] simp1511_0;
  wire [1:0] simp1521_0;
  wire [1:0] simp1531_0;
  wire [1:0] gfint6_0;
  wire [1:0] gfint6_1;
  wire [1:0] gtint6_0;
  wire [1:0] gtint6_1;
  wire selcomp6_0;
  wire selcomp6_1;
  wire sel6_0;
  wire sel6_1;
  wire selg6_0;
  wire selg6_1;
  wire icomplete6_0;
  wire scomplete6_0;
  wire [1:0] comp60_0;
  wire [1:0] comp61_0;
  wire [3:0] dcomp6_0;
  wire [1:0] simp1871_0;
  wire [3:0] match60_0;
  wire [1:0] simp2041_0;
  wire [1:0] simp2071_0;
  wire [1:0] simp2081_0;
  wire [1:0] match61_0;
  wire [1:0] simp2111_0;
  wire [1:0] simp2121_0;
  wire [31:0] gfint8_0;
  wire [31:0] gfint8_1;
  wire [31:0] gtint8_0;
  wire [31:0] gtint8_1;
  wire selcomp8_0;
  wire selcomp8_1;
  wire sel8_0;
  wire sel8_1;
  wire selg8_0;
  wire selg8_1;
  wire icomplete8_0;
  wire scomplete8_0;
  wire [31:0] comp80_0;
  wire [10:0] simp3221_0;
  wire [3:0] simp3222_0;
  wire [1:0] simp3223_0;
  wire [31:0] comp81_0;
  wire [10:0] simp3561_0;
  wire [3:0] simp3562_0;
  wire [1:0] simp3563_0;
  wire [1:0] dcomp8_0;
  wire match80_0;
  wire match81_0;
  wire [31:0] gfint10_0;
  wire [31:0] gfint10_1;
  wire [31:0] gtint10_0;
  wire [31:0] gtint10_1;
  wire selcomp10_0;
  wire selcomp10_1;
  wire sel10_0;
  wire sel10_1;
  wire selg10_0;
  wire selg10_1;
  wire icomplete10_0;
  wire scomplete10_0;
  wire [31:0] comp100_0;
  wire [10:0] simp6711_0;
  wire [3:0] simp6712_0;
  wire [1:0] simp6713_0;
  wire [31:0] comp101_0;
  wire [10:0] simp7051_0;
  wire [3:0] simp7052_0;
  wire [1:0] simp7053_0;
  wire [1:0] dcomp10_0;
  wire match100_0;
  wire match101_0;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I30 (gocomp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I31 (gocomp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I32 (gocomp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  OR2 I33 (gocomp_0[33:33], i_0r0[33:33], i_0r1[33:33]);
  OR2 I34 (gocomp_0[34:34], i_0r0[34:34], i_0r1[34:34]);
  OR2 I35 (gocomp_0[35:35], i_0r0[35:35], i_0r1[35:35]);
  OR2 I36 (gocomp_0[36:36], i_0r0[36:36], i_0r1[36:36]);
  OR2 I37 (gocomp_0[37:37], i_0r0[37:37], i_0r1[37:37]);
  OR2 I38 (gocomp_0[38:38], i_0r0[38:38], i_0r1[38:38]);
  OR2 I39 (gocomp_0[39:39], i_0r0[39:39], i_0r1[39:39]);
  OR2 I40 (gocomp_0[40:40], i_0r0[40:40], i_0r1[40:40]);
  OR2 I41 (gocomp_0[41:41], i_0r0[41:41], i_0r1[41:41]);
  OR2 I42 (gocomp_0[42:42], i_0r0[42:42], i_0r1[42:42]);
  OR2 I43 (gocomp_0[43:43], i_0r0[43:43], i_0r1[43:43]);
  OR2 I44 (gocomp_0[44:44], i_0r0[44:44], i_0r1[44:44]);
  OR2 I45 (gocomp_0[45:45], i_0r0[45:45], i_0r1[45:45]);
  OR2 I46 (gocomp_0[46:46], i_0r0[46:46], i_0r1[46:46]);
  OR2 I47 (gocomp_0[47:47], i_0r0[47:47], i_0r1[47:47]);
  OR2 I48 (gocomp_0[48:48], i_0r0[48:48], i_0r1[48:48]);
  OR2 I49 (gocomp_0[49:49], i_0r0[49:49], i_0r1[49:49]);
  OR2 I50 (gocomp_0[50:50], i_0r0[50:50], i_0r1[50:50]);
  OR2 I51 (gocomp_0[51:51], i_0r0[51:51], i_0r1[51:51]);
  OR2 I52 (gocomp_0[52:52], i_0r0[52:52], i_0r1[52:52]);
  OR2 I53 (gocomp_0[53:53], i_0r0[53:53], i_0r1[53:53]);
  OR2 I54 (gocomp_0[54:54], i_0r0[54:54], i_0r1[54:54]);
  OR2 I55 (gocomp_0[55:55], i_0r0[55:55], i_0r1[55:55]);
  OR2 I56 (gocomp_0[56:56], i_0r0[56:56], i_0r1[56:56]);
  OR2 I57 (gocomp_0[57:57], i_0r0[57:57], i_0r1[57:57]);
  OR2 I58 (gocomp_0[58:58], i_0r0[58:58], i_0r1[58:58]);
  OR2 I59 (gocomp_0[59:59], i_0r0[59:59], i_0r1[59:59]);
  OR2 I60 (gocomp_0[60:60], i_0r0[60:60], i_0r1[60:60]);
  OR2 I61 (gocomp_0[61:61], i_0r0[61:61], i_0r1[61:61]);
  OR2 I62 (gocomp_0[62:62], i_0r0[62:62], i_0r1[62:62]);
  OR2 I63 (gocomp_0[63:63], i_0r0[63:63], i_0r1[63:63]);
  OR2 I64 (gocomp_0[64:64], i_0r0[64:64], i_0r1[64:64]);
  OR2 I65 (gocomp_0[65:65], i_0r0[65:65], i_0r1[65:65]);
  OR2 I66 (gocomp_0[66:66], i_0r0[66:66], i_0r1[66:66]);
  OR2 I67 (gocomp_0[67:67], i_0r0[67:67], i_0r1[67:67]);
  OR2 I68 (gocomp_0[68:68], i_0r0[68:68], i_0r1[68:68]);
  C3 I69 (simp711_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  C3 I70 (simp711_0[1:1], gocomp_0[3:3], gocomp_0[4:4], gocomp_0[5:5]);
  C3 I71 (simp711_0[2:2], gocomp_0[6:6], gocomp_0[7:7], gocomp_0[8:8]);
  C3 I72 (simp711_0[3:3], gocomp_0[9:9], gocomp_0[10:10], gocomp_0[11:11]);
  C3 I73 (simp711_0[4:4], gocomp_0[12:12], gocomp_0[13:13], gocomp_0[14:14]);
  C3 I74 (simp711_0[5:5], gocomp_0[15:15], gocomp_0[16:16], gocomp_0[17:17]);
  C3 I75 (simp711_0[6:6], gocomp_0[18:18], gocomp_0[19:19], gocomp_0[20:20]);
  C3 I76 (simp711_0[7:7], gocomp_0[21:21], gocomp_0[22:22], gocomp_0[23:23]);
  C3 I77 (simp711_0[8:8], gocomp_0[24:24], gocomp_0[25:25], gocomp_0[26:26]);
  C3 I78 (simp711_0[9:9], gocomp_0[27:27], gocomp_0[28:28], gocomp_0[29:29]);
  C3 I79 (simp711_0[10:10], gocomp_0[30:30], gocomp_0[31:31], gocomp_0[32:32]);
  C3 I80 (simp711_0[11:11], gocomp_0[33:33], gocomp_0[34:34], gocomp_0[35:35]);
  C3 I81 (simp711_0[12:12], gocomp_0[36:36], gocomp_0[37:37], gocomp_0[38:38]);
  C3 I82 (simp711_0[13:13], gocomp_0[39:39], gocomp_0[40:40], gocomp_0[41:41]);
  C3 I83 (simp711_0[14:14], gocomp_0[42:42], gocomp_0[43:43], gocomp_0[44:44]);
  C3 I84 (simp711_0[15:15], gocomp_0[45:45], gocomp_0[46:46], gocomp_0[47:47]);
  C3 I85 (simp711_0[16:16], gocomp_0[48:48], gocomp_0[49:49], gocomp_0[50:50]);
  C3 I86 (simp711_0[17:17], gocomp_0[51:51], gocomp_0[52:52], gocomp_0[53:53]);
  C3 I87 (simp711_0[18:18], gocomp_0[54:54], gocomp_0[55:55], gocomp_0[56:56]);
  C3 I88 (simp711_0[19:19], gocomp_0[57:57], gocomp_0[58:58], gocomp_0[59:59]);
  C3 I89 (simp711_0[20:20], gocomp_0[60:60], gocomp_0[61:61], gocomp_0[62:62]);
  C3 I90 (simp711_0[21:21], gocomp_0[63:63], gocomp_0[64:64], gocomp_0[65:65]);
  C3 I91 (simp711_0[22:22], gocomp_0[66:66], gocomp_0[67:67], gocomp_0[68:68]);
  C3 I92 (simp712_0[0:0], simp711_0[0:0], simp711_0[1:1], simp711_0[2:2]);
  C3 I93 (simp712_0[1:1], simp711_0[3:3], simp711_0[4:4], simp711_0[5:5]);
  C3 I94 (simp712_0[2:2], simp711_0[6:6], simp711_0[7:7], simp711_0[8:8]);
  C3 I95 (simp712_0[3:3], simp711_0[9:9], simp711_0[10:10], simp711_0[11:11]);
  C3 I96 (simp712_0[4:4], simp711_0[12:12], simp711_0[13:13], simp711_0[14:14]);
  C3 I97 (simp712_0[5:5], simp711_0[15:15], simp711_0[16:16], simp711_0[17:17]);
  C3 I98 (simp712_0[6:6], simp711_0[18:18], simp711_0[19:19], simp711_0[20:20]);
  C2 I99 (simp712_0[7:7], simp711_0[21:21], simp711_0[22:22]);
  C3 I100 (simp713_0[0:0], simp712_0[0:0], simp712_0[1:1], simp712_0[2:2]);
  C3 I101 (simp713_0[1:1], simp712_0[3:3], simp712_0[4:4], simp712_0[5:5]);
  C2 I102 (simp713_0[2:2], simp712_0[6:6], simp712_0[7:7]);
  C3 I103 (go_0, simp713_0[0:0], simp713_0[1:1], simp713_0[2:2]);
  BUFF I104 (termt_1[0:0], go_0);
  GND I105 (termf_1[0:0]);
  BUFF I106 (termf_1[1:1], go_0);
  GND I107 (termt_1[1:1]);
  BUFF I108 (termt_2[1:1], go_0);
  GND I109 (termf_2[1:1]);
  BUFF I110 (termf_2[0:0], go_0);
  GND I111 (termt_2[0:0]);
  OR2 I112 (comp30_0[0:0], termf_1[0:0], termt_1[0:0]);
  OR2 I113 (comp30_0[1:1], termf_1[1:1], termt_1[1:1]);
  C2 I114 (selcomp3_0, comp30_0[0:0], comp30_0[1:1]);
  OR2 I115 (comp31_0[0:0], termf_2[0:0], termt_2[0:0]);
  OR2 I116 (comp31_0[1:1], termf_2[1:1], termt_2[1:1]);
  C2 I117 (selcomp3_1, comp31_0[0:0], comp31_0[1:1]);
  OR2 I118 (dcomp3_0[0:0], i_0r0[32:32], i_0r1[32:32]);
  OR2 I119 (dcomp3_0[1:1], i_0r0[33:33], i_0r1[33:33]);
  OR2 I120 (dcomp3_0[2:2], i_0r0[34:34], i_0r1[34:34]);
  OR2 I121 (dcomp3_0[3:3], i_0r0[35:35], i_0r1[35:35]);
  C3 I122 (simp1251_0[0:0], dcomp3_0[0:0], dcomp3_0[1:1], dcomp3_0[2:2]);
  BUFF I123 (simp1251_0[1:1], dcomp3_0[3:3]);
  C2 I124 (scomplete3_0, simp1251_0[0:0], simp1251_0[1:1]);
  C3 I125 (icomplete3_0, scomplete3_0, selcomp3_0, selcomp3_1);
  OR2 I126 (termf_3[0:0], gfint3_0[0:0], gfint3_1[0:0]);
  OR2 I127 (termf_3[1:1], gfint3_0[1:1], gfint3_1[1:1]);
  OR2 I128 (termt_3[0:0], gtint3_0[0:0], gtint3_1[0:0]);
  OR2 I129 (termt_3[1:1], gtint3_0[1:1], gtint3_1[1:1]);
  C2R I130 (sel3_0, selg3_0, icomplete3_0, reset);
  C2R I131 (sel3_1, selg3_1, icomplete3_0, reset);
  C2R I132 (gfint3_0[0:0], sel3_0, termf_1[0:0], reset);
  C2R I133 (gfint3_0[1:1], sel3_0, termf_1[1:1], reset);
  C2R I134 (gfint3_1[0:0], sel3_1, termf_2[0:0], reset);
  C2R I135 (gfint3_1[1:1], sel3_1, termf_2[1:1], reset);
  C2R I136 (gtint3_0[0:0], sel3_0, termt_1[0:0], reset);
  C2R I137 (gtint3_0[1:1], sel3_0, termt_1[1:1], reset);
  C2R I138 (gtint3_1[0:0], sel3_1, termt_2[0:0], reset);
  C2R I139 (gtint3_1[1:1], sel3_1, termt_2[1:1], reset);
  NOR3 I140 (simp1421_0[0:0], match30_0[0:0], match30_0[1:1], match30_0[2:2]);
  INV I141 (simp1421_0[1:1], match30_0[3:3]);
  NAND2 I142 (selg3_0, simp1421_0[0:0], simp1421_0[1:1]);
  C2 I143 (match30_0[0:0], i_0r0[32:32], i_0r0[33:33]);
  C2 I144 (match30_0[1:1], i_0r1[32:32], i_0r0[33:33]);
  C3 I145 (match30_0[2:2], i_0r1[32:32], i_0r1[33:33], i_0r0[34:34]);
  C3 I146 (simp1461_0[0:0], i_0r1[32:32], i_0r1[33:33], i_0r1[34:34]);
  BUFF I147 (simp1461_0[1:1], i_0r0[35:35]);
  C2 I148 (match30_0[3:3], simp1461_0[0:0], simp1461_0[1:1]);
  NOR3 I149 (simp1481_0[0:0], match31_0[0:0], match31_0[1:1], match31_0[2:2]);
  NOR2 I150 (simp1481_0[1:1], match31_0[3:3], match31_0[4:4]);
  NAND2 I151 (selg3_1, simp1481_0[0:0], simp1481_0[1:1]);
  C3 I152 (simp1491_0[0:0], i_0r0[32:32], i_0r1[33:33], i_0r0[34:34]);
  BUFF I153 (simp1491_0[1:1], i_0r0[35:35]);
  C2 I154 (match31_0[0:0], simp1491_0[0:0], simp1491_0[1:1]);
  C3 I155 (simp1501_0[0:0], i_0r0[32:32], i_0r1[33:33], i_0r1[34:34]);
  BUFF I156 (simp1501_0[1:1], i_0r0[35:35]);
  C2 I157 (match31_0[1:1], simp1501_0[0:0], simp1501_0[1:1]);
  C3 I158 (simp1511_0[0:0], i_0r0[32:32], i_0r1[33:33], i_0r0[34:34]);
  BUFF I159 (simp1511_0[1:1], i_0r1[35:35]);
  C2 I160 (match31_0[2:2], simp1511_0[0:0], simp1511_0[1:1]);
  C3 I161 (simp1521_0[0:0], i_0r0[32:32], i_0r1[33:33], i_0r1[34:34]);
  BUFF I162 (simp1521_0[1:1], i_0r1[35:35]);
  C2 I163 (match31_0[3:3], simp1521_0[0:0], simp1521_0[1:1]);
  C3 I164 (simp1531_0[0:0], i_0r1[32:32], i_0r1[33:33], i_0r1[34:34]);
  BUFF I165 (simp1531_0[1:1], i_0r1[35:35]);
  C2 I166 (match31_0[4:4], simp1531_0[0:0], simp1531_0[1:1]);
  BUFF I167 (termt_4[0:0], go_0);
  GND I168 (termf_4[0:0]);
  BUFF I169 (termf_4[1:1], go_0);
  GND I170 (termt_4[1:1]);
  BUFF I171 (termt_5[1:1], go_0);
  GND I172 (termf_5[1:1]);
  BUFF I173 (termf_5[0:0], go_0);
  GND I174 (termt_5[0:0]);
  OR2 I175 (comp60_0[0:0], termf_4[0:0], termt_4[0:0]);
  OR2 I176 (comp60_0[1:1], termf_4[1:1], termt_4[1:1]);
  C2 I177 (selcomp6_0, comp60_0[0:0], comp60_0[1:1]);
  OR2 I178 (comp61_0[0:0], termf_5[0:0], termt_5[0:0]);
  OR2 I179 (comp61_0[1:1], termf_5[1:1], termt_5[1:1]);
  C2 I180 (selcomp6_1, comp61_0[0:0], comp61_0[1:1]);
  OR2 I181 (dcomp6_0[0:0], i_0r0[32:32], i_0r1[32:32]);
  OR2 I182 (dcomp6_0[1:1], i_0r0[33:33], i_0r1[33:33]);
  OR2 I183 (dcomp6_0[2:2], i_0r0[34:34], i_0r1[34:34]);
  OR2 I184 (dcomp6_0[3:3], i_0r0[35:35], i_0r1[35:35]);
  C3 I185 (simp1871_0[0:0], dcomp6_0[0:0], dcomp6_0[1:1], dcomp6_0[2:2]);
  BUFF I186 (simp1871_0[1:1], dcomp6_0[3:3]);
  C2 I187 (scomplete6_0, simp1871_0[0:0], simp1871_0[1:1]);
  C3 I188 (icomplete6_0, scomplete6_0, selcomp6_0, selcomp6_1);
  OR2 I189 (termf_6[0:0], gfint6_0[0:0], gfint6_1[0:0]);
  OR2 I190 (termf_6[1:1], gfint6_0[1:1], gfint6_1[1:1]);
  OR2 I191 (termt_6[0:0], gtint6_0[0:0], gtint6_1[0:0]);
  OR2 I192 (termt_6[1:1], gtint6_0[1:1], gtint6_1[1:1]);
  C2R I193 (sel6_0, selg6_0, icomplete6_0, reset);
  C2R I194 (sel6_1, selg6_1, icomplete6_0, reset);
  C2R I195 (gfint6_0[0:0], sel6_0, termf_4[0:0], reset);
  C2R I196 (gfint6_0[1:1], sel6_0, termf_4[1:1], reset);
  C2R I197 (gfint6_1[0:0], sel6_1, termf_5[0:0], reset);
  C2R I198 (gfint6_1[1:1], sel6_1, termf_5[1:1], reset);
  C2R I199 (gtint6_0[0:0], sel6_0, termt_4[0:0], reset);
  C2R I200 (gtint6_0[1:1], sel6_0, termt_4[1:1], reset);
  C2R I201 (gtint6_1[0:0], sel6_1, termt_5[0:0], reset);
  C2R I202 (gtint6_1[1:1], sel6_1, termt_5[1:1], reset);
  NOR3 I203 (simp2041_0[0:0], match60_0[0:0], match60_0[1:1], match60_0[2:2]);
  INV I204 (simp2041_0[1:1], match60_0[3:3]);
  NAND2 I205 (selg6_0, simp2041_0[0:0], simp2041_0[1:1]);
  BUFF I206 (match60_0[0:0], i_0r0[32:32]);
  C2 I207 (match60_0[1:1], i_0r1[32:32], i_0r0[33:33]);
  C3 I208 (simp2071_0[0:0], i_0r1[32:32], i_0r1[33:33], i_0r0[34:34]);
  BUFF I209 (simp2071_0[1:1], i_0r1[35:35]);
  C2 I210 (match60_0[2:2], simp2071_0[0:0], simp2071_0[1:1]);
  C3 I211 (simp2081_0[0:0], i_0r1[32:32], i_0r1[33:33], i_0r1[34:34]);
  BUFF I212 (simp2081_0[1:1], i_0r1[35:35]);
  C2 I213 (match60_0[3:3], simp2081_0[0:0], simp2081_0[1:1]);
  OR2 I214 (selg6_1, match61_0[0:0], match61_0[1:1]);
  C3 I215 (simp2111_0[0:0], i_0r1[32:32], i_0r1[33:33], i_0r0[34:34]);
  BUFF I216 (simp2111_0[1:1], i_0r0[35:35]);
  C2 I217 (match61_0[0:0], simp2111_0[0:0], simp2111_0[1:1]);
  C3 I218 (simp2121_0[0:0], i_0r1[32:32], i_0r1[33:33], i_0r1[34:34]);
  BUFF I219 (simp2121_0[1:1], i_0r0[35:35]);
  C2 I220 (match61_0[1:1], simp2121_0[0:0], simp2121_0[1:1]);
  BUFF I221 (termt_7[0:0], i_0r0[36:36]);
  BUFF I222 (termf_7[0:0], i_0r1[36:36]);
  BUFF I223 (termt_7[1:1], i_0r0[37:37]);
  BUFF I224 (termf_7[1:1], i_0r1[37:37]);
  BUFF I225 (termt_7[2:2], i_0r0[38:38]);
  BUFF I226 (termf_7[2:2], i_0r1[38:38]);
  BUFF I227 (termt_7[3:3], i_0r0[39:39]);
  BUFF I228 (termf_7[3:3], i_0r1[39:39]);
  BUFF I229 (termt_7[4:4], i_0r0[40:40]);
  BUFF I230 (termf_7[4:4], i_0r1[40:40]);
  BUFF I231 (termt_7[5:5], i_0r0[41:41]);
  BUFF I232 (termf_7[5:5], i_0r1[41:41]);
  BUFF I233 (termt_7[6:6], i_0r0[42:42]);
  BUFF I234 (termf_7[6:6], i_0r1[42:42]);
  BUFF I235 (termt_7[7:7], i_0r0[43:43]);
  BUFF I236 (termf_7[7:7], i_0r1[43:43]);
  BUFF I237 (termt_7[8:8], i_0r0[44:44]);
  BUFF I238 (termf_7[8:8], i_0r1[44:44]);
  BUFF I239 (termt_7[9:9], i_0r0[45:45]);
  BUFF I240 (termf_7[9:9], i_0r1[45:45]);
  BUFF I241 (termt_7[10:10], i_0r0[46:46]);
  BUFF I242 (termf_7[10:10], i_0r1[46:46]);
  BUFF I243 (termt_7[11:11], i_0r0[47:47]);
  BUFF I244 (termf_7[11:11], i_0r1[47:47]);
  BUFF I245 (termt_7[12:12], i_0r0[48:48]);
  BUFF I246 (termf_7[12:12], i_0r1[48:48]);
  BUFF I247 (termt_7[13:13], i_0r0[49:49]);
  BUFF I248 (termf_7[13:13], i_0r1[49:49]);
  BUFF I249 (termt_7[14:14], i_0r0[50:50]);
  BUFF I250 (termf_7[14:14], i_0r1[50:50]);
  BUFF I251 (termt_7[15:15], i_0r0[51:51]);
  BUFF I252 (termf_7[15:15], i_0r1[51:51]);
  BUFF I253 (termt_7[16:16], i_0r0[52:52]);
  BUFF I254 (termf_7[16:16], i_0r1[52:52]);
  BUFF I255 (termt_7[17:17], i_0r0[53:53]);
  BUFF I256 (termf_7[17:17], i_0r1[53:53]);
  BUFF I257 (termt_7[18:18], i_0r0[54:54]);
  BUFF I258 (termf_7[18:18], i_0r1[54:54]);
  BUFF I259 (termt_7[19:19], i_0r0[55:55]);
  BUFF I260 (termf_7[19:19], i_0r1[55:55]);
  BUFF I261 (termt_7[20:20], i_0r0[56:56]);
  BUFF I262 (termf_7[20:20], i_0r1[56:56]);
  BUFF I263 (termt_7[21:21], i_0r0[57:57]);
  BUFF I264 (termf_7[21:21], i_0r1[57:57]);
  BUFF I265 (termt_7[22:22], i_0r0[58:58]);
  BUFF I266 (termf_7[22:22], i_0r1[58:58]);
  BUFF I267 (termt_7[23:23], i_0r0[59:59]);
  BUFF I268 (termf_7[23:23], i_0r1[59:59]);
  BUFF I269 (termt_7[24:24], i_0r0[60:60]);
  BUFF I270 (termf_7[24:24], i_0r1[60:60]);
  BUFF I271 (termt_7[25:25], i_0r0[61:61]);
  BUFF I272 (termf_7[25:25], i_0r1[61:61]);
  BUFF I273 (termt_7[26:26], i_0r0[62:62]);
  BUFF I274 (termf_7[26:26], i_0r1[62:62]);
  BUFF I275 (termt_7[27:27], i_0r0[63:63]);
  BUFF I276 (termf_7[27:27], i_0r1[63:63]);
  BUFF I277 (termt_7[28:28], i_0r0[64:64]);
  BUFF I278 (termf_7[28:28], i_0r1[64:64]);
  BUFF I279 (termt_7[29:29], i_0r0[65:65]);
  BUFF I280 (termf_7[29:29], i_0r1[65:65]);
  BUFF I281 (termt_7[30:30], i_0r0[66:66]);
  BUFF I282 (termf_7[30:30], i_0r1[66:66]);
  BUFF I283 (termt_7[31:31], i_0r0[67:67]);
  BUFF I284 (termf_7[31:31], i_0r1[67:67]);
  OR2 I285 (comp80_0[0:0], termf_7[0:0], termt_7[0:0]);
  OR2 I286 (comp80_0[1:1], termf_7[1:1], termt_7[1:1]);
  OR2 I287 (comp80_0[2:2], termf_7[2:2], termt_7[2:2]);
  OR2 I288 (comp80_0[3:3], termf_7[3:3], termt_7[3:3]);
  OR2 I289 (comp80_0[4:4], termf_7[4:4], termt_7[4:4]);
  OR2 I290 (comp80_0[5:5], termf_7[5:5], termt_7[5:5]);
  OR2 I291 (comp80_0[6:6], termf_7[6:6], termt_7[6:6]);
  OR2 I292 (comp80_0[7:7], termf_7[7:7], termt_7[7:7]);
  OR2 I293 (comp80_0[8:8], termf_7[8:8], termt_7[8:8]);
  OR2 I294 (comp80_0[9:9], termf_7[9:9], termt_7[9:9]);
  OR2 I295 (comp80_0[10:10], termf_7[10:10], termt_7[10:10]);
  OR2 I296 (comp80_0[11:11], termf_7[11:11], termt_7[11:11]);
  OR2 I297 (comp80_0[12:12], termf_7[12:12], termt_7[12:12]);
  OR2 I298 (comp80_0[13:13], termf_7[13:13], termt_7[13:13]);
  OR2 I299 (comp80_0[14:14], termf_7[14:14], termt_7[14:14]);
  OR2 I300 (comp80_0[15:15], termf_7[15:15], termt_7[15:15]);
  OR2 I301 (comp80_0[16:16], termf_7[16:16], termt_7[16:16]);
  OR2 I302 (comp80_0[17:17], termf_7[17:17], termt_7[17:17]);
  OR2 I303 (comp80_0[18:18], termf_7[18:18], termt_7[18:18]);
  OR2 I304 (comp80_0[19:19], termf_7[19:19], termt_7[19:19]);
  OR2 I305 (comp80_0[20:20], termf_7[20:20], termt_7[20:20]);
  OR2 I306 (comp80_0[21:21], termf_7[21:21], termt_7[21:21]);
  OR2 I307 (comp80_0[22:22], termf_7[22:22], termt_7[22:22]);
  OR2 I308 (comp80_0[23:23], termf_7[23:23], termt_7[23:23]);
  OR2 I309 (comp80_0[24:24], termf_7[24:24], termt_7[24:24]);
  OR2 I310 (comp80_0[25:25], termf_7[25:25], termt_7[25:25]);
  OR2 I311 (comp80_0[26:26], termf_7[26:26], termt_7[26:26]);
  OR2 I312 (comp80_0[27:27], termf_7[27:27], termt_7[27:27]);
  OR2 I313 (comp80_0[28:28], termf_7[28:28], termt_7[28:28]);
  OR2 I314 (comp80_0[29:29], termf_7[29:29], termt_7[29:29]);
  OR2 I315 (comp80_0[30:30], termf_7[30:30], termt_7[30:30]);
  OR2 I316 (comp80_0[31:31], termf_7[31:31], termt_7[31:31]);
  C3 I317 (simp3221_0[0:0], comp80_0[0:0], comp80_0[1:1], comp80_0[2:2]);
  C3 I318 (simp3221_0[1:1], comp80_0[3:3], comp80_0[4:4], comp80_0[5:5]);
  C3 I319 (simp3221_0[2:2], comp80_0[6:6], comp80_0[7:7], comp80_0[8:8]);
  C3 I320 (simp3221_0[3:3], comp80_0[9:9], comp80_0[10:10], comp80_0[11:11]);
  C3 I321 (simp3221_0[4:4], comp80_0[12:12], comp80_0[13:13], comp80_0[14:14]);
  C3 I322 (simp3221_0[5:5], comp80_0[15:15], comp80_0[16:16], comp80_0[17:17]);
  C3 I323 (simp3221_0[6:6], comp80_0[18:18], comp80_0[19:19], comp80_0[20:20]);
  C3 I324 (simp3221_0[7:7], comp80_0[21:21], comp80_0[22:22], comp80_0[23:23]);
  C3 I325 (simp3221_0[8:8], comp80_0[24:24], comp80_0[25:25], comp80_0[26:26]);
  C3 I326 (simp3221_0[9:9], comp80_0[27:27], comp80_0[28:28], comp80_0[29:29]);
  C2 I327 (simp3221_0[10:10], comp80_0[30:30], comp80_0[31:31]);
  C3 I328 (simp3222_0[0:0], simp3221_0[0:0], simp3221_0[1:1], simp3221_0[2:2]);
  C3 I329 (simp3222_0[1:1], simp3221_0[3:3], simp3221_0[4:4], simp3221_0[5:5]);
  C3 I330 (simp3222_0[2:2], simp3221_0[6:6], simp3221_0[7:7], simp3221_0[8:8]);
  C2 I331 (simp3222_0[3:3], simp3221_0[9:9], simp3221_0[10:10]);
  C3 I332 (simp3223_0[0:0], simp3222_0[0:0], simp3222_0[1:1], simp3222_0[2:2]);
  BUFF I333 (simp3223_0[1:1], simp3222_0[3:3]);
  C2 I334 (selcomp8_0, simp3223_0[0:0], simp3223_0[1:1]);
  OR2 I335 (comp81_0[0:0], i_0r0[36:36], i_0r1[36:36]);
  OR2 I336 (comp81_0[1:1], i_0r0[37:37], i_0r1[37:37]);
  OR2 I337 (comp81_0[2:2], i_0r0[38:38], i_0r1[38:38]);
  OR2 I338 (comp81_0[3:3], i_0r0[39:39], i_0r1[39:39]);
  OR2 I339 (comp81_0[4:4], i_0r0[40:40], i_0r1[40:40]);
  OR2 I340 (comp81_0[5:5], i_0r0[41:41], i_0r1[41:41]);
  OR2 I341 (comp81_0[6:6], i_0r0[42:42], i_0r1[42:42]);
  OR2 I342 (comp81_0[7:7], i_0r0[43:43], i_0r1[43:43]);
  OR2 I343 (comp81_0[8:8], i_0r0[44:44], i_0r1[44:44]);
  OR2 I344 (comp81_0[9:9], i_0r0[45:45], i_0r1[45:45]);
  OR2 I345 (comp81_0[10:10], i_0r0[46:46], i_0r1[46:46]);
  OR2 I346 (comp81_0[11:11], i_0r0[47:47], i_0r1[47:47]);
  OR2 I347 (comp81_0[12:12], i_0r0[48:48], i_0r1[48:48]);
  OR2 I348 (comp81_0[13:13], i_0r0[49:49], i_0r1[49:49]);
  OR2 I349 (comp81_0[14:14], i_0r0[50:50], i_0r1[50:50]);
  OR2 I350 (comp81_0[15:15], i_0r0[51:51], i_0r1[51:51]);
  OR2 I351 (comp81_0[16:16], i_0r0[52:52], i_0r1[52:52]);
  OR2 I352 (comp81_0[17:17], i_0r0[53:53], i_0r1[53:53]);
  OR2 I353 (comp81_0[18:18], i_0r0[54:54], i_0r1[54:54]);
  OR2 I354 (comp81_0[19:19], i_0r0[55:55], i_0r1[55:55]);
  OR2 I355 (comp81_0[20:20], i_0r0[56:56], i_0r1[56:56]);
  OR2 I356 (comp81_0[21:21], i_0r0[57:57], i_0r1[57:57]);
  OR2 I357 (comp81_0[22:22], i_0r0[58:58], i_0r1[58:58]);
  OR2 I358 (comp81_0[23:23], i_0r0[59:59], i_0r1[59:59]);
  OR2 I359 (comp81_0[24:24], i_0r0[60:60], i_0r1[60:60]);
  OR2 I360 (comp81_0[25:25], i_0r0[61:61], i_0r1[61:61]);
  OR2 I361 (comp81_0[26:26], i_0r0[62:62], i_0r1[62:62]);
  OR2 I362 (comp81_0[27:27], i_0r0[63:63], i_0r1[63:63]);
  OR2 I363 (comp81_0[28:28], i_0r0[64:64], i_0r1[64:64]);
  OR2 I364 (comp81_0[29:29], i_0r0[65:65], i_0r1[65:65]);
  OR2 I365 (comp81_0[30:30], i_0r0[66:66], i_0r1[66:66]);
  OR2 I366 (comp81_0[31:31], i_0r0[67:67], i_0r1[67:67]);
  C3 I367 (simp3561_0[0:0], comp81_0[0:0], comp81_0[1:1], comp81_0[2:2]);
  C3 I368 (simp3561_0[1:1], comp81_0[3:3], comp81_0[4:4], comp81_0[5:5]);
  C3 I369 (simp3561_0[2:2], comp81_0[6:6], comp81_0[7:7], comp81_0[8:8]);
  C3 I370 (simp3561_0[3:3], comp81_0[9:9], comp81_0[10:10], comp81_0[11:11]);
  C3 I371 (simp3561_0[4:4], comp81_0[12:12], comp81_0[13:13], comp81_0[14:14]);
  C3 I372 (simp3561_0[5:5], comp81_0[15:15], comp81_0[16:16], comp81_0[17:17]);
  C3 I373 (simp3561_0[6:6], comp81_0[18:18], comp81_0[19:19], comp81_0[20:20]);
  C3 I374 (simp3561_0[7:7], comp81_0[21:21], comp81_0[22:22], comp81_0[23:23]);
  C3 I375 (simp3561_0[8:8], comp81_0[24:24], comp81_0[25:25], comp81_0[26:26]);
  C3 I376 (simp3561_0[9:9], comp81_0[27:27], comp81_0[28:28], comp81_0[29:29]);
  C2 I377 (simp3561_0[10:10], comp81_0[30:30], comp81_0[31:31]);
  C3 I378 (simp3562_0[0:0], simp3561_0[0:0], simp3561_0[1:1], simp3561_0[2:2]);
  C3 I379 (simp3562_0[1:1], simp3561_0[3:3], simp3561_0[4:4], simp3561_0[5:5]);
  C3 I380 (simp3562_0[2:2], simp3561_0[6:6], simp3561_0[7:7], simp3561_0[8:8]);
  C2 I381 (simp3562_0[3:3], simp3561_0[9:9], simp3561_0[10:10]);
  C3 I382 (simp3563_0[0:0], simp3562_0[0:0], simp3562_0[1:1], simp3562_0[2:2]);
  BUFF I383 (simp3563_0[1:1], simp3562_0[3:3]);
  C2 I384 (selcomp8_1, simp3563_0[0:0], simp3563_0[1:1]);
  OR2 I385 (dcomp8_0[0:0], termf_3[0:0], termt_3[0:0]);
  OR2 I386 (dcomp8_0[1:1], termf_3[1:1], termt_3[1:1]);
  C2 I387 (scomplete8_0, dcomp8_0[0:0], dcomp8_0[1:1]);
  C3 I388 (icomplete8_0, scomplete8_0, selcomp8_0, selcomp8_1);
  OR2 I389 (termf_8[0:0], gfint8_0[0:0], gfint8_1[0:0]);
  OR2 I390 (termf_8[1:1], gfint8_0[1:1], gfint8_1[1:1]);
  OR2 I391 (termf_8[2:2], gfint8_0[2:2], gfint8_1[2:2]);
  OR2 I392 (termf_8[3:3], gfint8_0[3:3], gfint8_1[3:3]);
  OR2 I393 (termf_8[4:4], gfint8_0[4:4], gfint8_1[4:4]);
  OR2 I394 (termf_8[5:5], gfint8_0[5:5], gfint8_1[5:5]);
  OR2 I395 (termf_8[6:6], gfint8_0[6:6], gfint8_1[6:6]);
  OR2 I396 (termf_8[7:7], gfint8_0[7:7], gfint8_1[7:7]);
  OR2 I397 (termf_8[8:8], gfint8_0[8:8], gfint8_1[8:8]);
  OR2 I398 (termf_8[9:9], gfint8_0[9:9], gfint8_1[9:9]);
  OR2 I399 (termf_8[10:10], gfint8_0[10:10], gfint8_1[10:10]);
  OR2 I400 (termf_8[11:11], gfint8_0[11:11], gfint8_1[11:11]);
  OR2 I401 (termf_8[12:12], gfint8_0[12:12], gfint8_1[12:12]);
  OR2 I402 (termf_8[13:13], gfint8_0[13:13], gfint8_1[13:13]);
  OR2 I403 (termf_8[14:14], gfint8_0[14:14], gfint8_1[14:14]);
  OR2 I404 (termf_8[15:15], gfint8_0[15:15], gfint8_1[15:15]);
  OR2 I405 (termf_8[16:16], gfint8_0[16:16], gfint8_1[16:16]);
  OR2 I406 (termf_8[17:17], gfint8_0[17:17], gfint8_1[17:17]);
  OR2 I407 (termf_8[18:18], gfint8_0[18:18], gfint8_1[18:18]);
  OR2 I408 (termf_8[19:19], gfint8_0[19:19], gfint8_1[19:19]);
  OR2 I409 (termf_8[20:20], gfint8_0[20:20], gfint8_1[20:20]);
  OR2 I410 (termf_8[21:21], gfint8_0[21:21], gfint8_1[21:21]);
  OR2 I411 (termf_8[22:22], gfint8_0[22:22], gfint8_1[22:22]);
  OR2 I412 (termf_8[23:23], gfint8_0[23:23], gfint8_1[23:23]);
  OR2 I413 (termf_8[24:24], gfint8_0[24:24], gfint8_1[24:24]);
  OR2 I414 (termf_8[25:25], gfint8_0[25:25], gfint8_1[25:25]);
  OR2 I415 (termf_8[26:26], gfint8_0[26:26], gfint8_1[26:26]);
  OR2 I416 (termf_8[27:27], gfint8_0[27:27], gfint8_1[27:27]);
  OR2 I417 (termf_8[28:28], gfint8_0[28:28], gfint8_1[28:28]);
  OR2 I418 (termf_8[29:29], gfint8_0[29:29], gfint8_1[29:29]);
  OR2 I419 (termf_8[30:30], gfint8_0[30:30], gfint8_1[30:30]);
  OR2 I420 (termf_8[31:31], gfint8_0[31:31], gfint8_1[31:31]);
  OR2 I421 (termt_8[0:0], gtint8_0[0:0], gtint8_1[0:0]);
  OR2 I422 (termt_8[1:1], gtint8_0[1:1], gtint8_1[1:1]);
  OR2 I423 (termt_8[2:2], gtint8_0[2:2], gtint8_1[2:2]);
  OR2 I424 (termt_8[3:3], gtint8_0[3:3], gtint8_1[3:3]);
  OR2 I425 (termt_8[4:4], gtint8_0[4:4], gtint8_1[4:4]);
  OR2 I426 (termt_8[5:5], gtint8_0[5:5], gtint8_1[5:5]);
  OR2 I427 (termt_8[6:6], gtint8_0[6:6], gtint8_1[6:6]);
  OR2 I428 (termt_8[7:7], gtint8_0[7:7], gtint8_1[7:7]);
  OR2 I429 (termt_8[8:8], gtint8_0[8:8], gtint8_1[8:8]);
  OR2 I430 (termt_8[9:9], gtint8_0[9:9], gtint8_1[9:9]);
  OR2 I431 (termt_8[10:10], gtint8_0[10:10], gtint8_1[10:10]);
  OR2 I432 (termt_8[11:11], gtint8_0[11:11], gtint8_1[11:11]);
  OR2 I433 (termt_8[12:12], gtint8_0[12:12], gtint8_1[12:12]);
  OR2 I434 (termt_8[13:13], gtint8_0[13:13], gtint8_1[13:13]);
  OR2 I435 (termt_8[14:14], gtint8_0[14:14], gtint8_1[14:14]);
  OR2 I436 (termt_8[15:15], gtint8_0[15:15], gtint8_1[15:15]);
  OR2 I437 (termt_8[16:16], gtint8_0[16:16], gtint8_1[16:16]);
  OR2 I438 (termt_8[17:17], gtint8_0[17:17], gtint8_1[17:17]);
  OR2 I439 (termt_8[18:18], gtint8_0[18:18], gtint8_1[18:18]);
  OR2 I440 (termt_8[19:19], gtint8_0[19:19], gtint8_1[19:19]);
  OR2 I441 (termt_8[20:20], gtint8_0[20:20], gtint8_1[20:20]);
  OR2 I442 (termt_8[21:21], gtint8_0[21:21], gtint8_1[21:21]);
  OR2 I443 (termt_8[22:22], gtint8_0[22:22], gtint8_1[22:22]);
  OR2 I444 (termt_8[23:23], gtint8_0[23:23], gtint8_1[23:23]);
  OR2 I445 (termt_8[24:24], gtint8_0[24:24], gtint8_1[24:24]);
  OR2 I446 (termt_8[25:25], gtint8_0[25:25], gtint8_1[25:25]);
  OR2 I447 (termt_8[26:26], gtint8_0[26:26], gtint8_1[26:26]);
  OR2 I448 (termt_8[27:27], gtint8_0[27:27], gtint8_1[27:27]);
  OR2 I449 (termt_8[28:28], gtint8_0[28:28], gtint8_1[28:28]);
  OR2 I450 (termt_8[29:29], gtint8_0[29:29], gtint8_1[29:29]);
  OR2 I451 (termt_8[30:30], gtint8_0[30:30], gtint8_1[30:30]);
  OR2 I452 (termt_8[31:31], gtint8_0[31:31], gtint8_1[31:31]);
  C2R I453 (sel8_0, selg8_0, icomplete8_0, reset);
  C2R I454 (sel8_1, selg8_1, icomplete8_0, reset);
  C2R I455 (gfint8_0[0:0], sel8_0, termf_7[0:0], reset);
  C2R I456 (gfint8_0[1:1], sel8_0, termf_7[1:1], reset);
  C2R I457 (gfint8_0[2:2], sel8_0, termf_7[2:2], reset);
  C2R I458 (gfint8_0[3:3], sel8_0, termf_7[3:3], reset);
  C2R I459 (gfint8_0[4:4], sel8_0, termf_7[4:4], reset);
  C2R I460 (gfint8_0[5:5], sel8_0, termf_7[5:5], reset);
  C2R I461 (gfint8_0[6:6], sel8_0, termf_7[6:6], reset);
  C2R I462 (gfint8_0[7:7], sel8_0, termf_7[7:7], reset);
  C2R I463 (gfint8_0[8:8], sel8_0, termf_7[8:8], reset);
  C2R I464 (gfint8_0[9:9], sel8_0, termf_7[9:9], reset);
  C2R I465 (gfint8_0[10:10], sel8_0, termf_7[10:10], reset);
  C2R I466 (gfint8_0[11:11], sel8_0, termf_7[11:11], reset);
  C2R I467 (gfint8_0[12:12], sel8_0, termf_7[12:12], reset);
  C2R I468 (gfint8_0[13:13], sel8_0, termf_7[13:13], reset);
  C2R I469 (gfint8_0[14:14], sel8_0, termf_7[14:14], reset);
  C2R I470 (gfint8_0[15:15], sel8_0, termf_7[15:15], reset);
  C2R I471 (gfint8_0[16:16], sel8_0, termf_7[16:16], reset);
  C2R I472 (gfint8_0[17:17], sel8_0, termf_7[17:17], reset);
  C2R I473 (gfint8_0[18:18], sel8_0, termf_7[18:18], reset);
  C2R I474 (gfint8_0[19:19], sel8_0, termf_7[19:19], reset);
  C2R I475 (gfint8_0[20:20], sel8_0, termf_7[20:20], reset);
  C2R I476 (gfint8_0[21:21], sel8_0, termf_7[21:21], reset);
  C2R I477 (gfint8_0[22:22], sel8_0, termf_7[22:22], reset);
  C2R I478 (gfint8_0[23:23], sel8_0, termf_7[23:23], reset);
  C2R I479 (gfint8_0[24:24], sel8_0, termf_7[24:24], reset);
  C2R I480 (gfint8_0[25:25], sel8_0, termf_7[25:25], reset);
  C2R I481 (gfint8_0[26:26], sel8_0, termf_7[26:26], reset);
  C2R I482 (gfint8_0[27:27], sel8_0, termf_7[27:27], reset);
  C2R I483 (gfint8_0[28:28], sel8_0, termf_7[28:28], reset);
  C2R I484 (gfint8_0[29:29], sel8_0, termf_7[29:29], reset);
  C2R I485 (gfint8_0[30:30], sel8_0, termf_7[30:30], reset);
  C2R I486 (gfint8_0[31:31], sel8_0, termf_7[31:31], reset);
  C2R I487 (gfint8_1[0:0], sel8_1, i_0r0[36:36], reset);
  C2R I488 (gfint8_1[1:1], sel8_1, i_0r0[37:37], reset);
  C2R I489 (gfint8_1[2:2], sel8_1, i_0r0[38:38], reset);
  C2R I490 (gfint8_1[3:3], sel8_1, i_0r0[39:39], reset);
  C2R I491 (gfint8_1[4:4], sel8_1, i_0r0[40:40], reset);
  C2R I492 (gfint8_1[5:5], sel8_1, i_0r0[41:41], reset);
  C2R I493 (gfint8_1[6:6], sel8_1, i_0r0[42:42], reset);
  C2R I494 (gfint8_1[7:7], sel8_1, i_0r0[43:43], reset);
  C2R I495 (gfint8_1[8:8], sel8_1, i_0r0[44:44], reset);
  C2R I496 (gfint8_1[9:9], sel8_1, i_0r0[45:45], reset);
  C2R I497 (gfint8_1[10:10], sel8_1, i_0r0[46:46], reset);
  C2R I498 (gfint8_1[11:11], sel8_1, i_0r0[47:47], reset);
  C2R I499 (gfint8_1[12:12], sel8_1, i_0r0[48:48], reset);
  C2R I500 (gfint8_1[13:13], sel8_1, i_0r0[49:49], reset);
  C2R I501 (gfint8_1[14:14], sel8_1, i_0r0[50:50], reset);
  C2R I502 (gfint8_1[15:15], sel8_1, i_0r0[51:51], reset);
  C2R I503 (gfint8_1[16:16], sel8_1, i_0r0[52:52], reset);
  C2R I504 (gfint8_1[17:17], sel8_1, i_0r0[53:53], reset);
  C2R I505 (gfint8_1[18:18], sel8_1, i_0r0[54:54], reset);
  C2R I506 (gfint8_1[19:19], sel8_1, i_0r0[55:55], reset);
  C2R I507 (gfint8_1[20:20], sel8_1, i_0r0[56:56], reset);
  C2R I508 (gfint8_1[21:21], sel8_1, i_0r0[57:57], reset);
  C2R I509 (gfint8_1[22:22], sel8_1, i_0r0[58:58], reset);
  C2R I510 (gfint8_1[23:23], sel8_1, i_0r0[59:59], reset);
  C2R I511 (gfint8_1[24:24], sel8_1, i_0r0[60:60], reset);
  C2R I512 (gfint8_1[25:25], sel8_1, i_0r0[61:61], reset);
  C2R I513 (gfint8_1[26:26], sel8_1, i_0r0[62:62], reset);
  C2R I514 (gfint8_1[27:27], sel8_1, i_0r0[63:63], reset);
  C2R I515 (gfint8_1[28:28], sel8_1, i_0r0[64:64], reset);
  C2R I516 (gfint8_1[29:29], sel8_1, i_0r0[65:65], reset);
  C2R I517 (gfint8_1[30:30], sel8_1, i_0r0[66:66], reset);
  C2R I518 (gfint8_1[31:31], sel8_1, i_0r0[67:67], reset);
  C2R I519 (gtint8_0[0:0], sel8_0, termt_7[0:0], reset);
  C2R I520 (gtint8_0[1:1], sel8_0, termt_7[1:1], reset);
  C2R I521 (gtint8_0[2:2], sel8_0, termt_7[2:2], reset);
  C2R I522 (gtint8_0[3:3], sel8_0, termt_7[3:3], reset);
  C2R I523 (gtint8_0[4:4], sel8_0, termt_7[4:4], reset);
  C2R I524 (gtint8_0[5:5], sel8_0, termt_7[5:5], reset);
  C2R I525 (gtint8_0[6:6], sel8_0, termt_7[6:6], reset);
  C2R I526 (gtint8_0[7:7], sel8_0, termt_7[7:7], reset);
  C2R I527 (gtint8_0[8:8], sel8_0, termt_7[8:8], reset);
  C2R I528 (gtint8_0[9:9], sel8_0, termt_7[9:9], reset);
  C2R I529 (gtint8_0[10:10], sel8_0, termt_7[10:10], reset);
  C2R I530 (gtint8_0[11:11], sel8_0, termt_7[11:11], reset);
  C2R I531 (gtint8_0[12:12], sel8_0, termt_7[12:12], reset);
  C2R I532 (gtint8_0[13:13], sel8_0, termt_7[13:13], reset);
  C2R I533 (gtint8_0[14:14], sel8_0, termt_7[14:14], reset);
  C2R I534 (gtint8_0[15:15], sel8_0, termt_7[15:15], reset);
  C2R I535 (gtint8_0[16:16], sel8_0, termt_7[16:16], reset);
  C2R I536 (gtint8_0[17:17], sel8_0, termt_7[17:17], reset);
  C2R I537 (gtint8_0[18:18], sel8_0, termt_7[18:18], reset);
  C2R I538 (gtint8_0[19:19], sel8_0, termt_7[19:19], reset);
  C2R I539 (gtint8_0[20:20], sel8_0, termt_7[20:20], reset);
  C2R I540 (gtint8_0[21:21], sel8_0, termt_7[21:21], reset);
  C2R I541 (gtint8_0[22:22], sel8_0, termt_7[22:22], reset);
  C2R I542 (gtint8_0[23:23], sel8_0, termt_7[23:23], reset);
  C2R I543 (gtint8_0[24:24], sel8_0, termt_7[24:24], reset);
  C2R I544 (gtint8_0[25:25], sel8_0, termt_7[25:25], reset);
  C2R I545 (gtint8_0[26:26], sel8_0, termt_7[26:26], reset);
  C2R I546 (gtint8_0[27:27], sel8_0, termt_7[27:27], reset);
  C2R I547 (gtint8_0[28:28], sel8_0, termt_7[28:28], reset);
  C2R I548 (gtint8_0[29:29], sel8_0, termt_7[29:29], reset);
  C2R I549 (gtint8_0[30:30], sel8_0, termt_7[30:30], reset);
  C2R I550 (gtint8_0[31:31], sel8_0, termt_7[31:31], reset);
  C2R I551 (gtint8_1[0:0], sel8_1, i_0r1[36:36], reset);
  C2R I552 (gtint8_1[1:1], sel8_1, i_0r1[37:37], reset);
  C2R I553 (gtint8_1[2:2], sel8_1, i_0r1[38:38], reset);
  C2R I554 (gtint8_1[3:3], sel8_1, i_0r1[39:39], reset);
  C2R I555 (gtint8_1[4:4], sel8_1, i_0r1[40:40], reset);
  C2R I556 (gtint8_1[5:5], sel8_1, i_0r1[41:41], reset);
  C2R I557 (gtint8_1[6:6], sel8_1, i_0r1[42:42], reset);
  C2R I558 (gtint8_1[7:7], sel8_1, i_0r1[43:43], reset);
  C2R I559 (gtint8_1[8:8], sel8_1, i_0r1[44:44], reset);
  C2R I560 (gtint8_1[9:9], sel8_1, i_0r1[45:45], reset);
  C2R I561 (gtint8_1[10:10], sel8_1, i_0r1[46:46], reset);
  C2R I562 (gtint8_1[11:11], sel8_1, i_0r1[47:47], reset);
  C2R I563 (gtint8_1[12:12], sel8_1, i_0r1[48:48], reset);
  C2R I564 (gtint8_1[13:13], sel8_1, i_0r1[49:49], reset);
  C2R I565 (gtint8_1[14:14], sel8_1, i_0r1[50:50], reset);
  C2R I566 (gtint8_1[15:15], sel8_1, i_0r1[51:51], reset);
  C2R I567 (gtint8_1[16:16], sel8_1, i_0r1[52:52], reset);
  C2R I568 (gtint8_1[17:17], sel8_1, i_0r1[53:53], reset);
  C2R I569 (gtint8_1[18:18], sel8_1, i_0r1[54:54], reset);
  C2R I570 (gtint8_1[19:19], sel8_1, i_0r1[55:55], reset);
  C2R I571 (gtint8_1[20:20], sel8_1, i_0r1[56:56], reset);
  C2R I572 (gtint8_1[21:21], sel8_1, i_0r1[57:57], reset);
  C2R I573 (gtint8_1[22:22], sel8_1, i_0r1[58:58], reset);
  C2R I574 (gtint8_1[23:23], sel8_1, i_0r1[59:59], reset);
  C2R I575 (gtint8_1[24:24], sel8_1, i_0r1[60:60], reset);
  C2R I576 (gtint8_1[25:25], sel8_1, i_0r1[61:61], reset);
  C2R I577 (gtint8_1[26:26], sel8_1, i_0r1[62:62], reset);
  C2R I578 (gtint8_1[27:27], sel8_1, i_0r1[63:63], reset);
  C2R I579 (gtint8_1[28:28], sel8_1, i_0r1[64:64], reset);
  C2R I580 (gtint8_1[29:29], sel8_1, i_0r1[65:65], reset);
  C2R I581 (gtint8_1[30:30], sel8_1, i_0r1[66:66], reset);
  C2R I582 (gtint8_1[31:31], sel8_1, i_0r1[67:67], reset);
  BUFF I583 (selg8_0, match80_0);
  C2 I584 (match80_0, termf_3[0:0], termt_3[1:1]);
  BUFF I585 (selg8_1, match81_0);
  C2 I586 (match81_0, termt_3[0:0], termf_3[1:1]);
  BUFF I587 (termt_9[0:0], i_0r0[0:0]);
  BUFF I588 (termf_9[0:0], i_0r1[0:0]);
  BUFF I589 (termt_9[1:1], i_0r0[1:1]);
  BUFF I590 (termf_9[1:1], i_0r1[1:1]);
  BUFF I591 (termt_9[2:2], i_0r0[2:2]);
  BUFF I592 (termf_9[2:2], i_0r1[2:2]);
  BUFF I593 (termt_9[3:3], i_0r0[3:3]);
  BUFF I594 (termf_9[3:3], i_0r1[3:3]);
  BUFF I595 (termt_9[4:4], i_0r0[4:4]);
  BUFF I596 (termf_9[4:4], i_0r1[4:4]);
  BUFF I597 (termt_9[5:5], i_0r0[5:5]);
  BUFF I598 (termf_9[5:5], i_0r1[5:5]);
  BUFF I599 (termt_9[6:6], i_0r0[6:6]);
  BUFF I600 (termf_9[6:6], i_0r1[6:6]);
  BUFF I601 (termt_9[7:7], i_0r0[7:7]);
  BUFF I602 (termf_9[7:7], i_0r1[7:7]);
  BUFF I603 (termt_9[8:8], i_0r0[8:8]);
  BUFF I604 (termf_9[8:8], i_0r1[8:8]);
  BUFF I605 (termt_9[9:9], i_0r0[9:9]);
  BUFF I606 (termf_9[9:9], i_0r1[9:9]);
  BUFF I607 (termt_9[10:10], i_0r0[10:10]);
  BUFF I608 (termf_9[10:10], i_0r1[10:10]);
  BUFF I609 (termt_9[11:11], i_0r0[11:11]);
  BUFF I610 (termf_9[11:11], i_0r1[11:11]);
  BUFF I611 (termt_9[12:12], i_0r0[12:12]);
  BUFF I612 (termf_9[12:12], i_0r1[12:12]);
  BUFF I613 (termt_9[13:13], i_0r0[13:13]);
  BUFF I614 (termf_9[13:13], i_0r1[13:13]);
  BUFF I615 (termt_9[14:14], i_0r0[14:14]);
  BUFF I616 (termf_9[14:14], i_0r1[14:14]);
  BUFF I617 (termt_9[15:15], i_0r0[15:15]);
  BUFF I618 (termf_9[15:15], i_0r1[15:15]);
  BUFF I619 (termt_9[16:16], i_0r0[16:16]);
  BUFF I620 (termf_9[16:16], i_0r1[16:16]);
  BUFF I621 (termt_9[17:17], i_0r0[17:17]);
  BUFF I622 (termf_9[17:17], i_0r1[17:17]);
  BUFF I623 (termt_9[18:18], i_0r0[18:18]);
  BUFF I624 (termf_9[18:18], i_0r1[18:18]);
  BUFF I625 (termt_9[19:19], i_0r0[19:19]);
  BUFF I626 (termf_9[19:19], i_0r1[19:19]);
  BUFF I627 (termt_9[20:20], i_0r0[20:20]);
  BUFF I628 (termf_9[20:20], i_0r1[20:20]);
  BUFF I629 (termt_9[21:21], i_0r0[21:21]);
  BUFF I630 (termf_9[21:21], i_0r1[21:21]);
  BUFF I631 (termt_9[22:22], i_0r0[22:22]);
  BUFF I632 (termf_9[22:22], i_0r1[22:22]);
  BUFF I633 (termt_9[23:23], i_0r0[23:23]);
  BUFF I634 (termf_9[23:23], i_0r1[23:23]);
  BUFF I635 (termt_9[24:24], i_0r0[24:24]);
  BUFF I636 (termf_9[24:24], i_0r1[24:24]);
  BUFF I637 (termt_9[25:25], i_0r0[25:25]);
  BUFF I638 (termf_9[25:25], i_0r1[25:25]);
  BUFF I639 (termt_9[26:26], i_0r0[26:26]);
  BUFF I640 (termf_9[26:26], i_0r1[26:26]);
  BUFF I641 (termt_9[27:27], i_0r0[27:27]);
  BUFF I642 (termf_9[27:27], i_0r1[27:27]);
  BUFF I643 (termt_9[28:28], i_0r0[28:28]);
  BUFF I644 (termf_9[28:28], i_0r1[28:28]);
  BUFF I645 (termt_9[29:29], i_0r0[29:29]);
  BUFF I646 (termf_9[29:29], i_0r1[29:29]);
  BUFF I647 (termt_9[30:30], i_0r0[30:30]);
  BUFF I648 (termf_9[30:30], i_0r1[30:30]);
  BUFF I649 (termt_9[31:31], i_0r0[31:31]);
  BUFF I650 (termf_9[31:31], i_0r1[31:31]);
  OR2 I651 (comp100_0[0:0], termf_9[0:0], termt_9[0:0]);
  OR2 I652 (comp100_0[1:1], termf_9[1:1], termt_9[1:1]);
  OR2 I653 (comp100_0[2:2], termf_9[2:2], termt_9[2:2]);
  OR2 I654 (comp100_0[3:3], termf_9[3:3], termt_9[3:3]);
  OR2 I655 (comp100_0[4:4], termf_9[4:4], termt_9[4:4]);
  OR2 I656 (comp100_0[5:5], termf_9[5:5], termt_9[5:5]);
  OR2 I657 (comp100_0[6:6], termf_9[6:6], termt_9[6:6]);
  OR2 I658 (comp100_0[7:7], termf_9[7:7], termt_9[7:7]);
  OR2 I659 (comp100_0[8:8], termf_9[8:8], termt_9[8:8]);
  OR2 I660 (comp100_0[9:9], termf_9[9:9], termt_9[9:9]);
  OR2 I661 (comp100_0[10:10], termf_9[10:10], termt_9[10:10]);
  OR2 I662 (comp100_0[11:11], termf_9[11:11], termt_9[11:11]);
  OR2 I663 (comp100_0[12:12], termf_9[12:12], termt_9[12:12]);
  OR2 I664 (comp100_0[13:13], termf_9[13:13], termt_9[13:13]);
  OR2 I665 (comp100_0[14:14], termf_9[14:14], termt_9[14:14]);
  OR2 I666 (comp100_0[15:15], termf_9[15:15], termt_9[15:15]);
  OR2 I667 (comp100_0[16:16], termf_9[16:16], termt_9[16:16]);
  OR2 I668 (comp100_0[17:17], termf_9[17:17], termt_9[17:17]);
  OR2 I669 (comp100_0[18:18], termf_9[18:18], termt_9[18:18]);
  OR2 I670 (comp100_0[19:19], termf_9[19:19], termt_9[19:19]);
  OR2 I671 (comp100_0[20:20], termf_9[20:20], termt_9[20:20]);
  OR2 I672 (comp100_0[21:21], termf_9[21:21], termt_9[21:21]);
  OR2 I673 (comp100_0[22:22], termf_9[22:22], termt_9[22:22]);
  OR2 I674 (comp100_0[23:23], termf_9[23:23], termt_9[23:23]);
  OR2 I675 (comp100_0[24:24], termf_9[24:24], termt_9[24:24]);
  OR2 I676 (comp100_0[25:25], termf_9[25:25], termt_9[25:25]);
  OR2 I677 (comp100_0[26:26], termf_9[26:26], termt_9[26:26]);
  OR2 I678 (comp100_0[27:27], termf_9[27:27], termt_9[27:27]);
  OR2 I679 (comp100_0[28:28], termf_9[28:28], termt_9[28:28]);
  OR2 I680 (comp100_0[29:29], termf_9[29:29], termt_9[29:29]);
  OR2 I681 (comp100_0[30:30], termf_9[30:30], termt_9[30:30]);
  OR2 I682 (comp100_0[31:31], termf_9[31:31], termt_9[31:31]);
  C3 I683 (simp6711_0[0:0], comp100_0[0:0], comp100_0[1:1], comp100_0[2:2]);
  C3 I684 (simp6711_0[1:1], comp100_0[3:3], comp100_0[4:4], comp100_0[5:5]);
  C3 I685 (simp6711_0[2:2], comp100_0[6:6], comp100_0[7:7], comp100_0[8:8]);
  C3 I686 (simp6711_0[3:3], comp100_0[9:9], comp100_0[10:10], comp100_0[11:11]);
  C3 I687 (simp6711_0[4:4], comp100_0[12:12], comp100_0[13:13], comp100_0[14:14]);
  C3 I688 (simp6711_0[5:5], comp100_0[15:15], comp100_0[16:16], comp100_0[17:17]);
  C3 I689 (simp6711_0[6:6], comp100_0[18:18], comp100_0[19:19], comp100_0[20:20]);
  C3 I690 (simp6711_0[7:7], comp100_0[21:21], comp100_0[22:22], comp100_0[23:23]);
  C3 I691 (simp6711_0[8:8], comp100_0[24:24], comp100_0[25:25], comp100_0[26:26]);
  C3 I692 (simp6711_0[9:9], comp100_0[27:27], comp100_0[28:28], comp100_0[29:29]);
  C2 I693 (simp6711_0[10:10], comp100_0[30:30], comp100_0[31:31]);
  C3 I694 (simp6712_0[0:0], simp6711_0[0:0], simp6711_0[1:1], simp6711_0[2:2]);
  C3 I695 (simp6712_0[1:1], simp6711_0[3:3], simp6711_0[4:4], simp6711_0[5:5]);
  C3 I696 (simp6712_0[2:2], simp6711_0[6:6], simp6711_0[7:7], simp6711_0[8:8]);
  C2 I697 (simp6712_0[3:3], simp6711_0[9:9], simp6711_0[10:10]);
  C3 I698 (simp6713_0[0:0], simp6712_0[0:0], simp6712_0[1:1], simp6712_0[2:2]);
  BUFF I699 (simp6713_0[1:1], simp6712_0[3:3]);
  C2 I700 (selcomp10_0, simp6713_0[0:0], simp6713_0[1:1]);
  OR2 I701 (comp101_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I702 (comp101_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I703 (comp101_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I704 (comp101_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I705 (comp101_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I706 (comp101_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I707 (comp101_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I708 (comp101_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I709 (comp101_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I710 (comp101_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I711 (comp101_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I712 (comp101_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I713 (comp101_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I714 (comp101_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I715 (comp101_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I716 (comp101_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I717 (comp101_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I718 (comp101_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I719 (comp101_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I720 (comp101_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I721 (comp101_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I722 (comp101_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I723 (comp101_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I724 (comp101_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I725 (comp101_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I726 (comp101_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I727 (comp101_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I728 (comp101_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I729 (comp101_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I730 (comp101_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I731 (comp101_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I732 (comp101_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  C3 I733 (simp7051_0[0:0], comp101_0[0:0], comp101_0[1:1], comp101_0[2:2]);
  C3 I734 (simp7051_0[1:1], comp101_0[3:3], comp101_0[4:4], comp101_0[5:5]);
  C3 I735 (simp7051_0[2:2], comp101_0[6:6], comp101_0[7:7], comp101_0[8:8]);
  C3 I736 (simp7051_0[3:3], comp101_0[9:9], comp101_0[10:10], comp101_0[11:11]);
  C3 I737 (simp7051_0[4:4], comp101_0[12:12], comp101_0[13:13], comp101_0[14:14]);
  C3 I738 (simp7051_0[5:5], comp101_0[15:15], comp101_0[16:16], comp101_0[17:17]);
  C3 I739 (simp7051_0[6:6], comp101_0[18:18], comp101_0[19:19], comp101_0[20:20]);
  C3 I740 (simp7051_0[7:7], comp101_0[21:21], comp101_0[22:22], comp101_0[23:23]);
  C3 I741 (simp7051_0[8:8], comp101_0[24:24], comp101_0[25:25], comp101_0[26:26]);
  C3 I742 (simp7051_0[9:9], comp101_0[27:27], comp101_0[28:28], comp101_0[29:29]);
  C2 I743 (simp7051_0[10:10], comp101_0[30:30], comp101_0[31:31]);
  C3 I744 (simp7052_0[0:0], simp7051_0[0:0], simp7051_0[1:1], simp7051_0[2:2]);
  C3 I745 (simp7052_0[1:1], simp7051_0[3:3], simp7051_0[4:4], simp7051_0[5:5]);
  C3 I746 (simp7052_0[2:2], simp7051_0[6:6], simp7051_0[7:7], simp7051_0[8:8]);
  C2 I747 (simp7052_0[3:3], simp7051_0[9:9], simp7051_0[10:10]);
  C3 I748 (simp7053_0[0:0], simp7052_0[0:0], simp7052_0[1:1], simp7052_0[2:2]);
  BUFF I749 (simp7053_0[1:1], simp7052_0[3:3]);
  C2 I750 (selcomp10_1, simp7053_0[0:0], simp7053_0[1:1]);
  OR2 I751 (dcomp10_0[0:0], termf_6[0:0], termt_6[0:0]);
  OR2 I752 (dcomp10_0[1:1], termf_6[1:1], termt_6[1:1]);
  C2 I753 (scomplete10_0, dcomp10_0[0:0], dcomp10_0[1:1]);
  C3 I754 (icomplete10_0, scomplete10_0, selcomp10_0, selcomp10_1);
  OR2 I755 (termf_10[0:0], gfint10_0[0:0], gfint10_1[0:0]);
  OR2 I756 (termf_10[1:1], gfint10_0[1:1], gfint10_1[1:1]);
  OR2 I757 (termf_10[2:2], gfint10_0[2:2], gfint10_1[2:2]);
  OR2 I758 (termf_10[3:3], gfint10_0[3:3], gfint10_1[3:3]);
  OR2 I759 (termf_10[4:4], gfint10_0[4:4], gfint10_1[4:4]);
  OR2 I760 (termf_10[5:5], gfint10_0[5:5], gfint10_1[5:5]);
  OR2 I761 (termf_10[6:6], gfint10_0[6:6], gfint10_1[6:6]);
  OR2 I762 (termf_10[7:7], gfint10_0[7:7], gfint10_1[7:7]);
  OR2 I763 (termf_10[8:8], gfint10_0[8:8], gfint10_1[8:8]);
  OR2 I764 (termf_10[9:9], gfint10_0[9:9], gfint10_1[9:9]);
  OR2 I765 (termf_10[10:10], gfint10_0[10:10], gfint10_1[10:10]);
  OR2 I766 (termf_10[11:11], gfint10_0[11:11], gfint10_1[11:11]);
  OR2 I767 (termf_10[12:12], gfint10_0[12:12], gfint10_1[12:12]);
  OR2 I768 (termf_10[13:13], gfint10_0[13:13], gfint10_1[13:13]);
  OR2 I769 (termf_10[14:14], gfint10_0[14:14], gfint10_1[14:14]);
  OR2 I770 (termf_10[15:15], gfint10_0[15:15], gfint10_1[15:15]);
  OR2 I771 (termf_10[16:16], gfint10_0[16:16], gfint10_1[16:16]);
  OR2 I772 (termf_10[17:17], gfint10_0[17:17], gfint10_1[17:17]);
  OR2 I773 (termf_10[18:18], gfint10_0[18:18], gfint10_1[18:18]);
  OR2 I774 (termf_10[19:19], gfint10_0[19:19], gfint10_1[19:19]);
  OR2 I775 (termf_10[20:20], gfint10_0[20:20], gfint10_1[20:20]);
  OR2 I776 (termf_10[21:21], gfint10_0[21:21], gfint10_1[21:21]);
  OR2 I777 (termf_10[22:22], gfint10_0[22:22], gfint10_1[22:22]);
  OR2 I778 (termf_10[23:23], gfint10_0[23:23], gfint10_1[23:23]);
  OR2 I779 (termf_10[24:24], gfint10_0[24:24], gfint10_1[24:24]);
  OR2 I780 (termf_10[25:25], gfint10_0[25:25], gfint10_1[25:25]);
  OR2 I781 (termf_10[26:26], gfint10_0[26:26], gfint10_1[26:26]);
  OR2 I782 (termf_10[27:27], gfint10_0[27:27], gfint10_1[27:27]);
  OR2 I783 (termf_10[28:28], gfint10_0[28:28], gfint10_1[28:28]);
  OR2 I784 (termf_10[29:29], gfint10_0[29:29], gfint10_1[29:29]);
  OR2 I785 (termf_10[30:30], gfint10_0[30:30], gfint10_1[30:30]);
  OR2 I786 (termf_10[31:31], gfint10_0[31:31], gfint10_1[31:31]);
  OR2 I787 (termt_10[0:0], gtint10_0[0:0], gtint10_1[0:0]);
  OR2 I788 (termt_10[1:1], gtint10_0[1:1], gtint10_1[1:1]);
  OR2 I789 (termt_10[2:2], gtint10_0[2:2], gtint10_1[2:2]);
  OR2 I790 (termt_10[3:3], gtint10_0[3:3], gtint10_1[3:3]);
  OR2 I791 (termt_10[4:4], gtint10_0[4:4], gtint10_1[4:4]);
  OR2 I792 (termt_10[5:5], gtint10_0[5:5], gtint10_1[5:5]);
  OR2 I793 (termt_10[6:6], gtint10_0[6:6], gtint10_1[6:6]);
  OR2 I794 (termt_10[7:7], gtint10_0[7:7], gtint10_1[7:7]);
  OR2 I795 (termt_10[8:8], gtint10_0[8:8], gtint10_1[8:8]);
  OR2 I796 (termt_10[9:9], gtint10_0[9:9], gtint10_1[9:9]);
  OR2 I797 (termt_10[10:10], gtint10_0[10:10], gtint10_1[10:10]);
  OR2 I798 (termt_10[11:11], gtint10_0[11:11], gtint10_1[11:11]);
  OR2 I799 (termt_10[12:12], gtint10_0[12:12], gtint10_1[12:12]);
  OR2 I800 (termt_10[13:13], gtint10_0[13:13], gtint10_1[13:13]);
  OR2 I801 (termt_10[14:14], gtint10_0[14:14], gtint10_1[14:14]);
  OR2 I802 (termt_10[15:15], gtint10_0[15:15], gtint10_1[15:15]);
  OR2 I803 (termt_10[16:16], gtint10_0[16:16], gtint10_1[16:16]);
  OR2 I804 (termt_10[17:17], gtint10_0[17:17], gtint10_1[17:17]);
  OR2 I805 (termt_10[18:18], gtint10_0[18:18], gtint10_1[18:18]);
  OR2 I806 (termt_10[19:19], gtint10_0[19:19], gtint10_1[19:19]);
  OR2 I807 (termt_10[20:20], gtint10_0[20:20], gtint10_1[20:20]);
  OR2 I808 (termt_10[21:21], gtint10_0[21:21], gtint10_1[21:21]);
  OR2 I809 (termt_10[22:22], gtint10_0[22:22], gtint10_1[22:22]);
  OR2 I810 (termt_10[23:23], gtint10_0[23:23], gtint10_1[23:23]);
  OR2 I811 (termt_10[24:24], gtint10_0[24:24], gtint10_1[24:24]);
  OR2 I812 (termt_10[25:25], gtint10_0[25:25], gtint10_1[25:25]);
  OR2 I813 (termt_10[26:26], gtint10_0[26:26], gtint10_1[26:26]);
  OR2 I814 (termt_10[27:27], gtint10_0[27:27], gtint10_1[27:27]);
  OR2 I815 (termt_10[28:28], gtint10_0[28:28], gtint10_1[28:28]);
  OR2 I816 (termt_10[29:29], gtint10_0[29:29], gtint10_1[29:29]);
  OR2 I817 (termt_10[30:30], gtint10_0[30:30], gtint10_1[30:30]);
  OR2 I818 (termt_10[31:31], gtint10_0[31:31], gtint10_1[31:31]);
  C2R I819 (sel10_0, selg10_0, icomplete10_0, reset);
  C2R I820 (sel10_1, selg10_1, icomplete10_0, reset);
  C2R I821 (gfint10_0[0:0], sel10_0, termf_9[0:0], reset);
  C2R I822 (gfint10_0[1:1], sel10_0, termf_9[1:1], reset);
  C2R I823 (gfint10_0[2:2], sel10_0, termf_9[2:2], reset);
  C2R I824 (gfint10_0[3:3], sel10_0, termf_9[3:3], reset);
  C2R I825 (gfint10_0[4:4], sel10_0, termf_9[4:4], reset);
  C2R I826 (gfint10_0[5:5], sel10_0, termf_9[5:5], reset);
  C2R I827 (gfint10_0[6:6], sel10_0, termf_9[6:6], reset);
  C2R I828 (gfint10_0[7:7], sel10_0, termf_9[7:7], reset);
  C2R I829 (gfint10_0[8:8], sel10_0, termf_9[8:8], reset);
  C2R I830 (gfint10_0[9:9], sel10_0, termf_9[9:9], reset);
  C2R I831 (gfint10_0[10:10], sel10_0, termf_9[10:10], reset);
  C2R I832 (gfint10_0[11:11], sel10_0, termf_9[11:11], reset);
  C2R I833 (gfint10_0[12:12], sel10_0, termf_9[12:12], reset);
  C2R I834 (gfint10_0[13:13], sel10_0, termf_9[13:13], reset);
  C2R I835 (gfint10_0[14:14], sel10_0, termf_9[14:14], reset);
  C2R I836 (gfint10_0[15:15], sel10_0, termf_9[15:15], reset);
  C2R I837 (gfint10_0[16:16], sel10_0, termf_9[16:16], reset);
  C2R I838 (gfint10_0[17:17], sel10_0, termf_9[17:17], reset);
  C2R I839 (gfint10_0[18:18], sel10_0, termf_9[18:18], reset);
  C2R I840 (gfint10_0[19:19], sel10_0, termf_9[19:19], reset);
  C2R I841 (gfint10_0[20:20], sel10_0, termf_9[20:20], reset);
  C2R I842 (gfint10_0[21:21], sel10_0, termf_9[21:21], reset);
  C2R I843 (gfint10_0[22:22], sel10_0, termf_9[22:22], reset);
  C2R I844 (gfint10_0[23:23], sel10_0, termf_9[23:23], reset);
  C2R I845 (gfint10_0[24:24], sel10_0, termf_9[24:24], reset);
  C2R I846 (gfint10_0[25:25], sel10_0, termf_9[25:25], reset);
  C2R I847 (gfint10_0[26:26], sel10_0, termf_9[26:26], reset);
  C2R I848 (gfint10_0[27:27], sel10_0, termf_9[27:27], reset);
  C2R I849 (gfint10_0[28:28], sel10_0, termf_9[28:28], reset);
  C2R I850 (gfint10_0[29:29], sel10_0, termf_9[29:29], reset);
  C2R I851 (gfint10_0[30:30], sel10_0, termf_9[30:30], reset);
  C2R I852 (gfint10_0[31:31], sel10_0, termf_9[31:31], reset);
  C2R I853 (gfint10_1[0:0], sel10_1, i_0r0[0:0], reset);
  C2R I854 (gfint10_1[1:1], sel10_1, i_0r0[1:1], reset);
  C2R I855 (gfint10_1[2:2], sel10_1, i_0r0[2:2], reset);
  C2R I856 (gfint10_1[3:3], sel10_1, i_0r0[3:3], reset);
  C2R I857 (gfint10_1[4:4], sel10_1, i_0r0[4:4], reset);
  C2R I858 (gfint10_1[5:5], sel10_1, i_0r0[5:5], reset);
  C2R I859 (gfint10_1[6:6], sel10_1, i_0r0[6:6], reset);
  C2R I860 (gfint10_1[7:7], sel10_1, i_0r0[7:7], reset);
  C2R I861 (gfint10_1[8:8], sel10_1, i_0r0[8:8], reset);
  C2R I862 (gfint10_1[9:9], sel10_1, i_0r0[9:9], reset);
  C2R I863 (gfint10_1[10:10], sel10_1, i_0r0[10:10], reset);
  C2R I864 (gfint10_1[11:11], sel10_1, i_0r0[11:11], reset);
  C2R I865 (gfint10_1[12:12], sel10_1, i_0r0[12:12], reset);
  C2R I866 (gfint10_1[13:13], sel10_1, i_0r0[13:13], reset);
  C2R I867 (gfint10_1[14:14], sel10_1, i_0r0[14:14], reset);
  C2R I868 (gfint10_1[15:15], sel10_1, i_0r0[15:15], reset);
  C2R I869 (gfint10_1[16:16], sel10_1, i_0r0[16:16], reset);
  C2R I870 (gfint10_1[17:17], sel10_1, i_0r0[17:17], reset);
  C2R I871 (gfint10_1[18:18], sel10_1, i_0r0[18:18], reset);
  C2R I872 (gfint10_1[19:19], sel10_1, i_0r0[19:19], reset);
  C2R I873 (gfint10_1[20:20], sel10_1, i_0r0[20:20], reset);
  C2R I874 (gfint10_1[21:21], sel10_1, i_0r0[21:21], reset);
  C2R I875 (gfint10_1[22:22], sel10_1, i_0r0[22:22], reset);
  C2R I876 (gfint10_1[23:23], sel10_1, i_0r0[23:23], reset);
  C2R I877 (gfint10_1[24:24], sel10_1, i_0r0[24:24], reset);
  C2R I878 (gfint10_1[25:25], sel10_1, i_0r0[25:25], reset);
  C2R I879 (gfint10_1[26:26], sel10_1, i_0r0[26:26], reset);
  C2R I880 (gfint10_1[27:27], sel10_1, i_0r0[27:27], reset);
  C2R I881 (gfint10_1[28:28], sel10_1, i_0r0[28:28], reset);
  C2R I882 (gfint10_1[29:29], sel10_1, i_0r0[29:29], reset);
  C2R I883 (gfint10_1[30:30], sel10_1, i_0r0[30:30], reset);
  C2R I884 (gfint10_1[31:31], sel10_1, i_0r0[31:31], reset);
  C2R I885 (gtint10_0[0:0], sel10_0, termt_9[0:0], reset);
  C2R I886 (gtint10_0[1:1], sel10_0, termt_9[1:1], reset);
  C2R I887 (gtint10_0[2:2], sel10_0, termt_9[2:2], reset);
  C2R I888 (gtint10_0[3:3], sel10_0, termt_9[3:3], reset);
  C2R I889 (gtint10_0[4:4], sel10_0, termt_9[4:4], reset);
  C2R I890 (gtint10_0[5:5], sel10_0, termt_9[5:5], reset);
  C2R I891 (gtint10_0[6:6], sel10_0, termt_9[6:6], reset);
  C2R I892 (gtint10_0[7:7], sel10_0, termt_9[7:7], reset);
  C2R I893 (gtint10_0[8:8], sel10_0, termt_9[8:8], reset);
  C2R I894 (gtint10_0[9:9], sel10_0, termt_9[9:9], reset);
  C2R I895 (gtint10_0[10:10], sel10_0, termt_9[10:10], reset);
  C2R I896 (gtint10_0[11:11], sel10_0, termt_9[11:11], reset);
  C2R I897 (gtint10_0[12:12], sel10_0, termt_9[12:12], reset);
  C2R I898 (gtint10_0[13:13], sel10_0, termt_9[13:13], reset);
  C2R I899 (gtint10_0[14:14], sel10_0, termt_9[14:14], reset);
  C2R I900 (gtint10_0[15:15], sel10_0, termt_9[15:15], reset);
  C2R I901 (gtint10_0[16:16], sel10_0, termt_9[16:16], reset);
  C2R I902 (gtint10_0[17:17], sel10_0, termt_9[17:17], reset);
  C2R I903 (gtint10_0[18:18], sel10_0, termt_9[18:18], reset);
  C2R I904 (gtint10_0[19:19], sel10_0, termt_9[19:19], reset);
  C2R I905 (gtint10_0[20:20], sel10_0, termt_9[20:20], reset);
  C2R I906 (gtint10_0[21:21], sel10_0, termt_9[21:21], reset);
  C2R I907 (gtint10_0[22:22], sel10_0, termt_9[22:22], reset);
  C2R I908 (gtint10_0[23:23], sel10_0, termt_9[23:23], reset);
  C2R I909 (gtint10_0[24:24], sel10_0, termt_9[24:24], reset);
  C2R I910 (gtint10_0[25:25], sel10_0, termt_9[25:25], reset);
  C2R I911 (gtint10_0[26:26], sel10_0, termt_9[26:26], reset);
  C2R I912 (gtint10_0[27:27], sel10_0, termt_9[27:27], reset);
  C2R I913 (gtint10_0[28:28], sel10_0, termt_9[28:28], reset);
  C2R I914 (gtint10_0[29:29], sel10_0, termt_9[29:29], reset);
  C2R I915 (gtint10_0[30:30], sel10_0, termt_9[30:30], reset);
  C2R I916 (gtint10_0[31:31], sel10_0, termt_9[31:31], reset);
  C2R I917 (gtint10_1[0:0], sel10_1, i_0r1[0:0], reset);
  C2R I918 (gtint10_1[1:1], sel10_1, i_0r1[1:1], reset);
  C2R I919 (gtint10_1[2:2], sel10_1, i_0r1[2:2], reset);
  C2R I920 (gtint10_1[3:3], sel10_1, i_0r1[3:3], reset);
  C2R I921 (gtint10_1[4:4], sel10_1, i_0r1[4:4], reset);
  C2R I922 (gtint10_1[5:5], sel10_1, i_0r1[5:5], reset);
  C2R I923 (gtint10_1[6:6], sel10_1, i_0r1[6:6], reset);
  C2R I924 (gtint10_1[7:7], sel10_1, i_0r1[7:7], reset);
  C2R I925 (gtint10_1[8:8], sel10_1, i_0r1[8:8], reset);
  C2R I926 (gtint10_1[9:9], sel10_1, i_0r1[9:9], reset);
  C2R I927 (gtint10_1[10:10], sel10_1, i_0r1[10:10], reset);
  C2R I928 (gtint10_1[11:11], sel10_1, i_0r1[11:11], reset);
  C2R I929 (gtint10_1[12:12], sel10_1, i_0r1[12:12], reset);
  C2R I930 (gtint10_1[13:13], sel10_1, i_0r1[13:13], reset);
  C2R I931 (gtint10_1[14:14], sel10_1, i_0r1[14:14], reset);
  C2R I932 (gtint10_1[15:15], sel10_1, i_0r1[15:15], reset);
  C2R I933 (gtint10_1[16:16], sel10_1, i_0r1[16:16], reset);
  C2R I934 (gtint10_1[17:17], sel10_1, i_0r1[17:17], reset);
  C2R I935 (gtint10_1[18:18], sel10_1, i_0r1[18:18], reset);
  C2R I936 (gtint10_1[19:19], sel10_1, i_0r1[19:19], reset);
  C2R I937 (gtint10_1[20:20], sel10_1, i_0r1[20:20], reset);
  C2R I938 (gtint10_1[21:21], sel10_1, i_0r1[21:21], reset);
  C2R I939 (gtint10_1[22:22], sel10_1, i_0r1[22:22], reset);
  C2R I940 (gtint10_1[23:23], sel10_1, i_0r1[23:23], reset);
  C2R I941 (gtint10_1[24:24], sel10_1, i_0r1[24:24], reset);
  C2R I942 (gtint10_1[25:25], sel10_1, i_0r1[25:25], reset);
  C2R I943 (gtint10_1[26:26], sel10_1, i_0r1[26:26], reset);
  C2R I944 (gtint10_1[27:27], sel10_1, i_0r1[27:27], reset);
  C2R I945 (gtint10_1[28:28], sel10_1, i_0r1[28:28], reset);
  C2R I946 (gtint10_1[29:29], sel10_1, i_0r1[29:29], reset);
  C2R I947 (gtint10_1[30:30], sel10_1, i_0r1[30:30], reset);
  C2R I948 (gtint10_1[31:31], sel10_1, i_0r1[31:31], reset);
  BUFF I949 (selg10_0, match100_0);
  C2 I950 (match100_0, termf_6[0:0], termt_6[1:1]);
  BUFF I951 (selg10_1, match101_0);
  C2 I952 (match101_0, termt_6[0:0], termf_6[1:1]);
  BUFF I953 (o_0r0[0:0], termf_10[0:0]);
  BUFF I954 (o_0r0[1:1], termf_10[1:1]);
  BUFF I955 (o_0r0[2:2], termf_10[2:2]);
  BUFF I956 (o_0r0[3:3], termf_10[3:3]);
  BUFF I957 (o_0r0[4:4], termf_10[4:4]);
  BUFF I958 (o_0r0[5:5], termf_10[5:5]);
  BUFF I959 (o_0r0[6:6], termf_10[6:6]);
  BUFF I960 (o_0r0[7:7], termf_10[7:7]);
  BUFF I961 (o_0r0[8:8], termf_10[8:8]);
  BUFF I962 (o_0r0[9:9], termf_10[9:9]);
  BUFF I963 (o_0r0[10:10], termf_10[10:10]);
  BUFF I964 (o_0r0[11:11], termf_10[11:11]);
  BUFF I965 (o_0r0[12:12], termf_10[12:12]);
  BUFF I966 (o_0r0[13:13], termf_10[13:13]);
  BUFF I967 (o_0r0[14:14], termf_10[14:14]);
  BUFF I968 (o_0r0[15:15], termf_10[15:15]);
  BUFF I969 (o_0r0[16:16], termf_10[16:16]);
  BUFF I970 (o_0r0[17:17], termf_10[17:17]);
  BUFF I971 (o_0r0[18:18], termf_10[18:18]);
  BUFF I972 (o_0r0[19:19], termf_10[19:19]);
  BUFF I973 (o_0r0[20:20], termf_10[20:20]);
  BUFF I974 (o_0r0[21:21], termf_10[21:21]);
  BUFF I975 (o_0r0[22:22], termf_10[22:22]);
  BUFF I976 (o_0r0[23:23], termf_10[23:23]);
  BUFF I977 (o_0r0[24:24], termf_10[24:24]);
  BUFF I978 (o_0r0[25:25], termf_10[25:25]);
  BUFF I979 (o_0r0[26:26], termf_10[26:26]);
  BUFF I980 (o_0r0[27:27], termf_10[27:27]);
  BUFF I981 (o_0r0[28:28], termf_10[28:28]);
  BUFF I982 (o_0r0[29:29], termf_10[29:29]);
  BUFF I983 (o_0r0[30:30], termf_10[30:30]);
  BUFF I984 (o_0r0[31:31], termf_10[31:31]);
  BUFF I985 (o_0r0[32:32], termf_8[0:0]);
  BUFF I986 (o_0r0[33:33], termf_8[1:1]);
  BUFF I987 (o_0r0[34:34], termf_8[2:2]);
  BUFF I988 (o_0r0[35:35], termf_8[3:3]);
  BUFF I989 (o_0r0[36:36], termf_8[4:4]);
  BUFF I990 (o_0r0[37:37], termf_8[5:5]);
  BUFF I991 (o_0r0[38:38], termf_8[6:6]);
  BUFF I992 (o_0r0[39:39], termf_8[7:7]);
  BUFF I993 (o_0r0[40:40], termf_8[8:8]);
  BUFF I994 (o_0r0[41:41], termf_8[9:9]);
  BUFF I995 (o_0r0[42:42], termf_8[10:10]);
  BUFF I996 (o_0r0[43:43], termf_8[11:11]);
  BUFF I997 (o_0r0[44:44], termf_8[12:12]);
  BUFF I998 (o_0r0[45:45], termf_8[13:13]);
  BUFF I999 (o_0r0[46:46], termf_8[14:14]);
  BUFF I1000 (o_0r0[47:47], termf_8[15:15]);
  BUFF I1001 (o_0r0[48:48], termf_8[16:16]);
  BUFF I1002 (o_0r0[49:49], termf_8[17:17]);
  BUFF I1003 (o_0r0[50:50], termf_8[18:18]);
  BUFF I1004 (o_0r0[51:51], termf_8[19:19]);
  BUFF I1005 (o_0r0[52:52], termf_8[20:20]);
  BUFF I1006 (o_0r0[53:53], termf_8[21:21]);
  BUFF I1007 (o_0r0[54:54], termf_8[22:22]);
  BUFF I1008 (o_0r0[55:55], termf_8[23:23]);
  BUFF I1009 (o_0r0[56:56], termf_8[24:24]);
  BUFF I1010 (o_0r0[57:57], termf_8[25:25]);
  BUFF I1011 (o_0r0[58:58], termf_8[26:26]);
  BUFF I1012 (o_0r0[59:59], termf_8[27:27]);
  BUFF I1013 (o_0r0[60:60], termf_8[28:28]);
  BUFF I1014 (o_0r0[61:61], termf_8[29:29]);
  BUFF I1015 (o_0r0[62:62], termf_8[30:30]);
  BUFF I1016 (o_0r0[63:63], termf_8[31:31]);
  BUFF I1017 (o_0r0[64:64], i_0r0[68:68]);
  BUFF I1018 (o_0r1[0:0], termt_10[0:0]);
  BUFF I1019 (o_0r1[1:1], termt_10[1:1]);
  BUFF I1020 (o_0r1[2:2], termt_10[2:2]);
  BUFF I1021 (o_0r1[3:3], termt_10[3:3]);
  BUFF I1022 (o_0r1[4:4], termt_10[4:4]);
  BUFF I1023 (o_0r1[5:5], termt_10[5:5]);
  BUFF I1024 (o_0r1[6:6], termt_10[6:6]);
  BUFF I1025 (o_0r1[7:7], termt_10[7:7]);
  BUFF I1026 (o_0r1[8:8], termt_10[8:8]);
  BUFF I1027 (o_0r1[9:9], termt_10[9:9]);
  BUFF I1028 (o_0r1[10:10], termt_10[10:10]);
  BUFF I1029 (o_0r1[11:11], termt_10[11:11]);
  BUFF I1030 (o_0r1[12:12], termt_10[12:12]);
  BUFF I1031 (o_0r1[13:13], termt_10[13:13]);
  BUFF I1032 (o_0r1[14:14], termt_10[14:14]);
  BUFF I1033 (o_0r1[15:15], termt_10[15:15]);
  BUFF I1034 (o_0r1[16:16], termt_10[16:16]);
  BUFF I1035 (o_0r1[17:17], termt_10[17:17]);
  BUFF I1036 (o_0r1[18:18], termt_10[18:18]);
  BUFF I1037 (o_0r1[19:19], termt_10[19:19]);
  BUFF I1038 (o_0r1[20:20], termt_10[20:20]);
  BUFF I1039 (o_0r1[21:21], termt_10[21:21]);
  BUFF I1040 (o_0r1[22:22], termt_10[22:22]);
  BUFF I1041 (o_0r1[23:23], termt_10[23:23]);
  BUFF I1042 (o_0r1[24:24], termt_10[24:24]);
  BUFF I1043 (o_0r1[25:25], termt_10[25:25]);
  BUFF I1044 (o_0r1[26:26], termt_10[26:26]);
  BUFF I1045 (o_0r1[27:27], termt_10[27:27]);
  BUFF I1046 (o_0r1[28:28], termt_10[28:28]);
  BUFF I1047 (o_0r1[29:29], termt_10[29:29]);
  BUFF I1048 (o_0r1[30:30], termt_10[30:30]);
  BUFF I1049 (o_0r1[31:31], termt_10[31:31]);
  BUFF I1050 (o_0r1[32:32], termt_8[0:0]);
  BUFF I1051 (o_0r1[33:33], termt_8[1:1]);
  BUFF I1052 (o_0r1[34:34], termt_8[2:2]);
  BUFF I1053 (o_0r1[35:35], termt_8[3:3]);
  BUFF I1054 (o_0r1[36:36], termt_8[4:4]);
  BUFF I1055 (o_0r1[37:37], termt_8[5:5]);
  BUFF I1056 (o_0r1[38:38], termt_8[6:6]);
  BUFF I1057 (o_0r1[39:39], termt_8[7:7]);
  BUFF I1058 (o_0r1[40:40], termt_8[8:8]);
  BUFF I1059 (o_0r1[41:41], termt_8[9:9]);
  BUFF I1060 (o_0r1[42:42], termt_8[10:10]);
  BUFF I1061 (o_0r1[43:43], termt_8[11:11]);
  BUFF I1062 (o_0r1[44:44], termt_8[12:12]);
  BUFF I1063 (o_0r1[45:45], termt_8[13:13]);
  BUFF I1064 (o_0r1[46:46], termt_8[14:14]);
  BUFF I1065 (o_0r1[47:47], termt_8[15:15]);
  BUFF I1066 (o_0r1[48:48], termt_8[16:16]);
  BUFF I1067 (o_0r1[49:49], termt_8[17:17]);
  BUFF I1068 (o_0r1[50:50], termt_8[18:18]);
  BUFF I1069 (o_0r1[51:51], termt_8[19:19]);
  BUFF I1070 (o_0r1[52:52], termt_8[20:20]);
  BUFF I1071 (o_0r1[53:53], termt_8[21:21]);
  BUFF I1072 (o_0r1[54:54], termt_8[22:22]);
  BUFF I1073 (o_0r1[55:55], termt_8[23:23]);
  BUFF I1074 (o_0r1[56:56], termt_8[24:24]);
  BUFF I1075 (o_0r1[57:57], termt_8[25:25]);
  BUFF I1076 (o_0r1[58:58], termt_8[26:26]);
  BUFF I1077 (o_0r1[59:59], termt_8[27:27]);
  BUFF I1078 (o_0r1[60:60], termt_8[28:28]);
  BUFF I1079 (o_0r1[61:61], termt_8[29:29]);
  BUFF I1080 (o_0r1[62:62], termt_8[30:30]);
  BUFF I1081 (o_0r1[63:63], termt_8[31:31]);
  BUFF I1082 (o_0r1[64:64], i_0r1[68:68]);
  BUFF I1083 (i_0a, o_0a);
endmodule

// tki TeakI [One 0,One 0]
module tki (i_0r, i_0a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  input reset;
  wire nreset_0;
  wire firsthsa_0;
  wire nfirsthsa_0;
  wire firsthsd_0;
  wire noa_0;
  INV I0 (nreset_0, reset);
  INV I1 (nfirsthsa_0, firsthsa_0);
  INV I2 (noa_0, o_0a);
  AO22 I3 (o_0r, nreset_0, nfirsthsa_0, i_0r, firsthsd_0);
  AO22 I4 (firsthsa_0, nreset_0, o_0a, nreset_0, firsthsa_0);
  AO22 I5 (firsthsd_0, firsthsa_0, noa_0, firsthsa_0, firsthsd_0);
  AND2 I6 (i_0a, o_0a, firsthsd_0);
endmodule

module teak_nanoAlu (a_0r0, a_0r1, a_0a, b_0r0, b_0r1, b_0a, ctrl_0r0, ctrl_0r1, ctrl_0a, fi_0r0, fi_0r1, fi_0a, sfc_0r0, sfc_0r1, sfc_0a, o_0r0, o_0r1, o_0a, f_0r0, f_0r1, f_0a, reset);
  input [31:0] a_0r0;
  input [31:0] a_0r1;
  output a_0a;
  input [31:0] b_0r0;
  input [31:0] b_0r1;
  output b_0a;
  input [3:0] ctrl_0r0;
  input [3:0] ctrl_0r1;
  output ctrl_0a;
  input [3:0] fi_0r0;
  input [3:0] fi_0r1;
  output fi_0a;
  input sfc_0r0;
  input sfc_0r1;
  output sfc_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  output [3:0] f_0r0;
  output [3:0] f_0r1;
  input f_0a;
  input reset;
  wire L59_0r;
  wire L59_0a;
  wire [3:0] L60_0r0;
  wire [3:0] L60_0r1;
  wire L60_0a;
  wire L62_0r;
  wire L62_0a;
  wire L63_0r0;
  wire L63_0r1;
  wire L63_0a;
  wire L64_0r;
  wire L64_0a;
  wire [31:0] L65_0r0;
  wire [31:0] L65_0r1;
  wire L65_0a;
  wire L67_0r;
  wire L67_0a;
  wire L68_0r0;
  wire L68_0r1;
  wire L68_0a;
  wire L69_0r;
  wire L69_0a;
  wire [31:0] L70_0r0;
  wire [31:0] L70_0r1;
  wire L70_0a;
  wire [65:0] L72_0r0;
  wire [65:0] L72_0r1;
  wire L72_0a;
  wire L74_0r;
  wire L74_0a;
  wire L77_0r;
  wire L77_0a;
  wire [31:0] L78_0r0;
  wire [31:0] L78_0r1;
  wire L78_0a;
  wire L79_0r;
  wire L79_0a;
  wire L80_0r0;
  wire L80_0r1;
  wire L80_0a;
  wire L82_0r;
  wire L82_0a;
  wire L85_0r;
  wire L85_0a;
  wire [31:0] L86_0r0;
  wire [31:0] L86_0r1;
  wire L86_0a;
  wire L87_0r;
  wire L87_0a;
  wire [31:0] L88_0r0;
  wire [31:0] L88_0r1;
  wire L88_0a;
  wire L91_0r;
  wire L91_0a;
  wire L92_0r0;
  wire L92_0r1;
  wire L92_0a;
  wire L94_0r;
  wire L94_0a;
  wire L97_0r;
  wire L97_0a;
  wire [31:0] L98_0r0;
  wire [31:0] L98_0r1;
  wire L98_0a;
  wire L99_0r;
  wire L99_0a;
  wire [31:0] L100_0r0;
  wire [31:0] L100_0r1;
  wire L100_0a;
  wire L103_0r;
  wire L103_0a;
  wire L104_0r0;
  wire L104_0r1;
  wire L104_0a;
  wire L106_0r;
  wire L106_0a;
  wire L109_0r;
  wire L109_0a;
  wire [31:0] L110_0r0;
  wire [31:0] L110_0r1;
  wire L110_0a;
  wire L111_0r;
  wire L111_0a;
  wire [31:0] L112_0r0;
  wire [31:0] L112_0r1;
  wire L112_0a;
  wire L115_0r;
  wire L115_0a;
  wire L116_0r0;
  wire L116_0r1;
  wire L116_0a;
  wire L118_0r;
  wire L118_0a;
  wire L124_0r;
  wire L124_0a;
  wire L131_0r;
  wire L131_0a;
  wire L137_0r0;
  wire L137_0r1;
  wire L137_0a;
  wire L148_0r;
  wire L148_0a;
  wire [3:0] L149_0r0;
  wire [3:0] L149_0r1;
  wire L149_0a;
  wire L150_0r;
  wire L150_0a;
  wire L154_0r;
  wire L154_0a;
  wire L155_0r0;
  wire L155_0r1;
  wire L155_0a;
  wire L156_0r;
  wire L156_0a;
  wire L157_0r0;
  wire L157_0r1;
  wire L157_0a;
  wire L160_0r;
  wire L160_0a;
  wire L161_0r0;
  wire L161_0r1;
  wire L161_0a;
  wire L164_0r;
  wire L164_0a;
  wire L167_0r;
  wire L167_0a;
  wire L188_0r;
  wire L188_0a;
  wire L208_0r;
  wire L208_0a;
  wire L215_0r;
  wire L215_0a;
  wire [32:0] L220_0r0;
  wire [32:0] L220_0r1;
  wire L220_0a;
  wire [32:0] L222_0r0;
  wire [32:0] L222_0r1;
  wire L222_0a;
  wire [32:0] L224_0r0;
  wire [32:0] L224_0r1;
  wire L224_0a;
  wire [32:0] L226_0r0;
  wire [32:0] L226_0r1;
  wire L226_0a;
  wire [32:0] L228_0r0;
  wire [32:0] L228_0r1;
  wire L228_0a;
  wire [32:0] L231_0r0;
  wire [32:0] L231_0r1;
  wire L231_0a;
  wire L241_0r0;
  wire L241_0r1;
  wire L241_0a;
  wire L243_0r0;
  wire L243_0r1;
  wire L243_0a;
  wire L246_0r0;
  wire L246_0r1;
  wire L246_0a;
  wire L252_0r0;
  wire L252_0r1;
  wire L252_0a;
  wire L254_0r0;
  wire L254_0r1;
  wire L254_0a;
  wire L256_0r0;
  wire L256_0r1;
  wire L256_0a;
  wire [31:0] L290_0r0;
  wire [31:0] L290_0r1;
  wire L290_0a;
  wire [31:0] L295_0r0;
  wire [31:0] L295_0r1;
  wire L295_0a;
  wire [3:0] L300_0r0;
  wire [3:0] L300_0r1;
  wire L300_0a;
  wire [3:0] L301_0r0;
  wire [3:0] L301_0r1;
  wire L301_0a;
  wire L302_0r0;
  wire L302_0r1;
  wire L302_0a;
  wire [31:0] L303_0r0;
  wire [31:0] L303_0r1;
  wire L303_0a;
  wire [3:0] L304_0r0;
  wire [3:0] L304_0r1;
  wire L304_0a;
  wire [64:0] L317_0r0;
  wire [64:0] L317_0r1;
  wire L317_0a;
  wire [33:0] L321_0r0;
  wire [33:0] L321_0r1;
  wire L321_0a;
  wire [7:0] L323_0r0;
  wire [7:0] L323_0r1;
  wire L323_0a;
  wire [64:0] L325_0r0;
  wire [64:0] L325_0r1;
  wire L325_0a;
  wire [64:0] L326_0r0;
  wire [64:0] L326_0r1;
  wire L326_0a;
  wire [64:0] L327_0r0;
  wire [64:0] L327_0r1;
  wire L327_0a;
  wire [2:0] L329_0r0;
  wire [2:0] L329_0r1;
  wire L329_0a;
  wire [64:0] L336_0r0;
  wire [64:0] L336_0r1;
  wire L336_0a;
  wire [64:0] L337_0r0;
  wire [64:0] L337_0r1;
  wire L337_0a;
  wire [64:0] L338_0r0;
  wire [64:0] L338_0r1;
  wire L338_0a;
  wire L339_0r;
  wire L339_0a;
  wire L340_0r;
  wire L340_0a;
  wire L341_0r;
  wire L341_0a;
  wire [64:0] L350_0r0;
  wire [64:0] L350_0r1;
  wire L350_0a;
  wire [33:0] L360_0r0;
  wire [33:0] L360_0r1;
  wire L360_0a;
  wire [3:0] L367_0r0;
  wire [3:0] L367_0r1;
  wire L367_0a;
  wire [3:0] L369_0r0;
  wire [3:0] L369_0r1;
  wire L369_0a;
  wire [2:0] L371_0r0;
  wire [2:0] L371_0r1;
  wire L371_0a;
  wire L373_0r;
  wire L373_0a;
  wire L382_0r0;
  wire L382_0r1;
  wire L382_0a;
  wire [33:0] L383_0r0;
  wire [33:0] L383_0r1;
  wire L383_0a;
  wire L393_0r;
  wire L393_0a;
  wire L394_0r;
  wire L394_0a;
  wire L395_0r;
  wire L395_0a;
  wire L396_0r;
  wire L396_0a;
  wire L397_0r;
  wire L397_0a;
  wire [8:0] L406_0r0;
  wire [8:0] L406_0r1;
  wire L406_0a;
  wire L407_0r;
  wire L407_0a;
  wire [7:0] L410_0r0;
  wire [7:0] L410_0r1;
  wire L410_0a;
  wire [6:0] L413_0r0;
  wire [6:0] L413_0r1;
  wire L413_0a;
  wire [3:0] L421_0r0;
  wire [3:0] L421_0r1;
  wire L421_0a;
  wire [32:0] L429_0r0;
  wire [32:0] L429_0r1;
  wire L429_0a;
  wire L430_0r;
  wire L430_0a;
  wire [32:0] L431_0r0;
  wire [32:0] L431_0r1;
  wire L431_0a;
  wire [31:0] L432_0r0;
  wire [31:0] L432_0r1;
  wire L432_0a;
  wire [32:0] L433_0r0;
  wire [32:0] L433_0r1;
  wire L433_0a;
  wire [3:0] L437_0r0;
  wire [3:0] L437_0r1;
  wire L437_0a;
  wire [32:0] L442_0r0;
  wire [32:0] L442_0r1;
  wire L442_0a;
  wire [3:0] L445_0r0;
  wire [3:0] L445_0r1;
  wire L445_0a;
  wire [68:0] L446_0r0;
  wire [68:0] L446_0r1;
  wire L446_0a;
  tkj66m1_32_1_32 I0 (L63_0r0, L63_0r1, L63_0a, L65_0r0[31:0], L65_0r1[31:0], L65_0a, L68_0r0, L68_0r1, L68_0a, L70_0r0[31:0], L70_0r1[31:0], L70_0a, L72_0r0[65:0], L72_0r1[65:0], L72_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0 I1 (L74_0r, L74_0a, L62_0r, L62_0a, L64_0r, L64_0a, L67_0r, L67_0a, L69_0r, L69_0a, reset);
  tkj33m32_1 I2 (L78_0r0[31:0], L78_0r1[31:0], L78_0a, L80_0r0, L80_0r1, L80_0a, L222_0r0[32:0], L222_0r1[32:0], L222_0a, reset);
  tkf0mo0w0_o0w0 I3 (L82_0r, L82_0a, L77_0r, L77_0a, L79_0r, L79_0a, reset);
  tko65m33_1xori0w32bi32w32b_2apt1o0w32bi64w1b I4 (L336_0r0[64:0], L336_0r1[64:0], L336_0a, L224_0r0[32:0], L224_0r1[32:0], L224_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I5 (L94_0r, L94_0a, L85_0r, L85_0a, L87_0r, L87_0a, L91_0r, L91_0a, reset);
  tko65m33_1ori0w32bi32w32b_2apt1o0w32bi64w1b I6 (L337_0r0[64:0], L337_0r1[64:0], L337_0a, L226_0r0[32:0], L226_0r1[32:0], L226_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I7 (L106_0r, L106_0a, L97_0r, L97_0a, L99_0r, L99_0a, L103_0r, L103_0a, reset);
  tko65m33_1andi0w32bi32w32b_2apt1o0w32bi64w1b I8 (L338_0r0[64:0], L338_0r1[64:0], L338_0a, L228_0r0[32:0], L228_0r1[32:0], L228_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I9 (L118_0r, L118_0a, L109_0r, L109_0a, L111_0r, L111_0a, L115_0r, L115_0a, reset);
  tks4_o0w4_2m3m4m5m6m7mambo0w0_dmfo0w0_1m9o0w0_co0w0_0m8meo0w0 I10 (L60_0r0[3:0], L60_0r1[3:0], L60_0a, L74_0r, L74_0a, L82_0r, L82_0a, L94_0r, L94_0a, L106_0r, L106_0a, L118_0r, L118_0a, reset);
  tkf0mo0w0_o0w0 I11 (L131_0r, L131_0a, L124_0r, L124_0a, L59_0r, L59_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I12 (L164_0r, L164_0a, L154_0r, L154_0a, L156_0r, L156_0a, L160_0r, L160_0a, reset);
  tks4_o0w4_0c8m1c8mcmdmemfo0w0_2m3m4m5m6m7mambo0w0 I13 (L149_0r0[3:0], L149_0r1[3:0], L149_0a, L150_0r, L150_0a, L164_0r, L164_0a, reset);
  tkj0m0_0_0 I14 (L373_0r, L373_0a, L167_0r, L167_0a, L188_0r, L188_0a, L208_0r, L208_0a, reset);
  tkf65mo0w0_o0w65 I15 (L325_0r0[64:0], L325_0r1[64:0], L325_0a, L393_0r, L393_0a, L336_0r0[64:0], L336_0r1[64:0], L336_0a, reset);
  tkf65mo0w0_o0w65 I16 (L326_0r0[64:0], L326_0r1[64:0], L326_0a, L394_0r, L394_0a, L337_0r0[64:0], L337_0r1[64:0], L337_0a, reset);
  tkf65mo0w0_o0w65 I17 (L327_0r0[64:0], L327_0r1[64:0], L327_0a, L395_0r, L395_0a, L338_0r0[64:0], L338_0r1[64:0], L338_0a, reset);
  tkm4x33b I18 (L224_0r0[32:0], L224_0r1[32:0], L224_0a, L226_0r0[32:0], L226_0r1[32:0], L226_0a, L228_0r0[32:0], L228_0r1[32:0], L228_0a, L431_0r0[32:0], L431_0r1[32:0], L431_0a, L231_0r0[32:0], L231_0r1[32:0], L231_0a, reset);
  tkm4x0b I19 (L393_0r, L393_0a, L394_0r, L394_0a, L395_0r, L395_0a, L430_0r, L430_0a, L373_0r, L373_0a, reset);
  tkf3mo0w0_o0w3 I20 (L329_0r0[2:0], L329_0r1[2:0], L329_0a, L397_0r, L397_0a, L371_0r0[2:0], L371_0r1[2:0], L371_0a, reset);
  tkm2x1b I21 (L241_0r0, L241_0r1, L241_0a, L243_0r0, L243_0r1, L243_0a, L246_0r0, L246_0r1, L246_0a, reset);
  tkm2x0b I22 (L396_0r, L396_0a, L397_0r, L397_0a, L167_0r, L167_0a, reset);
  tkm3x1b I23 (L256_0r0, L256_0r1, L256_0a, L252_0r0, L252_0r1, L252_0a, L254_0r0, L254_0r1, L254_0a, L137_0r0, L137_0r1, L137_0a, reset);
  tkj8m1_7 I24 (sfc_0r0, sfc_0r1, sfc_0a, L413_0r0[6:0], L413_0r1[6:0], L413_0a, L410_0r0[7:0], L410_0r1[7:0], L410_0a, reset);
  tkf33mo0w0_o0w33 I25 (L433_0r0[32:0], L433_0r1[32:0], L433_0a, L188_0r, L188_0a, L442_0r0[32:0], L442_0r1[32:0], L442_0a, reset);
  tkvavbvciv65_wo0w65_ro0w32o0w32o0w32o0w32o32w32o32w32o32w32o32w32o32w32o64w1o64w1o64w1o64w1o64w1o64w1 I26 (L350_0r0[64:0], L350_0r1[64:0], L350_0a, L131_0r, L131_0a, L64_0r, L64_0a, L85_0r, L85_0a, L97_0r, L97_0a, L109_0r, L109_0a, L69_0r, L69_0a, L77_0r, L77_0a, L87_0r, L87_0a, L99_0r, L99_0a, L111_0r, L111_0a, L62_0r, L62_0a, L67_0r, L67_0a, L79_0r, L79_0a, L91_0r, L91_0a, L103_0r, L103_0a, L115_0r, L115_0a, L65_0r0[31:0], L65_0r1[31:0], L65_0a, L86_0r0[31:0], L86_0r1[31:0], L86_0a, L98_0r0[31:0], L98_0r1[31:0], L98_0a, L110_0r0[31:0], L110_0r1[31:0], L110_0a, L70_0r0[31:0], L70_0r1[31:0], L70_0a, L78_0r0[31:0], L78_0r1[31:0], L78_0a, L88_0r0[31:0], L88_0r1[31:0], L88_0a, L100_0r0[31:0], L100_0r1[31:0], L100_0a, L112_0r0[31:0], L112_0r1[31:0], L112_0a, L63_0r0, L63_0r1, L63_0a, L68_0r0, L68_0r1, L68_0a, L80_0r0, L80_0r1, L80_0a, L92_0r0, L92_0r1, L92_0a, L104_0r0, L104_0r1, L104_0a, L116_0r0, L116_0r1, L116_0a, reset);
  tkvaXORbresult34_wo0w34_ro0w1o33w1o32w1 I27 (L360_0r0[33:0], L360_0r1[33:0], L360_0a, L148_0r, L148_0a, L160_0r, L160_0a, L154_0r, L154_0a, L156_0r, L156_0a, L161_0r0, L161_0r1, L161_0a, L155_0r0, L155_0r1, L155_0a, L157_0r0, L157_0r1, L157_0a, reset);
  tkj8m4_4_0 I28 (ctrl_0r0[3:0], ctrl_0r1[3:0], ctrl_0a, fi_0r0[3:0], fi_0r1[3:0], fi_0a, L215_0r, L215_0a, L323_0r0[7:0], L323_0r1[7:0], L323_0a, reset);
  tkj65m32_32_1 I29 (L86_0r0[31:0], L86_0r1[31:0], L86_0a, L88_0r0[31:0], L88_0r1[31:0], L88_0a, L92_0r0, L92_0r1, L92_0a, L325_0r0[64:0], L325_0r1[64:0], L325_0a, reset);
  tkj65m32_32_1 I30 (L98_0r0[31:0], L98_0r1[31:0], L98_0a, L100_0r0[31:0], L100_0r1[31:0], L100_0a, L104_0r0, L104_0r1, L104_0a, L326_0r0[64:0], L326_0r1[64:0], L326_0a, reset);
  tkj65m32_32_1 I31 (L110_0r0[31:0], L110_0r1[31:0], L110_0a, L112_0r0[31:0], L112_0r1[31:0], L112_0a, L116_0r0, L116_0r1, L116_0a, L327_0r0[64:0], L327_0r1[64:0], L327_0a, reset);
  tkj34m1_0_33 I32 (L382_0r0, L382_0r1, L382_0a, L124_0r, L124_0a, L231_0r0[32:0], L231_0r1[32:0], L231_0a, L383_0r0[33:0], L383_0r1[33:0], L383_0a, reset);
  tkj3m1_1_1 I33 (L155_0r0, L155_0r1, L155_0a, L157_0r0, L157_0r1, L157_0a, L161_0r0, L161_0r1, L161_0a, L329_0r0[2:0], L329_0r1[2:0], L329_0a, reset);
  tko3m1_1xori0w1bi1w1b_2xort1o0w1bi2w1b I34 (L371_0r0[2:0], L371_0r1[2:0], L371_0a, L243_0r0, L243_0r1, L243_0a, reset);
  tkf0mo0w0_o0w0 I35 (L150_0r, L150_0a, L339_0r, L339_0a, L396_0r, L396_0a, reset);
  tkf65mo0w1_o0w65 I36 (L317_0r0[64:0], L317_0r1[64:0], L317_0a, L382_0r0, L382_0r1, L382_0a, L350_0r0[64:0], L350_0r1[64:0], L350_0a, reset);
  tkf34mo0w32_o0w34_o1w32 I37 (L321_0r0[33:0], L321_0r1[33:0], L321_0a, L432_0r0[31:0], L432_0r1[31:0], L432_0a, L360_0r0[33:0], L360_0r1[33:0], L360_0a, o_0r0[31:0], o_0r1[31:0], o_0a, reset);
  tkf8mo0w4_o0w7_o0w4_o0w4 I38 (L323_0r0[7:0], L323_0r1[7:0], L323_0a, L445_0r0[3:0], L445_0r1[3:0], L445_0a, L413_0r0[6:0], L413_0r1[6:0], L413_0a, L369_0r0[3:0], L369_0r1[3:0], L369_0a, L367_0r0[3:0], L367_0r1[3:0], L367_0a, reset);
  tkj4m0_4 I39 (L407_0r, L407_0a, L367_0r0[3:0], L367_0r1[3:0], L367_0a, L421_0r0[3:0], L421_0r1[3:0], L421_0a, reset);
  tkj4m4_0 I40 (L369_0r0[3:0], L369_0r1[3:0], L369_0a, L148_0r, L148_0a, L149_0r0[3:0], L149_0r1[3:0], L149_0a, reset);
  tkvctrlfisfc9_wo0w9_ro0w4o5w1o4w1o8w1 I41 (L406_0r0[8:0], L406_0r1[8:0], L406_0a, L407_0r, L407_0a, L59_0r, L59_0a, L341_0r, L341_0a, L339_0r, L339_0a, L340_0r, L340_0a, L60_0r0[3:0], L60_0r1[3:0], L60_0a, L254_0r0, L254_0r1, L254_0a, L241_0r0, L241_0r1, L241_0a, L252_0r0, L252_0r1, L252_0a, reset);
  tko34m34_1xori0w1bi0w1b_2apt1o0w1bi1w33b I42 (L383_0r0[33:0], L383_0r1[33:0], L383_0a, L321_0r0[33:0], L321_0r1[33:0], L321_0a, reset);
  tko8m9_1api0w8bi0w1b I43 (L410_0r0[7:0], L410_0r1[7:0], L410_0a, L406_0r0[8:0], L406_0r1[8:0], L406_0a, reset);
  tkj33m1_32 I44 (L246_0r0, L246_0r1, L246_0a, L432_0r0[31:0], L432_0r1[31:0], L432_0a, L433_0r0[32:0], L433_0r1[32:0], L433_0a, reset);
  tks4_o0w4_0c8m1c8mcmdmemfo0w0_5m6m7o0w0_2m3mam4mbo0w4 I45 (L421_0r0[3:0], L421_0r1[3:0], L421_0a, L340_0r, L340_0a, L341_0r, L341_0a, L437_0r0[3:0], L437_0r1[3:0], L437_0a, reset);
  tkm2x33b I46 (L220_0r0[32:0], L220_0r1[32:0], L220_0a, L222_0r0[32:0], L222_0r1[32:0], L222_0a, L429_0r0[32:0], L429_0r1[32:0], L429_0a, reset);
  tkf33mo0w0_o0w33 I47 (L429_0r0[32:0], L429_0r1[32:0], L429_0a, L430_0r, L430_0a, L431_0r0[32:0], L431_0r1[32:0], L431_0a, reset);
  tko4m1_1nm1b1_2nm1b0_3mx2o3o10_4o11_i0w4bt1o0w1bt2o0w1b I48 (L437_0r0[3:0], L437_0r1[3:0], L437_0a, L256_0r0, L256_0r1, L256_0a, reset);
  tko66m33_1nm1b0_2api0w33bt1o0w1b_3nm1b0_4api33w33bt3o0w1b_5addt2o0w34bt4o0w34b_6apt5o1w33b I49 (L72_0r0[65:0], L72_0r1[65:0], L72_0a, L220_0r0[32:0], L220_0r1[32:0], L220_0a, reset);
  tkj69m32_4_32_1 I50 (a_0r0[31:0], a_0r1[31:0], a_0a, L445_0r0[3:0], L445_0r1[3:0], L445_0a, b_0r0[31:0], b_0r1[31:0], b_0a, L137_0r0, L137_0r1, L137_0a, L446_0r0[68:0], L446_0r1[68:0], L446_0a, reset);
  tko33m4_1api0w2bi0w2b I51 (L442_0r0[32:0], L442_0r1[32:0], L442_0a, f_0r0[3:0], f_0r1[3:0], f_0a, reset);
  tko69m65_1nm2b1_2nm2b2_3mx0m12o1m12o3m8o7_2o6o10o14o15_i32w4bt1o0w2bt2o0w2b_4nm2b1_5nm2b2_6mx0m14o1m12o11o15_3o7_i32w4bt4o0w2bt5o0w2b_7noti36w32b_8mx2_1_t3o0w2bt7o0w32bi36w32b_9noti0w32b_10mx2_1_t6o0w2bt9o0w32bi0w32b_11apt10o0w32bt8o0w32bi68w1b I52 (L446_0r0[68:0], L446_0r1[68:0], L446_0a, L317_0r0[64:0], L317_0r1[64:0], L317_0a, reset);
  tki I53 (L208_0r, L208_0a, L215_0r, L215_0a, reset);
endmodule

