/*
    `nanoMultiplier.v'
    Balsa Verilog netlist file
    Created: Mon Nov  3 14:59:55 GMT 2008
    By: tarazonl@royaloak.cs.man.ac.uk (Linux)
    With net-verilog (balsa-netlist) version: 3.5gtk2
    Using technology: example/teak/Jbuf=1:Mbuf=1:Vbuf=0:Sbuf=1:Fbuf=1
    Command line : (balsa-netlist -Xexample/teak/Jbuf=1:Mbuf=1:Vbuf=0:Sbuf=1:Fbuf=1 -I /home/amulinks/balsa/linux/3.5gtk2/share/teak/ nanoMultiplier)

    Using `propagate-globals'
    The design contains the following global nets
		global-signal:  initialise input 1
*/

`timescale 1ns/1ps

module C2RI (
  o,
  i0,
  i1,
  initialise
);
  output o;
  input i0;
  input i1;
  input initialise;
  C2R I0 (o, i0, i1, initialise);
endmodule

module BrzF_0_l31__28_280_200_29_20_280_200_29_29 (
  i_0r, i_0a,
  o_0r, o_0a,
  o_1r, o_1a,
  initialise
);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input initialise;
  wire ifint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire ofint_1n;
  wire oaint_0n;
  wire oaint_1n;
  wire gate9_0n;
  wire gate6_0n;
  wire gate3_0n;
  assign oaint_1n = o_1r;
  INV I1 (gate9_0n, o_1a);
  C2RI I2 (o_1r, ofint_1n, gate9_0n, initialise);
  assign oaint_0n = o_0r;
  INV I4 (gate6_0n, o_0a);
  C2RI I5 (o_0r, ofint_0n, gate6_0n, initialise);
  assign i_0a = ifint_0n;
  INV I7 (gate3_0n, iaint_0n);
  C2RI I8 (ifint_0n, i_0r, gate3_0n, initialise);
  C2 I9 (iaint_0n, oaint_0n, oaint_1n);
  assign ofint_1n = ifint_0n;
  assign ofint_0n = ifint_0n;
endmodule

module BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m (
  i_0r, i_0a,
  o_0r, o_0a,
  o_1r, o_1a,
  o_2r, o_2a,
  initialise
);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  input initialise;
  wire ifint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire ofint_1n;
  wire ofint_2n;
  wire oaint_0n;
  wire oaint_1n;
  wire oaint_2n;
  wire gate21_0n;
  wire gate18_0n;
  wire gate15_0n;
  wire gate12_0n;
  assign oaint_2n = o_2r;
  INV I1 (gate21_0n, o_2a);
  C2RI I2 (o_2r, ofint_2n, gate21_0n, initialise);
  assign oaint_1n = o_1r;
  INV I4 (gate18_0n, o_1a);
  C2RI I5 (o_1r, ofint_1n, gate18_0n, initialise);
  assign oaint_0n = o_0r;
  INV I7 (gate15_0n, o_0a);
  C2RI I8 (o_0r, ofint_0n, gate15_0n, initialise);
  assign i_0a = ifint_0n;
  INV I10 (gate12_0n, iaint_0n);
  C2RI I11 (ifint_0n, i_0r, gate12_0n, initialise);
  C3 I12 (iaint_0n, oaint_0n, oaint_1n, oaint_2n);
  assign ofint_2n = ifint_0n;
  assign ofint_1n = ifint_0n;
  assign ofint_0n = ifint_0n;
endmodule

module BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m (
  i_0r, i_0a,
  o_0r, o_0a,
  o_1r, o_1a,
  o_2r, o_2a,
  o_3r, o_3a,
  initialise
);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  input initialise;
  wire [1:0] internal_0n;
  wire ifint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire ofint_1n;
  wire ofint_2n;
  wire ofint_3n;
  wire oaint_0n;
  wire oaint_1n;
  wire oaint_2n;
  wire oaint_3n;
  wire gate36_0n;
  wire gate33_0n;
  wire gate30_0n;
  wire gate27_0n;
  wire gate24_0n;
  assign oaint_3n = o_3r;
  INV I1 (gate36_0n, o_3a);
  C2RI I2 (o_3r, ofint_3n, gate36_0n, initialise);
  assign oaint_2n = o_2r;
  INV I4 (gate33_0n, o_2a);
  C2RI I5 (o_2r, ofint_2n, gate33_0n, initialise);
  assign oaint_1n = o_1r;
  INV I7 (gate30_0n, o_1a);
  C2RI I8 (o_1r, ofint_1n, gate30_0n, initialise);
  assign oaint_0n = o_0r;
  INV I10 (gate27_0n, o_0a);
  C2RI I11 (o_0r, ofint_0n, gate27_0n, initialise);
  assign i_0a = ifint_0n;
  INV I13 (gate24_0n, iaint_0n);
  C2RI I14 (ifint_0n, i_0r, gate24_0n, initialise);
  C2 I15 (internal_0n[0], oaint_0n, oaint_1n);
  C2 I16 (internal_0n[1], oaint_2n, oaint_3n);
  C2 I17 (iaint_0n, internal_0n[0], internal_0n[1]);
  assign ofint_3n = ifint_0n;
  assign ofint_2n = ifint_0n;
  assign ofint_1n = ifint_0n;
  assign ofint_0n = ifint_0n;
endmodule

module BrzF_0_l73__28_280_200_29_20_280_200_29_20_m35m (
  i_0r, i_0a,
  o_0r, o_0a,
  o_1r, o_1a,
  o_2r, o_2a,
  o_3r, o_3a,
  o_4r, o_4a,
  initialise
);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  input initialise;
  wire [1:0] internal_0n;
  wire ifint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire ofint_1n;
  wire ofint_2n;
  wire ofint_3n;
  wire ofint_4n;
  wire oaint_0n;
  wire oaint_1n;
  wire oaint_2n;
  wire oaint_3n;
  wire oaint_4n;
  wire gate54_0n;
  wire gate51_0n;
  wire gate48_0n;
  wire gate45_0n;
  wire gate42_0n;
  wire gate39_0n;
  assign oaint_4n = o_4r;
  INV I1 (gate54_0n, o_4a);
  C2RI I2 (o_4r, ofint_4n, gate54_0n, initialise);
  assign oaint_3n = o_3r;
  INV I4 (gate51_0n, o_3a);
  C2RI I5 (o_3r, ofint_3n, gate51_0n, initialise);
  assign oaint_2n = o_2r;
  INV I7 (gate48_0n, o_2a);
  C2RI I8 (o_2r, ofint_2n, gate48_0n, initialise);
  assign oaint_1n = o_1r;
  INV I10 (gate45_0n, o_1a);
  C2RI I11 (o_1r, ofint_1n, gate45_0n, initialise);
  assign oaint_0n = o_0r;
  INV I13 (gate42_0n, o_0a);
  C2RI I14 (o_0r, ofint_0n, gate42_0n, initialise);
  assign i_0a = ifint_0n;
  INV I16 (gate39_0n, iaint_0n);
  C2RI I17 (ifint_0n, i_0r, gate39_0n, initialise);
  C3 I18 (internal_0n[0], oaint_0n, oaint_1n, oaint_2n);
  C2 I19 (internal_0n[1], oaint_3n, oaint_4n);
  C2 I20 (iaint_0n, internal_0n[0], internal_0n[1]);
  assign ofint_4n = ifint_0n;
  assign ofint_3n = ifint_0n;
  assign ofint_2n = ifint_0n;
  assign ofint_1n = ifint_0n;
  assign ofint_0n = ifint_0n;
endmodule

module BrzF_0_l87__28_280_200_29_20_280_200_29_20_m36m (
  i_0r, i_0a,
  o_0r, o_0a,
  o_1r, o_1a,
  o_2r, o_2a,
  o_3r, o_3a,
  o_4r, o_4a,
  o_5r, o_5a,
  initialise
);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  input initialise;
  wire [1:0] internal_0n;
  wire ifint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire ofint_1n;
  wire ofint_2n;
  wire ofint_3n;
  wire ofint_4n;
  wire ofint_5n;
  wire oaint_0n;
  wire oaint_1n;
  wire oaint_2n;
  wire oaint_3n;
  wire oaint_4n;
  wire oaint_5n;
  wire gate75_0n;
  wire gate72_0n;
  wire gate69_0n;
  wire gate66_0n;
  wire gate63_0n;
  wire gate60_0n;
  wire gate57_0n;
  assign oaint_5n = o_5r;
  INV I1 (gate75_0n, o_5a);
  C2RI I2 (o_5r, ofint_5n, gate75_0n, initialise);
  assign oaint_4n = o_4r;
  INV I4 (gate72_0n, o_4a);
  C2RI I5 (o_4r, ofint_4n, gate72_0n, initialise);
  assign oaint_3n = o_3r;
  INV I7 (gate69_0n, o_3a);
  C2RI I8 (o_3r, ofint_3n, gate69_0n, initialise);
  assign oaint_2n = o_2r;
  INV I10 (gate66_0n, o_2a);
  C2RI I11 (o_2r, ofint_2n, gate66_0n, initialise);
  assign oaint_1n = o_1r;
  INV I13 (gate63_0n, o_1a);
  C2RI I14 (o_1r, ofint_1n, gate63_0n, initialise);
  assign oaint_0n = o_0r;
  INV I16 (gate60_0n, o_0a);
  C2RI I17 (o_0r, ofint_0n, gate60_0n, initialise);
  assign i_0a = ifint_0n;
  INV I19 (gate57_0n, iaint_0n);
  C2RI I20 (ifint_0n, i_0r, gate57_0n, initialise);
  C3 I21 (internal_0n[0], oaint_0n, oaint_1n, oaint_2n);
  C3 I22 (internal_0n[1], oaint_3n, oaint_4n, oaint_5n);
  C2 I23 (iaint_0n, internal_0n[0], internal_0n[1]);
  assign ofint_5n = ifint_0n;
  assign ofint_4n = ifint_0n;
  assign ofint_3n = ifint_0n;
  assign ofint_2n = ifint_0n;
  assign ofint_1n = ifint_0n;
  assign ofint_0n = ifint_0n;
endmodule

module BrzF_0_l101__28_280_200_29_20_280_200_29_2_m37m (
  i_0r, i_0a,
  o_0r, o_0a,
  o_1r, o_1a,
  o_2r, o_2a,
  o_3r, o_3a,
  o_4r, o_4a,
  o_5r, o_5a,
  o_6r, o_6a,
  initialise
);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  input initialise;
  wire [2:0] internal_0n;
  wire ifint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire ofint_1n;
  wire ofint_2n;
  wire ofint_3n;
  wire ofint_4n;
  wire ofint_5n;
  wire ofint_6n;
  wire oaint_0n;
  wire oaint_1n;
  wire oaint_2n;
  wire oaint_3n;
  wire oaint_4n;
  wire oaint_5n;
  wire oaint_6n;
  wire gate99_0n;
  wire gate96_0n;
  wire gate93_0n;
  wire gate90_0n;
  wire gate87_0n;
  wire gate84_0n;
  wire gate81_0n;
  wire gate78_0n;
  assign oaint_6n = o_6r;
  INV I1 (gate99_0n, o_6a);
  C2RI I2 (o_6r, ofint_6n, gate99_0n, initialise);
  assign oaint_5n = o_5r;
  INV I4 (gate96_0n, o_5a);
  C2RI I5 (o_5r, ofint_5n, gate96_0n, initialise);
  assign oaint_4n = o_4r;
  INV I7 (gate93_0n, o_4a);
  C2RI I8 (o_4r, ofint_4n, gate93_0n, initialise);
  assign oaint_3n = o_3r;
  INV I10 (gate90_0n, o_3a);
  C2RI I11 (o_3r, ofint_3n, gate90_0n, initialise);
  assign oaint_2n = o_2r;
  INV I13 (gate87_0n, o_2a);
  C2RI I14 (o_2r, ofint_2n, gate87_0n, initialise);
  assign oaint_1n = o_1r;
  INV I16 (gate84_0n, o_1a);
  C2RI I17 (o_1r, ofint_1n, gate84_0n, initialise);
  assign oaint_0n = o_0r;
  INV I19 (gate81_0n, o_0a);
  C2RI I20 (o_0r, ofint_0n, gate81_0n, initialise);
  assign i_0a = ifint_0n;
  INV I22 (gate78_0n, iaint_0n);
  C2RI I23 (ifint_0n, i_0r, gate78_0n, initialise);
  C3 I24 (internal_0n[0], oaint_0n, oaint_1n, oaint_2n);
  C2 I25 (internal_0n[1], oaint_3n, oaint_4n);
  C2 I26 (internal_0n[2], oaint_5n, oaint_6n);
  C3 I27 (iaint_0n, internal_0n[0], internal_0n[1], internal_0n[2]);
  assign ofint_6n = ifint_0n;
  assign ofint_5n = ifint_0n;
  assign ofint_4n = ifint_0n;
  assign ofint_3n = ifint_0n;
  assign ofint_2n = ifint_0n;
  assign ofint_1n = ifint_0n;
  assign ofint_0n = ifint_0n;
endmodule

module BrzF_0_l115__28_280_200_29_20_280_200_29_2_m38m (
  i_0r, i_0a,
  o_0r, o_0a,
  o_1r, o_1a,
  o_2r, o_2a,
  o_3r, o_3a,
  o_4r, o_4a,
  o_5r, o_5a,
  o_6r, o_6a,
  o_7r, o_7a,
  initialise
);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  output o_7r;
  input o_7a;
  input initialise;
  wire [2:0] internal_0n;
  wire ifint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire ofint_1n;
  wire ofint_2n;
  wire ofint_3n;
  wire ofint_4n;
  wire ofint_5n;
  wire ofint_6n;
  wire ofint_7n;
  wire oaint_0n;
  wire oaint_1n;
  wire oaint_2n;
  wire oaint_3n;
  wire oaint_4n;
  wire oaint_5n;
  wire oaint_6n;
  wire oaint_7n;
  wire gate126_0n;
  wire gate123_0n;
  wire gate120_0n;
  wire gate117_0n;
  wire gate114_0n;
  wire gate111_0n;
  wire gate108_0n;
  wire gate105_0n;
  wire gate102_0n;
  assign oaint_7n = o_7r;
  INV I1 (gate126_0n, o_7a);
  C2RI I2 (o_7r, ofint_7n, gate126_0n, initialise);
  assign oaint_6n = o_6r;
  INV I4 (gate123_0n, o_6a);
  C2RI I5 (o_6r, ofint_6n, gate123_0n, initialise);
  assign oaint_5n = o_5r;
  INV I7 (gate120_0n, o_5a);
  C2RI I8 (o_5r, ofint_5n, gate120_0n, initialise);
  assign oaint_4n = o_4r;
  INV I10 (gate117_0n, o_4a);
  C2RI I11 (o_4r, ofint_4n, gate117_0n, initialise);
  assign oaint_3n = o_3r;
  INV I13 (gate114_0n, o_3a);
  C2RI I14 (o_3r, ofint_3n, gate114_0n, initialise);
  assign oaint_2n = o_2r;
  INV I16 (gate111_0n, o_2a);
  C2RI I17 (o_2r, ofint_2n, gate111_0n, initialise);
  assign oaint_1n = o_1r;
  INV I19 (gate108_0n, o_1a);
  C2RI I20 (o_1r, ofint_1n, gate108_0n, initialise);
  assign oaint_0n = o_0r;
  INV I22 (gate105_0n, o_0a);
  C2RI I23 (o_0r, ofint_0n, gate105_0n, initialise);
  assign i_0a = ifint_0n;
  INV I25 (gate102_0n, iaint_0n);
  C2RI I26 (ifint_0n, i_0r, gate102_0n, initialise);
  C3 I27 (internal_0n[0], oaint_0n, oaint_1n, oaint_2n);
  C3 I28 (internal_0n[1], oaint_3n, oaint_4n, oaint_5n);
  C2 I29 (internal_0n[2], oaint_6n, oaint_7n);
  C3 I30 (iaint_0n, internal_0n[0], internal_0n[1], internal_0n[2]);
  assign ofint_7n = ifint_0n;
  assign ofint_6n = ifint_0n;
  assign ofint_5n = ifint_0n;
  assign ofint_4n = ifint_0n;
  assign ofint_3n = ifint_0n;
  assign ofint_2n = ifint_0n;
  assign ofint_1n = ifint_0n;
  assign ofint_0n = ifint_0n;
endmodule

module BrzF_0_l199__28_280_200_29_20_280_200_29_2_m39m (
  i_0r, i_0a,
  o_0r, o_0a,
  o_1r, o_1a,
  o_2r, o_2a,
  o_3r, o_3a,
  o_4r, o_4a,
  o_5r, o_5a,
  o_6r, o_6a,
  o_7r, o_7a,
  o_8r, o_8a,
  o_9r, o_9a,
  o_10r, o_10a,
  o_11r, o_11a,
  o_12r, o_12a,
  o_13r, o_13a,
  initialise
);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  output o_7r;
  input o_7a;
  output o_8r;
  input o_8a;
  output o_9r;
  input o_9a;
  output o_10r;
  input o_10a;
  output o_11r;
  input o_11a;
  output o_12r;
  input o_12a;
  output o_13r;
  input o_13a;
  input initialise;
  wire [6:0] internal_0n;
  wire ifint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire ofint_1n;
  wire ofint_2n;
  wire ofint_3n;
  wire ofint_4n;
  wire ofint_5n;
  wire ofint_6n;
  wire ofint_7n;
  wire ofint_8n;
  wire ofint_9n;
  wire ofint_10n;
  wire ofint_11n;
  wire ofint_12n;
  wire ofint_13n;
  wire oaint_0n;
  wire oaint_1n;
  wire oaint_2n;
  wire oaint_3n;
  wire oaint_4n;
  wire oaint_5n;
  wire oaint_6n;
  wire oaint_7n;
  wire oaint_8n;
  wire oaint_9n;
  wire oaint_10n;
  wire oaint_11n;
  wire oaint_12n;
  wire oaint_13n;
  wire gate171_0n;
  wire gate168_0n;
  wire gate165_0n;
  wire gate162_0n;
  wire gate159_0n;
  wire gate156_0n;
  wire gate153_0n;
  wire gate150_0n;
  wire gate147_0n;
  wire gate144_0n;
  wire gate141_0n;
  wire gate138_0n;
  wire gate135_0n;
  wire gate132_0n;
  wire gate129_0n;
  assign oaint_13n = o_13r;
  INV I1 (gate171_0n, o_13a);
  C2RI I2 (o_13r, ofint_13n, gate171_0n, initialise);
  assign oaint_12n = o_12r;
  INV I4 (gate168_0n, o_12a);
  C2RI I5 (o_12r, ofint_12n, gate168_0n, initialise);
  assign oaint_11n = o_11r;
  INV I7 (gate165_0n, o_11a);
  C2RI I8 (o_11r, ofint_11n, gate165_0n, initialise);
  assign oaint_10n = o_10r;
  INV I10 (gate162_0n, o_10a);
  C2RI I11 (o_10r, ofint_10n, gate162_0n, initialise);
  assign oaint_9n = o_9r;
  INV I13 (gate159_0n, o_9a);
  C2RI I14 (o_9r, ofint_9n, gate159_0n, initialise);
  assign oaint_8n = o_8r;
  INV I16 (gate156_0n, o_8a);
  C2RI I17 (o_8r, ofint_8n, gate156_0n, initialise);
  assign oaint_7n = o_7r;
  INV I19 (gate153_0n, o_7a);
  C2RI I20 (o_7r, ofint_7n, gate153_0n, initialise);
  assign oaint_6n = o_6r;
  INV I22 (gate150_0n, o_6a);
  C2RI I23 (o_6r, ofint_6n, gate150_0n, initialise);
  assign oaint_5n = o_5r;
  INV I25 (gate147_0n, o_5a);
  C2RI I26 (o_5r, ofint_5n, gate147_0n, initialise);
  assign oaint_4n = o_4r;
  INV I28 (gate144_0n, o_4a);
  C2RI I29 (o_4r, ofint_4n, gate144_0n, initialise);
  assign oaint_3n = o_3r;
  INV I31 (gate141_0n, o_3a);
  C2RI I32 (o_3r, ofint_3n, gate141_0n, initialise);
  assign oaint_2n = o_2r;
  INV I34 (gate138_0n, o_2a);
  C2RI I35 (o_2r, ofint_2n, gate138_0n, initialise);
  assign oaint_1n = o_1r;
  INV I37 (gate135_0n, o_1a);
  C2RI I38 (o_1r, ofint_1n, gate135_0n, initialise);
  assign oaint_0n = o_0r;
  INV I40 (gate132_0n, o_0a);
  C2RI I41 (o_0r, ofint_0n, gate132_0n, initialise);
  assign i_0a = ifint_0n;
  INV I43 (gate129_0n, iaint_0n);
  C2RI I44 (ifint_0n, i_0r, gate129_0n, initialise);
  C3 I45 (internal_0n[0], oaint_0n, oaint_1n, oaint_2n);
  C3 I46 (internal_0n[1], oaint_3n, oaint_4n, oaint_5n);
  C3 I47 (internal_0n[2], oaint_6n, oaint_7n, oaint_8n);
  C3 I48 (internal_0n[3], oaint_9n, oaint_10n, oaint_11n);
  C2 I49 (internal_0n[4], oaint_12n, oaint_13n);
  C3 I50 (internal_0n[5], internal_0n[0], internal_0n[1], internal_0n[2]);
  C2 I51 (internal_0n[6], internal_0n[3], internal_0n[4]);
  C2 I52 (iaint_0n, internal_0n[5], internal_0n[6]);
  assign ofint_13n = ifint_0n;
  assign ofint_12n = ifint_0n;
  assign ofint_11n = ifint_0n;
  assign ofint_10n = ifint_0n;
  assign ofint_9n = ifint_0n;
  assign ofint_8n = ifint_0n;
  assign ofint_7n = ifint_0n;
  assign ofint_6n = ifint_0n;
  assign ofint_5n = ifint_0n;
  assign ofint_4n = ifint_0n;
  assign ofint_3n = ifint_0n;
  assign ofint_2n = ifint_0n;
  assign ofint_1n = ifint_0n;
  assign ofint_0n = ifint_0n;
endmodule

module BrzF_1_l17__28_280_200_29_29 (
  i_0r0d, i_0r1d, i_0a,
  o_0r, o_0a,
  initialise
);
  input i_0r0d;
  input i_0r1d;
  output i_0a;
  output o_0r;
  input o_0a;
  input initialise;
  wire ifint_0n;
  wire itint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire oaint_0n;
  wire gate179_0n;
  wire complete176_0n;
  wire gate175_0n;
  wire complete172_0n;
  wire icomplete_0n;
  assign oaint_0n = o_0r;
  INV I1 (gate179_0n, o_0a);
  C2RI I2 (o_0r, ofint_0n, gate179_0n, initialise);
  assign i_0a = complete176_0n;
  OR2 I4 (complete176_0n, ifint_0n, itint_0n);
  INV I5 (gate175_0n, iaint_0n);
  C2RI I6 (itint_0n, i_0r1d, gate175_0n, initialise);
  C2RI I7 (ifint_0n, i_0r0d, gate175_0n, initialise);
  C2 I8 (iaint_0n, icomplete_0n, oaint_0n);
  assign ofint_0n = icomplete_0n;
  assign icomplete_0n = complete172_0n;
  OR2 I11 (complete172_0n, ifint_0n, itint_0n);
endmodule

module BrzF_1_l31__28_280_200_29_20_280_201_29_29 (
  i_0r0d, i_0r1d, i_0a,
  o_0r, o_0a,
  o_1r0d, o_1r1d, o_1a,
  initialise
);
  input i_0r0d;
  input i_0r1d;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r0d;
  output o_1r1d;
  input o_1a;
  input initialise;
  wire ifint_0n;
  wire itint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire ofint_1n;
  wire otint_1n;
  wire oaint_0n;
  wire oaint_1n;
  wire complete191_0n;
  wire gate190_0n;
  wire gate187_0n;
  wire complete184_0n;
  wire gate183_0n;
  wire complete180_0n;
  wire icomplete_0n;
  assign oaint_1n = complete191_0n;
  OR2 I1 (complete191_0n, o_1r0d, o_1r1d);
  INV I2 (gate190_0n, o_1a);
  C2RI I3 (o_1r1d, otint_1n, gate190_0n, initialise);
  C2RI I4 (o_1r0d, ofint_1n, gate190_0n, initialise);
  assign oaint_0n = o_0r;
  INV I6 (gate187_0n, o_0a);
  C2RI I7 (o_0r, ofint_0n, gate187_0n, initialise);
  assign i_0a = complete184_0n;
  OR2 I9 (complete184_0n, ifint_0n, itint_0n);
  INV I10 (gate183_0n, iaint_0n);
  C2RI I11 (itint_0n, i_0r1d, gate183_0n, initialise);
  C2RI I12 (ifint_0n, i_0r0d, gate183_0n, initialise);
  C3 I13 (iaint_0n, icomplete_0n, oaint_0n, oaint_1n);
  assign ofint_0n = icomplete_0n;
  assign otint_1n = itint_0n;
  assign ofint_1n = ifint_0n;
  assign icomplete_0n = complete180_0n;
  OR2 I18 (complete180_0n, ifint_0n, itint_0n);
endmodule

module BrzF_3_l31__28_280_200_29_20_280_203_29_29 (
  i_0r0d, i_0r1d, i_0a,
  o_0r, o_0a,
  o_1r0d, o_1r1d, o_1a,
  initialise
);
  input [2:0] i_0r0d;
  input [2:0] i_0r1d;
  output i_0a;
  output o_0r;
  input o_0a;
  output [2:0] o_1r0d;
  output [2:0] o_1r1d;
  input o_1a;
  input initialise;
  wire [2:0] ifint_0n;
  wire [2:0] itint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire [2:0] ofint_1n;
  wire [2:0] otint_1n;
  wire oaint_0n;
  wire oaint_1n;
  wire [2:0] complete203_0n;
  wire gate202_0n;
  wire gate199_0n;
  wire [2:0] complete196_0n;
  wire gate195_0n;
  wire [2:0] complete192_0n;
  wire icomplete_0n;
  C3 I0 (oaint_1n, complete203_0n[0], complete203_0n[1], complete203_0n[2]);
  OR2 I1 (complete203_0n[0], o_1r0d[0], o_1r1d[0]);
  OR2 I2 (complete203_0n[1], o_1r0d[1], o_1r1d[1]);
  OR2 I3 (complete203_0n[2], o_1r0d[2], o_1r1d[2]);
  INV I4 (gate202_0n, o_1a);
  C2RI I5 (o_1r1d[0], otint_1n[0], gate202_0n, initialise);
  C2RI I6 (o_1r1d[1], otint_1n[1], gate202_0n, initialise);
  C2RI I7 (o_1r1d[2], otint_1n[2], gate202_0n, initialise);
  C2RI I8 (o_1r0d[0], ofint_1n[0], gate202_0n, initialise);
  C2RI I9 (o_1r0d[1], ofint_1n[1], gate202_0n, initialise);
  C2RI I10 (o_1r0d[2], ofint_1n[2], gate202_0n, initialise);
  assign oaint_0n = o_0r;
  INV I12 (gate199_0n, o_0a);
  C2RI I13 (o_0r, ofint_0n, gate199_0n, initialise);
  C3 I14 (i_0a, complete196_0n[0], complete196_0n[1], complete196_0n[2]);
  OR2 I15 (complete196_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I16 (complete196_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I17 (complete196_0n[2], ifint_0n[2], itint_0n[2]);
  INV I18 (gate195_0n, iaint_0n);
  C2RI I19 (itint_0n[0], i_0r1d[0], gate195_0n, initialise);
  C2RI I20 (itint_0n[1], i_0r1d[1], gate195_0n, initialise);
  C2RI I21 (itint_0n[2], i_0r1d[2], gate195_0n, initialise);
  C2RI I22 (ifint_0n[0], i_0r0d[0], gate195_0n, initialise);
  C2RI I23 (ifint_0n[1], i_0r0d[1], gate195_0n, initialise);
  C2RI I24 (ifint_0n[2], i_0r0d[2], gate195_0n, initialise);
  C3 I25 (iaint_0n, icomplete_0n, oaint_0n, oaint_1n);
  assign ofint_0n = icomplete_0n;
  assign otint_1n[0] = itint_0n[0];
  assign otint_1n[1] = itint_0n[1];
  assign otint_1n[2] = itint_0n[2];
  assign ofint_1n[0] = ifint_0n[0];
  assign ofint_1n[1] = ifint_0n[1];
  assign ofint_1n[2] = ifint_0n[2];
  C3 I33 (icomplete_0n, complete192_0n[0], complete192_0n[1], complete192_0n[2]);
  OR2 I34 (complete192_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I35 (complete192_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I36 (complete192_0n[2], ifint_0n[2], itint_0n[2]);
endmodule

module BrzF_32_l17__28_280_200_29_29 (
  i_0r0d, i_0r1d, i_0a,
  o_0r, o_0a,
  initialise
);
  input [31:0] i_0r0d;
  input [31:0] i_0r1d;
  output i_0a;
  output o_0r;
  input o_0a;
  input initialise;
  wire [33:0] internal_0n;
  wire [31:0] ifint_0n;
  wire [31:0] itint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire oaint_0n;
  wire gate211_0n;
  wire [31:0] complete208_0n;
  wire gate207_0n;
  wire [31:0] complete204_0n;
  wire icomplete_0n;
  assign oaint_0n = o_0r;
  INV I1 (gate211_0n, o_0a);
  C2RI I2 (o_0r, ofint_0n, gate211_0n, initialise);
  C3 I3 (internal_0n[0], complete208_0n[0], complete208_0n[1], complete208_0n[2]);
  C3 I4 (internal_0n[1], complete208_0n[3], complete208_0n[4], complete208_0n[5]);
  C3 I5 (internal_0n[2], complete208_0n[6], complete208_0n[7], complete208_0n[8]);
  C3 I6 (internal_0n[3], complete208_0n[9], complete208_0n[10], complete208_0n[11]);
  C3 I7 (internal_0n[4], complete208_0n[12], complete208_0n[13], complete208_0n[14]);
  C3 I8 (internal_0n[5], complete208_0n[15], complete208_0n[16], complete208_0n[17]);
  C3 I9 (internal_0n[6], complete208_0n[18], complete208_0n[19], complete208_0n[20]);
  C3 I10 (internal_0n[7], complete208_0n[21], complete208_0n[22], complete208_0n[23]);
  C3 I11 (internal_0n[8], complete208_0n[24], complete208_0n[25], complete208_0n[26]);
  C3 I12 (internal_0n[9], complete208_0n[27], complete208_0n[28], complete208_0n[29]);
  C2 I13 (internal_0n[10], complete208_0n[30], complete208_0n[31]);
  C3 I14 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I15 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I16 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I17 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I18 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I19 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I20 (i_0a, internal_0n[15], internal_0n[16]);
  OR2 I21 (complete208_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I22 (complete208_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I23 (complete208_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I24 (complete208_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I25 (complete208_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I26 (complete208_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I27 (complete208_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I28 (complete208_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I29 (complete208_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I30 (complete208_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I31 (complete208_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I32 (complete208_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I33 (complete208_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I34 (complete208_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I35 (complete208_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I36 (complete208_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I37 (complete208_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I38 (complete208_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I39 (complete208_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I40 (complete208_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I41 (complete208_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I42 (complete208_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I43 (complete208_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I44 (complete208_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I45 (complete208_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I46 (complete208_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I47 (complete208_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I48 (complete208_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I49 (complete208_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I50 (complete208_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I51 (complete208_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I52 (complete208_0n[31], ifint_0n[31], itint_0n[31]);
  INV I53 (gate207_0n, iaint_0n);
  C2RI I54 (itint_0n[0], i_0r1d[0], gate207_0n, initialise);
  C2RI I55 (itint_0n[1], i_0r1d[1], gate207_0n, initialise);
  C2RI I56 (itint_0n[2], i_0r1d[2], gate207_0n, initialise);
  C2RI I57 (itint_0n[3], i_0r1d[3], gate207_0n, initialise);
  C2RI I58 (itint_0n[4], i_0r1d[4], gate207_0n, initialise);
  C2RI I59 (itint_0n[5], i_0r1d[5], gate207_0n, initialise);
  C2RI I60 (itint_0n[6], i_0r1d[6], gate207_0n, initialise);
  C2RI I61 (itint_0n[7], i_0r1d[7], gate207_0n, initialise);
  C2RI I62 (itint_0n[8], i_0r1d[8], gate207_0n, initialise);
  C2RI I63 (itint_0n[9], i_0r1d[9], gate207_0n, initialise);
  C2RI I64 (itint_0n[10], i_0r1d[10], gate207_0n, initialise);
  C2RI I65 (itint_0n[11], i_0r1d[11], gate207_0n, initialise);
  C2RI I66 (itint_0n[12], i_0r1d[12], gate207_0n, initialise);
  C2RI I67 (itint_0n[13], i_0r1d[13], gate207_0n, initialise);
  C2RI I68 (itint_0n[14], i_0r1d[14], gate207_0n, initialise);
  C2RI I69 (itint_0n[15], i_0r1d[15], gate207_0n, initialise);
  C2RI I70 (itint_0n[16], i_0r1d[16], gate207_0n, initialise);
  C2RI I71 (itint_0n[17], i_0r1d[17], gate207_0n, initialise);
  C2RI I72 (itint_0n[18], i_0r1d[18], gate207_0n, initialise);
  C2RI I73 (itint_0n[19], i_0r1d[19], gate207_0n, initialise);
  C2RI I74 (itint_0n[20], i_0r1d[20], gate207_0n, initialise);
  C2RI I75 (itint_0n[21], i_0r1d[21], gate207_0n, initialise);
  C2RI I76 (itint_0n[22], i_0r1d[22], gate207_0n, initialise);
  C2RI I77 (itint_0n[23], i_0r1d[23], gate207_0n, initialise);
  C2RI I78 (itint_0n[24], i_0r1d[24], gate207_0n, initialise);
  C2RI I79 (itint_0n[25], i_0r1d[25], gate207_0n, initialise);
  C2RI I80 (itint_0n[26], i_0r1d[26], gate207_0n, initialise);
  C2RI I81 (itint_0n[27], i_0r1d[27], gate207_0n, initialise);
  C2RI I82 (itint_0n[28], i_0r1d[28], gate207_0n, initialise);
  C2RI I83 (itint_0n[29], i_0r1d[29], gate207_0n, initialise);
  C2RI I84 (itint_0n[30], i_0r1d[30], gate207_0n, initialise);
  C2RI I85 (itint_0n[31], i_0r1d[31], gate207_0n, initialise);
  C2RI I86 (ifint_0n[0], i_0r0d[0], gate207_0n, initialise);
  C2RI I87 (ifint_0n[1], i_0r0d[1], gate207_0n, initialise);
  C2RI I88 (ifint_0n[2], i_0r0d[2], gate207_0n, initialise);
  C2RI I89 (ifint_0n[3], i_0r0d[3], gate207_0n, initialise);
  C2RI I90 (ifint_0n[4], i_0r0d[4], gate207_0n, initialise);
  C2RI I91 (ifint_0n[5], i_0r0d[5], gate207_0n, initialise);
  C2RI I92 (ifint_0n[6], i_0r0d[6], gate207_0n, initialise);
  C2RI I93 (ifint_0n[7], i_0r0d[7], gate207_0n, initialise);
  C2RI I94 (ifint_0n[8], i_0r0d[8], gate207_0n, initialise);
  C2RI I95 (ifint_0n[9], i_0r0d[9], gate207_0n, initialise);
  C2RI I96 (ifint_0n[10], i_0r0d[10], gate207_0n, initialise);
  C2RI I97 (ifint_0n[11], i_0r0d[11], gate207_0n, initialise);
  C2RI I98 (ifint_0n[12], i_0r0d[12], gate207_0n, initialise);
  C2RI I99 (ifint_0n[13], i_0r0d[13], gate207_0n, initialise);
  C2RI I100 (ifint_0n[14], i_0r0d[14], gate207_0n, initialise);
  C2RI I101 (ifint_0n[15], i_0r0d[15], gate207_0n, initialise);
  C2RI I102 (ifint_0n[16], i_0r0d[16], gate207_0n, initialise);
  C2RI I103 (ifint_0n[17], i_0r0d[17], gate207_0n, initialise);
  C2RI I104 (ifint_0n[18], i_0r0d[18], gate207_0n, initialise);
  C2RI I105 (ifint_0n[19], i_0r0d[19], gate207_0n, initialise);
  C2RI I106 (ifint_0n[20], i_0r0d[20], gate207_0n, initialise);
  C2RI I107 (ifint_0n[21], i_0r0d[21], gate207_0n, initialise);
  C2RI I108 (ifint_0n[22], i_0r0d[22], gate207_0n, initialise);
  C2RI I109 (ifint_0n[23], i_0r0d[23], gate207_0n, initialise);
  C2RI I110 (ifint_0n[24], i_0r0d[24], gate207_0n, initialise);
  C2RI I111 (ifint_0n[25], i_0r0d[25], gate207_0n, initialise);
  C2RI I112 (ifint_0n[26], i_0r0d[26], gate207_0n, initialise);
  C2RI I113 (ifint_0n[27], i_0r0d[27], gate207_0n, initialise);
  C2RI I114 (ifint_0n[28], i_0r0d[28], gate207_0n, initialise);
  C2RI I115 (ifint_0n[29], i_0r0d[29], gate207_0n, initialise);
  C2RI I116 (ifint_0n[30], i_0r0d[30], gate207_0n, initialise);
  C2RI I117 (ifint_0n[31], i_0r0d[31], gate207_0n, initialise);
  C2 I118 (iaint_0n, icomplete_0n, oaint_0n);
  assign ofint_0n = icomplete_0n;
  C3 I120 (internal_0n[17], complete204_0n[0], complete204_0n[1], complete204_0n[2]);
  C3 I121 (internal_0n[18], complete204_0n[3], complete204_0n[4], complete204_0n[5]);
  C3 I122 (internal_0n[19], complete204_0n[6], complete204_0n[7], complete204_0n[8]);
  C3 I123 (internal_0n[20], complete204_0n[9], complete204_0n[10], complete204_0n[11]);
  C3 I124 (internal_0n[21], complete204_0n[12], complete204_0n[13], complete204_0n[14]);
  C3 I125 (internal_0n[22], complete204_0n[15], complete204_0n[16], complete204_0n[17]);
  C3 I126 (internal_0n[23], complete204_0n[18], complete204_0n[19], complete204_0n[20]);
  C3 I127 (internal_0n[24], complete204_0n[21], complete204_0n[22], complete204_0n[23]);
  C3 I128 (internal_0n[25], complete204_0n[24], complete204_0n[25], complete204_0n[26]);
  C3 I129 (internal_0n[26], complete204_0n[27], complete204_0n[28], complete204_0n[29]);
  C2 I130 (internal_0n[27], complete204_0n[30], complete204_0n[31]);
  C3 I131 (internal_0n[28], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I132 (internal_0n[29], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I133 (internal_0n[30], internal_0n[23], internal_0n[24], internal_0n[25]);
  C2 I134 (internal_0n[31], internal_0n[26], internal_0n[27]);
  C2 I135 (internal_0n[32], internal_0n[28], internal_0n[29]);
  C2 I136 (internal_0n[33], internal_0n[30], internal_0n[31]);
  C2 I137 (icomplete_0n, internal_0n[32], internal_0n[33]);
  OR2 I138 (complete204_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I139 (complete204_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I140 (complete204_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I141 (complete204_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I142 (complete204_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I143 (complete204_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I144 (complete204_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I145 (complete204_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I146 (complete204_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I147 (complete204_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I148 (complete204_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I149 (complete204_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I150 (complete204_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I151 (complete204_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I152 (complete204_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I153 (complete204_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I154 (complete204_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I155 (complete204_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I156 (complete204_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I157 (complete204_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I158 (complete204_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I159 (complete204_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I160 (complete204_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I161 (complete204_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I162 (complete204_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I163 (complete204_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I164 (complete204_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I165 (complete204_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I166 (complete204_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I167 (complete204_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I168 (complete204_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I169 (complete204_0n[31], ifint_0n[31], itint_0n[31]);
endmodule

module BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m (
  i_0r0d, i_0r1d, i_0a,
  o_0r, o_0a,
  o_1r0d, o_1r1d, o_1a,
  initialise
);
  input [31:0] i_0r0d;
  input [31:0] i_0r1d;
  output i_0a;
  output o_0r;
  input o_0a;
  output [31:0] o_1r0d;
  output [31:0] o_1r1d;
  input o_1a;
  input initialise;
  wire [50:0] internal_0n;
  wire [31:0] ifint_0n;
  wire [31:0] itint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire [31:0] ofint_1n;
  wire [31:0] otint_1n;
  wire oaint_0n;
  wire oaint_1n;
  wire [31:0] complete223_0n;
  wire gate222_0n;
  wire gate219_0n;
  wire [31:0] complete216_0n;
  wire gate215_0n;
  wire [31:0] complete212_0n;
  wire icomplete_0n;
  C3 I0 (internal_0n[0], complete223_0n[0], complete223_0n[1], complete223_0n[2]);
  C3 I1 (internal_0n[1], complete223_0n[3], complete223_0n[4], complete223_0n[5]);
  C3 I2 (internal_0n[2], complete223_0n[6], complete223_0n[7], complete223_0n[8]);
  C3 I3 (internal_0n[3], complete223_0n[9], complete223_0n[10], complete223_0n[11]);
  C3 I4 (internal_0n[4], complete223_0n[12], complete223_0n[13], complete223_0n[14]);
  C3 I5 (internal_0n[5], complete223_0n[15], complete223_0n[16], complete223_0n[17]);
  C3 I6 (internal_0n[6], complete223_0n[18], complete223_0n[19], complete223_0n[20]);
  C3 I7 (internal_0n[7], complete223_0n[21], complete223_0n[22], complete223_0n[23]);
  C3 I8 (internal_0n[8], complete223_0n[24], complete223_0n[25], complete223_0n[26]);
  C3 I9 (internal_0n[9], complete223_0n[27], complete223_0n[28], complete223_0n[29]);
  C2 I10 (internal_0n[10], complete223_0n[30], complete223_0n[31]);
  C3 I11 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I12 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I13 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I14 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I15 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I16 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I17 (oaint_1n, internal_0n[15], internal_0n[16]);
  OR2 I18 (complete223_0n[0], o_1r0d[0], o_1r1d[0]);
  OR2 I19 (complete223_0n[1], o_1r0d[1], o_1r1d[1]);
  OR2 I20 (complete223_0n[2], o_1r0d[2], o_1r1d[2]);
  OR2 I21 (complete223_0n[3], o_1r0d[3], o_1r1d[3]);
  OR2 I22 (complete223_0n[4], o_1r0d[4], o_1r1d[4]);
  OR2 I23 (complete223_0n[5], o_1r0d[5], o_1r1d[5]);
  OR2 I24 (complete223_0n[6], o_1r0d[6], o_1r1d[6]);
  OR2 I25 (complete223_0n[7], o_1r0d[7], o_1r1d[7]);
  OR2 I26 (complete223_0n[8], o_1r0d[8], o_1r1d[8]);
  OR2 I27 (complete223_0n[9], o_1r0d[9], o_1r1d[9]);
  OR2 I28 (complete223_0n[10], o_1r0d[10], o_1r1d[10]);
  OR2 I29 (complete223_0n[11], o_1r0d[11], o_1r1d[11]);
  OR2 I30 (complete223_0n[12], o_1r0d[12], o_1r1d[12]);
  OR2 I31 (complete223_0n[13], o_1r0d[13], o_1r1d[13]);
  OR2 I32 (complete223_0n[14], o_1r0d[14], o_1r1d[14]);
  OR2 I33 (complete223_0n[15], o_1r0d[15], o_1r1d[15]);
  OR2 I34 (complete223_0n[16], o_1r0d[16], o_1r1d[16]);
  OR2 I35 (complete223_0n[17], o_1r0d[17], o_1r1d[17]);
  OR2 I36 (complete223_0n[18], o_1r0d[18], o_1r1d[18]);
  OR2 I37 (complete223_0n[19], o_1r0d[19], o_1r1d[19]);
  OR2 I38 (complete223_0n[20], o_1r0d[20], o_1r1d[20]);
  OR2 I39 (complete223_0n[21], o_1r0d[21], o_1r1d[21]);
  OR2 I40 (complete223_0n[22], o_1r0d[22], o_1r1d[22]);
  OR2 I41 (complete223_0n[23], o_1r0d[23], o_1r1d[23]);
  OR2 I42 (complete223_0n[24], o_1r0d[24], o_1r1d[24]);
  OR2 I43 (complete223_0n[25], o_1r0d[25], o_1r1d[25]);
  OR2 I44 (complete223_0n[26], o_1r0d[26], o_1r1d[26]);
  OR2 I45 (complete223_0n[27], o_1r0d[27], o_1r1d[27]);
  OR2 I46 (complete223_0n[28], o_1r0d[28], o_1r1d[28]);
  OR2 I47 (complete223_0n[29], o_1r0d[29], o_1r1d[29]);
  OR2 I48 (complete223_0n[30], o_1r0d[30], o_1r1d[30]);
  OR2 I49 (complete223_0n[31], o_1r0d[31], o_1r1d[31]);
  INV I50 (gate222_0n, o_1a);
  C2RI I51 (o_1r1d[0], otint_1n[0], gate222_0n, initialise);
  C2RI I52 (o_1r1d[1], otint_1n[1], gate222_0n, initialise);
  C2RI I53 (o_1r1d[2], otint_1n[2], gate222_0n, initialise);
  C2RI I54 (o_1r1d[3], otint_1n[3], gate222_0n, initialise);
  C2RI I55 (o_1r1d[4], otint_1n[4], gate222_0n, initialise);
  C2RI I56 (o_1r1d[5], otint_1n[5], gate222_0n, initialise);
  C2RI I57 (o_1r1d[6], otint_1n[6], gate222_0n, initialise);
  C2RI I58 (o_1r1d[7], otint_1n[7], gate222_0n, initialise);
  C2RI I59 (o_1r1d[8], otint_1n[8], gate222_0n, initialise);
  C2RI I60 (o_1r1d[9], otint_1n[9], gate222_0n, initialise);
  C2RI I61 (o_1r1d[10], otint_1n[10], gate222_0n, initialise);
  C2RI I62 (o_1r1d[11], otint_1n[11], gate222_0n, initialise);
  C2RI I63 (o_1r1d[12], otint_1n[12], gate222_0n, initialise);
  C2RI I64 (o_1r1d[13], otint_1n[13], gate222_0n, initialise);
  C2RI I65 (o_1r1d[14], otint_1n[14], gate222_0n, initialise);
  C2RI I66 (o_1r1d[15], otint_1n[15], gate222_0n, initialise);
  C2RI I67 (o_1r1d[16], otint_1n[16], gate222_0n, initialise);
  C2RI I68 (o_1r1d[17], otint_1n[17], gate222_0n, initialise);
  C2RI I69 (o_1r1d[18], otint_1n[18], gate222_0n, initialise);
  C2RI I70 (o_1r1d[19], otint_1n[19], gate222_0n, initialise);
  C2RI I71 (o_1r1d[20], otint_1n[20], gate222_0n, initialise);
  C2RI I72 (o_1r1d[21], otint_1n[21], gate222_0n, initialise);
  C2RI I73 (o_1r1d[22], otint_1n[22], gate222_0n, initialise);
  C2RI I74 (o_1r1d[23], otint_1n[23], gate222_0n, initialise);
  C2RI I75 (o_1r1d[24], otint_1n[24], gate222_0n, initialise);
  C2RI I76 (o_1r1d[25], otint_1n[25], gate222_0n, initialise);
  C2RI I77 (o_1r1d[26], otint_1n[26], gate222_0n, initialise);
  C2RI I78 (o_1r1d[27], otint_1n[27], gate222_0n, initialise);
  C2RI I79 (o_1r1d[28], otint_1n[28], gate222_0n, initialise);
  C2RI I80 (o_1r1d[29], otint_1n[29], gate222_0n, initialise);
  C2RI I81 (o_1r1d[30], otint_1n[30], gate222_0n, initialise);
  C2RI I82 (o_1r1d[31], otint_1n[31], gate222_0n, initialise);
  C2RI I83 (o_1r0d[0], ofint_1n[0], gate222_0n, initialise);
  C2RI I84 (o_1r0d[1], ofint_1n[1], gate222_0n, initialise);
  C2RI I85 (o_1r0d[2], ofint_1n[2], gate222_0n, initialise);
  C2RI I86 (o_1r0d[3], ofint_1n[3], gate222_0n, initialise);
  C2RI I87 (o_1r0d[4], ofint_1n[4], gate222_0n, initialise);
  C2RI I88 (o_1r0d[5], ofint_1n[5], gate222_0n, initialise);
  C2RI I89 (o_1r0d[6], ofint_1n[6], gate222_0n, initialise);
  C2RI I90 (o_1r0d[7], ofint_1n[7], gate222_0n, initialise);
  C2RI I91 (o_1r0d[8], ofint_1n[8], gate222_0n, initialise);
  C2RI I92 (o_1r0d[9], ofint_1n[9], gate222_0n, initialise);
  C2RI I93 (o_1r0d[10], ofint_1n[10], gate222_0n, initialise);
  C2RI I94 (o_1r0d[11], ofint_1n[11], gate222_0n, initialise);
  C2RI I95 (o_1r0d[12], ofint_1n[12], gate222_0n, initialise);
  C2RI I96 (o_1r0d[13], ofint_1n[13], gate222_0n, initialise);
  C2RI I97 (o_1r0d[14], ofint_1n[14], gate222_0n, initialise);
  C2RI I98 (o_1r0d[15], ofint_1n[15], gate222_0n, initialise);
  C2RI I99 (o_1r0d[16], ofint_1n[16], gate222_0n, initialise);
  C2RI I100 (o_1r0d[17], ofint_1n[17], gate222_0n, initialise);
  C2RI I101 (o_1r0d[18], ofint_1n[18], gate222_0n, initialise);
  C2RI I102 (o_1r0d[19], ofint_1n[19], gate222_0n, initialise);
  C2RI I103 (o_1r0d[20], ofint_1n[20], gate222_0n, initialise);
  C2RI I104 (o_1r0d[21], ofint_1n[21], gate222_0n, initialise);
  C2RI I105 (o_1r0d[22], ofint_1n[22], gate222_0n, initialise);
  C2RI I106 (o_1r0d[23], ofint_1n[23], gate222_0n, initialise);
  C2RI I107 (o_1r0d[24], ofint_1n[24], gate222_0n, initialise);
  C2RI I108 (o_1r0d[25], ofint_1n[25], gate222_0n, initialise);
  C2RI I109 (o_1r0d[26], ofint_1n[26], gate222_0n, initialise);
  C2RI I110 (o_1r0d[27], ofint_1n[27], gate222_0n, initialise);
  C2RI I111 (o_1r0d[28], ofint_1n[28], gate222_0n, initialise);
  C2RI I112 (o_1r0d[29], ofint_1n[29], gate222_0n, initialise);
  C2RI I113 (o_1r0d[30], ofint_1n[30], gate222_0n, initialise);
  C2RI I114 (o_1r0d[31], ofint_1n[31], gate222_0n, initialise);
  assign oaint_0n = o_0r;
  INV I116 (gate219_0n, o_0a);
  C2RI I117 (o_0r, ofint_0n, gate219_0n, initialise);
  C3 I118 (internal_0n[17], complete216_0n[0], complete216_0n[1], complete216_0n[2]);
  C3 I119 (internal_0n[18], complete216_0n[3], complete216_0n[4], complete216_0n[5]);
  C3 I120 (internal_0n[19], complete216_0n[6], complete216_0n[7], complete216_0n[8]);
  C3 I121 (internal_0n[20], complete216_0n[9], complete216_0n[10], complete216_0n[11]);
  C3 I122 (internal_0n[21], complete216_0n[12], complete216_0n[13], complete216_0n[14]);
  C3 I123 (internal_0n[22], complete216_0n[15], complete216_0n[16], complete216_0n[17]);
  C3 I124 (internal_0n[23], complete216_0n[18], complete216_0n[19], complete216_0n[20]);
  C3 I125 (internal_0n[24], complete216_0n[21], complete216_0n[22], complete216_0n[23]);
  C3 I126 (internal_0n[25], complete216_0n[24], complete216_0n[25], complete216_0n[26]);
  C3 I127 (internal_0n[26], complete216_0n[27], complete216_0n[28], complete216_0n[29]);
  C2 I128 (internal_0n[27], complete216_0n[30], complete216_0n[31]);
  C3 I129 (internal_0n[28], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I130 (internal_0n[29], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I131 (internal_0n[30], internal_0n[23], internal_0n[24], internal_0n[25]);
  C2 I132 (internal_0n[31], internal_0n[26], internal_0n[27]);
  C2 I133 (internal_0n[32], internal_0n[28], internal_0n[29]);
  C2 I134 (internal_0n[33], internal_0n[30], internal_0n[31]);
  C2 I135 (i_0a, internal_0n[32], internal_0n[33]);
  OR2 I136 (complete216_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I137 (complete216_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I138 (complete216_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I139 (complete216_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I140 (complete216_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I141 (complete216_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I142 (complete216_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I143 (complete216_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I144 (complete216_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I145 (complete216_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I146 (complete216_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I147 (complete216_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I148 (complete216_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I149 (complete216_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I150 (complete216_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I151 (complete216_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I152 (complete216_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I153 (complete216_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I154 (complete216_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I155 (complete216_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I156 (complete216_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I157 (complete216_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I158 (complete216_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I159 (complete216_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I160 (complete216_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I161 (complete216_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I162 (complete216_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I163 (complete216_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I164 (complete216_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I165 (complete216_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I166 (complete216_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I167 (complete216_0n[31], ifint_0n[31], itint_0n[31]);
  INV I168 (gate215_0n, iaint_0n);
  C2RI I169 (itint_0n[0], i_0r1d[0], gate215_0n, initialise);
  C2RI I170 (itint_0n[1], i_0r1d[1], gate215_0n, initialise);
  C2RI I171 (itint_0n[2], i_0r1d[2], gate215_0n, initialise);
  C2RI I172 (itint_0n[3], i_0r1d[3], gate215_0n, initialise);
  C2RI I173 (itint_0n[4], i_0r1d[4], gate215_0n, initialise);
  C2RI I174 (itint_0n[5], i_0r1d[5], gate215_0n, initialise);
  C2RI I175 (itint_0n[6], i_0r1d[6], gate215_0n, initialise);
  C2RI I176 (itint_0n[7], i_0r1d[7], gate215_0n, initialise);
  C2RI I177 (itint_0n[8], i_0r1d[8], gate215_0n, initialise);
  C2RI I178 (itint_0n[9], i_0r1d[9], gate215_0n, initialise);
  C2RI I179 (itint_0n[10], i_0r1d[10], gate215_0n, initialise);
  C2RI I180 (itint_0n[11], i_0r1d[11], gate215_0n, initialise);
  C2RI I181 (itint_0n[12], i_0r1d[12], gate215_0n, initialise);
  C2RI I182 (itint_0n[13], i_0r1d[13], gate215_0n, initialise);
  C2RI I183 (itint_0n[14], i_0r1d[14], gate215_0n, initialise);
  C2RI I184 (itint_0n[15], i_0r1d[15], gate215_0n, initialise);
  C2RI I185 (itint_0n[16], i_0r1d[16], gate215_0n, initialise);
  C2RI I186 (itint_0n[17], i_0r1d[17], gate215_0n, initialise);
  C2RI I187 (itint_0n[18], i_0r1d[18], gate215_0n, initialise);
  C2RI I188 (itint_0n[19], i_0r1d[19], gate215_0n, initialise);
  C2RI I189 (itint_0n[20], i_0r1d[20], gate215_0n, initialise);
  C2RI I190 (itint_0n[21], i_0r1d[21], gate215_0n, initialise);
  C2RI I191 (itint_0n[22], i_0r1d[22], gate215_0n, initialise);
  C2RI I192 (itint_0n[23], i_0r1d[23], gate215_0n, initialise);
  C2RI I193 (itint_0n[24], i_0r1d[24], gate215_0n, initialise);
  C2RI I194 (itint_0n[25], i_0r1d[25], gate215_0n, initialise);
  C2RI I195 (itint_0n[26], i_0r1d[26], gate215_0n, initialise);
  C2RI I196 (itint_0n[27], i_0r1d[27], gate215_0n, initialise);
  C2RI I197 (itint_0n[28], i_0r1d[28], gate215_0n, initialise);
  C2RI I198 (itint_0n[29], i_0r1d[29], gate215_0n, initialise);
  C2RI I199 (itint_0n[30], i_0r1d[30], gate215_0n, initialise);
  C2RI I200 (itint_0n[31], i_0r1d[31], gate215_0n, initialise);
  C2RI I201 (ifint_0n[0], i_0r0d[0], gate215_0n, initialise);
  C2RI I202 (ifint_0n[1], i_0r0d[1], gate215_0n, initialise);
  C2RI I203 (ifint_0n[2], i_0r0d[2], gate215_0n, initialise);
  C2RI I204 (ifint_0n[3], i_0r0d[3], gate215_0n, initialise);
  C2RI I205 (ifint_0n[4], i_0r0d[4], gate215_0n, initialise);
  C2RI I206 (ifint_0n[5], i_0r0d[5], gate215_0n, initialise);
  C2RI I207 (ifint_0n[6], i_0r0d[6], gate215_0n, initialise);
  C2RI I208 (ifint_0n[7], i_0r0d[7], gate215_0n, initialise);
  C2RI I209 (ifint_0n[8], i_0r0d[8], gate215_0n, initialise);
  C2RI I210 (ifint_0n[9], i_0r0d[9], gate215_0n, initialise);
  C2RI I211 (ifint_0n[10], i_0r0d[10], gate215_0n, initialise);
  C2RI I212 (ifint_0n[11], i_0r0d[11], gate215_0n, initialise);
  C2RI I213 (ifint_0n[12], i_0r0d[12], gate215_0n, initialise);
  C2RI I214 (ifint_0n[13], i_0r0d[13], gate215_0n, initialise);
  C2RI I215 (ifint_0n[14], i_0r0d[14], gate215_0n, initialise);
  C2RI I216 (ifint_0n[15], i_0r0d[15], gate215_0n, initialise);
  C2RI I217 (ifint_0n[16], i_0r0d[16], gate215_0n, initialise);
  C2RI I218 (ifint_0n[17], i_0r0d[17], gate215_0n, initialise);
  C2RI I219 (ifint_0n[18], i_0r0d[18], gate215_0n, initialise);
  C2RI I220 (ifint_0n[19], i_0r0d[19], gate215_0n, initialise);
  C2RI I221 (ifint_0n[20], i_0r0d[20], gate215_0n, initialise);
  C2RI I222 (ifint_0n[21], i_0r0d[21], gate215_0n, initialise);
  C2RI I223 (ifint_0n[22], i_0r0d[22], gate215_0n, initialise);
  C2RI I224 (ifint_0n[23], i_0r0d[23], gate215_0n, initialise);
  C2RI I225 (ifint_0n[24], i_0r0d[24], gate215_0n, initialise);
  C2RI I226 (ifint_0n[25], i_0r0d[25], gate215_0n, initialise);
  C2RI I227 (ifint_0n[26], i_0r0d[26], gate215_0n, initialise);
  C2RI I228 (ifint_0n[27], i_0r0d[27], gate215_0n, initialise);
  C2RI I229 (ifint_0n[28], i_0r0d[28], gate215_0n, initialise);
  C2RI I230 (ifint_0n[29], i_0r0d[29], gate215_0n, initialise);
  C2RI I231 (ifint_0n[30], i_0r0d[30], gate215_0n, initialise);
  C2RI I232 (ifint_0n[31], i_0r0d[31], gate215_0n, initialise);
  C3 I233 (iaint_0n, icomplete_0n, oaint_0n, oaint_1n);
  assign ofint_0n = icomplete_0n;
  assign otint_1n[0] = itint_0n[0];
  assign otint_1n[1] = itint_0n[1];
  assign otint_1n[2] = itint_0n[2];
  assign otint_1n[3] = itint_0n[3];
  assign otint_1n[4] = itint_0n[4];
  assign otint_1n[5] = itint_0n[5];
  assign otint_1n[6] = itint_0n[6];
  assign otint_1n[7] = itint_0n[7];
  assign otint_1n[8] = itint_0n[8];
  assign otint_1n[9] = itint_0n[9];
  assign otint_1n[10] = itint_0n[10];
  assign otint_1n[11] = itint_0n[11];
  assign otint_1n[12] = itint_0n[12];
  assign otint_1n[13] = itint_0n[13];
  assign otint_1n[14] = itint_0n[14];
  assign otint_1n[15] = itint_0n[15];
  assign otint_1n[16] = itint_0n[16];
  assign otint_1n[17] = itint_0n[17];
  assign otint_1n[18] = itint_0n[18];
  assign otint_1n[19] = itint_0n[19];
  assign otint_1n[20] = itint_0n[20];
  assign otint_1n[21] = itint_0n[21];
  assign otint_1n[22] = itint_0n[22];
  assign otint_1n[23] = itint_0n[23];
  assign otint_1n[24] = itint_0n[24];
  assign otint_1n[25] = itint_0n[25];
  assign otint_1n[26] = itint_0n[26];
  assign otint_1n[27] = itint_0n[27];
  assign otint_1n[28] = itint_0n[28];
  assign otint_1n[29] = itint_0n[29];
  assign otint_1n[30] = itint_0n[30];
  assign otint_1n[31] = itint_0n[31];
  assign ofint_1n[0] = ifint_0n[0];
  assign ofint_1n[1] = ifint_0n[1];
  assign ofint_1n[2] = ifint_0n[2];
  assign ofint_1n[3] = ifint_0n[3];
  assign ofint_1n[4] = ifint_0n[4];
  assign ofint_1n[5] = ifint_0n[5];
  assign ofint_1n[6] = ifint_0n[6];
  assign ofint_1n[7] = ifint_0n[7];
  assign ofint_1n[8] = ifint_0n[8];
  assign ofint_1n[9] = ifint_0n[9];
  assign ofint_1n[10] = ifint_0n[10];
  assign ofint_1n[11] = ifint_0n[11];
  assign ofint_1n[12] = ifint_0n[12];
  assign ofint_1n[13] = ifint_0n[13];
  assign ofint_1n[14] = ifint_0n[14];
  assign ofint_1n[15] = ifint_0n[15];
  assign ofint_1n[16] = ifint_0n[16];
  assign ofint_1n[17] = ifint_0n[17];
  assign ofint_1n[18] = ifint_0n[18];
  assign ofint_1n[19] = ifint_0n[19];
  assign ofint_1n[20] = ifint_0n[20];
  assign ofint_1n[21] = ifint_0n[21];
  assign ofint_1n[22] = ifint_0n[22];
  assign ofint_1n[23] = ifint_0n[23];
  assign ofint_1n[24] = ifint_0n[24];
  assign ofint_1n[25] = ifint_0n[25];
  assign ofint_1n[26] = ifint_0n[26];
  assign ofint_1n[27] = ifint_0n[27];
  assign ofint_1n[28] = ifint_0n[28];
  assign ofint_1n[29] = ifint_0n[29];
  assign ofint_1n[30] = ifint_0n[30];
  assign ofint_1n[31] = ifint_0n[31];
  C3 I299 (internal_0n[34], complete212_0n[0], complete212_0n[1], complete212_0n[2]);
  C3 I300 (internal_0n[35], complete212_0n[3], complete212_0n[4], complete212_0n[5]);
  C3 I301 (internal_0n[36], complete212_0n[6], complete212_0n[7], complete212_0n[8]);
  C3 I302 (internal_0n[37], complete212_0n[9], complete212_0n[10], complete212_0n[11]);
  C3 I303 (internal_0n[38], complete212_0n[12], complete212_0n[13], complete212_0n[14]);
  C3 I304 (internal_0n[39], complete212_0n[15], complete212_0n[16], complete212_0n[17]);
  C3 I305 (internal_0n[40], complete212_0n[18], complete212_0n[19], complete212_0n[20]);
  C3 I306 (internal_0n[41], complete212_0n[21], complete212_0n[22], complete212_0n[23]);
  C3 I307 (internal_0n[42], complete212_0n[24], complete212_0n[25], complete212_0n[26]);
  C3 I308 (internal_0n[43], complete212_0n[27], complete212_0n[28], complete212_0n[29]);
  C2 I309 (internal_0n[44], complete212_0n[30], complete212_0n[31]);
  C3 I310 (internal_0n[45], internal_0n[34], internal_0n[35], internal_0n[36]);
  C3 I311 (internal_0n[46], internal_0n[37], internal_0n[38], internal_0n[39]);
  C3 I312 (internal_0n[47], internal_0n[40], internal_0n[41], internal_0n[42]);
  C2 I313 (internal_0n[48], internal_0n[43], internal_0n[44]);
  C2 I314 (internal_0n[49], internal_0n[45], internal_0n[46]);
  C2 I315 (internal_0n[50], internal_0n[47], internal_0n[48]);
  C2 I316 (icomplete_0n, internal_0n[49], internal_0n[50]);
  OR2 I317 (complete212_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I318 (complete212_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I319 (complete212_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I320 (complete212_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I321 (complete212_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I322 (complete212_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I323 (complete212_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I324 (complete212_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I325 (complete212_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I326 (complete212_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I327 (complete212_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I328 (complete212_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I329 (complete212_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I330 (complete212_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I331 (complete212_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I332 (complete212_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I333 (complete212_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I334 (complete212_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I335 (complete212_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I336 (complete212_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I337 (complete212_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I338 (complete212_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I339 (complete212_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I340 (complete212_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I341 (complete212_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I342 (complete212_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I343 (complete212_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I344 (complete212_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I345 (complete212_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I346 (complete212_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I347 (complete212_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I348 (complete212_0n[31], ifint_0n[31], itint_0n[31]);
endmodule

module BrzF_33_l32__28_280_200_29_20_280_2033_29__m41m (
  i_0r0d, i_0r1d, i_0a,
  o_0r, o_0a,
  o_1r0d, o_1r1d, o_1a,
  initialise
);
  input [32:0] i_0r0d;
  input [32:0] i_0r1d;
  output i_0a;
  output o_0r;
  input o_0a;
  output [32:0] o_1r0d;
  output [32:0] o_1r1d;
  input o_1a;
  input initialise;
  wire [50:0] internal_0n;
  wire [32:0] ifint_0n;
  wire [32:0] itint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire [32:0] ofint_1n;
  wire [32:0] otint_1n;
  wire oaint_0n;
  wire oaint_1n;
  wire [32:0] complete235_0n;
  wire gate234_0n;
  wire gate231_0n;
  wire [32:0] complete228_0n;
  wire gate227_0n;
  wire [32:0] complete224_0n;
  wire icomplete_0n;
  C3 I0 (internal_0n[0], complete235_0n[0], complete235_0n[1], complete235_0n[2]);
  C3 I1 (internal_0n[1], complete235_0n[3], complete235_0n[4], complete235_0n[5]);
  C3 I2 (internal_0n[2], complete235_0n[6], complete235_0n[7], complete235_0n[8]);
  C3 I3 (internal_0n[3], complete235_0n[9], complete235_0n[10], complete235_0n[11]);
  C3 I4 (internal_0n[4], complete235_0n[12], complete235_0n[13], complete235_0n[14]);
  C3 I5 (internal_0n[5], complete235_0n[15], complete235_0n[16], complete235_0n[17]);
  C3 I6 (internal_0n[6], complete235_0n[18], complete235_0n[19], complete235_0n[20]);
  C3 I7 (internal_0n[7], complete235_0n[21], complete235_0n[22], complete235_0n[23]);
  C3 I8 (internal_0n[8], complete235_0n[24], complete235_0n[25], complete235_0n[26]);
  C3 I9 (internal_0n[9], complete235_0n[27], complete235_0n[28], complete235_0n[29]);
  C3 I10 (internal_0n[10], complete235_0n[30], complete235_0n[31], complete235_0n[32]);
  C3 I11 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I12 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I13 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I14 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I15 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I16 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I17 (oaint_1n, internal_0n[15], internal_0n[16]);
  OR2 I18 (complete235_0n[0], o_1r0d[0], o_1r1d[0]);
  OR2 I19 (complete235_0n[1], o_1r0d[1], o_1r1d[1]);
  OR2 I20 (complete235_0n[2], o_1r0d[2], o_1r1d[2]);
  OR2 I21 (complete235_0n[3], o_1r0d[3], o_1r1d[3]);
  OR2 I22 (complete235_0n[4], o_1r0d[4], o_1r1d[4]);
  OR2 I23 (complete235_0n[5], o_1r0d[5], o_1r1d[5]);
  OR2 I24 (complete235_0n[6], o_1r0d[6], o_1r1d[6]);
  OR2 I25 (complete235_0n[7], o_1r0d[7], o_1r1d[7]);
  OR2 I26 (complete235_0n[8], o_1r0d[8], o_1r1d[8]);
  OR2 I27 (complete235_0n[9], o_1r0d[9], o_1r1d[9]);
  OR2 I28 (complete235_0n[10], o_1r0d[10], o_1r1d[10]);
  OR2 I29 (complete235_0n[11], o_1r0d[11], o_1r1d[11]);
  OR2 I30 (complete235_0n[12], o_1r0d[12], o_1r1d[12]);
  OR2 I31 (complete235_0n[13], o_1r0d[13], o_1r1d[13]);
  OR2 I32 (complete235_0n[14], o_1r0d[14], o_1r1d[14]);
  OR2 I33 (complete235_0n[15], o_1r0d[15], o_1r1d[15]);
  OR2 I34 (complete235_0n[16], o_1r0d[16], o_1r1d[16]);
  OR2 I35 (complete235_0n[17], o_1r0d[17], o_1r1d[17]);
  OR2 I36 (complete235_0n[18], o_1r0d[18], o_1r1d[18]);
  OR2 I37 (complete235_0n[19], o_1r0d[19], o_1r1d[19]);
  OR2 I38 (complete235_0n[20], o_1r0d[20], o_1r1d[20]);
  OR2 I39 (complete235_0n[21], o_1r0d[21], o_1r1d[21]);
  OR2 I40 (complete235_0n[22], o_1r0d[22], o_1r1d[22]);
  OR2 I41 (complete235_0n[23], o_1r0d[23], o_1r1d[23]);
  OR2 I42 (complete235_0n[24], o_1r0d[24], o_1r1d[24]);
  OR2 I43 (complete235_0n[25], o_1r0d[25], o_1r1d[25]);
  OR2 I44 (complete235_0n[26], o_1r0d[26], o_1r1d[26]);
  OR2 I45 (complete235_0n[27], o_1r0d[27], o_1r1d[27]);
  OR2 I46 (complete235_0n[28], o_1r0d[28], o_1r1d[28]);
  OR2 I47 (complete235_0n[29], o_1r0d[29], o_1r1d[29]);
  OR2 I48 (complete235_0n[30], o_1r0d[30], o_1r1d[30]);
  OR2 I49 (complete235_0n[31], o_1r0d[31], o_1r1d[31]);
  OR2 I50 (complete235_0n[32], o_1r0d[32], o_1r1d[32]);
  INV I51 (gate234_0n, o_1a);
  C2RI I52 (o_1r1d[0], otint_1n[0], gate234_0n, initialise);
  C2RI I53 (o_1r1d[1], otint_1n[1], gate234_0n, initialise);
  C2RI I54 (o_1r1d[2], otint_1n[2], gate234_0n, initialise);
  C2RI I55 (o_1r1d[3], otint_1n[3], gate234_0n, initialise);
  C2RI I56 (o_1r1d[4], otint_1n[4], gate234_0n, initialise);
  C2RI I57 (o_1r1d[5], otint_1n[5], gate234_0n, initialise);
  C2RI I58 (o_1r1d[6], otint_1n[6], gate234_0n, initialise);
  C2RI I59 (o_1r1d[7], otint_1n[7], gate234_0n, initialise);
  C2RI I60 (o_1r1d[8], otint_1n[8], gate234_0n, initialise);
  C2RI I61 (o_1r1d[9], otint_1n[9], gate234_0n, initialise);
  C2RI I62 (o_1r1d[10], otint_1n[10], gate234_0n, initialise);
  C2RI I63 (o_1r1d[11], otint_1n[11], gate234_0n, initialise);
  C2RI I64 (o_1r1d[12], otint_1n[12], gate234_0n, initialise);
  C2RI I65 (o_1r1d[13], otint_1n[13], gate234_0n, initialise);
  C2RI I66 (o_1r1d[14], otint_1n[14], gate234_0n, initialise);
  C2RI I67 (o_1r1d[15], otint_1n[15], gate234_0n, initialise);
  C2RI I68 (o_1r1d[16], otint_1n[16], gate234_0n, initialise);
  C2RI I69 (o_1r1d[17], otint_1n[17], gate234_0n, initialise);
  C2RI I70 (o_1r1d[18], otint_1n[18], gate234_0n, initialise);
  C2RI I71 (o_1r1d[19], otint_1n[19], gate234_0n, initialise);
  C2RI I72 (o_1r1d[20], otint_1n[20], gate234_0n, initialise);
  C2RI I73 (o_1r1d[21], otint_1n[21], gate234_0n, initialise);
  C2RI I74 (o_1r1d[22], otint_1n[22], gate234_0n, initialise);
  C2RI I75 (o_1r1d[23], otint_1n[23], gate234_0n, initialise);
  C2RI I76 (o_1r1d[24], otint_1n[24], gate234_0n, initialise);
  C2RI I77 (o_1r1d[25], otint_1n[25], gate234_0n, initialise);
  C2RI I78 (o_1r1d[26], otint_1n[26], gate234_0n, initialise);
  C2RI I79 (o_1r1d[27], otint_1n[27], gate234_0n, initialise);
  C2RI I80 (o_1r1d[28], otint_1n[28], gate234_0n, initialise);
  C2RI I81 (o_1r1d[29], otint_1n[29], gate234_0n, initialise);
  C2RI I82 (o_1r1d[30], otint_1n[30], gate234_0n, initialise);
  C2RI I83 (o_1r1d[31], otint_1n[31], gate234_0n, initialise);
  C2RI I84 (o_1r1d[32], otint_1n[32], gate234_0n, initialise);
  C2RI I85 (o_1r0d[0], ofint_1n[0], gate234_0n, initialise);
  C2RI I86 (o_1r0d[1], ofint_1n[1], gate234_0n, initialise);
  C2RI I87 (o_1r0d[2], ofint_1n[2], gate234_0n, initialise);
  C2RI I88 (o_1r0d[3], ofint_1n[3], gate234_0n, initialise);
  C2RI I89 (o_1r0d[4], ofint_1n[4], gate234_0n, initialise);
  C2RI I90 (o_1r0d[5], ofint_1n[5], gate234_0n, initialise);
  C2RI I91 (o_1r0d[6], ofint_1n[6], gate234_0n, initialise);
  C2RI I92 (o_1r0d[7], ofint_1n[7], gate234_0n, initialise);
  C2RI I93 (o_1r0d[8], ofint_1n[8], gate234_0n, initialise);
  C2RI I94 (o_1r0d[9], ofint_1n[9], gate234_0n, initialise);
  C2RI I95 (o_1r0d[10], ofint_1n[10], gate234_0n, initialise);
  C2RI I96 (o_1r0d[11], ofint_1n[11], gate234_0n, initialise);
  C2RI I97 (o_1r0d[12], ofint_1n[12], gate234_0n, initialise);
  C2RI I98 (o_1r0d[13], ofint_1n[13], gate234_0n, initialise);
  C2RI I99 (o_1r0d[14], ofint_1n[14], gate234_0n, initialise);
  C2RI I100 (o_1r0d[15], ofint_1n[15], gate234_0n, initialise);
  C2RI I101 (o_1r0d[16], ofint_1n[16], gate234_0n, initialise);
  C2RI I102 (o_1r0d[17], ofint_1n[17], gate234_0n, initialise);
  C2RI I103 (o_1r0d[18], ofint_1n[18], gate234_0n, initialise);
  C2RI I104 (o_1r0d[19], ofint_1n[19], gate234_0n, initialise);
  C2RI I105 (o_1r0d[20], ofint_1n[20], gate234_0n, initialise);
  C2RI I106 (o_1r0d[21], ofint_1n[21], gate234_0n, initialise);
  C2RI I107 (o_1r0d[22], ofint_1n[22], gate234_0n, initialise);
  C2RI I108 (o_1r0d[23], ofint_1n[23], gate234_0n, initialise);
  C2RI I109 (o_1r0d[24], ofint_1n[24], gate234_0n, initialise);
  C2RI I110 (o_1r0d[25], ofint_1n[25], gate234_0n, initialise);
  C2RI I111 (o_1r0d[26], ofint_1n[26], gate234_0n, initialise);
  C2RI I112 (o_1r0d[27], ofint_1n[27], gate234_0n, initialise);
  C2RI I113 (o_1r0d[28], ofint_1n[28], gate234_0n, initialise);
  C2RI I114 (o_1r0d[29], ofint_1n[29], gate234_0n, initialise);
  C2RI I115 (o_1r0d[30], ofint_1n[30], gate234_0n, initialise);
  C2RI I116 (o_1r0d[31], ofint_1n[31], gate234_0n, initialise);
  C2RI I117 (o_1r0d[32], ofint_1n[32], gate234_0n, initialise);
  assign oaint_0n = o_0r;
  INV I119 (gate231_0n, o_0a);
  C2RI I120 (o_0r, ofint_0n, gate231_0n, initialise);
  C3 I121 (internal_0n[17], complete228_0n[0], complete228_0n[1], complete228_0n[2]);
  C3 I122 (internal_0n[18], complete228_0n[3], complete228_0n[4], complete228_0n[5]);
  C3 I123 (internal_0n[19], complete228_0n[6], complete228_0n[7], complete228_0n[8]);
  C3 I124 (internal_0n[20], complete228_0n[9], complete228_0n[10], complete228_0n[11]);
  C3 I125 (internal_0n[21], complete228_0n[12], complete228_0n[13], complete228_0n[14]);
  C3 I126 (internal_0n[22], complete228_0n[15], complete228_0n[16], complete228_0n[17]);
  C3 I127 (internal_0n[23], complete228_0n[18], complete228_0n[19], complete228_0n[20]);
  C3 I128 (internal_0n[24], complete228_0n[21], complete228_0n[22], complete228_0n[23]);
  C3 I129 (internal_0n[25], complete228_0n[24], complete228_0n[25], complete228_0n[26]);
  C3 I130 (internal_0n[26], complete228_0n[27], complete228_0n[28], complete228_0n[29]);
  C3 I131 (internal_0n[27], complete228_0n[30], complete228_0n[31], complete228_0n[32]);
  C3 I132 (internal_0n[28], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I133 (internal_0n[29], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I134 (internal_0n[30], internal_0n[23], internal_0n[24], internal_0n[25]);
  C2 I135 (internal_0n[31], internal_0n[26], internal_0n[27]);
  C2 I136 (internal_0n[32], internal_0n[28], internal_0n[29]);
  C2 I137 (internal_0n[33], internal_0n[30], internal_0n[31]);
  C2 I138 (i_0a, internal_0n[32], internal_0n[33]);
  OR2 I139 (complete228_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I140 (complete228_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I141 (complete228_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I142 (complete228_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I143 (complete228_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I144 (complete228_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I145 (complete228_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I146 (complete228_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I147 (complete228_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I148 (complete228_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I149 (complete228_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I150 (complete228_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I151 (complete228_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I152 (complete228_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I153 (complete228_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I154 (complete228_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I155 (complete228_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I156 (complete228_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I157 (complete228_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I158 (complete228_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I159 (complete228_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I160 (complete228_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I161 (complete228_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I162 (complete228_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I163 (complete228_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I164 (complete228_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I165 (complete228_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I166 (complete228_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I167 (complete228_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I168 (complete228_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I169 (complete228_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I170 (complete228_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I171 (complete228_0n[32], ifint_0n[32], itint_0n[32]);
  INV I172 (gate227_0n, iaint_0n);
  C2RI I173 (itint_0n[0], i_0r1d[0], gate227_0n, initialise);
  C2RI I174 (itint_0n[1], i_0r1d[1], gate227_0n, initialise);
  C2RI I175 (itint_0n[2], i_0r1d[2], gate227_0n, initialise);
  C2RI I176 (itint_0n[3], i_0r1d[3], gate227_0n, initialise);
  C2RI I177 (itint_0n[4], i_0r1d[4], gate227_0n, initialise);
  C2RI I178 (itint_0n[5], i_0r1d[5], gate227_0n, initialise);
  C2RI I179 (itint_0n[6], i_0r1d[6], gate227_0n, initialise);
  C2RI I180 (itint_0n[7], i_0r1d[7], gate227_0n, initialise);
  C2RI I181 (itint_0n[8], i_0r1d[8], gate227_0n, initialise);
  C2RI I182 (itint_0n[9], i_0r1d[9], gate227_0n, initialise);
  C2RI I183 (itint_0n[10], i_0r1d[10], gate227_0n, initialise);
  C2RI I184 (itint_0n[11], i_0r1d[11], gate227_0n, initialise);
  C2RI I185 (itint_0n[12], i_0r1d[12], gate227_0n, initialise);
  C2RI I186 (itint_0n[13], i_0r1d[13], gate227_0n, initialise);
  C2RI I187 (itint_0n[14], i_0r1d[14], gate227_0n, initialise);
  C2RI I188 (itint_0n[15], i_0r1d[15], gate227_0n, initialise);
  C2RI I189 (itint_0n[16], i_0r1d[16], gate227_0n, initialise);
  C2RI I190 (itint_0n[17], i_0r1d[17], gate227_0n, initialise);
  C2RI I191 (itint_0n[18], i_0r1d[18], gate227_0n, initialise);
  C2RI I192 (itint_0n[19], i_0r1d[19], gate227_0n, initialise);
  C2RI I193 (itint_0n[20], i_0r1d[20], gate227_0n, initialise);
  C2RI I194 (itint_0n[21], i_0r1d[21], gate227_0n, initialise);
  C2RI I195 (itint_0n[22], i_0r1d[22], gate227_0n, initialise);
  C2RI I196 (itint_0n[23], i_0r1d[23], gate227_0n, initialise);
  C2RI I197 (itint_0n[24], i_0r1d[24], gate227_0n, initialise);
  C2RI I198 (itint_0n[25], i_0r1d[25], gate227_0n, initialise);
  C2RI I199 (itint_0n[26], i_0r1d[26], gate227_0n, initialise);
  C2RI I200 (itint_0n[27], i_0r1d[27], gate227_0n, initialise);
  C2RI I201 (itint_0n[28], i_0r1d[28], gate227_0n, initialise);
  C2RI I202 (itint_0n[29], i_0r1d[29], gate227_0n, initialise);
  C2RI I203 (itint_0n[30], i_0r1d[30], gate227_0n, initialise);
  C2RI I204 (itint_0n[31], i_0r1d[31], gate227_0n, initialise);
  C2RI I205 (itint_0n[32], i_0r1d[32], gate227_0n, initialise);
  C2RI I206 (ifint_0n[0], i_0r0d[0], gate227_0n, initialise);
  C2RI I207 (ifint_0n[1], i_0r0d[1], gate227_0n, initialise);
  C2RI I208 (ifint_0n[2], i_0r0d[2], gate227_0n, initialise);
  C2RI I209 (ifint_0n[3], i_0r0d[3], gate227_0n, initialise);
  C2RI I210 (ifint_0n[4], i_0r0d[4], gate227_0n, initialise);
  C2RI I211 (ifint_0n[5], i_0r0d[5], gate227_0n, initialise);
  C2RI I212 (ifint_0n[6], i_0r0d[6], gate227_0n, initialise);
  C2RI I213 (ifint_0n[7], i_0r0d[7], gate227_0n, initialise);
  C2RI I214 (ifint_0n[8], i_0r0d[8], gate227_0n, initialise);
  C2RI I215 (ifint_0n[9], i_0r0d[9], gate227_0n, initialise);
  C2RI I216 (ifint_0n[10], i_0r0d[10], gate227_0n, initialise);
  C2RI I217 (ifint_0n[11], i_0r0d[11], gate227_0n, initialise);
  C2RI I218 (ifint_0n[12], i_0r0d[12], gate227_0n, initialise);
  C2RI I219 (ifint_0n[13], i_0r0d[13], gate227_0n, initialise);
  C2RI I220 (ifint_0n[14], i_0r0d[14], gate227_0n, initialise);
  C2RI I221 (ifint_0n[15], i_0r0d[15], gate227_0n, initialise);
  C2RI I222 (ifint_0n[16], i_0r0d[16], gate227_0n, initialise);
  C2RI I223 (ifint_0n[17], i_0r0d[17], gate227_0n, initialise);
  C2RI I224 (ifint_0n[18], i_0r0d[18], gate227_0n, initialise);
  C2RI I225 (ifint_0n[19], i_0r0d[19], gate227_0n, initialise);
  C2RI I226 (ifint_0n[20], i_0r0d[20], gate227_0n, initialise);
  C2RI I227 (ifint_0n[21], i_0r0d[21], gate227_0n, initialise);
  C2RI I228 (ifint_0n[22], i_0r0d[22], gate227_0n, initialise);
  C2RI I229 (ifint_0n[23], i_0r0d[23], gate227_0n, initialise);
  C2RI I230 (ifint_0n[24], i_0r0d[24], gate227_0n, initialise);
  C2RI I231 (ifint_0n[25], i_0r0d[25], gate227_0n, initialise);
  C2RI I232 (ifint_0n[26], i_0r0d[26], gate227_0n, initialise);
  C2RI I233 (ifint_0n[27], i_0r0d[27], gate227_0n, initialise);
  C2RI I234 (ifint_0n[28], i_0r0d[28], gate227_0n, initialise);
  C2RI I235 (ifint_0n[29], i_0r0d[29], gate227_0n, initialise);
  C2RI I236 (ifint_0n[30], i_0r0d[30], gate227_0n, initialise);
  C2RI I237 (ifint_0n[31], i_0r0d[31], gate227_0n, initialise);
  C2RI I238 (ifint_0n[32], i_0r0d[32], gate227_0n, initialise);
  C3 I239 (iaint_0n, icomplete_0n, oaint_0n, oaint_1n);
  assign ofint_0n = icomplete_0n;
  assign otint_1n[0] = itint_0n[0];
  assign otint_1n[1] = itint_0n[1];
  assign otint_1n[2] = itint_0n[2];
  assign otint_1n[3] = itint_0n[3];
  assign otint_1n[4] = itint_0n[4];
  assign otint_1n[5] = itint_0n[5];
  assign otint_1n[6] = itint_0n[6];
  assign otint_1n[7] = itint_0n[7];
  assign otint_1n[8] = itint_0n[8];
  assign otint_1n[9] = itint_0n[9];
  assign otint_1n[10] = itint_0n[10];
  assign otint_1n[11] = itint_0n[11];
  assign otint_1n[12] = itint_0n[12];
  assign otint_1n[13] = itint_0n[13];
  assign otint_1n[14] = itint_0n[14];
  assign otint_1n[15] = itint_0n[15];
  assign otint_1n[16] = itint_0n[16];
  assign otint_1n[17] = itint_0n[17];
  assign otint_1n[18] = itint_0n[18];
  assign otint_1n[19] = itint_0n[19];
  assign otint_1n[20] = itint_0n[20];
  assign otint_1n[21] = itint_0n[21];
  assign otint_1n[22] = itint_0n[22];
  assign otint_1n[23] = itint_0n[23];
  assign otint_1n[24] = itint_0n[24];
  assign otint_1n[25] = itint_0n[25];
  assign otint_1n[26] = itint_0n[26];
  assign otint_1n[27] = itint_0n[27];
  assign otint_1n[28] = itint_0n[28];
  assign otint_1n[29] = itint_0n[29];
  assign otint_1n[30] = itint_0n[30];
  assign otint_1n[31] = itint_0n[31];
  assign otint_1n[32] = itint_0n[32];
  assign ofint_1n[0] = ifint_0n[0];
  assign ofint_1n[1] = ifint_0n[1];
  assign ofint_1n[2] = ifint_0n[2];
  assign ofint_1n[3] = ifint_0n[3];
  assign ofint_1n[4] = ifint_0n[4];
  assign ofint_1n[5] = ifint_0n[5];
  assign ofint_1n[6] = ifint_0n[6];
  assign ofint_1n[7] = ifint_0n[7];
  assign ofint_1n[8] = ifint_0n[8];
  assign ofint_1n[9] = ifint_0n[9];
  assign ofint_1n[10] = ifint_0n[10];
  assign ofint_1n[11] = ifint_0n[11];
  assign ofint_1n[12] = ifint_0n[12];
  assign ofint_1n[13] = ifint_0n[13];
  assign ofint_1n[14] = ifint_0n[14];
  assign ofint_1n[15] = ifint_0n[15];
  assign ofint_1n[16] = ifint_0n[16];
  assign ofint_1n[17] = ifint_0n[17];
  assign ofint_1n[18] = ifint_0n[18];
  assign ofint_1n[19] = ifint_0n[19];
  assign ofint_1n[20] = ifint_0n[20];
  assign ofint_1n[21] = ifint_0n[21];
  assign ofint_1n[22] = ifint_0n[22];
  assign ofint_1n[23] = ifint_0n[23];
  assign ofint_1n[24] = ifint_0n[24];
  assign ofint_1n[25] = ifint_0n[25];
  assign ofint_1n[26] = ifint_0n[26];
  assign ofint_1n[27] = ifint_0n[27];
  assign ofint_1n[28] = ifint_0n[28];
  assign ofint_1n[29] = ifint_0n[29];
  assign ofint_1n[30] = ifint_0n[30];
  assign ofint_1n[31] = ifint_0n[31];
  assign ofint_1n[32] = ifint_0n[32];
  C3 I307 (internal_0n[34], complete224_0n[0], complete224_0n[1], complete224_0n[2]);
  C3 I308 (internal_0n[35], complete224_0n[3], complete224_0n[4], complete224_0n[5]);
  C3 I309 (internal_0n[36], complete224_0n[6], complete224_0n[7], complete224_0n[8]);
  C3 I310 (internal_0n[37], complete224_0n[9], complete224_0n[10], complete224_0n[11]);
  C3 I311 (internal_0n[38], complete224_0n[12], complete224_0n[13], complete224_0n[14]);
  C3 I312 (internal_0n[39], complete224_0n[15], complete224_0n[16], complete224_0n[17]);
  C3 I313 (internal_0n[40], complete224_0n[18], complete224_0n[19], complete224_0n[20]);
  C3 I314 (internal_0n[41], complete224_0n[21], complete224_0n[22], complete224_0n[23]);
  C3 I315 (internal_0n[42], complete224_0n[24], complete224_0n[25], complete224_0n[26]);
  C3 I316 (internal_0n[43], complete224_0n[27], complete224_0n[28], complete224_0n[29]);
  C3 I317 (internal_0n[44], complete224_0n[30], complete224_0n[31], complete224_0n[32]);
  C3 I318 (internal_0n[45], internal_0n[34], internal_0n[35], internal_0n[36]);
  C3 I319 (internal_0n[46], internal_0n[37], internal_0n[38], internal_0n[39]);
  C3 I320 (internal_0n[47], internal_0n[40], internal_0n[41], internal_0n[42]);
  C2 I321 (internal_0n[48], internal_0n[43], internal_0n[44]);
  C2 I322 (internal_0n[49], internal_0n[45], internal_0n[46]);
  C2 I323 (internal_0n[50], internal_0n[47], internal_0n[48]);
  C2 I324 (icomplete_0n, internal_0n[49], internal_0n[50]);
  OR2 I325 (complete224_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I326 (complete224_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I327 (complete224_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I328 (complete224_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I329 (complete224_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I330 (complete224_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I331 (complete224_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I332 (complete224_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I333 (complete224_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I334 (complete224_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I335 (complete224_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I336 (complete224_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I337 (complete224_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I338 (complete224_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I339 (complete224_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I340 (complete224_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I341 (complete224_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I342 (complete224_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I343 (complete224_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I344 (complete224_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I345 (complete224_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I346 (complete224_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I347 (complete224_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I348 (complete224_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I349 (complete224_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I350 (complete224_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I351 (complete224_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I352 (complete224_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I353 (complete224_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I354 (complete224_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I355 (complete224_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I356 (complete224_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I357 (complete224_0n[32], ifint_0n[32], itint_0n[32]);
endmodule

module BrzF_34_l32__28_280_200_29_20_280_2034_29__m42m (
  i_0r0d, i_0r1d, i_0a,
  o_0r, o_0a,
  o_1r0d, o_1r1d, o_1a,
  initialise
);
  input [33:0] i_0r0d;
  input [33:0] i_0r1d;
  output i_0a;
  output o_0r;
  input o_0a;
  output [33:0] o_1r0d;
  output [33:0] o_1r1d;
  input o_1a;
  input initialise;
  wire [53:0] internal_0n;
  wire [33:0] ifint_0n;
  wire [33:0] itint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire [33:0] ofint_1n;
  wire [33:0] otint_1n;
  wire oaint_0n;
  wire oaint_1n;
  wire [33:0] complete247_0n;
  wire gate246_0n;
  wire gate243_0n;
  wire [33:0] complete240_0n;
  wire gate239_0n;
  wire [33:0] complete236_0n;
  wire icomplete_0n;
  C3 I0 (internal_0n[0], complete247_0n[0], complete247_0n[1], complete247_0n[2]);
  C3 I1 (internal_0n[1], complete247_0n[3], complete247_0n[4], complete247_0n[5]);
  C3 I2 (internal_0n[2], complete247_0n[6], complete247_0n[7], complete247_0n[8]);
  C3 I3 (internal_0n[3], complete247_0n[9], complete247_0n[10], complete247_0n[11]);
  C3 I4 (internal_0n[4], complete247_0n[12], complete247_0n[13], complete247_0n[14]);
  C3 I5 (internal_0n[5], complete247_0n[15], complete247_0n[16], complete247_0n[17]);
  C3 I6 (internal_0n[6], complete247_0n[18], complete247_0n[19], complete247_0n[20]);
  C3 I7 (internal_0n[7], complete247_0n[21], complete247_0n[22], complete247_0n[23]);
  C3 I8 (internal_0n[8], complete247_0n[24], complete247_0n[25], complete247_0n[26]);
  C3 I9 (internal_0n[9], complete247_0n[27], complete247_0n[28], complete247_0n[29]);
  C2 I10 (internal_0n[10], complete247_0n[30], complete247_0n[31]);
  C2 I11 (internal_0n[11], complete247_0n[32], complete247_0n[33]);
  C3 I12 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I13 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I14 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I15 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I16 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I17 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I18 (oaint_1n, internal_0n[16], internal_0n[17]);
  OR2 I19 (complete247_0n[0], o_1r0d[0], o_1r1d[0]);
  OR2 I20 (complete247_0n[1], o_1r0d[1], o_1r1d[1]);
  OR2 I21 (complete247_0n[2], o_1r0d[2], o_1r1d[2]);
  OR2 I22 (complete247_0n[3], o_1r0d[3], o_1r1d[3]);
  OR2 I23 (complete247_0n[4], o_1r0d[4], o_1r1d[4]);
  OR2 I24 (complete247_0n[5], o_1r0d[5], o_1r1d[5]);
  OR2 I25 (complete247_0n[6], o_1r0d[6], o_1r1d[6]);
  OR2 I26 (complete247_0n[7], o_1r0d[7], o_1r1d[7]);
  OR2 I27 (complete247_0n[8], o_1r0d[8], o_1r1d[8]);
  OR2 I28 (complete247_0n[9], o_1r0d[9], o_1r1d[9]);
  OR2 I29 (complete247_0n[10], o_1r0d[10], o_1r1d[10]);
  OR2 I30 (complete247_0n[11], o_1r0d[11], o_1r1d[11]);
  OR2 I31 (complete247_0n[12], o_1r0d[12], o_1r1d[12]);
  OR2 I32 (complete247_0n[13], o_1r0d[13], o_1r1d[13]);
  OR2 I33 (complete247_0n[14], o_1r0d[14], o_1r1d[14]);
  OR2 I34 (complete247_0n[15], o_1r0d[15], o_1r1d[15]);
  OR2 I35 (complete247_0n[16], o_1r0d[16], o_1r1d[16]);
  OR2 I36 (complete247_0n[17], o_1r0d[17], o_1r1d[17]);
  OR2 I37 (complete247_0n[18], o_1r0d[18], o_1r1d[18]);
  OR2 I38 (complete247_0n[19], o_1r0d[19], o_1r1d[19]);
  OR2 I39 (complete247_0n[20], o_1r0d[20], o_1r1d[20]);
  OR2 I40 (complete247_0n[21], o_1r0d[21], o_1r1d[21]);
  OR2 I41 (complete247_0n[22], o_1r0d[22], o_1r1d[22]);
  OR2 I42 (complete247_0n[23], o_1r0d[23], o_1r1d[23]);
  OR2 I43 (complete247_0n[24], o_1r0d[24], o_1r1d[24]);
  OR2 I44 (complete247_0n[25], o_1r0d[25], o_1r1d[25]);
  OR2 I45 (complete247_0n[26], o_1r0d[26], o_1r1d[26]);
  OR2 I46 (complete247_0n[27], o_1r0d[27], o_1r1d[27]);
  OR2 I47 (complete247_0n[28], o_1r0d[28], o_1r1d[28]);
  OR2 I48 (complete247_0n[29], o_1r0d[29], o_1r1d[29]);
  OR2 I49 (complete247_0n[30], o_1r0d[30], o_1r1d[30]);
  OR2 I50 (complete247_0n[31], o_1r0d[31], o_1r1d[31]);
  OR2 I51 (complete247_0n[32], o_1r0d[32], o_1r1d[32]);
  OR2 I52 (complete247_0n[33], o_1r0d[33], o_1r1d[33]);
  INV I53 (gate246_0n, o_1a);
  C2RI I54 (o_1r1d[0], otint_1n[0], gate246_0n, initialise);
  C2RI I55 (o_1r1d[1], otint_1n[1], gate246_0n, initialise);
  C2RI I56 (o_1r1d[2], otint_1n[2], gate246_0n, initialise);
  C2RI I57 (o_1r1d[3], otint_1n[3], gate246_0n, initialise);
  C2RI I58 (o_1r1d[4], otint_1n[4], gate246_0n, initialise);
  C2RI I59 (o_1r1d[5], otint_1n[5], gate246_0n, initialise);
  C2RI I60 (o_1r1d[6], otint_1n[6], gate246_0n, initialise);
  C2RI I61 (o_1r1d[7], otint_1n[7], gate246_0n, initialise);
  C2RI I62 (o_1r1d[8], otint_1n[8], gate246_0n, initialise);
  C2RI I63 (o_1r1d[9], otint_1n[9], gate246_0n, initialise);
  C2RI I64 (o_1r1d[10], otint_1n[10], gate246_0n, initialise);
  C2RI I65 (o_1r1d[11], otint_1n[11], gate246_0n, initialise);
  C2RI I66 (o_1r1d[12], otint_1n[12], gate246_0n, initialise);
  C2RI I67 (o_1r1d[13], otint_1n[13], gate246_0n, initialise);
  C2RI I68 (o_1r1d[14], otint_1n[14], gate246_0n, initialise);
  C2RI I69 (o_1r1d[15], otint_1n[15], gate246_0n, initialise);
  C2RI I70 (o_1r1d[16], otint_1n[16], gate246_0n, initialise);
  C2RI I71 (o_1r1d[17], otint_1n[17], gate246_0n, initialise);
  C2RI I72 (o_1r1d[18], otint_1n[18], gate246_0n, initialise);
  C2RI I73 (o_1r1d[19], otint_1n[19], gate246_0n, initialise);
  C2RI I74 (o_1r1d[20], otint_1n[20], gate246_0n, initialise);
  C2RI I75 (o_1r1d[21], otint_1n[21], gate246_0n, initialise);
  C2RI I76 (o_1r1d[22], otint_1n[22], gate246_0n, initialise);
  C2RI I77 (o_1r1d[23], otint_1n[23], gate246_0n, initialise);
  C2RI I78 (o_1r1d[24], otint_1n[24], gate246_0n, initialise);
  C2RI I79 (o_1r1d[25], otint_1n[25], gate246_0n, initialise);
  C2RI I80 (o_1r1d[26], otint_1n[26], gate246_0n, initialise);
  C2RI I81 (o_1r1d[27], otint_1n[27], gate246_0n, initialise);
  C2RI I82 (o_1r1d[28], otint_1n[28], gate246_0n, initialise);
  C2RI I83 (o_1r1d[29], otint_1n[29], gate246_0n, initialise);
  C2RI I84 (o_1r1d[30], otint_1n[30], gate246_0n, initialise);
  C2RI I85 (o_1r1d[31], otint_1n[31], gate246_0n, initialise);
  C2RI I86 (o_1r1d[32], otint_1n[32], gate246_0n, initialise);
  C2RI I87 (o_1r1d[33], otint_1n[33], gate246_0n, initialise);
  C2RI I88 (o_1r0d[0], ofint_1n[0], gate246_0n, initialise);
  C2RI I89 (o_1r0d[1], ofint_1n[1], gate246_0n, initialise);
  C2RI I90 (o_1r0d[2], ofint_1n[2], gate246_0n, initialise);
  C2RI I91 (o_1r0d[3], ofint_1n[3], gate246_0n, initialise);
  C2RI I92 (o_1r0d[4], ofint_1n[4], gate246_0n, initialise);
  C2RI I93 (o_1r0d[5], ofint_1n[5], gate246_0n, initialise);
  C2RI I94 (o_1r0d[6], ofint_1n[6], gate246_0n, initialise);
  C2RI I95 (o_1r0d[7], ofint_1n[7], gate246_0n, initialise);
  C2RI I96 (o_1r0d[8], ofint_1n[8], gate246_0n, initialise);
  C2RI I97 (o_1r0d[9], ofint_1n[9], gate246_0n, initialise);
  C2RI I98 (o_1r0d[10], ofint_1n[10], gate246_0n, initialise);
  C2RI I99 (o_1r0d[11], ofint_1n[11], gate246_0n, initialise);
  C2RI I100 (o_1r0d[12], ofint_1n[12], gate246_0n, initialise);
  C2RI I101 (o_1r0d[13], ofint_1n[13], gate246_0n, initialise);
  C2RI I102 (o_1r0d[14], ofint_1n[14], gate246_0n, initialise);
  C2RI I103 (o_1r0d[15], ofint_1n[15], gate246_0n, initialise);
  C2RI I104 (o_1r0d[16], ofint_1n[16], gate246_0n, initialise);
  C2RI I105 (o_1r0d[17], ofint_1n[17], gate246_0n, initialise);
  C2RI I106 (o_1r0d[18], ofint_1n[18], gate246_0n, initialise);
  C2RI I107 (o_1r0d[19], ofint_1n[19], gate246_0n, initialise);
  C2RI I108 (o_1r0d[20], ofint_1n[20], gate246_0n, initialise);
  C2RI I109 (o_1r0d[21], ofint_1n[21], gate246_0n, initialise);
  C2RI I110 (o_1r0d[22], ofint_1n[22], gate246_0n, initialise);
  C2RI I111 (o_1r0d[23], ofint_1n[23], gate246_0n, initialise);
  C2RI I112 (o_1r0d[24], ofint_1n[24], gate246_0n, initialise);
  C2RI I113 (o_1r0d[25], ofint_1n[25], gate246_0n, initialise);
  C2RI I114 (o_1r0d[26], ofint_1n[26], gate246_0n, initialise);
  C2RI I115 (o_1r0d[27], ofint_1n[27], gate246_0n, initialise);
  C2RI I116 (o_1r0d[28], ofint_1n[28], gate246_0n, initialise);
  C2RI I117 (o_1r0d[29], ofint_1n[29], gate246_0n, initialise);
  C2RI I118 (o_1r0d[30], ofint_1n[30], gate246_0n, initialise);
  C2RI I119 (o_1r0d[31], ofint_1n[31], gate246_0n, initialise);
  C2RI I120 (o_1r0d[32], ofint_1n[32], gate246_0n, initialise);
  C2RI I121 (o_1r0d[33], ofint_1n[33], gate246_0n, initialise);
  assign oaint_0n = o_0r;
  INV I123 (gate243_0n, o_0a);
  C2RI I124 (o_0r, ofint_0n, gate243_0n, initialise);
  C3 I125 (internal_0n[18], complete240_0n[0], complete240_0n[1], complete240_0n[2]);
  C3 I126 (internal_0n[19], complete240_0n[3], complete240_0n[4], complete240_0n[5]);
  C3 I127 (internal_0n[20], complete240_0n[6], complete240_0n[7], complete240_0n[8]);
  C3 I128 (internal_0n[21], complete240_0n[9], complete240_0n[10], complete240_0n[11]);
  C3 I129 (internal_0n[22], complete240_0n[12], complete240_0n[13], complete240_0n[14]);
  C3 I130 (internal_0n[23], complete240_0n[15], complete240_0n[16], complete240_0n[17]);
  C3 I131 (internal_0n[24], complete240_0n[18], complete240_0n[19], complete240_0n[20]);
  C3 I132 (internal_0n[25], complete240_0n[21], complete240_0n[22], complete240_0n[23]);
  C3 I133 (internal_0n[26], complete240_0n[24], complete240_0n[25], complete240_0n[26]);
  C3 I134 (internal_0n[27], complete240_0n[27], complete240_0n[28], complete240_0n[29]);
  C2 I135 (internal_0n[28], complete240_0n[30], complete240_0n[31]);
  C2 I136 (internal_0n[29], complete240_0n[32], complete240_0n[33]);
  C3 I137 (internal_0n[30], internal_0n[18], internal_0n[19], internal_0n[20]);
  C3 I138 (internal_0n[31], internal_0n[21], internal_0n[22], internal_0n[23]);
  C3 I139 (internal_0n[32], internal_0n[24], internal_0n[25], internal_0n[26]);
  C3 I140 (internal_0n[33], internal_0n[27], internal_0n[28], internal_0n[29]);
  C2 I141 (internal_0n[34], internal_0n[30], internal_0n[31]);
  C2 I142 (internal_0n[35], internal_0n[32], internal_0n[33]);
  C2 I143 (i_0a, internal_0n[34], internal_0n[35]);
  OR2 I144 (complete240_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I145 (complete240_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I146 (complete240_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I147 (complete240_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I148 (complete240_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I149 (complete240_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I150 (complete240_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I151 (complete240_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I152 (complete240_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I153 (complete240_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I154 (complete240_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I155 (complete240_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I156 (complete240_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I157 (complete240_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I158 (complete240_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I159 (complete240_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I160 (complete240_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I161 (complete240_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I162 (complete240_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I163 (complete240_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I164 (complete240_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I165 (complete240_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I166 (complete240_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I167 (complete240_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I168 (complete240_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I169 (complete240_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I170 (complete240_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I171 (complete240_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I172 (complete240_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I173 (complete240_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I174 (complete240_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I175 (complete240_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I176 (complete240_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I177 (complete240_0n[33], ifint_0n[33], itint_0n[33]);
  INV I178 (gate239_0n, iaint_0n);
  C2RI I179 (itint_0n[0], i_0r1d[0], gate239_0n, initialise);
  C2RI I180 (itint_0n[1], i_0r1d[1], gate239_0n, initialise);
  C2RI I181 (itint_0n[2], i_0r1d[2], gate239_0n, initialise);
  C2RI I182 (itint_0n[3], i_0r1d[3], gate239_0n, initialise);
  C2RI I183 (itint_0n[4], i_0r1d[4], gate239_0n, initialise);
  C2RI I184 (itint_0n[5], i_0r1d[5], gate239_0n, initialise);
  C2RI I185 (itint_0n[6], i_0r1d[6], gate239_0n, initialise);
  C2RI I186 (itint_0n[7], i_0r1d[7], gate239_0n, initialise);
  C2RI I187 (itint_0n[8], i_0r1d[8], gate239_0n, initialise);
  C2RI I188 (itint_0n[9], i_0r1d[9], gate239_0n, initialise);
  C2RI I189 (itint_0n[10], i_0r1d[10], gate239_0n, initialise);
  C2RI I190 (itint_0n[11], i_0r1d[11], gate239_0n, initialise);
  C2RI I191 (itint_0n[12], i_0r1d[12], gate239_0n, initialise);
  C2RI I192 (itint_0n[13], i_0r1d[13], gate239_0n, initialise);
  C2RI I193 (itint_0n[14], i_0r1d[14], gate239_0n, initialise);
  C2RI I194 (itint_0n[15], i_0r1d[15], gate239_0n, initialise);
  C2RI I195 (itint_0n[16], i_0r1d[16], gate239_0n, initialise);
  C2RI I196 (itint_0n[17], i_0r1d[17], gate239_0n, initialise);
  C2RI I197 (itint_0n[18], i_0r1d[18], gate239_0n, initialise);
  C2RI I198 (itint_0n[19], i_0r1d[19], gate239_0n, initialise);
  C2RI I199 (itint_0n[20], i_0r1d[20], gate239_0n, initialise);
  C2RI I200 (itint_0n[21], i_0r1d[21], gate239_0n, initialise);
  C2RI I201 (itint_0n[22], i_0r1d[22], gate239_0n, initialise);
  C2RI I202 (itint_0n[23], i_0r1d[23], gate239_0n, initialise);
  C2RI I203 (itint_0n[24], i_0r1d[24], gate239_0n, initialise);
  C2RI I204 (itint_0n[25], i_0r1d[25], gate239_0n, initialise);
  C2RI I205 (itint_0n[26], i_0r1d[26], gate239_0n, initialise);
  C2RI I206 (itint_0n[27], i_0r1d[27], gate239_0n, initialise);
  C2RI I207 (itint_0n[28], i_0r1d[28], gate239_0n, initialise);
  C2RI I208 (itint_0n[29], i_0r1d[29], gate239_0n, initialise);
  C2RI I209 (itint_0n[30], i_0r1d[30], gate239_0n, initialise);
  C2RI I210 (itint_0n[31], i_0r1d[31], gate239_0n, initialise);
  C2RI I211 (itint_0n[32], i_0r1d[32], gate239_0n, initialise);
  C2RI I212 (itint_0n[33], i_0r1d[33], gate239_0n, initialise);
  C2RI I213 (ifint_0n[0], i_0r0d[0], gate239_0n, initialise);
  C2RI I214 (ifint_0n[1], i_0r0d[1], gate239_0n, initialise);
  C2RI I215 (ifint_0n[2], i_0r0d[2], gate239_0n, initialise);
  C2RI I216 (ifint_0n[3], i_0r0d[3], gate239_0n, initialise);
  C2RI I217 (ifint_0n[4], i_0r0d[4], gate239_0n, initialise);
  C2RI I218 (ifint_0n[5], i_0r0d[5], gate239_0n, initialise);
  C2RI I219 (ifint_0n[6], i_0r0d[6], gate239_0n, initialise);
  C2RI I220 (ifint_0n[7], i_0r0d[7], gate239_0n, initialise);
  C2RI I221 (ifint_0n[8], i_0r0d[8], gate239_0n, initialise);
  C2RI I222 (ifint_0n[9], i_0r0d[9], gate239_0n, initialise);
  C2RI I223 (ifint_0n[10], i_0r0d[10], gate239_0n, initialise);
  C2RI I224 (ifint_0n[11], i_0r0d[11], gate239_0n, initialise);
  C2RI I225 (ifint_0n[12], i_0r0d[12], gate239_0n, initialise);
  C2RI I226 (ifint_0n[13], i_0r0d[13], gate239_0n, initialise);
  C2RI I227 (ifint_0n[14], i_0r0d[14], gate239_0n, initialise);
  C2RI I228 (ifint_0n[15], i_0r0d[15], gate239_0n, initialise);
  C2RI I229 (ifint_0n[16], i_0r0d[16], gate239_0n, initialise);
  C2RI I230 (ifint_0n[17], i_0r0d[17], gate239_0n, initialise);
  C2RI I231 (ifint_0n[18], i_0r0d[18], gate239_0n, initialise);
  C2RI I232 (ifint_0n[19], i_0r0d[19], gate239_0n, initialise);
  C2RI I233 (ifint_0n[20], i_0r0d[20], gate239_0n, initialise);
  C2RI I234 (ifint_0n[21], i_0r0d[21], gate239_0n, initialise);
  C2RI I235 (ifint_0n[22], i_0r0d[22], gate239_0n, initialise);
  C2RI I236 (ifint_0n[23], i_0r0d[23], gate239_0n, initialise);
  C2RI I237 (ifint_0n[24], i_0r0d[24], gate239_0n, initialise);
  C2RI I238 (ifint_0n[25], i_0r0d[25], gate239_0n, initialise);
  C2RI I239 (ifint_0n[26], i_0r0d[26], gate239_0n, initialise);
  C2RI I240 (ifint_0n[27], i_0r0d[27], gate239_0n, initialise);
  C2RI I241 (ifint_0n[28], i_0r0d[28], gate239_0n, initialise);
  C2RI I242 (ifint_0n[29], i_0r0d[29], gate239_0n, initialise);
  C2RI I243 (ifint_0n[30], i_0r0d[30], gate239_0n, initialise);
  C2RI I244 (ifint_0n[31], i_0r0d[31], gate239_0n, initialise);
  C2RI I245 (ifint_0n[32], i_0r0d[32], gate239_0n, initialise);
  C2RI I246 (ifint_0n[33], i_0r0d[33], gate239_0n, initialise);
  C3 I247 (iaint_0n, icomplete_0n, oaint_0n, oaint_1n);
  assign ofint_0n = icomplete_0n;
  assign otint_1n[0] = itint_0n[0];
  assign otint_1n[1] = itint_0n[1];
  assign otint_1n[2] = itint_0n[2];
  assign otint_1n[3] = itint_0n[3];
  assign otint_1n[4] = itint_0n[4];
  assign otint_1n[5] = itint_0n[5];
  assign otint_1n[6] = itint_0n[6];
  assign otint_1n[7] = itint_0n[7];
  assign otint_1n[8] = itint_0n[8];
  assign otint_1n[9] = itint_0n[9];
  assign otint_1n[10] = itint_0n[10];
  assign otint_1n[11] = itint_0n[11];
  assign otint_1n[12] = itint_0n[12];
  assign otint_1n[13] = itint_0n[13];
  assign otint_1n[14] = itint_0n[14];
  assign otint_1n[15] = itint_0n[15];
  assign otint_1n[16] = itint_0n[16];
  assign otint_1n[17] = itint_0n[17];
  assign otint_1n[18] = itint_0n[18];
  assign otint_1n[19] = itint_0n[19];
  assign otint_1n[20] = itint_0n[20];
  assign otint_1n[21] = itint_0n[21];
  assign otint_1n[22] = itint_0n[22];
  assign otint_1n[23] = itint_0n[23];
  assign otint_1n[24] = itint_0n[24];
  assign otint_1n[25] = itint_0n[25];
  assign otint_1n[26] = itint_0n[26];
  assign otint_1n[27] = itint_0n[27];
  assign otint_1n[28] = itint_0n[28];
  assign otint_1n[29] = itint_0n[29];
  assign otint_1n[30] = itint_0n[30];
  assign otint_1n[31] = itint_0n[31];
  assign otint_1n[32] = itint_0n[32];
  assign otint_1n[33] = itint_0n[33];
  assign ofint_1n[0] = ifint_0n[0];
  assign ofint_1n[1] = ifint_0n[1];
  assign ofint_1n[2] = ifint_0n[2];
  assign ofint_1n[3] = ifint_0n[3];
  assign ofint_1n[4] = ifint_0n[4];
  assign ofint_1n[5] = ifint_0n[5];
  assign ofint_1n[6] = ifint_0n[6];
  assign ofint_1n[7] = ifint_0n[7];
  assign ofint_1n[8] = ifint_0n[8];
  assign ofint_1n[9] = ifint_0n[9];
  assign ofint_1n[10] = ifint_0n[10];
  assign ofint_1n[11] = ifint_0n[11];
  assign ofint_1n[12] = ifint_0n[12];
  assign ofint_1n[13] = ifint_0n[13];
  assign ofint_1n[14] = ifint_0n[14];
  assign ofint_1n[15] = ifint_0n[15];
  assign ofint_1n[16] = ifint_0n[16];
  assign ofint_1n[17] = ifint_0n[17];
  assign ofint_1n[18] = ifint_0n[18];
  assign ofint_1n[19] = ifint_0n[19];
  assign ofint_1n[20] = ifint_0n[20];
  assign ofint_1n[21] = ifint_0n[21];
  assign ofint_1n[22] = ifint_0n[22];
  assign ofint_1n[23] = ifint_0n[23];
  assign ofint_1n[24] = ifint_0n[24];
  assign ofint_1n[25] = ifint_0n[25];
  assign ofint_1n[26] = ifint_0n[26];
  assign ofint_1n[27] = ifint_0n[27];
  assign ofint_1n[28] = ifint_0n[28];
  assign ofint_1n[29] = ifint_0n[29];
  assign ofint_1n[30] = ifint_0n[30];
  assign ofint_1n[31] = ifint_0n[31];
  assign ofint_1n[32] = ifint_0n[32];
  assign ofint_1n[33] = ifint_0n[33];
  C3 I317 (internal_0n[36], complete236_0n[0], complete236_0n[1], complete236_0n[2]);
  C3 I318 (internal_0n[37], complete236_0n[3], complete236_0n[4], complete236_0n[5]);
  C3 I319 (internal_0n[38], complete236_0n[6], complete236_0n[7], complete236_0n[8]);
  C3 I320 (internal_0n[39], complete236_0n[9], complete236_0n[10], complete236_0n[11]);
  C3 I321 (internal_0n[40], complete236_0n[12], complete236_0n[13], complete236_0n[14]);
  C3 I322 (internal_0n[41], complete236_0n[15], complete236_0n[16], complete236_0n[17]);
  C3 I323 (internal_0n[42], complete236_0n[18], complete236_0n[19], complete236_0n[20]);
  C3 I324 (internal_0n[43], complete236_0n[21], complete236_0n[22], complete236_0n[23]);
  C3 I325 (internal_0n[44], complete236_0n[24], complete236_0n[25], complete236_0n[26]);
  C3 I326 (internal_0n[45], complete236_0n[27], complete236_0n[28], complete236_0n[29]);
  C2 I327 (internal_0n[46], complete236_0n[30], complete236_0n[31]);
  C2 I328 (internal_0n[47], complete236_0n[32], complete236_0n[33]);
  C3 I329 (internal_0n[48], internal_0n[36], internal_0n[37], internal_0n[38]);
  C3 I330 (internal_0n[49], internal_0n[39], internal_0n[40], internal_0n[41]);
  C3 I331 (internal_0n[50], internal_0n[42], internal_0n[43], internal_0n[44]);
  C3 I332 (internal_0n[51], internal_0n[45], internal_0n[46], internal_0n[47]);
  C2 I333 (internal_0n[52], internal_0n[48], internal_0n[49]);
  C2 I334 (internal_0n[53], internal_0n[50], internal_0n[51]);
  C2 I335 (icomplete_0n, internal_0n[52], internal_0n[53]);
  OR2 I336 (complete236_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I337 (complete236_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I338 (complete236_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I339 (complete236_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I340 (complete236_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I341 (complete236_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I342 (complete236_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I343 (complete236_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I344 (complete236_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I345 (complete236_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I346 (complete236_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I347 (complete236_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I348 (complete236_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I349 (complete236_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I350 (complete236_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I351 (complete236_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I352 (complete236_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I353 (complete236_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I354 (complete236_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I355 (complete236_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I356 (complete236_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I357 (complete236_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I358 (complete236_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I359 (complete236_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I360 (complete236_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I361 (complete236_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I362 (complete236_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I363 (complete236_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I364 (complete236_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I365 (complete236_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I366 (complete236_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I367 (complete236_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I368 (complete236_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I369 (complete236_0n[33], ifint_0n[33], itint_0n[33]);
endmodule

module BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m (
  i_0r0d, i_0r1d, i_0a,
  o_0r, o_0a,
  o_1r0d, o_1r1d, o_1a,
  initialise
);
  input [34:0] i_0r0d;
  input [34:0] i_0r1d;
  output i_0a;
  output o_0r;
  input o_0a;
  output [34:0] o_1r0d;
  output [34:0] o_1r1d;
  input o_1a;
  input initialise;
  wire [53:0] internal_0n;
  wire [34:0] ifint_0n;
  wire [34:0] itint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire [34:0] ofint_1n;
  wire [34:0] otint_1n;
  wire oaint_0n;
  wire oaint_1n;
  wire [34:0] complete259_0n;
  wire gate258_0n;
  wire gate255_0n;
  wire [34:0] complete252_0n;
  wire gate251_0n;
  wire [34:0] complete248_0n;
  wire icomplete_0n;
  C3 I0 (internal_0n[0], complete259_0n[0], complete259_0n[1], complete259_0n[2]);
  C3 I1 (internal_0n[1], complete259_0n[3], complete259_0n[4], complete259_0n[5]);
  C3 I2 (internal_0n[2], complete259_0n[6], complete259_0n[7], complete259_0n[8]);
  C3 I3 (internal_0n[3], complete259_0n[9], complete259_0n[10], complete259_0n[11]);
  C3 I4 (internal_0n[4], complete259_0n[12], complete259_0n[13], complete259_0n[14]);
  C3 I5 (internal_0n[5], complete259_0n[15], complete259_0n[16], complete259_0n[17]);
  C3 I6 (internal_0n[6], complete259_0n[18], complete259_0n[19], complete259_0n[20]);
  C3 I7 (internal_0n[7], complete259_0n[21], complete259_0n[22], complete259_0n[23]);
  C3 I8 (internal_0n[8], complete259_0n[24], complete259_0n[25], complete259_0n[26]);
  C3 I9 (internal_0n[9], complete259_0n[27], complete259_0n[28], complete259_0n[29]);
  C3 I10 (internal_0n[10], complete259_0n[30], complete259_0n[31], complete259_0n[32]);
  C2 I11 (internal_0n[11], complete259_0n[33], complete259_0n[34]);
  C3 I12 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I13 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I14 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I15 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I16 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I17 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I18 (oaint_1n, internal_0n[16], internal_0n[17]);
  OR2 I19 (complete259_0n[0], o_1r0d[0], o_1r1d[0]);
  OR2 I20 (complete259_0n[1], o_1r0d[1], o_1r1d[1]);
  OR2 I21 (complete259_0n[2], o_1r0d[2], o_1r1d[2]);
  OR2 I22 (complete259_0n[3], o_1r0d[3], o_1r1d[3]);
  OR2 I23 (complete259_0n[4], o_1r0d[4], o_1r1d[4]);
  OR2 I24 (complete259_0n[5], o_1r0d[5], o_1r1d[5]);
  OR2 I25 (complete259_0n[6], o_1r0d[6], o_1r1d[6]);
  OR2 I26 (complete259_0n[7], o_1r0d[7], o_1r1d[7]);
  OR2 I27 (complete259_0n[8], o_1r0d[8], o_1r1d[8]);
  OR2 I28 (complete259_0n[9], o_1r0d[9], o_1r1d[9]);
  OR2 I29 (complete259_0n[10], o_1r0d[10], o_1r1d[10]);
  OR2 I30 (complete259_0n[11], o_1r0d[11], o_1r1d[11]);
  OR2 I31 (complete259_0n[12], o_1r0d[12], o_1r1d[12]);
  OR2 I32 (complete259_0n[13], o_1r0d[13], o_1r1d[13]);
  OR2 I33 (complete259_0n[14], o_1r0d[14], o_1r1d[14]);
  OR2 I34 (complete259_0n[15], o_1r0d[15], o_1r1d[15]);
  OR2 I35 (complete259_0n[16], o_1r0d[16], o_1r1d[16]);
  OR2 I36 (complete259_0n[17], o_1r0d[17], o_1r1d[17]);
  OR2 I37 (complete259_0n[18], o_1r0d[18], o_1r1d[18]);
  OR2 I38 (complete259_0n[19], o_1r0d[19], o_1r1d[19]);
  OR2 I39 (complete259_0n[20], o_1r0d[20], o_1r1d[20]);
  OR2 I40 (complete259_0n[21], o_1r0d[21], o_1r1d[21]);
  OR2 I41 (complete259_0n[22], o_1r0d[22], o_1r1d[22]);
  OR2 I42 (complete259_0n[23], o_1r0d[23], o_1r1d[23]);
  OR2 I43 (complete259_0n[24], o_1r0d[24], o_1r1d[24]);
  OR2 I44 (complete259_0n[25], o_1r0d[25], o_1r1d[25]);
  OR2 I45 (complete259_0n[26], o_1r0d[26], o_1r1d[26]);
  OR2 I46 (complete259_0n[27], o_1r0d[27], o_1r1d[27]);
  OR2 I47 (complete259_0n[28], o_1r0d[28], o_1r1d[28]);
  OR2 I48 (complete259_0n[29], o_1r0d[29], o_1r1d[29]);
  OR2 I49 (complete259_0n[30], o_1r0d[30], o_1r1d[30]);
  OR2 I50 (complete259_0n[31], o_1r0d[31], o_1r1d[31]);
  OR2 I51 (complete259_0n[32], o_1r0d[32], o_1r1d[32]);
  OR2 I52 (complete259_0n[33], o_1r0d[33], o_1r1d[33]);
  OR2 I53 (complete259_0n[34], o_1r0d[34], o_1r1d[34]);
  INV I54 (gate258_0n, o_1a);
  C2RI I55 (o_1r1d[0], otint_1n[0], gate258_0n, initialise);
  C2RI I56 (o_1r1d[1], otint_1n[1], gate258_0n, initialise);
  C2RI I57 (o_1r1d[2], otint_1n[2], gate258_0n, initialise);
  C2RI I58 (o_1r1d[3], otint_1n[3], gate258_0n, initialise);
  C2RI I59 (o_1r1d[4], otint_1n[4], gate258_0n, initialise);
  C2RI I60 (o_1r1d[5], otint_1n[5], gate258_0n, initialise);
  C2RI I61 (o_1r1d[6], otint_1n[6], gate258_0n, initialise);
  C2RI I62 (o_1r1d[7], otint_1n[7], gate258_0n, initialise);
  C2RI I63 (o_1r1d[8], otint_1n[8], gate258_0n, initialise);
  C2RI I64 (o_1r1d[9], otint_1n[9], gate258_0n, initialise);
  C2RI I65 (o_1r1d[10], otint_1n[10], gate258_0n, initialise);
  C2RI I66 (o_1r1d[11], otint_1n[11], gate258_0n, initialise);
  C2RI I67 (o_1r1d[12], otint_1n[12], gate258_0n, initialise);
  C2RI I68 (o_1r1d[13], otint_1n[13], gate258_0n, initialise);
  C2RI I69 (o_1r1d[14], otint_1n[14], gate258_0n, initialise);
  C2RI I70 (o_1r1d[15], otint_1n[15], gate258_0n, initialise);
  C2RI I71 (o_1r1d[16], otint_1n[16], gate258_0n, initialise);
  C2RI I72 (o_1r1d[17], otint_1n[17], gate258_0n, initialise);
  C2RI I73 (o_1r1d[18], otint_1n[18], gate258_0n, initialise);
  C2RI I74 (o_1r1d[19], otint_1n[19], gate258_0n, initialise);
  C2RI I75 (o_1r1d[20], otint_1n[20], gate258_0n, initialise);
  C2RI I76 (o_1r1d[21], otint_1n[21], gate258_0n, initialise);
  C2RI I77 (o_1r1d[22], otint_1n[22], gate258_0n, initialise);
  C2RI I78 (o_1r1d[23], otint_1n[23], gate258_0n, initialise);
  C2RI I79 (o_1r1d[24], otint_1n[24], gate258_0n, initialise);
  C2RI I80 (o_1r1d[25], otint_1n[25], gate258_0n, initialise);
  C2RI I81 (o_1r1d[26], otint_1n[26], gate258_0n, initialise);
  C2RI I82 (o_1r1d[27], otint_1n[27], gate258_0n, initialise);
  C2RI I83 (o_1r1d[28], otint_1n[28], gate258_0n, initialise);
  C2RI I84 (o_1r1d[29], otint_1n[29], gate258_0n, initialise);
  C2RI I85 (o_1r1d[30], otint_1n[30], gate258_0n, initialise);
  C2RI I86 (o_1r1d[31], otint_1n[31], gate258_0n, initialise);
  C2RI I87 (o_1r1d[32], otint_1n[32], gate258_0n, initialise);
  C2RI I88 (o_1r1d[33], otint_1n[33], gate258_0n, initialise);
  C2RI I89 (o_1r1d[34], otint_1n[34], gate258_0n, initialise);
  C2RI I90 (o_1r0d[0], ofint_1n[0], gate258_0n, initialise);
  C2RI I91 (o_1r0d[1], ofint_1n[1], gate258_0n, initialise);
  C2RI I92 (o_1r0d[2], ofint_1n[2], gate258_0n, initialise);
  C2RI I93 (o_1r0d[3], ofint_1n[3], gate258_0n, initialise);
  C2RI I94 (o_1r0d[4], ofint_1n[4], gate258_0n, initialise);
  C2RI I95 (o_1r0d[5], ofint_1n[5], gate258_0n, initialise);
  C2RI I96 (o_1r0d[6], ofint_1n[6], gate258_0n, initialise);
  C2RI I97 (o_1r0d[7], ofint_1n[7], gate258_0n, initialise);
  C2RI I98 (o_1r0d[8], ofint_1n[8], gate258_0n, initialise);
  C2RI I99 (o_1r0d[9], ofint_1n[9], gate258_0n, initialise);
  C2RI I100 (o_1r0d[10], ofint_1n[10], gate258_0n, initialise);
  C2RI I101 (o_1r0d[11], ofint_1n[11], gate258_0n, initialise);
  C2RI I102 (o_1r0d[12], ofint_1n[12], gate258_0n, initialise);
  C2RI I103 (o_1r0d[13], ofint_1n[13], gate258_0n, initialise);
  C2RI I104 (o_1r0d[14], ofint_1n[14], gate258_0n, initialise);
  C2RI I105 (o_1r0d[15], ofint_1n[15], gate258_0n, initialise);
  C2RI I106 (o_1r0d[16], ofint_1n[16], gate258_0n, initialise);
  C2RI I107 (o_1r0d[17], ofint_1n[17], gate258_0n, initialise);
  C2RI I108 (o_1r0d[18], ofint_1n[18], gate258_0n, initialise);
  C2RI I109 (o_1r0d[19], ofint_1n[19], gate258_0n, initialise);
  C2RI I110 (o_1r0d[20], ofint_1n[20], gate258_0n, initialise);
  C2RI I111 (o_1r0d[21], ofint_1n[21], gate258_0n, initialise);
  C2RI I112 (o_1r0d[22], ofint_1n[22], gate258_0n, initialise);
  C2RI I113 (o_1r0d[23], ofint_1n[23], gate258_0n, initialise);
  C2RI I114 (o_1r0d[24], ofint_1n[24], gate258_0n, initialise);
  C2RI I115 (o_1r0d[25], ofint_1n[25], gate258_0n, initialise);
  C2RI I116 (o_1r0d[26], ofint_1n[26], gate258_0n, initialise);
  C2RI I117 (o_1r0d[27], ofint_1n[27], gate258_0n, initialise);
  C2RI I118 (o_1r0d[28], ofint_1n[28], gate258_0n, initialise);
  C2RI I119 (o_1r0d[29], ofint_1n[29], gate258_0n, initialise);
  C2RI I120 (o_1r0d[30], ofint_1n[30], gate258_0n, initialise);
  C2RI I121 (o_1r0d[31], ofint_1n[31], gate258_0n, initialise);
  C2RI I122 (o_1r0d[32], ofint_1n[32], gate258_0n, initialise);
  C2RI I123 (o_1r0d[33], ofint_1n[33], gate258_0n, initialise);
  C2RI I124 (o_1r0d[34], ofint_1n[34], gate258_0n, initialise);
  assign oaint_0n = o_0r;
  INV I126 (gate255_0n, o_0a);
  C2RI I127 (o_0r, ofint_0n, gate255_0n, initialise);
  C3 I128 (internal_0n[18], complete252_0n[0], complete252_0n[1], complete252_0n[2]);
  C3 I129 (internal_0n[19], complete252_0n[3], complete252_0n[4], complete252_0n[5]);
  C3 I130 (internal_0n[20], complete252_0n[6], complete252_0n[7], complete252_0n[8]);
  C3 I131 (internal_0n[21], complete252_0n[9], complete252_0n[10], complete252_0n[11]);
  C3 I132 (internal_0n[22], complete252_0n[12], complete252_0n[13], complete252_0n[14]);
  C3 I133 (internal_0n[23], complete252_0n[15], complete252_0n[16], complete252_0n[17]);
  C3 I134 (internal_0n[24], complete252_0n[18], complete252_0n[19], complete252_0n[20]);
  C3 I135 (internal_0n[25], complete252_0n[21], complete252_0n[22], complete252_0n[23]);
  C3 I136 (internal_0n[26], complete252_0n[24], complete252_0n[25], complete252_0n[26]);
  C3 I137 (internal_0n[27], complete252_0n[27], complete252_0n[28], complete252_0n[29]);
  C3 I138 (internal_0n[28], complete252_0n[30], complete252_0n[31], complete252_0n[32]);
  C2 I139 (internal_0n[29], complete252_0n[33], complete252_0n[34]);
  C3 I140 (internal_0n[30], internal_0n[18], internal_0n[19], internal_0n[20]);
  C3 I141 (internal_0n[31], internal_0n[21], internal_0n[22], internal_0n[23]);
  C3 I142 (internal_0n[32], internal_0n[24], internal_0n[25], internal_0n[26]);
  C3 I143 (internal_0n[33], internal_0n[27], internal_0n[28], internal_0n[29]);
  C2 I144 (internal_0n[34], internal_0n[30], internal_0n[31]);
  C2 I145 (internal_0n[35], internal_0n[32], internal_0n[33]);
  C2 I146 (i_0a, internal_0n[34], internal_0n[35]);
  OR2 I147 (complete252_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I148 (complete252_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I149 (complete252_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I150 (complete252_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I151 (complete252_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I152 (complete252_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I153 (complete252_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I154 (complete252_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I155 (complete252_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I156 (complete252_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I157 (complete252_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I158 (complete252_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I159 (complete252_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I160 (complete252_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I161 (complete252_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I162 (complete252_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I163 (complete252_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I164 (complete252_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I165 (complete252_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I166 (complete252_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I167 (complete252_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I168 (complete252_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I169 (complete252_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I170 (complete252_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I171 (complete252_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I172 (complete252_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I173 (complete252_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I174 (complete252_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I175 (complete252_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I176 (complete252_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I177 (complete252_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I178 (complete252_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I179 (complete252_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I180 (complete252_0n[33], ifint_0n[33], itint_0n[33]);
  OR2 I181 (complete252_0n[34], ifint_0n[34], itint_0n[34]);
  INV I182 (gate251_0n, iaint_0n);
  C2RI I183 (itint_0n[0], i_0r1d[0], gate251_0n, initialise);
  C2RI I184 (itint_0n[1], i_0r1d[1], gate251_0n, initialise);
  C2RI I185 (itint_0n[2], i_0r1d[2], gate251_0n, initialise);
  C2RI I186 (itint_0n[3], i_0r1d[3], gate251_0n, initialise);
  C2RI I187 (itint_0n[4], i_0r1d[4], gate251_0n, initialise);
  C2RI I188 (itint_0n[5], i_0r1d[5], gate251_0n, initialise);
  C2RI I189 (itint_0n[6], i_0r1d[6], gate251_0n, initialise);
  C2RI I190 (itint_0n[7], i_0r1d[7], gate251_0n, initialise);
  C2RI I191 (itint_0n[8], i_0r1d[8], gate251_0n, initialise);
  C2RI I192 (itint_0n[9], i_0r1d[9], gate251_0n, initialise);
  C2RI I193 (itint_0n[10], i_0r1d[10], gate251_0n, initialise);
  C2RI I194 (itint_0n[11], i_0r1d[11], gate251_0n, initialise);
  C2RI I195 (itint_0n[12], i_0r1d[12], gate251_0n, initialise);
  C2RI I196 (itint_0n[13], i_0r1d[13], gate251_0n, initialise);
  C2RI I197 (itint_0n[14], i_0r1d[14], gate251_0n, initialise);
  C2RI I198 (itint_0n[15], i_0r1d[15], gate251_0n, initialise);
  C2RI I199 (itint_0n[16], i_0r1d[16], gate251_0n, initialise);
  C2RI I200 (itint_0n[17], i_0r1d[17], gate251_0n, initialise);
  C2RI I201 (itint_0n[18], i_0r1d[18], gate251_0n, initialise);
  C2RI I202 (itint_0n[19], i_0r1d[19], gate251_0n, initialise);
  C2RI I203 (itint_0n[20], i_0r1d[20], gate251_0n, initialise);
  C2RI I204 (itint_0n[21], i_0r1d[21], gate251_0n, initialise);
  C2RI I205 (itint_0n[22], i_0r1d[22], gate251_0n, initialise);
  C2RI I206 (itint_0n[23], i_0r1d[23], gate251_0n, initialise);
  C2RI I207 (itint_0n[24], i_0r1d[24], gate251_0n, initialise);
  C2RI I208 (itint_0n[25], i_0r1d[25], gate251_0n, initialise);
  C2RI I209 (itint_0n[26], i_0r1d[26], gate251_0n, initialise);
  C2RI I210 (itint_0n[27], i_0r1d[27], gate251_0n, initialise);
  C2RI I211 (itint_0n[28], i_0r1d[28], gate251_0n, initialise);
  C2RI I212 (itint_0n[29], i_0r1d[29], gate251_0n, initialise);
  C2RI I213 (itint_0n[30], i_0r1d[30], gate251_0n, initialise);
  C2RI I214 (itint_0n[31], i_0r1d[31], gate251_0n, initialise);
  C2RI I215 (itint_0n[32], i_0r1d[32], gate251_0n, initialise);
  C2RI I216 (itint_0n[33], i_0r1d[33], gate251_0n, initialise);
  C2RI I217 (itint_0n[34], i_0r1d[34], gate251_0n, initialise);
  C2RI I218 (ifint_0n[0], i_0r0d[0], gate251_0n, initialise);
  C2RI I219 (ifint_0n[1], i_0r0d[1], gate251_0n, initialise);
  C2RI I220 (ifint_0n[2], i_0r0d[2], gate251_0n, initialise);
  C2RI I221 (ifint_0n[3], i_0r0d[3], gate251_0n, initialise);
  C2RI I222 (ifint_0n[4], i_0r0d[4], gate251_0n, initialise);
  C2RI I223 (ifint_0n[5], i_0r0d[5], gate251_0n, initialise);
  C2RI I224 (ifint_0n[6], i_0r0d[6], gate251_0n, initialise);
  C2RI I225 (ifint_0n[7], i_0r0d[7], gate251_0n, initialise);
  C2RI I226 (ifint_0n[8], i_0r0d[8], gate251_0n, initialise);
  C2RI I227 (ifint_0n[9], i_0r0d[9], gate251_0n, initialise);
  C2RI I228 (ifint_0n[10], i_0r0d[10], gate251_0n, initialise);
  C2RI I229 (ifint_0n[11], i_0r0d[11], gate251_0n, initialise);
  C2RI I230 (ifint_0n[12], i_0r0d[12], gate251_0n, initialise);
  C2RI I231 (ifint_0n[13], i_0r0d[13], gate251_0n, initialise);
  C2RI I232 (ifint_0n[14], i_0r0d[14], gate251_0n, initialise);
  C2RI I233 (ifint_0n[15], i_0r0d[15], gate251_0n, initialise);
  C2RI I234 (ifint_0n[16], i_0r0d[16], gate251_0n, initialise);
  C2RI I235 (ifint_0n[17], i_0r0d[17], gate251_0n, initialise);
  C2RI I236 (ifint_0n[18], i_0r0d[18], gate251_0n, initialise);
  C2RI I237 (ifint_0n[19], i_0r0d[19], gate251_0n, initialise);
  C2RI I238 (ifint_0n[20], i_0r0d[20], gate251_0n, initialise);
  C2RI I239 (ifint_0n[21], i_0r0d[21], gate251_0n, initialise);
  C2RI I240 (ifint_0n[22], i_0r0d[22], gate251_0n, initialise);
  C2RI I241 (ifint_0n[23], i_0r0d[23], gate251_0n, initialise);
  C2RI I242 (ifint_0n[24], i_0r0d[24], gate251_0n, initialise);
  C2RI I243 (ifint_0n[25], i_0r0d[25], gate251_0n, initialise);
  C2RI I244 (ifint_0n[26], i_0r0d[26], gate251_0n, initialise);
  C2RI I245 (ifint_0n[27], i_0r0d[27], gate251_0n, initialise);
  C2RI I246 (ifint_0n[28], i_0r0d[28], gate251_0n, initialise);
  C2RI I247 (ifint_0n[29], i_0r0d[29], gate251_0n, initialise);
  C2RI I248 (ifint_0n[30], i_0r0d[30], gate251_0n, initialise);
  C2RI I249 (ifint_0n[31], i_0r0d[31], gate251_0n, initialise);
  C2RI I250 (ifint_0n[32], i_0r0d[32], gate251_0n, initialise);
  C2RI I251 (ifint_0n[33], i_0r0d[33], gate251_0n, initialise);
  C2RI I252 (ifint_0n[34], i_0r0d[34], gate251_0n, initialise);
  C3 I253 (iaint_0n, icomplete_0n, oaint_0n, oaint_1n);
  assign ofint_0n = icomplete_0n;
  assign otint_1n[0] = itint_0n[0];
  assign otint_1n[1] = itint_0n[1];
  assign otint_1n[2] = itint_0n[2];
  assign otint_1n[3] = itint_0n[3];
  assign otint_1n[4] = itint_0n[4];
  assign otint_1n[5] = itint_0n[5];
  assign otint_1n[6] = itint_0n[6];
  assign otint_1n[7] = itint_0n[7];
  assign otint_1n[8] = itint_0n[8];
  assign otint_1n[9] = itint_0n[9];
  assign otint_1n[10] = itint_0n[10];
  assign otint_1n[11] = itint_0n[11];
  assign otint_1n[12] = itint_0n[12];
  assign otint_1n[13] = itint_0n[13];
  assign otint_1n[14] = itint_0n[14];
  assign otint_1n[15] = itint_0n[15];
  assign otint_1n[16] = itint_0n[16];
  assign otint_1n[17] = itint_0n[17];
  assign otint_1n[18] = itint_0n[18];
  assign otint_1n[19] = itint_0n[19];
  assign otint_1n[20] = itint_0n[20];
  assign otint_1n[21] = itint_0n[21];
  assign otint_1n[22] = itint_0n[22];
  assign otint_1n[23] = itint_0n[23];
  assign otint_1n[24] = itint_0n[24];
  assign otint_1n[25] = itint_0n[25];
  assign otint_1n[26] = itint_0n[26];
  assign otint_1n[27] = itint_0n[27];
  assign otint_1n[28] = itint_0n[28];
  assign otint_1n[29] = itint_0n[29];
  assign otint_1n[30] = itint_0n[30];
  assign otint_1n[31] = itint_0n[31];
  assign otint_1n[32] = itint_0n[32];
  assign otint_1n[33] = itint_0n[33];
  assign otint_1n[34] = itint_0n[34];
  assign ofint_1n[0] = ifint_0n[0];
  assign ofint_1n[1] = ifint_0n[1];
  assign ofint_1n[2] = ifint_0n[2];
  assign ofint_1n[3] = ifint_0n[3];
  assign ofint_1n[4] = ifint_0n[4];
  assign ofint_1n[5] = ifint_0n[5];
  assign ofint_1n[6] = ifint_0n[6];
  assign ofint_1n[7] = ifint_0n[7];
  assign ofint_1n[8] = ifint_0n[8];
  assign ofint_1n[9] = ifint_0n[9];
  assign ofint_1n[10] = ifint_0n[10];
  assign ofint_1n[11] = ifint_0n[11];
  assign ofint_1n[12] = ifint_0n[12];
  assign ofint_1n[13] = ifint_0n[13];
  assign ofint_1n[14] = ifint_0n[14];
  assign ofint_1n[15] = ifint_0n[15];
  assign ofint_1n[16] = ifint_0n[16];
  assign ofint_1n[17] = ifint_0n[17];
  assign ofint_1n[18] = ifint_0n[18];
  assign ofint_1n[19] = ifint_0n[19];
  assign ofint_1n[20] = ifint_0n[20];
  assign ofint_1n[21] = ifint_0n[21];
  assign ofint_1n[22] = ifint_0n[22];
  assign ofint_1n[23] = ifint_0n[23];
  assign ofint_1n[24] = ifint_0n[24];
  assign ofint_1n[25] = ifint_0n[25];
  assign ofint_1n[26] = ifint_0n[26];
  assign ofint_1n[27] = ifint_0n[27];
  assign ofint_1n[28] = ifint_0n[28];
  assign ofint_1n[29] = ifint_0n[29];
  assign ofint_1n[30] = ifint_0n[30];
  assign ofint_1n[31] = ifint_0n[31];
  assign ofint_1n[32] = ifint_0n[32];
  assign ofint_1n[33] = ifint_0n[33];
  assign ofint_1n[34] = ifint_0n[34];
  C3 I325 (internal_0n[36], complete248_0n[0], complete248_0n[1], complete248_0n[2]);
  C3 I326 (internal_0n[37], complete248_0n[3], complete248_0n[4], complete248_0n[5]);
  C3 I327 (internal_0n[38], complete248_0n[6], complete248_0n[7], complete248_0n[8]);
  C3 I328 (internal_0n[39], complete248_0n[9], complete248_0n[10], complete248_0n[11]);
  C3 I329 (internal_0n[40], complete248_0n[12], complete248_0n[13], complete248_0n[14]);
  C3 I330 (internal_0n[41], complete248_0n[15], complete248_0n[16], complete248_0n[17]);
  C3 I331 (internal_0n[42], complete248_0n[18], complete248_0n[19], complete248_0n[20]);
  C3 I332 (internal_0n[43], complete248_0n[21], complete248_0n[22], complete248_0n[23]);
  C3 I333 (internal_0n[44], complete248_0n[24], complete248_0n[25], complete248_0n[26]);
  C3 I334 (internal_0n[45], complete248_0n[27], complete248_0n[28], complete248_0n[29]);
  C3 I335 (internal_0n[46], complete248_0n[30], complete248_0n[31], complete248_0n[32]);
  C2 I336 (internal_0n[47], complete248_0n[33], complete248_0n[34]);
  C3 I337 (internal_0n[48], internal_0n[36], internal_0n[37], internal_0n[38]);
  C3 I338 (internal_0n[49], internal_0n[39], internal_0n[40], internal_0n[41]);
  C3 I339 (internal_0n[50], internal_0n[42], internal_0n[43], internal_0n[44]);
  C3 I340 (internal_0n[51], internal_0n[45], internal_0n[46], internal_0n[47]);
  C2 I341 (internal_0n[52], internal_0n[48], internal_0n[49]);
  C2 I342 (internal_0n[53], internal_0n[50], internal_0n[51]);
  C2 I343 (icomplete_0n, internal_0n[52], internal_0n[53]);
  OR2 I344 (complete248_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I345 (complete248_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I346 (complete248_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I347 (complete248_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I348 (complete248_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I349 (complete248_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I350 (complete248_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I351 (complete248_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I352 (complete248_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I353 (complete248_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I354 (complete248_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I355 (complete248_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I356 (complete248_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I357 (complete248_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I358 (complete248_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I359 (complete248_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I360 (complete248_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I361 (complete248_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I362 (complete248_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I363 (complete248_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I364 (complete248_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I365 (complete248_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I366 (complete248_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I367 (complete248_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I368 (complete248_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I369 (complete248_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I370 (complete248_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I371 (complete248_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I372 (complete248_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I373 (complete248_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I374 (complete248_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I375 (complete248_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I376 (complete248_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I377 (complete248_0n[33], ifint_0n[33], itint_0n[33]);
  OR2 I378 (complete248_0n[34], ifint_0n[34], itint_0n[34]);
endmodule

module BrzF_36_l32__28_280_200_29_20_280_2036_29__m44m (
  i_0r0d, i_0r1d, i_0a,
  o_0r, o_0a,
  o_1r0d, o_1r1d, o_1a,
  initialise
);
  input [35:0] i_0r0d;
  input [35:0] i_0r1d;
  output i_0a;
  output o_0r;
  input o_0a;
  output [35:0] o_1r0d;
  output [35:0] o_1r1d;
  input o_1a;
  input initialise;
  wire [53:0] internal_0n;
  wire [35:0] ifint_0n;
  wire [35:0] itint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire [35:0] ofint_1n;
  wire [35:0] otint_1n;
  wire oaint_0n;
  wire oaint_1n;
  wire [35:0] complete271_0n;
  wire gate270_0n;
  wire gate267_0n;
  wire [35:0] complete264_0n;
  wire gate263_0n;
  wire [35:0] complete260_0n;
  wire icomplete_0n;
  C3 I0 (internal_0n[0], complete271_0n[0], complete271_0n[1], complete271_0n[2]);
  C3 I1 (internal_0n[1], complete271_0n[3], complete271_0n[4], complete271_0n[5]);
  C3 I2 (internal_0n[2], complete271_0n[6], complete271_0n[7], complete271_0n[8]);
  C3 I3 (internal_0n[3], complete271_0n[9], complete271_0n[10], complete271_0n[11]);
  C3 I4 (internal_0n[4], complete271_0n[12], complete271_0n[13], complete271_0n[14]);
  C3 I5 (internal_0n[5], complete271_0n[15], complete271_0n[16], complete271_0n[17]);
  C3 I6 (internal_0n[6], complete271_0n[18], complete271_0n[19], complete271_0n[20]);
  C3 I7 (internal_0n[7], complete271_0n[21], complete271_0n[22], complete271_0n[23]);
  C3 I8 (internal_0n[8], complete271_0n[24], complete271_0n[25], complete271_0n[26]);
  C3 I9 (internal_0n[9], complete271_0n[27], complete271_0n[28], complete271_0n[29]);
  C3 I10 (internal_0n[10], complete271_0n[30], complete271_0n[31], complete271_0n[32]);
  C3 I11 (internal_0n[11], complete271_0n[33], complete271_0n[34], complete271_0n[35]);
  C3 I12 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I13 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I14 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I15 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I16 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I17 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I18 (oaint_1n, internal_0n[16], internal_0n[17]);
  OR2 I19 (complete271_0n[0], o_1r0d[0], o_1r1d[0]);
  OR2 I20 (complete271_0n[1], o_1r0d[1], o_1r1d[1]);
  OR2 I21 (complete271_0n[2], o_1r0d[2], o_1r1d[2]);
  OR2 I22 (complete271_0n[3], o_1r0d[3], o_1r1d[3]);
  OR2 I23 (complete271_0n[4], o_1r0d[4], o_1r1d[4]);
  OR2 I24 (complete271_0n[5], o_1r0d[5], o_1r1d[5]);
  OR2 I25 (complete271_0n[6], o_1r0d[6], o_1r1d[6]);
  OR2 I26 (complete271_0n[7], o_1r0d[7], o_1r1d[7]);
  OR2 I27 (complete271_0n[8], o_1r0d[8], o_1r1d[8]);
  OR2 I28 (complete271_0n[9], o_1r0d[9], o_1r1d[9]);
  OR2 I29 (complete271_0n[10], o_1r0d[10], o_1r1d[10]);
  OR2 I30 (complete271_0n[11], o_1r0d[11], o_1r1d[11]);
  OR2 I31 (complete271_0n[12], o_1r0d[12], o_1r1d[12]);
  OR2 I32 (complete271_0n[13], o_1r0d[13], o_1r1d[13]);
  OR2 I33 (complete271_0n[14], o_1r0d[14], o_1r1d[14]);
  OR2 I34 (complete271_0n[15], o_1r0d[15], o_1r1d[15]);
  OR2 I35 (complete271_0n[16], o_1r0d[16], o_1r1d[16]);
  OR2 I36 (complete271_0n[17], o_1r0d[17], o_1r1d[17]);
  OR2 I37 (complete271_0n[18], o_1r0d[18], o_1r1d[18]);
  OR2 I38 (complete271_0n[19], o_1r0d[19], o_1r1d[19]);
  OR2 I39 (complete271_0n[20], o_1r0d[20], o_1r1d[20]);
  OR2 I40 (complete271_0n[21], o_1r0d[21], o_1r1d[21]);
  OR2 I41 (complete271_0n[22], o_1r0d[22], o_1r1d[22]);
  OR2 I42 (complete271_0n[23], o_1r0d[23], o_1r1d[23]);
  OR2 I43 (complete271_0n[24], o_1r0d[24], o_1r1d[24]);
  OR2 I44 (complete271_0n[25], o_1r0d[25], o_1r1d[25]);
  OR2 I45 (complete271_0n[26], o_1r0d[26], o_1r1d[26]);
  OR2 I46 (complete271_0n[27], o_1r0d[27], o_1r1d[27]);
  OR2 I47 (complete271_0n[28], o_1r0d[28], o_1r1d[28]);
  OR2 I48 (complete271_0n[29], o_1r0d[29], o_1r1d[29]);
  OR2 I49 (complete271_0n[30], o_1r0d[30], o_1r1d[30]);
  OR2 I50 (complete271_0n[31], o_1r0d[31], o_1r1d[31]);
  OR2 I51 (complete271_0n[32], o_1r0d[32], o_1r1d[32]);
  OR2 I52 (complete271_0n[33], o_1r0d[33], o_1r1d[33]);
  OR2 I53 (complete271_0n[34], o_1r0d[34], o_1r1d[34]);
  OR2 I54 (complete271_0n[35], o_1r0d[35], o_1r1d[35]);
  INV I55 (gate270_0n, o_1a);
  C2RI I56 (o_1r1d[0], otint_1n[0], gate270_0n, initialise);
  C2RI I57 (o_1r1d[1], otint_1n[1], gate270_0n, initialise);
  C2RI I58 (o_1r1d[2], otint_1n[2], gate270_0n, initialise);
  C2RI I59 (o_1r1d[3], otint_1n[3], gate270_0n, initialise);
  C2RI I60 (o_1r1d[4], otint_1n[4], gate270_0n, initialise);
  C2RI I61 (o_1r1d[5], otint_1n[5], gate270_0n, initialise);
  C2RI I62 (o_1r1d[6], otint_1n[6], gate270_0n, initialise);
  C2RI I63 (o_1r1d[7], otint_1n[7], gate270_0n, initialise);
  C2RI I64 (o_1r1d[8], otint_1n[8], gate270_0n, initialise);
  C2RI I65 (o_1r1d[9], otint_1n[9], gate270_0n, initialise);
  C2RI I66 (o_1r1d[10], otint_1n[10], gate270_0n, initialise);
  C2RI I67 (o_1r1d[11], otint_1n[11], gate270_0n, initialise);
  C2RI I68 (o_1r1d[12], otint_1n[12], gate270_0n, initialise);
  C2RI I69 (o_1r1d[13], otint_1n[13], gate270_0n, initialise);
  C2RI I70 (o_1r1d[14], otint_1n[14], gate270_0n, initialise);
  C2RI I71 (o_1r1d[15], otint_1n[15], gate270_0n, initialise);
  C2RI I72 (o_1r1d[16], otint_1n[16], gate270_0n, initialise);
  C2RI I73 (o_1r1d[17], otint_1n[17], gate270_0n, initialise);
  C2RI I74 (o_1r1d[18], otint_1n[18], gate270_0n, initialise);
  C2RI I75 (o_1r1d[19], otint_1n[19], gate270_0n, initialise);
  C2RI I76 (o_1r1d[20], otint_1n[20], gate270_0n, initialise);
  C2RI I77 (o_1r1d[21], otint_1n[21], gate270_0n, initialise);
  C2RI I78 (o_1r1d[22], otint_1n[22], gate270_0n, initialise);
  C2RI I79 (o_1r1d[23], otint_1n[23], gate270_0n, initialise);
  C2RI I80 (o_1r1d[24], otint_1n[24], gate270_0n, initialise);
  C2RI I81 (o_1r1d[25], otint_1n[25], gate270_0n, initialise);
  C2RI I82 (o_1r1d[26], otint_1n[26], gate270_0n, initialise);
  C2RI I83 (o_1r1d[27], otint_1n[27], gate270_0n, initialise);
  C2RI I84 (o_1r1d[28], otint_1n[28], gate270_0n, initialise);
  C2RI I85 (o_1r1d[29], otint_1n[29], gate270_0n, initialise);
  C2RI I86 (o_1r1d[30], otint_1n[30], gate270_0n, initialise);
  C2RI I87 (o_1r1d[31], otint_1n[31], gate270_0n, initialise);
  C2RI I88 (o_1r1d[32], otint_1n[32], gate270_0n, initialise);
  C2RI I89 (o_1r1d[33], otint_1n[33], gate270_0n, initialise);
  C2RI I90 (o_1r1d[34], otint_1n[34], gate270_0n, initialise);
  C2RI I91 (o_1r1d[35], otint_1n[35], gate270_0n, initialise);
  C2RI I92 (o_1r0d[0], ofint_1n[0], gate270_0n, initialise);
  C2RI I93 (o_1r0d[1], ofint_1n[1], gate270_0n, initialise);
  C2RI I94 (o_1r0d[2], ofint_1n[2], gate270_0n, initialise);
  C2RI I95 (o_1r0d[3], ofint_1n[3], gate270_0n, initialise);
  C2RI I96 (o_1r0d[4], ofint_1n[4], gate270_0n, initialise);
  C2RI I97 (o_1r0d[5], ofint_1n[5], gate270_0n, initialise);
  C2RI I98 (o_1r0d[6], ofint_1n[6], gate270_0n, initialise);
  C2RI I99 (o_1r0d[7], ofint_1n[7], gate270_0n, initialise);
  C2RI I100 (o_1r0d[8], ofint_1n[8], gate270_0n, initialise);
  C2RI I101 (o_1r0d[9], ofint_1n[9], gate270_0n, initialise);
  C2RI I102 (o_1r0d[10], ofint_1n[10], gate270_0n, initialise);
  C2RI I103 (o_1r0d[11], ofint_1n[11], gate270_0n, initialise);
  C2RI I104 (o_1r0d[12], ofint_1n[12], gate270_0n, initialise);
  C2RI I105 (o_1r0d[13], ofint_1n[13], gate270_0n, initialise);
  C2RI I106 (o_1r0d[14], ofint_1n[14], gate270_0n, initialise);
  C2RI I107 (o_1r0d[15], ofint_1n[15], gate270_0n, initialise);
  C2RI I108 (o_1r0d[16], ofint_1n[16], gate270_0n, initialise);
  C2RI I109 (o_1r0d[17], ofint_1n[17], gate270_0n, initialise);
  C2RI I110 (o_1r0d[18], ofint_1n[18], gate270_0n, initialise);
  C2RI I111 (o_1r0d[19], ofint_1n[19], gate270_0n, initialise);
  C2RI I112 (o_1r0d[20], ofint_1n[20], gate270_0n, initialise);
  C2RI I113 (o_1r0d[21], ofint_1n[21], gate270_0n, initialise);
  C2RI I114 (o_1r0d[22], ofint_1n[22], gate270_0n, initialise);
  C2RI I115 (o_1r0d[23], ofint_1n[23], gate270_0n, initialise);
  C2RI I116 (o_1r0d[24], ofint_1n[24], gate270_0n, initialise);
  C2RI I117 (o_1r0d[25], ofint_1n[25], gate270_0n, initialise);
  C2RI I118 (o_1r0d[26], ofint_1n[26], gate270_0n, initialise);
  C2RI I119 (o_1r0d[27], ofint_1n[27], gate270_0n, initialise);
  C2RI I120 (o_1r0d[28], ofint_1n[28], gate270_0n, initialise);
  C2RI I121 (o_1r0d[29], ofint_1n[29], gate270_0n, initialise);
  C2RI I122 (o_1r0d[30], ofint_1n[30], gate270_0n, initialise);
  C2RI I123 (o_1r0d[31], ofint_1n[31], gate270_0n, initialise);
  C2RI I124 (o_1r0d[32], ofint_1n[32], gate270_0n, initialise);
  C2RI I125 (o_1r0d[33], ofint_1n[33], gate270_0n, initialise);
  C2RI I126 (o_1r0d[34], ofint_1n[34], gate270_0n, initialise);
  C2RI I127 (o_1r0d[35], ofint_1n[35], gate270_0n, initialise);
  assign oaint_0n = o_0r;
  INV I129 (gate267_0n, o_0a);
  C2RI I130 (o_0r, ofint_0n, gate267_0n, initialise);
  C3 I131 (internal_0n[18], complete264_0n[0], complete264_0n[1], complete264_0n[2]);
  C3 I132 (internal_0n[19], complete264_0n[3], complete264_0n[4], complete264_0n[5]);
  C3 I133 (internal_0n[20], complete264_0n[6], complete264_0n[7], complete264_0n[8]);
  C3 I134 (internal_0n[21], complete264_0n[9], complete264_0n[10], complete264_0n[11]);
  C3 I135 (internal_0n[22], complete264_0n[12], complete264_0n[13], complete264_0n[14]);
  C3 I136 (internal_0n[23], complete264_0n[15], complete264_0n[16], complete264_0n[17]);
  C3 I137 (internal_0n[24], complete264_0n[18], complete264_0n[19], complete264_0n[20]);
  C3 I138 (internal_0n[25], complete264_0n[21], complete264_0n[22], complete264_0n[23]);
  C3 I139 (internal_0n[26], complete264_0n[24], complete264_0n[25], complete264_0n[26]);
  C3 I140 (internal_0n[27], complete264_0n[27], complete264_0n[28], complete264_0n[29]);
  C3 I141 (internal_0n[28], complete264_0n[30], complete264_0n[31], complete264_0n[32]);
  C3 I142 (internal_0n[29], complete264_0n[33], complete264_0n[34], complete264_0n[35]);
  C3 I143 (internal_0n[30], internal_0n[18], internal_0n[19], internal_0n[20]);
  C3 I144 (internal_0n[31], internal_0n[21], internal_0n[22], internal_0n[23]);
  C3 I145 (internal_0n[32], internal_0n[24], internal_0n[25], internal_0n[26]);
  C3 I146 (internal_0n[33], internal_0n[27], internal_0n[28], internal_0n[29]);
  C2 I147 (internal_0n[34], internal_0n[30], internal_0n[31]);
  C2 I148 (internal_0n[35], internal_0n[32], internal_0n[33]);
  C2 I149 (i_0a, internal_0n[34], internal_0n[35]);
  OR2 I150 (complete264_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I151 (complete264_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I152 (complete264_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I153 (complete264_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I154 (complete264_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I155 (complete264_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I156 (complete264_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I157 (complete264_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I158 (complete264_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I159 (complete264_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I160 (complete264_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I161 (complete264_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I162 (complete264_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I163 (complete264_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I164 (complete264_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I165 (complete264_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I166 (complete264_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I167 (complete264_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I168 (complete264_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I169 (complete264_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I170 (complete264_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I171 (complete264_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I172 (complete264_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I173 (complete264_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I174 (complete264_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I175 (complete264_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I176 (complete264_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I177 (complete264_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I178 (complete264_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I179 (complete264_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I180 (complete264_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I181 (complete264_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I182 (complete264_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I183 (complete264_0n[33], ifint_0n[33], itint_0n[33]);
  OR2 I184 (complete264_0n[34], ifint_0n[34], itint_0n[34]);
  OR2 I185 (complete264_0n[35], ifint_0n[35], itint_0n[35]);
  INV I186 (gate263_0n, iaint_0n);
  C2RI I187 (itint_0n[0], i_0r1d[0], gate263_0n, initialise);
  C2RI I188 (itint_0n[1], i_0r1d[1], gate263_0n, initialise);
  C2RI I189 (itint_0n[2], i_0r1d[2], gate263_0n, initialise);
  C2RI I190 (itint_0n[3], i_0r1d[3], gate263_0n, initialise);
  C2RI I191 (itint_0n[4], i_0r1d[4], gate263_0n, initialise);
  C2RI I192 (itint_0n[5], i_0r1d[5], gate263_0n, initialise);
  C2RI I193 (itint_0n[6], i_0r1d[6], gate263_0n, initialise);
  C2RI I194 (itint_0n[7], i_0r1d[7], gate263_0n, initialise);
  C2RI I195 (itint_0n[8], i_0r1d[8], gate263_0n, initialise);
  C2RI I196 (itint_0n[9], i_0r1d[9], gate263_0n, initialise);
  C2RI I197 (itint_0n[10], i_0r1d[10], gate263_0n, initialise);
  C2RI I198 (itint_0n[11], i_0r1d[11], gate263_0n, initialise);
  C2RI I199 (itint_0n[12], i_0r1d[12], gate263_0n, initialise);
  C2RI I200 (itint_0n[13], i_0r1d[13], gate263_0n, initialise);
  C2RI I201 (itint_0n[14], i_0r1d[14], gate263_0n, initialise);
  C2RI I202 (itint_0n[15], i_0r1d[15], gate263_0n, initialise);
  C2RI I203 (itint_0n[16], i_0r1d[16], gate263_0n, initialise);
  C2RI I204 (itint_0n[17], i_0r1d[17], gate263_0n, initialise);
  C2RI I205 (itint_0n[18], i_0r1d[18], gate263_0n, initialise);
  C2RI I206 (itint_0n[19], i_0r1d[19], gate263_0n, initialise);
  C2RI I207 (itint_0n[20], i_0r1d[20], gate263_0n, initialise);
  C2RI I208 (itint_0n[21], i_0r1d[21], gate263_0n, initialise);
  C2RI I209 (itint_0n[22], i_0r1d[22], gate263_0n, initialise);
  C2RI I210 (itint_0n[23], i_0r1d[23], gate263_0n, initialise);
  C2RI I211 (itint_0n[24], i_0r1d[24], gate263_0n, initialise);
  C2RI I212 (itint_0n[25], i_0r1d[25], gate263_0n, initialise);
  C2RI I213 (itint_0n[26], i_0r1d[26], gate263_0n, initialise);
  C2RI I214 (itint_0n[27], i_0r1d[27], gate263_0n, initialise);
  C2RI I215 (itint_0n[28], i_0r1d[28], gate263_0n, initialise);
  C2RI I216 (itint_0n[29], i_0r1d[29], gate263_0n, initialise);
  C2RI I217 (itint_0n[30], i_0r1d[30], gate263_0n, initialise);
  C2RI I218 (itint_0n[31], i_0r1d[31], gate263_0n, initialise);
  C2RI I219 (itint_0n[32], i_0r1d[32], gate263_0n, initialise);
  C2RI I220 (itint_0n[33], i_0r1d[33], gate263_0n, initialise);
  C2RI I221 (itint_0n[34], i_0r1d[34], gate263_0n, initialise);
  C2RI I222 (itint_0n[35], i_0r1d[35], gate263_0n, initialise);
  C2RI I223 (ifint_0n[0], i_0r0d[0], gate263_0n, initialise);
  C2RI I224 (ifint_0n[1], i_0r0d[1], gate263_0n, initialise);
  C2RI I225 (ifint_0n[2], i_0r0d[2], gate263_0n, initialise);
  C2RI I226 (ifint_0n[3], i_0r0d[3], gate263_0n, initialise);
  C2RI I227 (ifint_0n[4], i_0r0d[4], gate263_0n, initialise);
  C2RI I228 (ifint_0n[5], i_0r0d[5], gate263_0n, initialise);
  C2RI I229 (ifint_0n[6], i_0r0d[6], gate263_0n, initialise);
  C2RI I230 (ifint_0n[7], i_0r0d[7], gate263_0n, initialise);
  C2RI I231 (ifint_0n[8], i_0r0d[8], gate263_0n, initialise);
  C2RI I232 (ifint_0n[9], i_0r0d[9], gate263_0n, initialise);
  C2RI I233 (ifint_0n[10], i_0r0d[10], gate263_0n, initialise);
  C2RI I234 (ifint_0n[11], i_0r0d[11], gate263_0n, initialise);
  C2RI I235 (ifint_0n[12], i_0r0d[12], gate263_0n, initialise);
  C2RI I236 (ifint_0n[13], i_0r0d[13], gate263_0n, initialise);
  C2RI I237 (ifint_0n[14], i_0r0d[14], gate263_0n, initialise);
  C2RI I238 (ifint_0n[15], i_0r0d[15], gate263_0n, initialise);
  C2RI I239 (ifint_0n[16], i_0r0d[16], gate263_0n, initialise);
  C2RI I240 (ifint_0n[17], i_0r0d[17], gate263_0n, initialise);
  C2RI I241 (ifint_0n[18], i_0r0d[18], gate263_0n, initialise);
  C2RI I242 (ifint_0n[19], i_0r0d[19], gate263_0n, initialise);
  C2RI I243 (ifint_0n[20], i_0r0d[20], gate263_0n, initialise);
  C2RI I244 (ifint_0n[21], i_0r0d[21], gate263_0n, initialise);
  C2RI I245 (ifint_0n[22], i_0r0d[22], gate263_0n, initialise);
  C2RI I246 (ifint_0n[23], i_0r0d[23], gate263_0n, initialise);
  C2RI I247 (ifint_0n[24], i_0r0d[24], gate263_0n, initialise);
  C2RI I248 (ifint_0n[25], i_0r0d[25], gate263_0n, initialise);
  C2RI I249 (ifint_0n[26], i_0r0d[26], gate263_0n, initialise);
  C2RI I250 (ifint_0n[27], i_0r0d[27], gate263_0n, initialise);
  C2RI I251 (ifint_0n[28], i_0r0d[28], gate263_0n, initialise);
  C2RI I252 (ifint_0n[29], i_0r0d[29], gate263_0n, initialise);
  C2RI I253 (ifint_0n[30], i_0r0d[30], gate263_0n, initialise);
  C2RI I254 (ifint_0n[31], i_0r0d[31], gate263_0n, initialise);
  C2RI I255 (ifint_0n[32], i_0r0d[32], gate263_0n, initialise);
  C2RI I256 (ifint_0n[33], i_0r0d[33], gate263_0n, initialise);
  C2RI I257 (ifint_0n[34], i_0r0d[34], gate263_0n, initialise);
  C2RI I258 (ifint_0n[35], i_0r0d[35], gate263_0n, initialise);
  C3 I259 (iaint_0n, icomplete_0n, oaint_0n, oaint_1n);
  assign ofint_0n = icomplete_0n;
  assign otint_1n[0] = itint_0n[0];
  assign otint_1n[1] = itint_0n[1];
  assign otint_1n[2] = itint_0n[2];
  assign otint_1n[3] = itint_0n[3];
  assign otint_1n[4] = itint_0n[4];
  assign otint_1n[5] = itint_0n[5];
  assign otint_1n[6] = itint_0n[6];
  assign otint_1n[7] = itint_0n[7];
  assign otint_1n[8] = itint_0n[8];
  assign otint_1n[9] = itint_0n[9];
  assign otint_1n[10] = itint_0n[10];
  assign otint_1n[11] = itint_0n[11];
  assign otint_1n[12] = itint_0n[12];
  assign otint_1n[13] = itint_0n[13];
  assign otint_1n[14] = itint_0n[14];
  assign otint_1n[15] = itint_0n[15];
  assign otint_1n[16] = itint_0n[16];
  assign otint_1n[17] = itint_0n[17];
  assign otint_1n[18] = itint_0n[18];
  assign otint_1n[19] = itint_0n[19];
  assign otint_1n[20] = itint_0n[20];
  assign otint_1n[21] = itint_0n[21];
  assign otint_1n[22] = itint_0n[22];
  assign otint_1n[23] = itint_0n[23];
  assign otint_1n[24] = itint_0n[24];
  assign otint_1n[25] = itint_0n[25];
  assign otint_1n[26] = itint_0n[26];
  assign otint_1n[27] = itint_0n[27];
  assign otint_1n[28] = itint_0n[28];
  assign otint_1n[29] = itint_0n[29];
  assign otint_1n[30] = itint_0n[30];
  assign otint_1n[31] = itint_0n[31];
  assign otint_1n[32] = itint_0n[32];
  assign otint_1n[33] = itint_0n[33];
  assign otint_1n[34] = itint_0n[34];
  assign otint_1n[35] = itint_0n[35];
  assign ofint_1n[0] = ifint_0n[0];
  assign ofint_1n[1] = ifint_0n[1];
  assign ofint_1n[2] = ifint_0n[2];
  assign ofint_1n[3] = ifint_0n[3];
  assign ofint_1n[4] = ifint_0n[4];
  assign ofint_1n[5] = ifint_0n[5];
  assign ofint_1n[6] = ifint_0n[6];
  assign ofint_1n[7] = ifint_0n[7];
  assign ofint_1n[8] = ifint_0n[8];
  assign ofint_1n[9] = ifint_0n[9];
  assign ofint_1n[10] = ifint_0n[10];
  assign ofint_1n[11] = ifint_0n[11];
  assign ofint_1n[12] = ifint_0n[12];
  assign ofint_1n[13] = ifint_0n[13];
  assign ofint_1n[14] = ifint_0n[14];
  assign ofint_1n[15] = ifint_0n[15];
  assign ofint_1n[16] = ifint_0n[16];
  assign ofint_1n[17] = ifint_0n[17];
  assign ofint_1n[18] = ifint_0n[18];
  assign ofint_1n[19] = ifint_0n[19];
  assign ofint_1n[20] = ifint_0n[20];
  assign ofint_1n[21] = ifint_0n[21];
  assign ofint_1n[22] = ifint_0n[22];
  assign ofint_1n[23] = ifint_0n[23];
  assign ofint_1n[24] = ifint_0n[24];
  assign ofint_1n[25] = ifint_0n[25];
  assign ofint_1n[26] = ifint_0n[26];
  assign ofint_1n[27] = ifint_0n[27];
  assign ofint_1n[28] = ifint_0n[28];
  assign ofint_1n[29] = ifint_0n[29];
  assign ofint_1n[30] = ifint_0n[30];
  assign ofint_1n[31] = ifint_0n[31];
  assign ofint_1n[32] = ifint_0n[32];
  assign ofint_1n[33] = ifint_0n[33];
  assign ofint_1n[34] = ifint_0n[34];
  assign ofint_1n[35] = ifint_0n[35];
  C3 I333 (internal_0n[36], complete260_0n[0], complete260_0n[1], complete260_0n[2]);
  C3 I334 (internal_0n[37], complete260_0n[3], complete260_0n[4], complete260_0n[5]);
  C3 I335 (internal_0n[38], complete260_0n[6], complete260_0n[7], complete260_0n[8]);
  C3 I336 (internal_0n[39], complete260_0n[9], complete260_0n[10], complete260_0n[11]);
  C3 I337 (internal_0n[40], complete260_0n[12], complete260_0n[13], complete260_0n[14]);
  C3 I338 (internal_0n[41], complete260_0n[15], complete260_0n[16], complete260_0n[17]);
  C3 I339 (internal_0n[42], complete260_0n[18], complete260_0n[19], complete260_0n[20]);
  C3 I340 (internal_0n[43], complete260_0n[21], complete260_0n[22], complete260_0n[23]);
  C3 I341 (internal_0n[44], complete260_0n[24], complete260_0n[25], complete260_0n[26]);
  C3 I342 (internal_0n[45], complete260_0n[27], complete260_0n[28], complete260_0n[29]);
  C3 I343 (internal_0n[46], complete260_0n[30], complete260_0n[31], complete260_0n[32]);
  C3 I344 (internal_0n[47], complete260_0n[33], complete260_0n[34], complete260_0n[35]);
  C3 I345 (internal_0n[48], internal_0n[36], internal_0n[37], internal_0n[38]);
  C3 I346 (internal_0n[49], internal_0n[39], internal_0n[40], internal_0n[41]);
  C3 I347 (internal_0n[50], internal_0n[42], internal_0n[43], internal_0n[44]);
  C3 I348 (internal_0n[51], internal_0n[45], internal_0n[46], internal_0n[47]);
  C2 I349 (internal_0n[52], internal_0n[48], internal_0n[49]);
  C2 I350 (internal_0n[53], internal_0n[50], internal_0n[51]);
  C2 I351 (icomplete_0n, internal_0n[52], internal_0n[53]);
  OR2 I352 (complete260_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I353 (complete260_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I354 (complete260_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I355 (complete260_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I356 (complete260_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I357 (complete260_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I358 (complete260_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I359 (complete260_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I360 (complete260_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I361 (complete260_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I362 (complete260_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I363 (complete260_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I364 (complete260_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I365 (complete260_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I366 (complete260_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I367 (complete260_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I368 (complete260_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I369 (complete260_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I370 (complete260_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I371 (complete260_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I372 (complete260_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I373 (complete260_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I374 (complete260_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I375 (complete260_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I376 (complete260_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I377 (complete260_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I378 (complete260_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I379 (complete260_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I380 (complete260_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I381 (complete260_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I382 (complete260_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I383 (complete260_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I384 (complete260_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I385 (complete260_0n[33], ifint_0n[33], itint_0n[33]);
  OR2 I386 (complete260_0n[34], ifint_0n[34], itint_0n[34]);
  OR2 I387 (complete260_0n[35], ifint_0n[35], itint_0n[35]);
endmodule

module BrzJ_l11__280_200_29 (
  i_0r, i_0a,
  i_1r, i_1a,
  o_0r, o_0a,
  initialise
);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  output o_0r;
  input o_0a;
  input initialise;
  wire ofint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire ifint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire gate280_0n;
  wire gate277_0n;
  wire gate274_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign i_1a = ifint_1n;
  INV I3 (gate280_0n, iaint_1n);
  C2RI I4 (ifint_1n, i_1r, gate280_0n, initialise);
  assign i_0a = ifint_0n;
  INV I6 (gate277_0n, iaint_0n);
  C2RI I7 (ifint_0n, i_0r, gate277_0n, initialise);
  assign oaint_0n = o_0r;
  INV I9 (gate274_0n, o_0a);
  C2RI I10 (o_0r, ofint_0n, gate274_0n, initialise);
  C2 I11 (ofint_0n, ifint_0n, ifint_1n);
endmodule

module BrzJ_l15__280_200_200_29 (
  i_0r, i_0a,
  i_1r, i_1a,
  i_2r, i_2a,
  o_0r, o_0a,
  initialise
);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  output o_0r;
  input o_0a;
  input initialise;
  wire ofint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire ifint_1n;
  wire ifint_2n;
  wire iaint_0n;
  wire iaint_1n;
  wire iaint_2n;
  wire gate292_0n;
  wire gate289_0n;
  wire gate286_0n;
  wire gate283_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign iaint_2n = oaint_0n;
  assign i_2a = ifint_2n;
  INV I4 (gate292_0n, iaint_2n);
  C2RI I5 (ifint_2n, i_2r, gate292_0n, initialise);
  assign i_1a = ifint_1n;
  INV I7 (gate289_0n, iaint_1n);
  C2RI I8 (ifint_1n, i_1r, gate289_0n, initialise);
  assign i_0a = ifint_0n;
  INV I10 (gate286_0n, iaint_0n);
  C2RI I11 (ifint_0n, i_0r, gate286_0n, initialise);
  assign oaint_0n = o_0r;
  INV I13 (gate283_0n, o_0a);
  C2RI I14 (o_0r, ofint_0n, gate283_0n, initialise);
  C3 I15 (ofint_0n, ifint_0n, ifint_1n, ifint_2n);
endmodule

module BrzJ_l19__280_200_200_200_29 (
  i_0r, i_0a,
  i_1r, i_1a,
  i_2r, i_2a,
  i_3r, i_3a,
  o_0r, o_0a,
  initialise
);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  output o_0r;
  input o_0a;
  input initialise;
  wire [1:0] internal_0n;
  wire ofint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire ifint_1n;
  wire ifint_2n;
  wire ifint_3n;
  wire iaint_0n;
  wire iaint_1n;
  wire iaint_2n;
  wire iaint_3n;
  wire gate307_0n;
  wire gate304_0n;
  wire gate301_0n;
  wire gate298_0n;
  wire gate295_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign iaint_2n = oaint_0n;
  assign iaint_3n = oaint_0n;
  assign i_3a = ifint_3n;
  INV I5 (gate307_0n, iaint_3n);
  C2RI I6 (ifint_3n, i_3r, gate307_0n, initialise);
  assign i_2a = ifint_2n;
  INV I8 (gate304_0n, iaint_2n);
  C2RI I9 (ifint_2n, i_2r, gate304_0n, initialise);
  assign i_1a = ifint_1n;
  INV I11 (gate301_0n, iaint_1n);
  C2RI I12 (ifint_1n, i_1r, gate301_0n, initialise);
  assign i_0a = ifint_0n;
  INV I14 (gate298_0n, iaint_0n);
  C2RI I15 (ifint_0n, i_0r, gate298_0n, initialise);
  assign oaint_0n = o_0r;
  INV I17 (gate295_0n, o_0a);
  C2RI I18 (o_0r, ofint_0n, gate295_0n, initialise);
  C2 I19 (internal_0n[0], ifint_0n, ifint_1n);
  C2 I20 (internal_0n[1], ifint_2n, ifint_3n);
  C2 I21 (ofint_0n, internal_0n[0], internal_0n[1]);
endmodule

module BrzJ_l23__280_200_200_200_200_29 (
  i_0r, i_0a,
  i_1r, i_1a,
  i_2r, i_2a,
  i_3r, i_3a,
  i_4r, i_4a,
  o_0r, o_0a,
  initialise
);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  input i_4r;
  output i_4a;
  output o_0r;
  input o_0a;
  input initialise;
  wire [1:0] internal_0n;
  wire ofint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire ifint_1n;
  wire ifint_2n;
  wire ifint_3n;
  wire ifint_4n;
  wire iaint_0n;
  wire iaint_1n;
  wire iaint_2n;
  wire iaint_3n;
  wire iaint_4n;
  wire gate325_0n;
  wire gate322_0n;
  wire gate319_0n;
  wire gate316_0n;
  wire gate313_0n;
  wire gate310_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign iaint_2n = oaint_0n;
  assign iaint_3n = oaint_0n;
  assign iaint_4n = oaint_0n;
  assign i_4a = ifint_4n;
  INV I6 (gate325_0n, iaint_4n);
  C2RI I7 (ifint_4n, i_4r, gate325_0n, initialise);
  assign i_3a = ifint_3n;
  INV I9 (gate322_0n, iaint_3n);
  C2RI I10 (ifint_3n, i_3r, gate322_0n, initialise);
  assign i_2a = ifint_2n;
  INV I12 (gate319_0n, iaint_2n);
  C2RI I13 (ifint_2n, i_2r, gate319_0n, initialise);
  assign i_1a = ifint_1n;
  INV I15 (gate316_0n, iaint_1n);
  C2RI I16 (ifint_1n, i_1r, gate316_0n, initialise);
  assign i_0a = ifint_0n;
  INV I18 (gate313_0n, iaint_0n);
  C2RI I19 (ifint_0n, i_0r, gate313_0n, initialise);
  assign oaint_0n = o_0r;
  INV I21 (gate310_0n, o_0a);
  C2RI I22 (o_0r, ofint_0n, gate310_0n, initialise);
  C3 I23 (internal_0n[0], ifint_0n, ifint_1n, ifint_2n);
  C2 I24 (internal_0n[1], ifint_3n, ifint_4n);
  C2 I25 (ofint_0n, internal_0n[0], internal_0n[1]);
endmodule

module BrzJ_l27__280_200_200_200_200_200_29 (
  i_0r, i_0a,
  i_1r, i_1a,
  i_2r, i_2a,
  i_3r, i_3a,
  i_4r, i_4a,
  i_5r, i_5a,
  o_0r, o_0a,
  initialise
);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  input i_4r;
  output i_4a;
  input i_5r;
  output i_5a;
  output o_0r;
  input o_0a;
  input initialise;
  wire [1:0] internal_0n;
  wire ofint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire ifint_1n;
  wire ifint_2n;
  wire ifint_3n;
  wire ifint_4n;
  wire ifint_5n;
  wire iaint_0n;
  wire iaint_1n;
  wire iaint_2n;
  wire iaint_3n;
  wire iaint_4n;
  wire iaint_5n;
  wire gate346_0n;
  wire gate343_0n;
  wire gate340_0n;
  wire gate337_0n;
  wire gate334_0n;
  wire gate331_0n;
  wire gate328_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign iaint_2n = oaint_0n;
  assign iaint_3n = oaint_0n;
  assign iaint_4n = oaint_0n;
  assign iaint_5n = oaint_0n;
  assign i_5a = ifint_5n;
  INV I7 (gate346_0n, iaint_5n);
  C2RI I8 (ifint_5n, i_5r, gate346_0n, initialise);
  assign i_4a = ifint_4n;
  INV I10 (gate343_0n, iaint_4n);
  C2RI I11 (ifint_4n, i_4r, gate343_0n, initialise);
  assign i_3a = ifint_3n;
  INV I13 (gate340_0n, iaint_3n);
  C2RI I14 (ifint_3n, i_3r, gate340_0n, initialise);
  assign i_2a = ifint_2n;
  INV I16 (gate337_0n, iaint_2n);
  C2RI I17 (ifint_2n, i_2r, gate337_0n, initialise);
  assign i_1a = ifint_1n;
  INV I19 (gate334_0n, iaint_1n);
  C2RI I20 (ifint_1n, i_1r, gate334_0n, initialise);
  assign i_0a = ifint_0n;
  INV I22 (gate331_0n, iaint_0n);
  C2RI I23 (ifint_0n, i_0r, gate331_0n, initialise);
  assign oaint_0n = o_0r;
  INV I25 (gate328_0n, o_0a);
  C2RI I26 (o_0r, ofint_0n, gate328_0n, initialise);
  C3 I27 (internal_0n[0], ifint_0n, ifint_1n, ifint_2n);
  C3 I28 (internal_0n[1], ifint_3n, ifint_4n, ifint_5n);
  C2 I29 (ofint_0n, internal_0n[0], internal_0n[1]);
endmodule

module BrzJ_l35__280_200_200_200_200_200_200_200__m45m (
  i_0r, i_0a,
  i_1r, i_1a,
  i_2r, i_2a,
  i_3r, i_3a,
  i_4r, i_4a,
  i_5r, i_5a,
  i_6r, i_6a,
  i_7r, i_7a,
  o_0r, o_0a,
  initialise
);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  input i_4r;
  output i_4a;
  input i_5r;
  output i_5a;
  input i_6r;
  output i_6a;
  input i_7r;
  output i_7a;
  output o_0r;
  input o_0a;
  input initialise;
  wire [2:0] internal_0n;
  wire ofint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire ifint_1n;
  wire ifint_2n;
  wire ifint_3n;
  wire ifint_4n;
  wire ifint_5n;
  wire ifint_6n;
  wire ifint_7n;
  wire iaint_0n;
  wire iaint_1n;
  wire iaint_2n;
  wire iaint_3n;
  wire iaint_4n;
  wire iaint_5n;
  wire iaint_6n;
  wire iaint_7n;
  wire gate373_0n;
  wire gate370_0n;
  wire gate367_0n;
  wire gate364_0n;
  wire gate361_0n;
  wire gate358_0n;
  wire gate355_0n;
  wire gate352_0n;
  wire gate349_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign iaint_2n = oaint_0n;
  assign iaint_3n = oaint_0n;
  assign iaint_4n = oaint_0n;
  assign iaint_5n = oaint_0n;
  assign iaint_6n = oaint_0n;
  assign iaint_7n = oaint_0n;
  assign i_7a = ifint_7n;
  INV I9 (gate373_0n, iaint_7n);
  C2RI I10 (ifint_7n, i_7r, gate373_0n, initialise);
  assign i_6a = ifint_6n;
  INV I12 (gate370_0n, iaint_6n);
  C2RI I13 (ifint_6n, i_6r, gate370_0n, initialise);
  assign i_5a = ifint_5n;
  INV I15 (gate367_0n, iaint_5n);
  C2RI I16 (ifint_5n, i_5r, gate367_0n, initialise);
  assign i_4a = ifint_4n;
  INV I18 (gate364_0n, iaint_4n);
  C2RI I19 (ifint_4n, i_4r, gate364_0n, initialise);
  assign i_3a = ifint_3n;
  INV I21 (gate361_0n, iaint_3n);
  C2RI I22 (ifint_3n, i_3r, gate361_0n, initialise);
  assign i_2a = ifint_2n;
  INV I24 (gate358_0n, iaint_2n);
  C2RI I25 (ifint_2n, i_2r, gate358_0n, initialise);
  assign i_1a = ifint_1n;
  INV I27 (gate355_0n, iaint_1n);
  C2RI I28 (ifint_1n, i_1r, gate355_0n, initialise);
  assign i_0a = ifint_0n;
  INV I30 (gate352_0n, iaint_0n);
  C2RI I31 (ifint_0n, i_0r, gate352_0n, initialise);
  assign oaint_0n = o_0r;
  INV I33 (gate349_0n, o_0a);
  C2RI I34 (o_0r, ofint_0n, gate349_0n, initialise);
  C3 I35 (internal_0n[0], ifint_0n, ifint_1n, ifint_2n);
  C3 I36 (internal_0n[1], ifint_3n, ifint_4n, ifint_5n);
  C2 I37 (internal_0n[2], ifint_6n, ifint_7n);
  C3 I38 (ofint_0n, internal_0n[0], internal_0n[1], internal_0n[2]);
endmodule

module BrzJ_l59__280_200_200_200_200_200_200_200__m46m (
  i_0r, i_0a,
  i_1r, i_1a,
  i_2r, i_2a,
  i_3r, i_3a,
  i_4r, i_4a,
  i_5r, i_5a,
  i_6r, i_6a,
  i_7r, i_7a,
  i_8r, i_8a,
  i_9r, i_9a,
  i_10r, i_10a,
  i_11r, i_11a,
  i_12r, i_12a,
  i_13r, i_13a,
  o_0r, o_0a,
  initialise
);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  input i_4r;
  output i_4a;
  input i_5r;
  output i_5a;
  input i_6r;
  output i_6a;
  input i_7r;
  output i_7a;
  input i_8r;
  output i_8a;
  input i_9r;
  output i_9a;
  input i_10r;
  output i_10a;
  input i_11r;
  output i_11a;
  input i_12r;
  output i_12a;
  input i_13r;
  output i_13a;
  output o_0r;
  input o_0a;
  input initialise;
  wire [6:0] internal_0n;
  wire ofint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire ifint_1n;
  wire ifint_2n;
  wire ifint_3n;
  wire ifint_4n;
  wire ifint_5n;
  wire ifint_6n;
  wire ifint_7n;
  wire ifint_8n;
  wire ifint_9n;
  wire ifint_10n;
  wire ifint_11n;
  wire ifint_12n;
  wire ifint_13n;
  wire iaint_0n;
  wire iaint_1n;
  wire iaint_2n;
  wire iaint_3n;
  wire iaint_4n;
  wire iaint_5n;
  wire iaint_6n;
  wire iaint_7n;
  wire iaint_8n;
  wire iaint_9n;
  wire iaint_10n;
  wire iaint_11n;
  wire iaint_12n;
  wire iaint_13n;
  wire gate418_0n;
  wire gate415_0n;
  wire gate412_0n;
  wire gate409_0n;
  wire gate406_0n;
  wire gate403_0n;
  wire gate400_0n;
  wire gate397_0n;
  wire gate394_0n;
  wire gate391_0n;
  wire gate388_0n;
  wire gate385_0n;
  wire gate382_0n;
  wire gate379_0n;
  wire gate376_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign iaint_2n = oaint_0n;
  assign iaint_3n = oaint_0n;
  assign iaint_4n = oaint_0n;
  assign iaint_5n = oaint_0n;
  assign iaint_6n = oaint_0n;
  assign iaint_7n = oaint_0n;
  assign iaint_8n = oaint_0n;
  assign iaint_9n = oaint_0n;
  assign iaint_10n = oaint_0n;
  assign iaint_11n = oaint_0n;
  assign iaint_12n = oaint_0n;
  assign iaint_13n = oaint_0n;
  assign i_13a = ifint_13n;
  INV I15 (gate418_0n, iaint_13n);
  C2RI I16 (ifint_13n, i_13r, gate418_0n, initialise);
  assign i_12a = ifint_12n;
  INV I18 (gate415_0n, iaint_12n);
  C2RI I19 (ifint_12n, i_12r, gate415_0n, initialise);
  assign i_11a = ifint_11n;
  INV I21 (gate412_0n, iaint_11n);
  C2RI I22 (ifint_11n, i_11r, gate412_0n, initialise);
  assign i_10a = ifint_10n;
  INV I24 (gate409_0n, iaint_10n);
  C2RI I25 (ifint_10n, i_10r, gate409_0n, initialise);
  assign i_9a = ifint_9n;
  INV I27 (gate406_0n, iaint_9n);
  C2RI I28 (ifint_9n, i_9r, gate406_0n, initialise);
  assign i_8a = ifint_8n;
  INV I30 (gate403_0n, iaint_8n);
  C2RI I31 (ifint_8n, i_8r, gate403_0n, initialise);
  assign i_7a = ifint_7n;
  INV I33 (gate400_0n, iaint_7n);
  C2RI I34 (ifint_7n, i_7r, gate400_0n, initialise);
  assign i_6a = ifint_6n;
  INV I36 (gate397_0n, iaint_6n);
  C2RI I37 (ifint_6n, i_6r, gate397_0n, initialise);
  assign i_5a = ifint_5n;
  INV I39 (gate394_0n, iaint_5n);
  C2RI I40 (ifint_5n, i_5r, gate394_0n, initialise);
  assign i_4a = ifint_4n;
  INV I42 (gate391_0n, iaint_4n);
  C2RI I43 (ifint_4n, i_4r, gate391_0n, initialise);
  assign i_3a = ifint_3n;
  INV I45 (gate388_0n, iaint_3n);
  C2RI I46 (ifint_3n, i_3r, gate388_0n, initialise);
  assign i_2a = ifint_2n;
  INV I48 (gate385_0n, iaint_2n);
  C2RI I49 (ifint_2n, i_2r, gate385_0n, initialise);
  assign i_1a = ifint_1n;
  INV I51 (gate382_0n, iaint_1n);
  C2RI I52 (ifint_1n, i_1r, gate382_0n, initialise);
  assign i_0a = ifint_0n;
  INV I54 (gate379_0n, iaint_0n);
  C2RI I55 (ifint_0n, i_0r, gate379_0n, initialise);
  assign oaint_0n = o_0r;
  INV I57 (gate376_0n, o_0a);
  C2RI I58 (o_0r, ofint_0n, gate376_0n, initialise);
  C3 I59 (internal_0n[0], ifint_0n, ifint_1n, ifint_2n);
  C3 I60 (internal_0n[1], ifint_3n, ifint_4n, ifint_5n);
  C3 I61 (internal_0n[2], ifint_6n, ifint_7n, ifint_8n);
  C3 I62 (internal_0n[3], ifint_9n, ifint_10n, ifint_11n);
  C2 I63 (internal_0n[4], ifint_12n, ifint_13n);
  C3 I64 (internal_0n[5], internal_0n[0], internal_0n[1], internal_0n[2]);
  C2 I65 (internal_0n[6], internal_0n[3], internal_0n[4]);
  C2 I66 (ofint_0n, internal_0n[5], internal_0n[6]);
endmodule

module BrzJ_l11__280_202_29 (
  i_0r, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input i_0r;
  output i_0a;
  input [1:0] i_1r0d;
  input [1:0] i_1r1d;
  output i_1a;
  output [1:0] o_0r0d;
  output [1:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [1:0] ofint_0n;
  wire [1:0] otint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire [1:0] ifint_1n;
  wire [1:0] itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [1:0] complete429_0n;
  wire gate428_0n;
  wire gate425_0n;
  wire [1:0] complete422_0n;
  wire gate421_0n;
  wire [1:0] joint_0n;
  wire [1:0] joinf_0n;
  wire icomplete_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  C2 I2 (i_1a, complete429_0n[0], complete429_0n[1]);
  OR2 I3 (complete429_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I4 (complete429_0n[1], ifint_1n[1], itint_1n[1]);
  INV I5 (gate428_0n, iaint_1n);
  C2RI I6 (itint_1n[0], i_1r1d[0], gate428_0n, initialise);
  C2RI I7 (itint_1n[1], i_1r1d[1], gate428_0n, initialise);
  C2RI I8 (ifint_1n[0], i_1r0d[0], gate428_0n, initialise);
  C2RI I9 (ifint_1n[1], i_1r0d[1], gate428_0n, initialise);
  assign i_0a = ifint_0n;
  INV I11 (gate425_0n, iaint_0n);
  C2RI I12 (ifint_0n, i_0r, gate425_0n, initialise);
  C2 I13 (oaint_0n, complete422_0n[0], complete422_0n[1]);
  OR2 I14 (complete422_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I15 (complete422_0n[1], o_0r0d[1], o_0r1d[1]);
  INV I16 (gate421_0n, o_0a);
  C2RI I17 (o_0r1d[0], otint_0n[0], gate421_0n, initialise);
  C2RI I18 (o_0r1d[1], otint_0n[1], gate421_0n, initialise);
  C2RI I19 (o_0r0d[0], ofint_0n[0], gate421_0n, initialise);
  C2RI I20 (o_0r0d[1], ofint_0n[1], gate421_0n, initialise);
  assign otint_0n[1] = joint_0n[1];
  assign ofint_0n[1] = joinf_0n[1];
  C2 I23 (otint_0n[0], joint_0n[0], icomplete_0n);
  C2 I24 (ofint_0n[0], joinf_0n[0], icomplete_0n);
  assign icomplete_0n = ifint_0n;
  assign joint_0n[0] = itint_1n[0];
  assign joint_0n[1] = itint_1n[1];
  assign joinf_0n[0] = ifint_1n[0];
  assign joinf_0n[1] = ifint_1n[1];
endmodule

module BrzJ_l11__280_203_29 (
  i_0r, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input i_0r;
  output i_0a;
  input [2:0] i_1r0d;
  input [2:0] i_1r1d;
  output i_1a;
  output [2:0] o_0r0d;
  output [2:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [2:0] ofint_0n;
  wire [2:0] otint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire [2:0] ifint_1n;
  wire [2:0] itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [2:0] complete440_0n;
  wire gate439_0n;
  wire gate436_0n;
  wire [2:0] complete433_0n;
  wire gate432_0n;
  wire [2:0] joint_0n;
  wire [2:0] joinf_0n;
  wire icomplete_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  C3 I2 (i_1a, complete440_0n[0], complete440_0n[1], complete440_0n[2]);
  OR2 I3 (complete440_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I4 (complete440_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I5 (complete440_0n[2], ifint_1n[2], itint_1n[2]);
  INV I6 (gate439_0n, iaint_1n);
  C2RI I7 (itint_1n[0], i_1r1d[0], gate439_0n, initialise);
  C2RI I8 (itint_1n[1], i_1r1d[1], gate439_0n, initialise);
  C2RI I9 (itint_1n[2], i_1r1d[2], gate439_0n, initialise);
  C2RI I10 (ifint_1n[0], i_1r0d[0], gate439_0n, initialise);
  C2RI I11 (ifint_1n[1], i_1r0d[1], gate439_0n, initialise);
  C2RI I12 (ifint_1n[2], i_1r0d[2], gate439_0n, initialise);
  assign i_0a = ifint_0n;
  INV I14 (gate436_0n, iaint_0n);
  C2RI I15 (ifint_0n, i_0r, gate436_0n, initialise);
  C3 I16 (oaint_0n, complete433_0n[0], complete433_0n[1], complete433_0n[2]);
  OR2 I17 (complete433_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I18 (complete433_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I19 (complete433_0n[2], o_0r0d[2], o_0r1d[2]);
  INV I20 (gate432_0n, o_0a);
  C2RI I21 (o_0r1d[0], otint_0n[0], gate432_0n, initialise);
  C2RI I22 (o_0r1d[1], otint_0n[1], gate432_0n, initialise);
  C2RI I23 (o_0r1d[2], otint_0n[2], gate432_0n, initialise);
  C2RI I24 (o_0r0d[0], ofint_0n[0], gate432_0n, initialise);
  C2RI I25 (o_0r0d[1], ofint_0n[1], gate432_0n, initialise);
  C2RI I26 (o_0r0d[2], ofint_0n[2], gate432_0n, initialise);
  assign otint_0n[1] = joint_0n[1];
  assign otint_0n[2] = joint_0n[2];
  assign ofint_0n[1] = joinf_0n[1];
  assign ofint_0n[2] = joinf_0n[2];
  C2 I31 (otint_0n[0], joint_0n[0], icomplete_0n);
  C2 I32 (ofint_0n[0], joinf_0n[0], icomplete_0n);
  assign icomplete_0n = ifint_0n;
  assign joint_0n[0] = itint_1n[0];
  assign joint_0n[1] = itint_1n[1];
  assign joint_0n[2] = itint_1n[2];
  assign joinf_0n[0] = ifint_1n[0];
  assign joinf_0n[1] = ifint_1n[1];
  assign joinf_0n[2] = ifint_1n[2];
endmodule

module BrzJ_l11__280_209_29 (
  i_0r, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input i_0r;
  output i_0a;
  input [8:0] i_1r0d;
  input [8:0] i_1r1d;
  output i_1a;
  output [8:0] o_0r0d;
  output [8:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [5:0] internal_0n;
  wire [8:0] ofint_0n;
  wire [8:0] otint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire [8:0] ifint_1n;
  wire [8:0] itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [8:0] complete451_0n;
  wire gate450_0n;
  wire gate447_0n;
  wire [8:0] complete444_0n;
  wire gate443_0n;
  wire [8:0] joint_0n;
  wire [8:0] joinf_0n;
  wire icomplete_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  C3 I2 (internal_0n[0], complete451_0n[0], complete451_0n[1], complete451_0n[2]);
  C3 I3 (internal_0n[1], complete451_0n[3], complete451_0n[4], complete451_0n[5]);
  C3 I4 (internal_0n[2], complete451_0n[6], complete451_0n[7], complete451_0n[8]);
  C3 I5 (i_1a, internal_0n[0], internal_0n[1], internal_0n[2]);
  OR2 I6 (complete451_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I7 (complete451_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I8 (complete451_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I9 (complete451_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I10 (complete451_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I11 (complete451_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I12 (complete451_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I13 (complete451_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I14 (complete451_0n[8], ifint_1n[8], itint_1n[8]);
  INV I15 (gate450_0n, iaint_1n);
  C2RI I16 (itint_1n[0], i_1r1d[0], gate450_0n, initialise);
  C2RI I17 (itint_1n[1], i_1r1d[1], gate450_0n, initialise);
  C2RI I18 (itint_1n[2], i_1r1d[2], gate450_0n, initialise);
  C2RI I19 (itint_1n[3], i_1r1d[3], gate450_0n, initialise);
  C2RI I20 (itint_1n[4], i_1r1d[4], gate450_0n, initialise);
  C2RI I21 (itint_1n[5], i_1r1d[5], gate450_0n, initialise);
  C2RI I22 (itint_1n[6], i_1r1d[6], gate450_0n, initialise);
  C2RI I23 (itint_1n[7], i_1r1d[7], gate450_0n, initialise);
  C2RI I24 (itint_1n[8], i_1r1d[8], gate450_0n, initialise);
  C2RI I25 (ifint_1n[0], i_1r0d[0], gate450_0n, initialise);
  C2RI I26 (ifint_1n[1], i_1r0d[1], gate450_0n, initialise);
  C2RI I27 (ifint_1n[2], i_1r0d[2], gate450_0n, initialise);
  C2RI I28 (ifint_1n[3], i_1r0d[3], gate450_0n, initialise);
  C2RI I29 (ifint_1n[4], i_1r0d[4], gate450_0n, initialise);
  C2RI I30 (ifint_1n[5], i_1r0d[5], gate450_0n, initialise);
  C2RI I31 (ifint_1n[6], i_1r0d[6], gate450_0n, initialise);
  C2RI I32 (ifint_1n[7], i_1r0d[7], gate450_0n, initialise);
  C2RI I33 (ifint_1n[8], i_1r0d[8], gate450_0n, initialise);
  assign i_0a = ifint_0n;
  INV I35 (gate447_0n, iaint_0n);
  C2RI I36 (ifint_0n, i_0r, gate447_0n, initialise);
  C3 I37 (internal_0n[3], complete444_0n[0], complete444_0n[1], complete444_0n[2]);
  C3 I38 (internal_0n[4], complete444_0n[3], complete444_0n[4], complete444_0n[5]);
  C3 I39 (internal_0n[5], complete444_0n[6], complete444_0n[7], complete444_0n[8]);
  C3 I40 (oaint_0n, internal_0n[3], internal_0n[4], internal_0n[5]);
  OR2 I41 (complete444_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I42 (complete444_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I43 (complete444_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I44 (complete444_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I45 (complete444_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I46 (complete444_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I47 (complete444_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I48 (complete444_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I49 (complete444_0n[8], o_0r0d[8], o_0r1d[8]);
  INV I50 (gate443_0n, o_0a);
  C2RI I51 (o_0r1d[0], otint_0n[0], gate443_0n, initialise);
  C2RI I52 (o_0r1d[1], otint_0n[1], gate443_0n, initialise);
  C2RI I53 (o_0r1d[2], otint_0n[2], gate443_0n, initialise);
  C2RI I54 (o_0r1d[3], otint_0n[3], gate443_0n, initialise);
  C2RI I55 (o_0r1d[4], otint_0n[4], gate443_0n, initialise);
  C2RI I56 (o_0r1d[5], otint_0n[5], gate443_0n, initialise);
  C2RI I57 (o_0r1d[6], otint_0n[6], gate443_0n, initialise);
  C2RI I58 (o_0r1d[7], otint_0n[7], gate443_0n, initialise);
  C2RI I59 (o_0r1d[8], otint_0n[8], gate443_0n, initialise);
  C2RI I60 (o_0r0d[0], ofint_0n[0], gate443_0n, initialise);
  C2RI I61 (o_0r0d[1], ofint_0n[1], gate443_0n, initialise);
  C2RI I62 (o_0r0d[2], ofint_0n[2], gate443_0n, initialise);
  C2RI I63 (o_0r0d[3], ofint_0n[3], gate443_0n, initialise);
  C2RI I64 (o_0r0d[4], ofint_0n[4], gate443_0n, initialise);
  C2RI I65 (o_0r0d[5], ofint_0n[5], gate443_0n, initialise);
  C2RI I66 (o_0r0d[6], ofint_0n[6], gate443_0n, initialise);
  C2RI I67 (o_0r0d[7], ofint_0n[7], gate443_0n, initialise);
  C2RI I68 (o_0r0d[8], ofint_0n[8], gate443_0n, initialise);
  assign otint_0n[1] = joint_0n[1];
  assign otint_0n[2] = joint_0n[2];
  assign otint_0n[3] = joint_0n[3];
  assign otint_0n[4] = joint_0n[4];
  assign otint_0n[5] = joint_0n[5];
  assign otint_0n[6] = joint_0n[6];
  assign otint_0n[7] = joint_0n[7];
  assign otint_0n[8] = joint_0n[8];
  assign ofint_0n[1] = joinf_0n[1];
  assign ofint_0n[2] = joinf_0n[2];
  assign ofint_0n[3] = joinf_0n[3];
  assign ofint_0n[4] = joinf_0n[4];
  assign ofint_0n[5] = joinf_0n[5];
  assign ofint_0n[6] = joinf_0n[6];
  assign ofint_0n[7] = joinf_0n[7];
  assign ofint_0n[8] = joinf_0n[8];
  C2 I85 (otint_0n[0], joint_0n[0], icomplete_0n);
  C2 I86 (ofint_0n[0], joinf_0n[0], icomplete_0n);
  assign icomplete_0n = ifint_0n;
  assign joint_0n[0] = itint_1n[0];
  assign joint_0n[1] = itint_1n[1];
  assign joint_0n[2] = itint_1n[2];
  assign joint_0n[3] = itint_1n[3];
  assign joint_0n[4] = itint_1n[4];
  assign joint_0n[5] = itint_1n[5];
  assign joint_0n[6] = itint_1n[6];
  assign joint_0n[7] = itint_1n[7];
  assign joint_0n[8] = itint_1n[8];
  assign joinf_0n[0] = ifint_1n[0];
  assign joinf_0n[1] = ifint_1n[1];
  assign joinf_0n[2] = ifint_1n[2];
  assign joinf_0n[3] = ifint_1n[3];
  assign joinf_0n[4] = ifint_1n[4];
  assign joinf_0n[5] = ifint_1n[5];
  assign joinf_0n[6] = ifint_1n[6];
  assign joinf_0n[7] = ifint_1n[7];
  assign joinf_0n[8] = ifint_1n[8];
endmodule

module BrzJ_l11__281_200_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input i_0r0d;
  input i_0r1d;
  output i_0a;
  input i_1r;
  output i_1a;
  output o_0r0d;
  output o_0r1d;
  input o_0a;
  input initialise;
  wire ofint_0n;
  wire otint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire ifint_1n;
  wire itint_0n;
  wire iaint_0n;
  wire iaint_1n;
  wire gate462_0n;
  wire complete459_0n;
  wire gate458_0n;
  wire complete455_0n;
  wire gate454_0n;
  wire joint_0n;
  wire joinf_0n;
  wire icomplete_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign i_1a = ifint_1n;
  INV I3 (gate462_0n, iaint_1n);
  C2RI I4 (ifint_1n, i_1r, gate462_0n, initialise);
  assign i_0a = complete459_0n;
  OR2 I6 (complete459_0n, ifint_0n, itint_0n);
  INV I7 (gate458_0n, iaint_0n);
  C2RI I8 (itint_0n, i_0r1d, gate458_0n, initialise);
  C2RI I9 (ifint_0n, i_0r0d, gate458_0n, initialise);
  assign oaint_0n = complete455_0n;
  OR2 I11 (complete455_0n, o_0r0d, o_0r1d);
  INV I12 (gate454_0n, o_0a);
  C2RI I13 (o_0r1d, otint_0n, gate454_0n, initialise);
  C2RI I14 (o_0r0d, ofint_0n, gate454_0n, initialise);
  C2 I15 (otint_0n, joint_0n, icomplete_0n);
  C2 I16 (ofint_0n, joinf_0n, icomplete_0n);
  assign icomplete_0n = ifint_1n;
  assign joint_0n = itint_0n;
  assign joinf_0n = ifint_0n;
endmodule

module BrzJ_l11__281_201_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input i_0r0d;
  input i_0r1d;
  output i_0a;
  input i_1r0d;
  input i_1r1d;
  output i_1a;
  output [1:0] o_0r0d;
  output [1:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [1:0] ofint_0n;
  wire [1:0] otint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire ifint_1n;
  wire itint_0n;
  wire itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire complete474_0n;
  wire gate473_0n;
  wire complete470_0n;
  wire gate469_0n;
  wire [1:0] complete466_0n;
  wire gate465_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign i_1a = complete474_0n;
  OR2 I3 (complete474_0n, ifint_1n, itint_1n);
  INV I4 (gate473_0n, iaint_1n);
  C2RI I5 (itint_1n, i_1r1d, gate473_0n, initialise);
  C2RI I6 (ifint_1n, i_1r0d, gate473_0n, initialise);
  assign i_0a = complete470_0n;
  OR2 I8 (complete470_0n, ifint_0n, itint_0n);
  INV I9 (gate469_0n, iaint_0n);
  C2RI I10 (itint_0n, i_0r1d, gate469_0n, initialise);
  C2RI I11 (ifint_0n, i_0r0d, gate469_0n, initialise);
  C2 I12 (oaint_0n, complete466_0n[0], complete466_0n[1]);
  OR2 I13 (complete466_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I14 (complete466_0n[1], o_0r0d[1], o_0r1d[1]);
  INV I15 (gate465_0n, o_0a);
  C2RI I16 (o_0r1d[0], otint_0n[0], gate465_0n, initialise);
  C2RI I17 (o_0r1d[1], otint_0n[1], gate465_0n, initialise);
  C2RI I18 (o_0r0d[0], ofint_0n[0], gate465_0n, initialise);
  C2RI I19 (o_0r0d[1], ofint_0n[1], gate465_0n, initialise);
  assign otint_0n[0] = itint_0n;
  assign otint_0n[1] = itint_1n;
  assign ofint_0n[0] = ifint_0n;
  assign ofint_0n[1] = ifint_1n;
endmodule

module BrzJ_l11__281_203_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input i_0r0d;
  input i_0r1d;
  output i_0a;
  input [2:0] i_1r0d;
  input [2:0] i_1r1d;
  output i_1a;
  output [3:0] o_0r0d;
  output [3:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [1:0] internal_0n;
  wire [3:0] ofint_0n;
  wire [3:0] otint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire [2:0] ifint_1n;
  wire itint_0n;
  wire [2:0] itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [2:0] complete486_0n;
  wire gate485_0n;
  wire complete482_0n;
  wire gate481_0n;
  wire [3:0] complete478_0n;
  wire gate477_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  C3 I2 (i_1a, complete486_0n[0], complete486_0n[1], complete486_0n[2]);
  OR2 I3 (complete486_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I4 (complete486_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I5 (complete486_0n[2], ifint_1n[2], itint_1n[2]);
  INV I6 (gate485_0n, iaint_1n);
  C2RI I7 (itint_1n[0], i_1r1d[0], gate485_0n, initialise);
  C2RI I8 (itint_1n[1], i_1r1d[1], gate485_0n, initialise);
  C2RI I9 (itint_1n[2], i_1r1d[2], gate485_0n, initialise);
  C2RI I10 (ifint_1n[0], i_1r0d[0], gate485_0n, initialise);
  C2RI I11 (ifint_1n[1], i_1r0d[1], gate485_0n, initialise);
  C2RI I12 (ifint_1n[2], i_1r0d[2], gate485_0n, initialise);
  assign i_0a = complete482_0n;
  OR2 I14 (complete482_0n, ifint_0n, itint_0n);
  INV I15 (gate481_0n, iaint_0n);
  C2RI I16 (itint_0n, i_0r1d, gate481_0n, initialise);
  C2RI I17 (ifint_0n, i_0r0d, gate481_0n, initialise);
  C2 I18 (internal_0n[0], complete478_0n[0], complete478_0n[1]);
  C2 I19 (internal_0n[1], complete478_0n[2], complete478_0n[3]);
  C2 I20 (oaint_0n, internal_0n[0], internal_0n[1]);
  OR2 I21 (complete478_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I22 (complete478_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I23 (complete478_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I24 (complete478_0n[3], o_0r0d[3], o_0r1d[3]);
  INV I25 (gate477_0n, o_0a);
  C2RI I26 (o_0r1d[0], otint_0n[0], gate477_0n, initialise);
  C2RI I27 (o_0r1d[1], otint_0n[1], gate477_0n, initialise);
  C2RI I28 (o_0r1d[2], otint_0n[2], gate477_0n, initialise);
  C2RI I29 (o_0r1d[3], otint_0n[3], gate477_0n, initialise);
  C2RI I30 (o_0r0d[0], ofint_0n[0], gate477_0n, initialise);
  C2RI I31 (o_0r0d[1], ofint_0n[1], gate477_0n, initialise);
  C2RI I32 (o_0r0d[2], ofint_0n[2], gate477_0n, initialise);
  C2RI I33 (o_0r0d[3], ofint_0n[3], gate477_0n, initialise);
  assign otint_0n[0] = itint_0n;
  assign otint_0n[1] = itint_1n[0];
  assign otint_0n[2] = itint_1n[1];
  assign otint_0n[3] = itint_1n[2];
  assign ofint_0n[0] = ifint_0n;
  assign ofint_0n[1] = ifint_1n[0];
  assign ofint_0n[2] = ifint_1n[1];
  assign ofint_0n[3] = ifint_1n[2];
endmodule

module BrzJ_l12__281_2031_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input i_0r0d;
  input i_0r1d;
  output i_0a;
  input [30:0] i_1r0d;
  input [30:0] i_1r1d;
  output i_1a;
  output [31:0] o_0r0d;
  output [31:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [33:0] internal_0n;
  wire [31:0] ofint_0n;
  wire [31:0] otint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire [30:0] ifint_1n;
  wire itint_0n;
  wire [30:0] itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [30:0] complete498_0n;
  wire gate497_0n;
  wire complete494_0n;
  wire gate493_0n;
  wire [31:0] complete490_0n;
  wire gate489_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  C3 I2 (internal_0n[0], complete498_0n[0], complete498_0n[1], complete498_0n[2]);
  C3 I3 (internal_0n[1], complete498_0n[3], complete498_0n[4], complete498_0n[5]);
  C3 I4 (internal_0n[2], complete498_0n[6], complete498_0n[7], complete498_0n[8]);
  C3 I5 (internal_0n[3], complete498_0n[9], complete498_0n[10], complete498_0n[11]);
  C3 I6 (internal_0n[4], complete498_0n[12], complete498_0n[13], complete498_0n[14]);
  C3 I7 (internal_0n[5], complete498_0n[15], complete498_0n[16], complete498_0n[17]);
  C3 I8 (internal_0n[6], complete498_0n[18], complete498_0n[19], complete498_0n[20]);
  C3 I9 (internal_0n[7], complete498_0n[21], complete498_0n[22], complete498_0n[23]);
  C3 I10 (internal_0n[8], complete498_0n[24], complete498_0n[25], complete498_0n[26]);
  C2 I11 (internal_0n[9], complete498_0n[27], complete498_0n[28]);
  C2 I12 (internal_0n[10], complete498_0n[29], complete498_0n[30]);
  C3 I13 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I14 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I15 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I16 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I17 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I18 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I19 (i_1a, internal_0n[15], internal_0n[16]);
  OR2 I20 (complete498_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I21 (complete498_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I22 (complete498_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I23 (complete498_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I24 (complete498_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I25 (complete498_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I26 (complete498_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I27 (complete498_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I28 (complete498_0n[8], ifint_1n[8], itint_1n[8]);
  OR2 I29 (complete498_0n[9], ifint_1n[9], itint_1n[9]);
  OR2 I30 (complete498_0n[10], ifint_1n[10], itint_1n[10]);
  OR2 I31 (complete498_0n[11], ifint_1n[11], itint_1n[11]);
  OR2 I32 (complete498_0n[12], ifint_1n[12], itint_1n[12]);
  OR2 I33 (complete498_0n[13], ifint_1n[13], itint_1n[13]);
  OR2 I34 (complete498_0n[14], ifint_1n[14], itint_1n[14]);
  OR2 I35 (complete498_0n[15], ifint_1n[15], itint_1n[15]);
  OR2 I36 (complete498_0n[16], ifint_1n[16], itint_1n[16]);
  OR2 I37 (complete498_0n[17], ifint_1n[17], itint_1n[17]);
  OR2 I38 (complete498_0n[18], ifint_1n[18], itint_1n[18]);
  OR2 I39 (complete498_0n[19], ifint_1n[19], itint_1n[19]);
  OR2 I40 (complete498_0n[20], ifint_1n[20], itint_1n[20]);
  OR2 I41 (complete498_0n[21], ifint_1n[21], itint_1n[21]);
  OR2 I42 (complete498_0n[22], ifint_1n[22], itint_1n[22]);
  OR2 I43 (complete498_0n[23], ifint_1n[23], itint_1n[23]);
  OR2 I44 (complete498_0n[24], ifint_1n[24], itint_1n[24]);
  OR2 I45 (complete498_0n[25], ifint_1n[25], itint_1n[25]);
  OR2 I46 (complete498_0n[26], ifint_1n[26], itint_1n[26]);
  OR2 I47 (complete498_0n[27], ifint_1n[27], itint_1n[27]);
  OR2 I48 (complete498_0n[28], ifint_1n[28], itint_1n[28]);
  OR2 I49 (complete498_0n[29], ifint_1n[29], itint_1n[29]);
  OR2 I50 (complete498_0n[30], ifint_1n[30], itint_1n[30]);
  INV I51 (gate497_0n, iaint_1n);
  C2RI I52 (itint_1n[0], i_1r1d[0], gate497_0n, initialise);
  C2RI I53 (itint_1n[1], i_1r1d[1], gate497_0n, initialise);
  C2RI I54 (itint_1n[2], i_1r1d[2], gate497_0n, initialise);
  C2RI I55 (itint_1n[3], i_1r1d[3], gate497_0n, initialise);
  C2RI I56 (itint_1n[4], i_1r1d[4], gate497_0n, initialise);
  C2RI I57 (itint_1n[5], i_1r1d[5], gate497_0n, initialise);
  C2RI I58 (itint_1n[6], i_1r1d[6], gate497_0n, initialise);
  C2RI I59 (itint_1n[7], i_1r1d[7], gate497_0n, initialise);
  C2RI I60 (itint_1n[8], i_1r1d[8], gate497_0n, initialise);
  C2RI I61 (itint_1n[9], i_1r1d[9], gate497_0n, initialise);
  C2RI I62 (itint_1n[10], i_1r1d[10], gate497_0n, initialise);
  C2RI I63 (itint_1n[11], i_1r1d[11], gate497_0n, initialise);
  C2RI I64 (itint_1n[12], i_1r1d[12], gate497_0n, initialise);
  C2RI I65 (itint_1n[13], i_1r1d[13], gate497_0n, initialise);
  C2RI I66 (itint_1n[14], i_1r1d[14], gate497_0n, initialise);
  C2RI I67 (itint_1n[15], i_1r1d[15], gate497_0n, initialise);
  C2RI I68 (itint_1n[16], i_1r1d[16], gate497_0n, initialise);
  C2RI I69 (itint_1n[17], i_1r1d[17], gate497_0n, initialise);
  C2RI I70 (itint_1n[18], i_1r1d[18], gate497_0n, initialise);
  C2RI I71 (itint_1n[19], i_1r1d[19], gate497_0n, initialise);
  C2RI I72 (itint_1n[20], i_1r1d[20], gate497_0n, initialise);
  C2RI I73 (itint_1n[21], i_1r1d[21], gate497_0n, initialise);
  C2RI I74 (itint_1n[22], i_1r1d[22], gate497_0n, initialise);
  C2RI I75 (itint_1n[23], i_1r1d[23], gate497_0n, initialise);
  C2RI I76 (itint_1n[24], i_1r1d[24], gate497_0n, initialise);
  C2RI I77 (itint_1n[25], i_1r1d[25], gate497_0n, initialise);
  C2RI I78 (itint_1n[26], i_1r1d[26], gate497_0n, initialise);
  C2RI I79 (itint_1n[27], i_1r1d[27], gate497_0n, initialise);
  C2RI I80 (itint_1n[28], i_1r1d[28], gate497_0n, initialise);
  C2RI I81 (itint_1n[29], i_1r1d[29], gate497_0n, initialise);
  C2RI I82 (itint_1n[30], i_1r1d[30], gate497_0n, initialise);
  C2RI I83 (ifint_1n[0], i_1r0d[0], gate497_0n, initialise);
  C2RI I84 (ifint_1n[1], i_1r0d[1], gate497_0n, initialise);
  C2RI I85 (ifint_1n[2], i_1r0d[2], gate497_0n, initialise);
  C2RI I86 (ifint_1n[3], i_1r0d[3], gate497_0n, initialise);
  C2RI I87 (ifint_1n[4], i_1r0d[4], gate497_0n, initialise);
  C2RI I88 (ifint_1n[5], i_1r0d[5], gate497_0n, initialise);
  C2RI I89 (ifint_1n[6], i_1r0d[6], gate497_0n, initialise);
  C2RI I90 (ifint_1n[7], i_1r0d[7], gate497_0n, initialise);
  C2RI I91 (ifint_1n[8], i_1r0d[8], gate497_0n, initialise);
  C2RI I92 (ifint_1n[9], i_1r0d[9], gate497_0n, initialise);
  C2RI I93 (ifint_1n[10], i_1r0d[10], gate497_0n, initialise);
  C2RI I94 (ifint_1n[11], i_1r0d[11], gate497_0n, initialise);
  C2RI I95 (ifint_1n[12], i_1r0d[12], gate497_0n, initialise);
  C2RI I96 (ifint_1n[13], i_1r0d[13], gate497_0n, initialise);
  C2RI I97 (ifint_1n[14], i_1r0d[14], gate497_0n, initialise);
  C2RI I98 (ifint_1n[15], i_1r0d[15], gate497_0n, initialise);
  C2RI I99 (ifint_1n[16], i_1r0d[16], gate497_0n, initialise);
  C2RI I100 (ifint_1n[17], i_1r0d[17], gate497_0n, initialise);
  C2RI I101 (ifint_1n[18], i_1r0d[18], gate497_0n, initialise);
  C2RI I102 (ifint_1n[19], i_1r0d[19], gate497_0n, initialise);
  C2RI I103 (ifint_1n[20], i_1r0d[20], gate497_0n, initialise);
  C2RI I104 (ifint_1n[21], i_1r0d[21], gate497_0n, initialise);
  C2RI I105 (ifint_1n[22], i_1r0d[22], gate497_0n, initialise);
  C2RI I106 (ifint_1n[23], i_1r0d[23], gate497_0n, initialise);
  C2RI I107 (ifint_1n[24], i_1r0d[24], gate497_0n, initialise);
  C2RI I108 (ifint_1n[25], i_1r0d[25], gate497_0n, initialise);
  C2RI I109 (ifint_1n[26], i_1r0d[26], gate497_0n, initialise);
  C2RI I110 (ifint_1n[27], i_1r0d[27], gate497_0n, initialise);
  C2RI I111 (ifint_1n[28], i_1r0d[28], gate497_0n, initialise);
  C2RI I112 (ifint_1n[29], i_1r0d[29], gate497_0n, initialise);
  C2RI I113 (ifint_1n[30], i_1r0d[30], gate497_0n, initialise);
  assign i_0a = complete494_0n;
  OR2 I115 (complete494_0n, ifint_0n, itint_0n);
  INV I116 (gate493_0n, iaint_0n);
  C2RI I117 (itint_0n, i_0r1d, gate493_0n, initialise);
  C2RI I118 (ifint_0n, i_0r0d, gate493_0n, initialise);
  C3 I119 (internal_0n[17], complete490_0n[0], complete490_0n[1], complete490_0n[2]);
  C3 I120 (internal_0n[18], complete490_0n[3], complete490_0n[4], complete490_0n[5]);
  C3 I121 (internal_0n[19], complete490_0n[6], complete490_0n[7], complete490_0n[8]);
  C3 I122 (internal_0n[20], complete490_0n[9], complete490_0n[10], complete490_0n[11]);
  C3 I123 (internal_0n[21], complete490_0n[12], complete490_0n[13], complete490_0n[14]);
  C3 I124 (internal_0n[22], complete490_0n[15], complete490_0n[16], complete490_0n[17]);
  C3 I125 (internal_0n[23], complete490_0n[18], complete490_0n[19], complete490_0n[20]);
  C3 I126 (internal_0n[24], complete490_0n[21], complete490_0n[22], complete490_0n[23]);
  C3 I127 (internal_0n[25], complete490_0n[24], complete490_0n[25], complete490_0n[26]);
  C3 I128 (internal_0n[26], complete490_0n[27], complete490_0n[28], complete490_0n[29]);
  C2 I129 (internal_0n[27], complete490_0n[30], complete490_0n[31]);
  C3 I130 (internal_0n[28], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I131 (internal_0n[29], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I132 (internal_0n[30], internal_0n[23], internal_0n[24], internal_0n[25]);
  C2 I133 (internal_0n[31], internal_0n[26], internal_0n[27]);
  C2 I134 (internal_0n[32], internal_0n[28], internal_0n[29]);
  C2 I135 (internal_0n[33], internal_0n[30], internal_0n[31]);
  C2 I136 (oaint_0n, internal_0n[32], internal_0n[33]);
  OR2 I137 (complete490_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I138 (complete490_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I139 (complete490_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I140 (complete490_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I141 (complete490_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I142 (complete490_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I143 (complete490_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I144 (complete490_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I145 (complete490_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I146 (complete490_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I147 (complete490_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I148 (complete490_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I149 (complete490_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I150 (complete490_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I151 (complete490_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I152 (complete490_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I153 (complete490_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I154 (complete490_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I155 (complete490_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I156 (complete490_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I157 (complete490_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I158 (complete490_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I159 (complete490_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I160 (complete490_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I161 (complete490_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I162 (complete490_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I163 (complete490_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I164 (complete490_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I165 (complete490_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I166 (complete490_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I167 (complete490_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I168 (complete490_0n[31], o_0r0d[31], o_0r1d[31]);
  INV I169 (gate489_0n, o_0a);
  C2RI I170 (o_0r1d[0], otint_0n[0], gate489_0n, initialise);
  C2RI I171 (o_0r1d[1], otint_0n[1], gate489_0n, initialise);
  C2RI I172 (o_0r1d[2], otint_0n[2], gate489_0n, initialise);
  C2RI I173 (o_0r1d[3], otint_0n[3], gate489_0n, initialise);
  C2RI I174 (o_0r1d[4], otint_0n[4], gate489_0n, initialise);
  C2RI I175 (o_0r1d[5], otint_0n[5], gate489_0n, initialise);
  C2RI I176 (o_0r1d[6], otint_0n[6], gate489_0n, initialise);
  C2RI I177 (o_0r1d[7], otint_0n[7], gate489_0n, initialise);
  C2RI I178 (o_0r1d[8], otint_0n[8], gate489_0n, initialise);
  C2RI I179 (o_0r1d[9], otint_0n[9], gate489_0n, initialise);
  C2RI I180 (o_0r1d[10], otint_0n[10], gate489_0n, initialise);
  C2RI I181 (o_0r1d[11], otint_0n[11], gate489_0n, initialise);
  C2RI I182 (o_0r1d[12], otint_0n[12], gate489_0n, initialise);
  C2RI I183 (o_0r1d[13], otint_0n[13], gate489_0n, initialise);
  C2RI I184 (o_0r1d[14], otint_0n[14], gate489_0n, initialise);
  C2RI I185 (o_0r1d[15], otint_0n[15], gate489_0n, initialise);
  C2RI I186 (o_0r1d[16], otint_0n[16], gate489_0n, initialise);
  C2RI I187 (o_0r1d[17], otint_0n[17], gate489_0n, initialise);
  C2RI I188 (o_0r1d[18], otint_0n[18], gate489_0n, initialise);
  C2RI I189 (o_0r1d[19], otint_0n[19], gate489_0n, initialise);
  C2RI I190 (o_0r1d[20], otint_0n[20], gate489_0n, initialise);
  C2RI I191 (o_0r1d[21], otint_0n[21], gate489_0n, initialise);
  C2RI I192 (o_0r1d[22], otint_0n[22], gate489_0n, initialise);
  C2RI I193 (o_0r1d[23], otint_0n[23], gate489_0n, initialise);
  C2RI I194 (o_0r1d[24], otint_0n[24], gate489_0n, initialise);
  C2RI I195 (o_0r1d[25], otint_0n[25], gate489_0n, initialise);
  C2RI I196 (o_0r1d[26], otint_0n[26], gate489_0n, initialise);
  C2RI I197 (o_0r1d[27], otint_0n[27], gate489_0n, initialise);
  C2RI I198 (o_0r1d[28], otint_0n[28], gate489_0n, initialise);
  C2RI I199 (o_0r1d[29], otint_0n[29], gate489_0n, initialise);
  C2RI I200 (o_0r1d[30], otint_0n[30], gate489_0n, initialise);
  C2RI I201 (o_0r1d[31], otint_0n[31], gate489_0n, initialise);
  C2RI I202 (o_0r0d[0], ofint_0n[0], gate489_0n, initialise);
  C2RI I203 (o_0r0d[1], ofint_0n[1], gate489_0n, initialise);
  C2RI I204 (o_0r0d[2], ofint_0n[2], gate489_0n, initialise);
  C2RI I205 (o_0r0d[3], ofint_0n[3], gate489_0n, initialise);
  C2RI I206 (o_0r0d[4], ofint_0n[4], gate489_0n, initialise);
  C2RI I207 (o_0r0d[5], ofint_0n[5], gate489_0n, initialise);
  C2RI I208 (o_0r0d[6], ofint_0n[6], gate489_0n, initialise);
  C2RI I209 (o_0r0d[7], ofint_0n[7], gate489_0n, initialise);
  C2RI I210 (o_0r0d[8], ofint_0n[8], gate489_0n, initialise);
  C2RI I211 (o_0r0d[9], ofint_0n[9], gate489_0n, initialise);
  C2RI I212 (o_0r0d[10], ofint_0n[10], gate489_0n, initialise);
  C2RI I213 (o_0r0d[11], ofint_0n[11], gate489_0n, initialise);
  C2RI I214 (o_0r0d[12], ofint_0n[12], gate489_0n, initialise);
  C2RI I215 (o_0r0d[13], ofint_0n[13], gate489_0n, initialise);
  C2RI I216 (o_0r0d[14], ofint_0n[14], gate489_0n, initialise);
  C2RI I217 (o_0r0d[15], ofint_0n[15], gate489_0n, initialise);
  C2RI I218 (o_0r0d[16], ofint_0n[16], gate489_0n, initialise);
  C2RI I219 (o_0r0d[17], ofint_0n[17], gate489_0n, initialise);
  C2RI I220 (o_0r0d[18], ofint_0n[18], gate489_0n, initialise);
  C2RI I221 (o_0r0d[19], ofint_0n[19], gate489_0n, initialise);
  C2RI I222 (o_0r0d[20], ofint_0n[20], gate489_0n, initialise);
  C2RI I223 (o_0r0d[21], ofint_0n[21], gate489_0n, initialise);
  C2RI I224 (o_0r0d[22], ofint_0n[22], gate489_0n, initialise);
  C2RI I225 (o_0r0d[23], ofint_0n[23], gate489_0n, initialise);
  C2RI I226 (o_0r0d[24], ofint_0n[24], gate489_0n, initialise);
  C2RI I227 (o_0r0d[25], ofint_0n[25], gate489_0n, initialise);
  C2RI I228 (o_0r0d[26], ofint_0n[26], gate489_0n, initialise);
  C2RI I229 (o_0r0d[27], ofint_0n[27], gate489_0n, initialise);
  C2RI I230 (o_0r0d[28], ofint_0n[28], gate489_0n, initialise);
  C2RI I231 (o_0r0d[29], ofint_0n[29], gate489_0n, initialise);
  C2RI I232 (o_0r0d[30], ofint_0n[30], gate489_0n, initialise);
  C2RI I233 (o_0r0d[31], ofint_0n[31], gate489_0n, initialise);
  assign otint_0n[0] = itint_0n;
  assign otint_0n[1] = itint_1n[0];
  assign otint_0n[2] = itint_1n[1];
  assign otint_0n[3] = itint_1n[2];
  assign otint_0n[4] = itint_1n[3];
  assign otint_0n[5] = itint_1n[4];
  assign otint_0n[6] = itint_1n[5];
  assign otint_0n[7] = itint_1n[6];
  assign otint_0n[8] = itint_1n[7];
  assign otint_0n[9] = itint_1n[8];
  assign otint_0n[10] = itint_1n[9];
  assign otint_0n[11] = itint_1n[10];
  assign otint_0n[12] = itint_1n[11];
  assign otint_0n[13] = itint_1n[12];
  assign otint_0n[14] = itint_1n[13];
  assign otint_0n[15] = itint_1n[14];
  assign otint_0n[16] = itint_1n[15];
  assign otint_0n[17] = itint_1n[16];
  assign otint_0n[18] = itint_1n[17];
  assign otint_0n[19] = itint_1n[18];
  assign otint_0n[20] = itint_1n[19];
  assign otint_0n[21] = itint_1n[20];
  assign otint_0n[22] = itint_1n[21];
  assign otint_0n[23] = itint_1n[22];
  assign otint_0n[24] = itint_1n[23];
  assign otint_0n[25] = itint_1n[24];
  assign otint_0n[26] = itint_1n[25];
  assign otint_0n[27] = itint_1n[26];
  assign otint_0n[28] = itint_1n[27];
  assign otint_0n[29] = itint_1n[28];
  assign otint_0n[30] = itint_1n[29];
  assign otint_0n[31] = itint_1n[30];
  assign ofint_0n[0] = ifint_0n;
  assign ofint_0n[1] = ifint_1n[0];
  assign ofint_0n[2] = ifint_1n[1];
  assign ofint_0n[3] = ifint_1n[2];
  assign ofint_0n[4] = ifint_1n[3];
  assign ofint_0n[5] = ifint_1n[4];
  assign ofint_0n[6] = ifint_1n[5];
  assign ofint_0n[7] = ifint_1n[6];
  assign ofint_0n[8] = ifint_1n[7];
  assign ofint_0n[9] = ifint_1n[8];
  assign ofint_0n[10] = ifint_1n[9];
  assign ofint_0n[11] = ifint_1n[10];
  assign ofint_0n[12] = ifint_1n[11];
  assign ofint_0n[13] = ifint_1n[12];
  assign ofint_0n[14] = ifint_1n[13];
  assign ofint_0n[15] = ifint_1n[14];
  assign ofint_0n[16] = ifint_1n[15];
  assign ofint_0n[17] = ifint_1n[16];
  assign ofint_0n[18] = ifint_1n[17];
  assign ofint_0n[19] = ifint_1n[18];
  assign ofint_0n[20] = ifint_1n[19];
  assign ofint_0n[21] = ifint_1n[20];
  assign ofint_0n[22] = ifint_1n[21];
  assign ofint_0n[23] = ifint_1n[22];
  assign ofint_0n[24] = ifint_1n[23];
  assign ofint_0n[25] = ifint_1n[24];
  assign ofint_0n[26] = ifint_1n[25];
  assign ofint_0n[27] = ifint_1n[26];
  assign ofint_0n[28] = ifint_1n[27];
  assign ofint_0n[29] = ifint_1n[28];
  assign ofint_0n[30] = ifint_1n[29];
  assign ofint_0n[31] = ifint_1n[30];
endmodule

module BrzJ_l12__281_2032_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input i_0r0d;
  input i_0r1d;
  output i_0a;
  input [31:0] i_1r0d;
  input [31:0] i_1r1d;
  output i_1a;
  output [32:0] o_0r0d;
  output [32:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [33:0] internal_0n;
  wire [32:0] ofint_0n;
  wire [32:0] otint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire [31:0] ifint_1n;
  wire itint_0n;
  wire [31:0] itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [31:0] complete510_0n;
  wire gate509_0n;
  wire complete506_0n;
  wire gate505_0n;
  wire [32:0] complete502_0n;
  wire gate501_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  C3 I2 (internal_0n[0], complete510_0n[0], complete510_0n[1], complete510_0n[2]);
  C3 I3 (internal_0n[1], complete510_0n[3], complete510_0n[4], complete510_0n[5]);
  C3 I4 (internal_0n[2], complete510_0n[6], complete510_0n[7], complete510_0n[8]);
  C3 I5 (internal_0n[3], complete510_0n[9], complete510_0n[10], complete510_0n[11]);
  C3 I6 (internal_0n[4], complete510_0n[12], complete510_0n[13], complete510_0n[14]);
  C3 I7 (internal_0n[5], complete510_0n[15], complete510_0n[16], complete510_0n[17]);
  C3 I8 (internal_0n[6], complete510_0n[18], complete510_0n[19], complete510_0n[20]);
  C3 I9 (internal_0n[7], complete510_0n[21], complete510_0n[22], complete510_0n[23]);
  C3 I10 (internal_0n[8], complete510_0n[24], complete510_0n[25], complete510_0n[26]);
  C3 I11 (internal_0n[9], complete510_0n[27], complete510_0n[28], complete510_0n[29]);
  C2 I12 (internal_0n[10], complete510_0n[30], complete510_0n[31]);
  C3 I13 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I14 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I15 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I16 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I17 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I18 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I19 (i_1a, internal_0n[15], internal_0n[16]);
  OR2 I20 (complete510_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I21 (complete510_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I22 (complete510_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I23 (complete510_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I24 (complete510_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I25 (complete510_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I26 (complete510_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I27 (complete510_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I28 (complete510_0n[8], ifint_1n[8], itint_1n[8]);
  OR2 I29 (complete510_0n[9], ifint_1n[9], itint_1n[9]);
  OR2 I30 (complete510_0n[10], ifint_1n[10], itint_1n[10]);
  OR2 I31 (complete510_0n[11], ifint_1n[11], itint_1n[11]);
  OR2 I32 (complete510_0n[12], ifint_1n[12], itint_1n[12]);
  OR2 I33 (complete510_0n[13], ifint_1n[13], itint_1n[13]);
  OR2 I34 (complete510_0n[14], ifint_1n[14], itint_1n[14]);
  OR2 I35 (complete510_0n[15], ifint_1n[15], itint_1n[15]);
  OR2 I36 (complete510_0n[16], ifint_1n[16], itint_1n[16]);
  OR2 I37 (complete510_0n[17], ifint_1n[17], itint_1n[17]);
  OR2 I38 (complete510_0n[18], ifint_1n[18], itint_1n[18]);
  OR2 I39 (complete510_0n[19], ifint_1n[19], itint_1n[19]);
  OR2 I40 (complete510_0n[20], ifint_1n[20], itint_1n[20]);
  OR2 I41 (complete510_0n[21], ifint_1n[21], itint_1n[21]);
  OR2 I42 (complete510_0n[22], ifint_1n[22], itint_1n[22]);
  OR2 I43 (complete510_0n[23], ifint_1n[23], itint_1n[23]);
  OR2 I44 (complete510_0n[24], ifint_1n[24], itint_1n[24]);
  OR2 I45 (complete510_0n[25], ifint_1n[25], itint_1n[25]);
  OR2 I46 (complete510_0n[26], ifint_1n[26], itint_1n[26]);
  OR2 I47 (complete510_0n[27], ifint_1n[27], itint_1n[27]);
  OR2 I48 (complete510_0n[28], ifint_1n[28], itint_1n[28]);
  OR2 I49 (complete510_0n[29], ifint_1n[29], itint_1n[29]);
  OR2 I50 (complete510_0n[30], ifint_1n[30], itint_1n[30]);
  OR2 I51 (complete510_0n[31], ifint_1n[31], itint_1n[31]);
  INV I52 (gate509_0n, iaint_1n);
  C2RI I53 (itint_1n[0], i_1r1d[0], gate509_0n, initialise);
  C2RI I54 (itint_1n[1], i_1r1d[1], gate509_0n, initialise);
  C2RI I55 (itint_1n[2], i_1r1d[2], gate509_0n, initialise);
  C2RI I56 (itint_1n[3], i_1r1d[3], gate509_0n, initialise);
  C2RI I57 (itint_1n[4], i_1r1d[4], gate509_0n, initialise);
  C2RI I58 (itint_1n[5], i_1r1d[5], gate509_0n, initialise);
  C2RI I59 (itint_1n[6], i_1r1d[6], gate509_0n, initialise);
  C2RI I60 (itint_1n[7], i_1r1d[7], gate509_0n, initialise);
  C2RI I61 (itint_1n[8], i_1r1d[8], gate509_0n, initialise);
  C2RI I62 (itint_1n[9], i_1r1d[9], gate509_0n, initialise);
  C2RI I63 (itint_1n[10], i_1r1d[10], gate509_0n, initialise);
  C2RI I64 (itint_1n[11], i_1r1d[11], gate509_0n, initialise);
  C2RI I65 (itint_1n[12], i_1r1d[12], gate509_0n, initialise);
  C2RI I66 (itint_1n[13], i_1r1d[13], gate509_0n, initialise);
  C2RI I67 (itint_1n[14], i_1r1d[14], gate509_0n, initialise);
  C2RI I68 (itint_1n[15], i_1r1d[15], gate509_0n, initialise);
  C2RI I69 (itint_1n[16], i_1r1d[16], gate509_0n, initialise);
  C2RI I70 (itint_1n[17], i_1r1d[17], gate509_0n, initialise);
  C2RI I71 (itint_1n[18], i_1r1d[18], gate509_0n, initialise);
  C2RI I72 (itint_1n[19], i_1r1d[19], gate509_0n, initialise);
  C2RI I73 (itint_1n[20], i_1r1d[20], gate509_0n, initialise);
  C2RI I74 (itint_1n[21], i_1r1d[21], gate509_0n, initialise);
  C2RI I75 (itint_1n[22], i_1r1d[22], gate509_0n, initialise);
  C2RI I76 (itint_1n[23], i_1r1d[23], gate509_0n, initialise);
  C2RI I77 (itint_1n[24], i_1r1d[24], gate509_0n, initialise);
  C2RI I78 (itint_1n[25], i_1r1d[25], gate509_0n, initialise);
  C2RI I79 (itint_1n[26], i_1r1d[26], gate509_0n, initialise);
  C2RI I80 (itint_1n[27], i_1r1d[27], gate509_0n, initialise);
  C2RI I81 (itint_1n[28], i_1r1d[28], gate509_0n, initialise);
  C2RI I82 (itint_1n[29], i_1r1d[29], gate509_0n, initialise);
  C2RI I83 (itint_1n[30], i_1r1d[30], gate509_0n, initialise);
  C2RI I84 (itint_1n[31], i_1r1d[31], gate509_0n, initialise);
  C2RI I85 (ifint_1n[0], i_1r0d[0], gate509_0n, initialise);
  C2RI I86 (ifint_1n[1], i_1r0d[1], gate509_0n, initialise);
  C2RI I87 (ifint_1n[2], i_1r0d[2], gate509_0n, initialise);
  C2RI I88 (ifint_1n[3], i_1r0d[3], gate509_0n, initialise);
  C2RI I89 (ifint_1n[4], i_1r0d[4], gate509_0n, initialise);
  C2RI I90 (ifint_1n[5], i_1r0d[5], gate509_0n, initialise);
  C2RI I91 (ifint_1n[6], i_1r0d[6], gate509_0n, initialise);
  C2RI I92 (ifint_1n[7], i_1r0d[7], gate509_0n, initialise);
  C2RI I93 (ifint_1n[8], i_1r0d[8], gate509_0n, initialise);
  C2RI I94 (ifint_1n[9], i_1r0d[9], gate509_0n, initialise);
  C2RI I95 (ifint_1n[10], i_1r0d[10], gate509_0n, initialise);
  C2RI I96 (ifint_1n[11], i_1r0d[11], gate509_0n, initialise);
  C2RI I97 (ifint_1n[12], i_1r0d[12], gate509_0n, initialise);
  C2RI I98 (ifint_1n[13], i_1r0d[13], gate509_0n, initialise);
  C2RI I99 (ifint_1n[14], i_1r0d[14], gate509_0n, initialise);
  C2RI I100 (ifint_1n[15], i_1r0d[15], gate509_0n, initialise);
  C2RI I101 (ifint_1n[16], i_1r0d[16], gate509_0n, initialise);
  C2RI I102 (ifint_1n[17], i_1r0d[17], gate509_0n, initialise);
  C2RI I103 (ifint_1n[18], i_1r0d[18], gate509_0n, initialise);
  C2RI I104 (ifint_1n[19], i_1r0d[19], gate509_0n, initialise);
  C2RI I105 (ifint_1n[20], i_1r0d[20], gate509_0n, initialise);
  C2RI I106 (ifint_1n[21], i_1r0d[21], gate509_0n, initialise);
  C2RI I107 (ifint_1n[22], i_1r0d[22], gate509_0n, initialise);
  C2RI I108 (ifint_1n[23], i_1r0d[23], gate509_0n, initialise);
  C2RI I109 (ifint_1n[24], i_1r0d[24], gate509_0n, initialise);
  C2RI I110 (ifint_1n[25], i_1r0d[25], gate509_0n, initialise);
  C2RI I111 (ifint_1n[26], i_1r0d[26], gate509_0n, initialise);
  C2RI I112 (ifint_1n[27], i_1r0d[27], gate509_0n, initialise);
  C2RI I113 (ifint_1n[28], i_1r0d[28], gate509_0n, initialise);
  C2RI I114 (ifint_1n[29], i_1r0d[29], gate509_0n, initialise);
  C2RI I115 (ifint_1n[30], i_1r0d[30], gate509_0n, initialise);
  C2RI I116 (ifint_1n[31], i_1r0d[31], gate509_0n, initialise);
  assign i_0a = complete506_0n;
  OR2 I118 (complete506_0n, ifint_0n, itint_0n);
  INV I119 (gate505_0n, iaint_0n);
  C2RI I120 (itint_0n, i_0r1d, gate505_0n, initialise);
  C2RI I121 (ifint_0n, i_0r0d, gate505_0n, initialise);
  C3 I122 (internal_0n[17], complete502_0n[0], complete502_0n[1], complete502_0n[2]);
  C3 I123 (internal_0n[18], complete502_0n[3], complete502_0n[4], complete502_0n[5]);
  C3 I124 (internal_0n[19], complete502_0n[6], complete502_0n[7], complete502_0n[8]);
  C3 I125 (internal_0n[20], complete502_0n[9], complete502_0n[10], complete502_0n[11]);
  C3 I126 (internal_0n[21], complete502_0n[12], complete502_0n[13], complete502_0n[14]);
  C3 I127 (internal_0n[22], complete502_0n[15], complete502_0n[16], complete502_0n[17]);
  C3 I128 (internal_0n[23], complete502_0n[18], complete502_0n[19], complete502_0n[20]);
  C3 I129 (internal_0n[24], complete502_0n[21], complete502_0n[22], complete502_0n[23]);
  C3 I130 (internal_0n[25], complete502_0n[24], complete502_0n[25], complete502_0n[26]);
  C3 I131 (internal_0n[26], complete502_0n[27], complete502_0n[28], complete502_0n[29]);
  C3 I132 (internal_0n[27], complete502_0n[30], complete502_0n[31], complete502_0n[32]);
  C3 I133 (internal_0n[28], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I134 (internal_0n[29], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I135 (internal_0n[30], internal_0n[23], internal_0n[24], internal_0n[25]);
  C2 I136 (internal_0n[31], internal_0n[26], internal_0n[27]);
  C2 I137 (internal_0n[32], internal_0n[28], internal_0n[29]);
  C2 I138 (internal_0n[33], internal_0n[30], internal_0n[31]);
  C2 I139 (oaint_0n, internal_0n[32], internal_0n[33]);
  OR2 I140 (complete502_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I141 (complete502_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I142 (complete502_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I143 (complete502_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I144 (complete502_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I145 (complete502_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I146 (complete502_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I147 (complete502_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I148 (complete502_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I149 (complete502_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I150 (complete502_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I151 (complete502_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I152 (complete502_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I153 (complete502_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I154 (complete502_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I155 (complete502_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I156 (complete502_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I157 (complete502_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I158 (complete502_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I159 (complete502_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I160 (complete502_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I161 (complete502_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I162 (complete502_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I163 (complete502_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I164 (complete502_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I165 (complete502_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I166 (complete502_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I167 (complete502_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I168 (complete502_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I169 (complete502_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I170 (complete502_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I171 (complete502_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I172 (complete502_0n[32], o_0r0d[32], o_0r1d[32]);
  INV I173 (gate501_0n, o_0a);
  C2RI I174 (o_0r1d[0], otint_0n[0], gate501_0n, initialise);
  C2RI I175 (o_0r1d[1], otint_0n[1], gate501_0n, initialise);
  C2RI I176 (o_0r1d[2], otint_0n[2], gate501_0n, initialise);
  C2RI I177 (o_0r1d[3], otint_0n[3], gate501_0n, initialise);
  C2RI I178 (o_0r1d[4], otint_0n[4], gate501_0n, initialise);
  C2RI I179 (o_0r1d[5], otint_0n[5], gate501_0n, initialise);
  C2RI I180 (o_0r1d[6], otint_0n[6], gate501_0n, initialise);
  C2RI I181 (o_0r1d[7], otint_0n[7], gate501_0n, initialise);
  C2RI I182 (o_0r1d[8], otint_0n[8], gate501_0n, initialise);
  C2RI I183 (o_0r1d[9], otint_0n[9], gate501_0n, initialise);
  C2RI I184 (o_0r1d[10], otint_0n[10], gate501_0n, initialise);
  C2RI I185 (o_0r1d[11], otint_0n[11], gate501_0n, initialise);
  C2RI I186 (o_0r1d[12], otint_0n[12], gate501_0n, initialise);
  C2RI I187 (o_0r1d[13], otint_0n[13], gate501_0n, initialise);
  C2RI I188 (o_0r1d[14], otint_0n[14], gate501_0n, initialise);
  C2RI I189 (o_0r1d[15], otint_0n[15], gate501_0n, initialise);
  C2RI I190 (o_0r1d[16], otint_0n[16], gate501_0n, initialise);
  C2RI I191 (o_0r1d[17], otint_0n[17], gate501_0n, initialise);
  C2RI I192 (o_0r1d[18], otint_0n[18], gate501_0n, initialise);
  C2RI I193 (o_0r1d[19], otint_0n[19], gate501_0n, initialise);
  C2RI I194 (o_0r1d[20], otint_0n[20], gate501_0n, initialise);
  C2RI I195 (o_0r1d[21], otint_0n[21], gate501_0n, initialise);
  C2RI I196 (o_0r1d[22], otint_0n[22], gate501_0n, initialise);
  C2RI I197 (o_0r1d[23], otint_0n[23], gate501_0n, initialise);
  C2RI I198 (o_0r1d[24], otint_0n[24], gate501_0n, initialise);
  C2RI I199 (o_0r1d[25], otint_0n[25], gate501_0n, initialise);
  C2RI I200 (o_0r1d[26], otint_0n[26], gate501_0n, initialise);
  C2RI I201 (o_0r1d[27], otint_0n[27], gate501_0n, initialise);
  C2RI I202 (o_0r1d[28], otint_0n[28], gate501_0n, initialise);
  C2RI I203 (o_0r1d[29], otint_0n[29], gate501_0n, initialise);
  C2RI I204 (o_0r1d[30], otint_0n[30], gate501_0n, initialise);
  C2RI I205 (o_0r1d[31], otint_0n[31], gate501_0n, initialise);
  C2RI I206 (o_0r1d[32], otint_0n[32], gate501_0n, initialise);
  C2RI I207 (o_0r0d[0], ofint_0n[0], gate501_0n, initialise);
  C2RI I208 (o_0r0d[1], ofint_0n[1], gate501_0n, initialise);
  C2RI I209 (o_0r0d[2], ofint_0n[2], gate501_0n, initialise);
  C2RI I210 (o_0r0d[3], ofint_0n[3], gate501_0n, initialise);
  C2RI I211 (o_0r0d[4], ofint_0n[4], gate501_0n, initialise);
  C2RI I212 (o_0r0d[5], ofint_0n[5], gate501_0n, initialise);
  C2RI I213 (o_0r0d[6], ofint_0n[6], gate501_0n, initialise);
  C2RI I214 (o_0r0d[7], ofint_0n[7], gate501_0n, initialise);
  C2RI I215 (o_0r0d[8], ofint_0n[8], gate501_0n, initialise);
  C2RI I216 (o_0r0d[9], ofint_0n[9], gate501_0n, initialise);
  C2RI I217 (o_0r0d[10], ofint_0n[10], gate501_0n, initialise);
  C2RI I218 (o_0r0d[11], ofint_0n[11], gate501_0n, initialise);
  C2RI I219 (o_0r0d[12], ofint_0n[12], gate501_0n, initialise);
  C2RI I220 (o_0r0d[13], ofint_0n[13], gate501_0n, initialise);
  C2RI I221 (o_0r0d[14], ofint_0n[14], gate501_0n, initialise);
  C2RI I222 (o_0r0d[15], ofint_0n[15], gate501_0n, initialise);
  C2RI I223 (o_0r0d[16], ofint_0n[16], gate501_0n, initialise);
  C2RI I224 (o_0r0d[17], ofint_0n[17], gate501_0n, initialise);
  C2RI I225 (o_0r0d[18], ofint_0n[18], gate501_0n, initialise);
  C2RI I226 (o_0r0d[19], ofint_0n[19], gate501_0n, initialise);
  C2RI I227 (o_0r0d[20], ofint_0n[20], gate501_0n, initialise);
  C2RI I228 (o_0r0d[21], ofint_0n[21], gate501_0n, initialise);
  C2RI I229 (o_0r0d[22], ofint_0n[22], gate501_0n, initialise);
  C2RI I230 (o_0r0d[23], ofint_0n[23], gate501_0n, initialise);
  C2RI I231 (o_0r0d[24], ofint_0n[24], gate501_0n, initialise);
  C2RI I232 (o_0r0d[25], ofint_0n[25], gate501_0n, initialise);
  C2RI I233 (o_0r0d[26], ofint_0n[26], gate501_0n, initialise);
  C2RI I234 (o_0r0d[27], ofint_0n[27], gate501_0n, initialise);
  C2RI I235 (o_0r0d[28], ofint_0n[28], gate501_0n, initialise);
  C2RI I236 (o_0r0d[29], ofint_0n[29], gate501_0n, initialise);
  C2RI I237 (o_0r0d[30], ofint_0n[30], gate501_0n, initialise);
  C2RI I238 (o_0r0d[31], ofint_0n[31], gate501_0n, initialise);
  C2RI I239 (o_0r0d[32], ofint_0n[32], gate501_0n, initialise);
  assign otint_0n[0] = itint_0n;
  assign otint_0n[1] = itint_1n[0];
  assign otint_0n[2] = itint_1n[1];
  assign otint_0n[3] = itint_1n[2];
  assign otint_0n[4] = itint_1n[3];
  assign otint_0n[5] = itint_1n[4];
  assign otint_0n[6] = itint_1n[5];
  assign otint_0n[7] = itint_1n[6];
  assign otint_0n[8] = itint_1n[7];
  assign otint_0n[9] = itint_1n[8];
  assign otint_0n[10] = itint_1n[9];
  assign otint_0n[11] = itint_1n[10];
  assign otint_0n[12] = itint_1n[11];
  assign otint_0n[13] = itint_1n[12];
  assign otint_0n[14] = itint_1n[13];
  assign otint_0n[15] = itint_1n[14];
  assign otint_0n[16] = itint_1n[15];
  assign otint_0n[17] = itint_1n[16];
  assign otint_0n[18] = itint_1n[17];
  assign otint_0n[19] = itint_1n[18];
  assign otint_0n[20] = itint_1n[19];
  assign otint_0n[21] = itint_1n[20];
  assign otint_0n[22] = itint_1n[21];
  assign otint_0n[23] = itint_1n[22];
  assign otint_0n[24] = itint_1n[23];
  assign otint_0n[25] = itint_1n[24];
  assign otint_0n[26] = itint_1n[25];
  assign otint_0n[27] = itint_1n[26];
  assign otint_0n[28] = itint_1n[27];
  assign otint_0n[29] = itint_1n[28];
  assign otint_0n[30] = itint_1n[29];
  assign otint_0n[31] = itint_1n[30];
  assign otint_0n[32] = itint_1n[31];
  assign ofint_0n[0] = ifint_0n;
  assign ofint_0n[1] = ifint_1n[0];
  assign ofint_0n[2] = ifint_1n[1];
  assign ofint_0n[3] = ifint_1n[2];
  assign ofint_0n[4] = ifint_1n[3];
  assign ofint_0n[5] = ifint_1n[4];
  assign ofint_0n[6] = ifint_1n[5];
  assign ofint_0n[7] = ifint_1n[6];
  assign ofint_0n[8] = ifint_1n[7];
  assign ofint_0n[9] = ifint_1n[8];
  assign ofint_0n[10] = ifint_1n[9];
  assign ofint_0n[11] = ifint_1n[10];
  assign ofint_0n[12] = ifint_1n[11];
  assign ofint_0n[13] = ifint_1n[12];
  assign ofint_0n[14] = ifint_1n[13];
  assign ofint_0n[15] = ifint_1n[14];
  assign ofint_0n[16] = ifint_1n[15];
  assign ofint_0n[17] = ifint_1n[16];
  assign ofint_0n[18] = ifint_1n[17];
  assign ofint_0n[19] = ifint_1n[18];
  assign ofint_0n[20] = ifint_1n[19];
  assign ofint_0n[21] = ifint_1n[20];
  assign ofint_0n[22] = ifint_1n[21];
  assign ofint_0n[23] = ifint_1n[22];
  assign ofint_0n[24] = ifint_1n[23];
  assign ofint_0n[25] = ifint_1n[24];
  assign ofint_0n[26] = ifint_1n[25];
  assign ofint_0n[27] = ifint_1n[26];
  assign ofint_0n[28] = ifint_1n[27];
  assign ofint_0n[29] = ifint_1n[28];
  assign ofint_0n[30] = ifint_1n[29];
  assign ofint_0n[31] = ifint_1n[30];
  assign ofint_0n[32] = ifint_1n[31];
endmodule

module BrzJ_l12__281_2034_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input i_0r0d;
  input i_0r1d;
  output i_0a;
  input [33:0] i_1r0d;
  input [33:0] i_1r1d;
  output i_1a;
  output [34:0] o_0r0d;
  output [34:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [35:0] internal_0n;
  wire [34:0] ofint_0n;
  wire [34:0] otint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire [33:0] ifint_1n;
  wire itint_0n;
  wire [33:0] itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [33:0] complete522_0n;
  wire gate521_0n;
  wire complete518_0n;
  wire gate517_0n;
  wire [34:0] complete514_0n;
  wire gate513_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  C3 I2 (internal_0n[0], complete522_0n[0], complete522_0n[1], complete522_0n[2]);
  C3 I3 (internal_0n[1], complete522_0n[3], complete522_0n[4], complete522_0n[5]);
  C3 I4 (internal_0n[2], complete522_0n[6], complete522_0n[7], complete522_0n[8]);
  C3 I5 (internal_0n[3], complete522_0n[9], complete522_0n[10], complete522_0n[11]);
  C3 I6 (internal_0n[4], complete522_0n[12], complete522_0n[13], complete522_0n[14]);
  C3 I7 (internal_0n[5], complete522_0n[15], complete522_0n[16], complete522_0n[17]);
  C3 I8 (internal_0n[6], complete522_0n[18], complete522_0n[19], complete522_0n[20]);
  C3 I9 (internal_0n[7], complete522_0n[21], complete522_0n[22], complete522_0n[23]);
  C3 I10 (internal_0n[8], complete522_0n[24], complete522_0n[25], complete522_0n[26]);
  C3 I11 (internal_0n[9], complete522_0n[27], complete522_0n[28], complete522_0n[29]);
  C2 I12 (internal_0n[10], complete522_0n[30], complete522_0n[31]);
  C2 I13 (internal_0n[11], complete522_0n[32], complete522_0n[33]);
  C3 I14 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I15 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I16 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I17 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I18 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I19 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I20 (i_1a, internal_0n[16], internal_0n[17]);
  OR2 I21 (complete522_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I22 (complete522_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I23 (complete522_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I24 (complete522_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I25 (complete522_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I26 (complete522_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I27 (complete522_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I28 (complete522_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I29 (complete522_0n[8], ifint_1n[8], itint_1n[8]);
  OR2 I30 (complete522_0n[9], ifint_1n[9], itint_1n[9]);
  OR2 I31 (complete522_0n[10], ifint_1n[10], itint_1n[10]);
  OR2 I32 (complete522_0n[11], ifint_1n[11], itint_1n[11]);
  OR2 I33 (complete522_0n[12], ifint_1n[12], itint_1n[12]);
  OR2 I34 (complete522_0n[13], ifint_1n[13], itint_1n[13]);
  OR2 I35 (complete522_0n[14], ifint_1n[14], itint_1n[14]);
  OR2 I36 (complete522_0n[15], ifint_1n[15], itint_1n[15]);
  OR2 I37 (complete522_0n[16], ifint_1n[16], itint_1n[16]);
  OR2 I38 (complete522_0n[17], ifint_1n[17], itint_1n[17]);
  OR2 I39 (complete522_0n[18], ifint_1n[18], itint_1n[18]);
  OR2 I40 (complete522_0n[19], ifint_1n[19], itint_1n[19]);
  OR2 I41 (complete522_0n[20], ifint_1n[20], itint_1n[20]);
  OR2 I42 (complete522_0n[21], ifint_1n[21], itint_1n[21]);
  OR2 I43 (complete522_0n[22], ifint_1n[22], itint_1n[22]);
  OR2 I44 (complete522_0n[23], ifint_1n[23], itint_1n[23]);
  OR2 I45 (complete522_0n[24], ifint_1n[24], itint_1n[24]);
  OR2 I46 (complete522_0n[25], ifint_1n[25], itint_1n[25]);
  OR2 I47 (complete522_0n[26], ifint_1n[26], itint_1n[26]);
  OR2 I48 (complete522_0n[27], ifint_1n[27], itint_1n[27]);
  OR2 I49 (complete522_0n[28], ifint_1n[28], itint_1n[28]);
  OR2 I50 (complete522_0n[29], ifint_1n[29], itint_1n[29]);
  OR2 I51 (complete522_0n[30], ifint_1n[30], itint_1n[30]);
  OR2 I52 (complete522_0n[31], ifint_1n[31], itint_1n[31]);
  OR2 I53 (complete522_0n[32], ifint_1n[32], itint_1n[32]);
  OR2 I54 (complete522_0n[33], ifint_1n[33], itint_1n[33]);
  INV I55 (gate521_0n, iaint_1n);
  C2RI I56 (itint_1n[0], i_1r1d[0], gate521_0n, initialise);
  C2RI I57 (itint_1n[1], i_1r1d[1], gate521_0n, initialise);
  C2RI I58 (itint_1n[2], i_1r1d[2], gate521_0n, initialise);
  C2RI I59 (itint_1n[3], i_1r1d[3], gate521_0n, initialise);
  C2RI I60 (itint_1n[4], i_1r1d[4], gate521_0n, initialise);
  C2RI I61 (itint_1n[5], i_1r1d[5], gate521_0n, initialise);
  C2RI I62 (itint_1n[6], i_1r1d[6], gate521_0n, initialise);
  C2RI I63 (itint_1n[7], i_1r1d[7], gate521_0n, initialise);
  C2RI I64 (itint_1n[8], i_1r1d[8], gate521_0n, initialise);
  C2RI I65 (itint_1n[9], i_1r1d[9], gate521_0n, initialise);
  C2RI I66 (itint_1n[10], i_1r1d[10], gate521_0n, initialise);
  C2RI I67 (itint_1n[11], i_1r1d[11], gate521_0n, initialise);
  C2RI I68 (itint_1n[12], i_1r1d[12], gate521_0n, initialise);
  C2RI I69 (itint_1n[13], i_1r1d[13], gate521_0n, initialise);
  C2RI I70 (itint_1n[14], i_1r1d[14], gate521_0n, initialise);
  C2RI I71 (itint_1n[15], i_1r1d[15], gate521_0n, initialise);
  C2RI I72 (itint_1n[16], i_1r1d[16], gate521_0n, initialise);
  C2RI I73 (itint_1n[17], i_1r1d[17], gate521_0n, initialise);
  C2RI I74 (itint_1n[18], i_1r1d[18], gate521_0n, initialise);
  C2RI I75 (itint_1n[19], i_1r1d[19], gate521_0n, initialise);
  C2RI I76 (itint_1n[20], i_1r1d[20], gate521_0n, initialise);
  C2RI I77 (itint_1n[21], i_1r1d[21], gate521_0n, initialise);
  C2RI I78 (itint_1n[22], i_1r1d[22], gate521_0n, initialise);
  C2RI I79 (itint_1n[23], i_1r1d[23], gate521_0n, initialise);
  C2RI I80 (itint_1n[24], i_1r1d[24], gate521_0n, initialise);
  C2RI I81 (itint_1n[25], i_1r1d[25], gate521_0n, initialise);
  C2RI I82 (itint_1n[26], i_1r1d[26], gate521_0n, initialise);
  C2RI I83 (itint_1n[27], i_1r1d[27], gate521_0n, initialise);
  C2RI I84 (itint_1n[28], i_1r1d[28], gate521_0n, initialise);
  C2RI I85 (itint_1n[29], i_1r1d[29], gate521_0n, initialise);
  C2RI I86 (itint_1n[30], i_1r1d[30], gate521_0n, initialise);
  C2RI I87 (itint_1n[31], i_1r1d[31], gate521_0n, initialise);
  C2RI I88 (itint_1n[32], i_1r1d[32], gate521_0n, initialise);
  C2RI I89 (itint_1n[33], i_1r1d[33], gate521_0n, initialise);
  C2RI I90 (ifint_1n[0], i_1r0d[0], gate521_0n, initialise);
  C2RI I91 (ifint_1n[1], i_1r0d[1], gate521_0n, initialise);
  C2RI I92 (ifint_1n[2], i_1r0d[2], gate521_0n, initialise);
  C2RI I93 (ifint_1n[3], i_1r0d[3], gate521_0n, initialise);
  C2RI I94 (ifint_1n[4], i_1r0d[4], gate521_0n, initialise);
  C2RI I95 (ifint_1n[5], i_1r0d[5], gate521_0n, initialise);
  C2RI I96 (ifint_1n[6], i_1r0d[6], gate521_0n, initialise);
  C2RI I97 (ifint_1n[7], i_1r0d[7], gate521_0n, initialise);
  C2RI I98 (ifint_1n[8], i_1r0d[8], gate521_0n, initialise);
  C2RI I99 (ifint_1n[9], i_1r0d[9], gate521_0n, initialise);
  C2RI I100 (ifint_1n[10], i_1r0d[10], gate521_0n, initialise);
  C2RI I101 (ifint_1n[11], i_1r0d[11], gate521_0n, initialise);
  C2RI I102 (ifint_1n[12], i_1r0d[12], gate521_0n, initialise);
  C2RI I103 (ifint_1n[13], i_1r0d[13], gate521_0n, initialise);
  C2RI I104 (ifint_1n[14], i_1r0d[14], gate521_0n, initialise);
  C2RI I105 (ifint_1n[15], i_1r0d[15], gate521_0n, initialise);
  C2RI I106 (ifint_1n[16], i_1r0d[16], gate521_0n, initialise);
  C2RI I107 (ifint_1n[17], i_1r0d[17], gate521_0n, initialise);
  C2RI I108 (ifint_1n[18], i_1r0d[18], gate521_0n, initialise);
  C2RI I109 (ifint_1n[19], i_1r0d[19], gate521_0n, initialise);
  C2RI I110 (ifint_1n[20], i_1r0d[20], gate521_0n, initialise);
  C2RI I111 (ifint_1n[21], i_1r0d[21], gate521_0n, initialise);
  C2RI I112 (ifint_1n[22], i_1r0d[22], gate521_0n, initialise);
  C2RI I113 (ifint_1n[23], i_1r0d[23], gate521_0n, initialise);
  C2RI I114 (ifint_1n[24], i_1r0d[24], gate521_0n, initialise);
  C2RI I115 (ifint_1n[25], i_1r0d[25], gate521_0n, initialise);
  C2RI I116 (ifint_1n[26], i_1r0d[26], gate521_0n, initialise);
  C2RI I117 (ifint_1n[27], i_1r0d[27], gate521_0n, initialise);
  C2RI I118 (ifint_1n[28], i_1r0d[28], gate521_0n, initialise);
  C2RI I119 (ifint_1n[29], i_1r0d[29], gate521_0n, initialise);
  C2RI I120 (ifint_1n[30], i_1r0d[30], gate521_0n, initialise);
  C2RI I121 (ifint_1n[31], i_1r0d[31], gate521_0n, initialise);
  C2RI I122 (ifint_1n[32], i_1r0d[32], gate521_0n, initialise);
  C2RI I123 (ifint_1n[33], i_1r0d[33], gate521_0n, initialise);
  assign i_0a = complete518_0n;
  OR2 I125 (complete518_0n, ifint_0n, itint_0n);
  INV I126 (gate517_0n, iaint_0n);
  C2RI I127 (itint_0n, i_0r1d, gate517_0n, initialise);
  C2RI I128 (ifint_0n, i_0r0d, gate517_0n, initialise);
  C3 I129 (internal_0n[18], complete514_0n[0], complete514_0n[1], complete514_0n[2]);
  C3 I130 (internal_0n[19], complete514_0n[3], complete514_0n[4], complete514_0n[5]);
  C3 I131 (internal_0n[20], complete514_0n[6], complete514_0n[7], complete514_0n[8]);
  C3 I132 (internal_0n[21], complete514_0n[9], complete514_0n[10], complete514_0n[11]);
  C3 I133 (internal_0n[22], complete514_0n[12], complete514_0n[13], complete514_0n[14]);
  C3 I134 (internal_0n[23], complete514_0n[15], complete514_0n[16], complete514_0n[17]);
  C3 I135 (internal_0n[24], complete514_0n[18], complete514_0n[19], complete514_0n[20]);
  C3 I136 (internal_0n[25], complete514_0n[21], complete514_0n[22], complete514_0n[23]);
  C3 I137 (internal_0n[26], complete514_0n[24], complete514_0n[25], complete514_0n[26]);
  C3 I138 (internal_0n[27], complete514_0n[27], complete514_0n[28], complete514_0n[29]);
  C3 I139 (internal_0n[28], complete514_0n[30], complete514_0n[31], complete514_0n[32]);
  C2 I140 (internal_0n[29], complete514_0n[33], complete514_0n[34]);
  C3 I141 (internal_0n[30], internal_0n[18], internal_0n[19], internal_0n[20]);
  C3 I142 (internal_0n[31], internal_0n[21], internal_0n[22], internal_0n[23]);
  C3 I143 (internal_0n[32], internal_0n[24], internal_0n[25], internal_0n[26]);
  C3 I144 (internal_0n[33], internal_0n[27], internal_0n[28], internal_0n[29]);
  C2 I145 (internal_0n[34], internal_0n[30], internal_0n[31]);
  C2 I146 (internal_0n[35], internal_0n[32], internal_0n[33]);
  C2 I147 (oaint_0n, internal_0n[34], internal_0n[35]);
  OR2 I148 (complete514_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I149 (complete514_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I150 (complete514_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I151 (complete514_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I152 (complete514_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I153 (complete514_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I154 (complete514_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I155 (complete514_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I156 (complete514_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I157 (complete514_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I158 (complete514_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I159 (complete514_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I160 (complete514_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I161 (complete514_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I162 (complete514_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I163 (complete514_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I164 (complete514_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I165 (complete514_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I166 (complete514_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I167 (complete514_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I168 (complete514_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I169 (complete514_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I170 (complete514_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I171 (complete514_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I172 (complete514_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I173 (complete514_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I174 (complete514_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I175 (complete514_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I176 (complete514_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I177 (complete514_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I178 (complete514_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I179 (complete514_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I180 (complete514_0n[32], o_0r0d[32], o_0r1d[32]);
  OR2 I181 (complete514_0n[33], o_0r0d[33], o_0r1d[33]);
  OR2 I182 (complete514_0n[34], o_0r0d[34], o_0r1d[34]);
  INV I183 (gate513_0n, o_0a);
  C2RI I184 (o_0r1d[0], otint_0n[0], gate513_0n, initialise);
  C2RI I185 (o_0r1d[1], otint_0n[1], gate513_0n, initialise);
  C2RI I186 (o_0r1d[2], otint_0n[2], gate513_0n, initialise);
  C2RI I187 (o_0r1d[3], otint_0n[3], gate513_0n, initialise);
  C2RI I188 (o_0r1d[4], otint_0n[4], gate513_0n, initialise);
  C2RI I189 (o_0r1d[5], otint_0n[5], gate513_0n, initialise);
  C2RI I190 (o_0r1d[6], otint_0n[6], gate513_0n, initialise);
  C2RI I191 (o_0r1d[7], otint_0n[7], gate513_0n, initialise);
  C2RI I192 (o_0r1d[8], otint_0n[8], gate513_0n, initialise);
  C2RI I193 (o_0r1d[9], otint_0n[9], gate513_0n, initialise);
  C2RI I194 (o_0r1d[10], otint_0n[10], gate513_0n, initialise);
  C2RI I195 (o_0r1d[11], otint_0n[11], gate513_0n, initialise);
  C2RI I196 (o_0r1d[12], otint_0n[12], gate513_0n, initialise);
  C2RI I197 (o_0r1d[13], otint_0n[13], gate513_0n, initialise);
  C2RI I198 (o_0r1d[14], otint_0n[14], gate513_0n, initialise);
  C2RI I199 (o_0r1d[15], otint_0n[15], gate513_0n, initialise);
  C2RI I200 (o_0r1d[16], otint_0n[16], gate513_0n, initialise);
  C2RI I201 (o_0r1d[17], otint_0n[17], gate513_0n, initialise);
  C2RI I202 (o_0r1d[18], otint_0n[18], gate513_0n, initialise);
  C2RI I203 (o_0r1d[19], otint_0n[19], gate513_0n, initialise);
  C2RI I204 (o_0r1d[20], otint_0n[20], gate513_0n, initialise);
  C2RI I205 (o_0r1d[21], otint_0n[21], gate513_0n, initialise);
  C2RI I206 (o_0r1d[22], otint_0n[22], gate513_0n, initialise);
  C2RI I207 (o_0r1d[23], otint_0n[23], gate513_0n, initialise);
  C2RI I208 (o_0r1d[24], otint_0n[24], gate513_0n, initialise);
  C2RI I209 (o_0r1d[25], otint_0n[25], gate513_0n, initialise);
  C2RI I210 (o_0r1d[26], otint_0n[26], gate513_0n, initialise);
  C2RI I211 (o_0r1d[27], otint_0n[27], gate513_0n, initialise);
  C2RI I212 (o_0r1d[28], otint_0n[28], gate513_0n, initialise);
  C2RI I213 (o_0r1d[29], otint_0n[29], gate513_0n, initialise);
  C2RI I214 (o_0r1d[30], otint_0n[30], gate513_0n, initialise);
  C2RI I215 (o_0r1d[31], otint_0n[31], gate513_0n, initialise);
  C2RI I216 (o_0r1d[32], otint_0n[32], gate513_0n, initialise);
  C2RI I217 (o_0r1d[33], otint_0n[33], gate513_0n, initialise);
  C2RI I218 (o_0r1d[34], otint_0n[34], gate513_0n, initialise);
  C2RI I219 (o_0r0d[0], ofint_0n[0], gate513_0n, initialise);
  C2RI I220 (o_0r0d[1], ofint_0n[1], gate513_0n, initialise);
  C2RI I221 (o_0r0d[2], ofint_0n[2], gate513_0n, initialise);
  C2RI I222 (o_0r0d[3], ofint_0n[3], gate513_0n, initialise);
  C2RI I223 (o_0r0d[4], ofint_0n[4], gate513_0n, initialise);
  C2RI I224 (o_0r0d[5], ofint_0n[5], gate513_0n, initialise);
  C2RI I225 (o_0r0d[6], ofint_0n[6], gate513_0n, initialise);
  C2RI I226 (o_0r0d[7], ofint_0n[7], gate513_0n, initialise);
  C2RI I227 (o_0r0d[8], ofint_0n[8], gate513_0n, initialise);
  C2RI I228 (o_0r0d[9], ofint_0n[9], gate513_0n, initialise);
  C2RI I229 (o_0r0d[10], ofint_0n[10], gate513_0n, initialise);
  C2RI I230 (o_0r0d[11], ofint_0n[11], gate513_0n, initialise);
  C2RI I231 (o_0r0d[12], ofint_0n[12], gate513_0n, initialise);
  C2RI I232 (o_0r0d[13], ofint_0n[13], gate513_0n, initialise);
  C2RI I233 (o_0r0d[14], ofint_0n[14], gate513_0n, initialise);
  C2RI I234 (o_0r0d[15], ofint_0n[15], gate513_0n, initialise);
  C2RI I235 (o_0r0d[16], ofint_0n[16], gate513_0n, initialise);
  C2RI I236 (o_0r0d[17], ofint_0n[17], gate513_0n, initialise);
  C2RI I237 (o_0r0d[18], ofint_0n[18], gate513_0n, initialise);
  C2RI I238 (o_0r0d[19], ofint_0n[19], gate513_0n, initialise);
  C2RI I239 (o_0r0d[20], ofint_0n[20], gate513_0n, initialise);
  C2RI I240 (o_0r0d[21], ofint_0n[21], gate513_0n, initialise);
  C2RI I241 (o_0r0d[22], ofint_0n[22], gate513_0n, initialise);
  C2RI I242 (o_0r0d[23], ofint_0n[23], gate513_0n, initialise);
  C2RI I243 (o_0r0d[24], ofint_0n[24], gate513_0n, initialise);
  C2RI I244 (o_0r0d[25], ofint_0n[25], gate513_0n, initialise);
  C2RI I245 (o_0r0d[26], ofint_0n[26], gate513_0n, initialise);
  C2RI I246 (o_0r0d[27], ofint_0n[27], gate513_0n, initialise);
  C2RI I247 (o_0r0d[28], ofint_0n[28], gate513_0n, initialise);
  C2RI I248 (o_0r0d[29], ofint_0n[29], gate513_0n, initialise);
  C2RI I249 (o_0r0d[30], ofint_0n[30], gate513_0n, initialise);
  C2RI I250 (o_0r0d[31], ofint_0n[31], gate513_0n, initialise);
  C2RI I251 (o_0r0d[32], ofint_0n[32], gate513_0n, initialise);
  C2RI I252 (o_0r0d[33], ofint_0n[33], gate513_0n, initialise);
  C2RI I253 (o_0r0d[34], ofint_0n[34], gate513_0n, initialise);
  assign otint_0n[0] = itint_0n;
  assign otint_0n[1] = itint_1n[0];
  assign otint_0n[2] = itint_1n[1];
  assign otint_0n[3] = itint_1n[2];
  assign otint_0n[4] = itint_1n[3];
  assign otint_0n[5] = itint_1n[4];
  assign otint_0n[6] = itint_1n[5];
  assign otint_0n[7] = itint_1n[6];
  assign otint_0n[8] = itint_1n[7];
  assign otint_0n[9] = itint_1n[8];
  assign otint_0n[10] = itint_1n[9];
  assign otint_0n[11] = itint_1n[10];
  assign otint_0n[12] = itint_1n[11];
  assign otint_0n[13] = itint_1n[12];
  assign otint_0n[14] = itint_1n[13];
  assign otint_0n[15] = itint_1n[14];
  assign otint_0n[16] = itint_1n[15];
  assign otint_0n[17] = itint_1n[16];
  assign otint_0n[18] = itint_1n[17];
  assign otint_0n[19] = itint_1n[18];
  assign otint_0n[20] = itint_1n[19];
  assign otint_0n[21] = itint_1n[20];
  assign otint_0n[22] = itint_1n[21];
  assign otint_0n[23] = itint_1n[22];
  assign otint_0n[24] = itint_1n[23];
  assign otint_0n[25] = itint_1n[24];
  assign otint_0n[26] = itint_1n[25];
  assign otint_0n[27] = itint_1n[26];
  assign otint_0n[28] = itint_1n[27];
  assign otint_0n[29] = itint_1n[28];
  assign otint_0n[30] = itint_1n[29];
  assign otint_0n[31] = itint_1n[30];
  assign otint_0n[32] = itint_1n[31];
  assign otint_0n[33] = itint_1n[32];
  assign otint_0n[34] = itint_1n[33];
  assign ofint_0n[0] = ifint_0n;
  assign ofint_0n[1] = ifint_1n[0];
  assign ofint_0n[2] = ifint_1n[1];
  assign ofint_0n[3] = ifint_1n[2];
  assign ofint_0n[4] = ifint_1n[3];
  assign ofint_0n[5] = ifint_1n[4];
  assign ofint_0n[6] = ifint_1n[5];
  assign ofint_0n[7] = ifint_1n[6];
  assign ofint_0n[8] = ifint_1n[7];
  assign ofint_0n[9] = ifint_1n[8];
  assign ofint_0n[10] = ifint_1n[9];
  assign ofint_0n[11] = ifint_1n[10];
  assign ofint_0n[12] = ifint_1n[11];
  assign ofint_0n[13] = ifint_1n[12];
  assign ofint_0n[14] = ifint_1n[13];
  assign ofint_0n[15] = ifint_1n[14];
  assign ofint_0n[16] = ifint_1n[15];
  assign ofint_0n[17] = ifint_1n[16];
  assign ofint_0n[18] = ifint_1n[17];
  assign ofint_0n[19] = ifint_1n[18];
  assign ofint_0n[20] = ifint_1n[19];
  assign ofint_0n[21] = ifint_1n[20];
  assign ofint_0n[22] = ifint_1n[21];
  assign ofint_0n[23] = ifint_1n[22];
  assign ofint_0n[24] = ifint_1n[23];
  assign ofint_0n[25] = ifint_1n[24];
  assign ofint_0n[26] = ifint_1n[25];
  assign ofint_0n[27] = ifint_1n[26];
  assign ofint_0n[28] = ifint_1n[27];
  assign ofint_0n[29] = ifint_1n[28];
  assign ofint_0n[30] = ifint_1n[29];
  assign ofint_0n[31] = ifint_1n[30];
  assign ofint_0n[32] = ifint_1n[31];
  assign ofint_0n[33] = ifint_1n[32];
  assign ofint_0n[34] = ifint_1n[33];
endmodule

module BrzJ_l12__282_2033_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [1:0] i_0r0d;
  input [1:0] i_0r1d;
  output i_0a;
  input [32:0] i_1r0d;
  input [32:0] i_1r1d;
  output i_1a;
  output [34:0] o_0r0d;
  output [34:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [34:0] internal_0n;
  wire [34:0] ofint_0n;
  wire [34:0] otint_0n;
  wire oaint_0n;
  wire [1:0] ifint_0n;
  wire [32:0] ifint_1n;
  wire [1:0] itint_0n;
  wire [32:0] itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [32:0] complete534_0n;
  wire gate533_0n;
  wire [1:0] complete530_0n;
  wire gate529_0n;
  wire [34:0] complete526_0n;
  wire gate525_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  C3 I2 (internal_0n[0], complete534_0n[0], complete534_0n[1], complete534_0n[2]);
  C3 I3 (internal_0n[1], complete534_0n[3], complete534_0n[4], complete534_0n[5]);
  C3 I4 (internal_0n[2], complete534_0n[6], complete534_0n[7], complete534_0n[8]);
  C3 I5 (internal_0n[3], complete534_0n[9], complete534_0n[10], complete534_0n[11]);
  C3 I6 (internal_0n[4], complete534_0n[12], complete534_0n[13], complete534_0n[14]);
  C3 I7 (internal_0n[5], complete534_0n[15], complete534_0n[16], complete534_0n[17]);
  C3 I8 (internal_0n[6], complete534_0n[18], complete534_0n[19], complete534_0n[20]);
  C3 I9 (internal_0n[7], complete534_0n[21], complete534_0n[22], complete534_0n[23]);
  C3 I10 (internal_0n[8], complete534_0n[24], complete534_0n[25], complete534_0n[26]);
  C3 I11 (internal_0n[9], complete534_0n[27], complete534_0n[28], complete534_0n[29]);
  C3 I12 (internal_0n[10], complete534_0n[30], complete534_0n[31], complete534_0n[32]);
  C3 I13 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I14 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I15 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I16 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I17 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I18 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I19 (i_1a, internal_0n[15], internal_0n[16]);
  OR2 I20 (complete534_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I21 (complete534_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I22 (complete534_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I23 (complete534_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I24 (complete534_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I25 (complete534_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I26 (complete534_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I27 (complete534_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I28 (complete534_0n[8], ifint_1n[8], itint_1n[8]);
  OR2 I29 (complete534_0n[9], ifint_1n[9], itint_1n[9]);
  OR2 I30 (complete534_0n[10], ifint_1n[10], itint_1n[10]);
  OR2 I31 (complete534_0n[11], ifint_1n[11], itint_1n[11]);
  OR2 I32 (complete534_0n[12], ifint_1n[12], itint_1n[12]);
  OR2 I33 (complete534_0n[13], ifint_1n[13], itint_1n[13]);
  OR2 I34 (complete534_0n[14], ifint_1n[14], itint_1n[14]);
  OR2 I35 (complete534_0n[15], ifint_1n[15], itint_1n[15]);
  OR2 I36 (complete534_0n[16], ifint_1n[16], itint_1n[16]);
  OR2 I37 (complete534_0n[17], ifint_1n[17], itint_1n[17]);
  OR2 I38 (complete534_0n[18], ifint_1n[18], itint_1n[18]);
  OR2 I39 (complete534_0n[19], ifint_1n[19], itint_1n[19]);
  OR2 I40 (complete534_0n[20], ifint_1n[20], itint_1n[20]);
  OR2 I41 (complete534_0n[21], ifint_1n[21], itint_1n[21]);
  OR2 I42 (complete534_0n[22], ifint_1n[22], itint_1n[22]);
  OR2 I43 (complete534_0n[23], ifint_1n[23], itint_1n[23]);
  OR2 I44 (complete534_0n[24], ifint_1n[24], itint_1n[24]);
  OR2 I45 (complete534_0n[25], ifint_1n[25], itint_1n[25]);
  OR2 I46 (complete534_0n[26], ifint_1n[26], itint_1n[26]);
  OR2 I47 (complete534_0n[27], ifint_1n[27], itint_1n[27]);
  OR2 I48 (complete534_0n[28], ifint_1n[28], itint_1n[28]);
  OR2 I49 (complete534_0n[29], ifint_1n[29], itint_1n[29]);
  OR2 I50 (complete534_0n[30], ifint_1n[30], itint_1n[30]);
  OR2 I51 (complete534_0n[31], ifint_1n[31], itint_1n[31]);
  OR2 I52 (complete534_0n[32], ifint_1n[32], itint_1n[32]);
  INV I53 (gate533_0n, iaint_1n);
  C2RI I54 (itint_1n[0], i_1r1d[0], gate533_0n, initialise);
  C2RI I55 (itint_1n[1], i_1r1d[1], gate533_0n, initialise);
  C2RI I56 (itint_1n[2], i_1r1d[2], gate533_0n, initialise);
  C2RI I57 (itint_1n[3], i_1r1d[3], gate533_0n, initialise);
  C2RI I58 (itint_1n[4], i_1r1d[4], gate533_0n, initialise);
  C2RI I59 (itint_1n[5], i_1r1d[5], gate533_0n, initialise);
  C2RI I60 (itint_1n[6], i_1r1d[6], gate533_0n, initialise);
  C2RI I61 (itint_1n[7], i_1r1d[7], gate533_0n, initialise);
  C2RI I62 (itint_1n[8], i_1r1d[8], gate533_0n, initialise);
  C2RI I63 (itint_1n[9], i_1r1d[9], gate533_0n, initialise);
  C2RI I64 (itint_1n[10], i_1r1d[10], gate533_0n, initialise);
  C2RI I65 (itint_1n[11], i_1r1d[11], gate533_0n, initialise);
  C2RI I66 (itint_1n[12], i_1r1d[12], gate533_0n, initialise);
  C2RI I67 (itint_1n[13], i_1r1d[13], gate533_0n, initialise);
  C2RI I68 (itint_1n[14], i_1r1d[14], gate533_0n, initialise);
  C2RI I69 (itint_1n[15], i_1r1d[15], gate533_0n, initialise);
  C2RI I70 (itint_1n[16], i_1r1d[16], gate533_0n, initialise);
  C2RI I71 (itint_1n[17], i_1r1d[17], gate533_0n, initialise);
  C2RI I72 (itint_1n[18], i_1r1d[18], gate533_0n, initialise);
  C2RI I73 (itint_1n[19], i_1r1d[19], gate533_0n, initialise);
  C2RI I74 (itint_1n[20], i_1r1d[20], gate533_0n, initialise);
  C2RI I75 (itint_1n[21], i_1r1d[21], gate533_0n, initialise);
  C2RI I76 (itint_1n[22], i_1r1d[22], gate533_0n, initialise);
  C2RI I77 (itint_1n[23], i_1r1d[23], gate533_0n, initialise);
  C2RI I78 (itint_1n[24], i_1r1d[24], gate533_0n, initialise);
  C2RI I79 (itint_1n[25], i_1r1d[25], gate533_0n, initialise);
  C2RI I80 (itint_1n[26], i_1r1d[26], gate533_0n, initialise);
  C2RI I81 (itint_1n[27], i_1r1d[27], gate533_0n, initialise);
  C2RI I82 (itint_1n[28], i_1r1d[28], gate533_0n, initialise);
  C2RI I83 (itint_1n[29], i_1r1d[29], gate533_0n, initialise);
  C2RI I84 (itint_1n[30], i_1r1d[30], gate533_0n, initialise);
  C2RI I85 (itint_1n[31], i_1r1d[31], gate533_0n, initialise);
  C2RI I86 (itint_1n[32], i_1r1d[32], gate533_0n, initialise);
  C2RI I87 (ifint_1n[0], i_1r0d[0], gate533_0n, initialise);
  C2RI I88 (ifint_1n[1], i_1r0d[1], gate533_0n, initialise);
  C2RI I89 (ifint_1n[2], i_1r0d[2], gate533_0n, initialise);
  C2RI I90 (ifint_1n[3], i_1r0d[3], gate533_0n, initialise);
  C2RI I91 (ifint_1n[4], i_1r0d[4], gate533_0n, initialise);
  C2RI I92 (ifint_1n[5], i_1r0d[5], gate533_0n, initialise);
  C2RI I93 (ifint_1n[6], i_1r0d[6], gate533_0n, initialise);
  C2RI I94 (ifint_1n[7], i_1r0d[7], gate533_0n, initialise);
  C2RI I95 (ifint_1n[8], i_1r0d[8], gate533_0n, initialise);
  C2RI I96 (ifint_1n[9], i_1r0d[9], gate533_0n, initialise);
  C2RI I97 (ifint_1n[10], i_1r0d[10], gate533_0n, initialise);
  C2RI I98 (ifint_1n[11], i_1r0d[11], gate533_0n, initialise);
  C2RI I99 (ifint_1n[12], i_1r0d[12], gate533_0n, initialise);
  C2RI I100 (ifint_1n[13], i_1r0d[13], gate533_0n, initialise);
  C2RI I101 (ifint_1n[14], i_1r0d[14], gate533_0n, initialise);
  C2RI I102 (ifint_1n[15], i_1r0d[15], gate533_0n, initialise);
  C2RI I103 (ifint_1n[16], i_1r0d[16], gate533_0n, initialise);
  C2RI I104 (ifint_1n[17], i_1r0d[17], gate533_0n, initialise);
  C2RI I105 (ifint_1n[18], i_1r0d[18], gate533_0n, initialise);
  C2RI I106 (ifint_1n[19], i_1r0d[19], gate533_0n, initialise);
  C2RI I107 (ifint_1n[20], i_1r0d[20], gate533_0n, initialise);
  C2RI I108 (ifint_1n[21], i_1r0d[21], gate533_0n, initialise);
  C2RI I109 (ifint_1n[22], i_1r0d[22], gate533_0n, initialise);
  C2RI I110 (ifint_1n[23], i_1r0d[23], gate533_0n, initialise);
  C2RI I111 (ifint_1n[24], i_1r0d[24], gate533_0n, initialise);
  C2RI I112 (ifint_1n[25], i_1r0d[25], gate533_0n, initialise);
  C2RI I113 (ifint_1n[26], i_1r0d[26], gate533_0n, initialise);
  C2RI I114 (ifint_1n[27], i_1r0d[27], gate533_0n, initialise);
  C2RI I115 (ifint_1n[28], i_1r0d[28], gate533_0n, initialise);
  C2RI I116 (ifint_1n[29], i_1r0d[29], gate533_0n, initialise);
  C2RI I117 (ifint_1n[30], i_1r0d[30], gate533_0n, initialise);
  C2RI I118 (ifint_1n[31], i_1r0d[31], gate533_0n, initialise);
  C2RI I119 (ifint_1n[32], i_1r0d[32], gate533_0n, initialise);
  C2 I120 (i_0a, complete530_0n[0], complete530_0n[1]);
  OR2 I121 (complete530_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I122 (complete530_0n[1], ifint_0n[1], itint_0n[1]);
  INV I123 (gate529_0n, iaint_0n);
  C2RI I124 (itint_0n[0], i_0r1d[0], gate529_0n, initialise);
  C2RI I125 (itint_0n[1], i_0r1d[1], gate529_0n, initialise);
  C2RI I126 (ifint_0n[0], i_0r0d[0], gate529_0n, initialise);
  C2RI I127 (ifint_0n[1], i_0r0d[1], gate529_0n, initialise);
  C3 I128 (internal_0n[17], complete526_0n[0], complete526_0n[1], complete526_0n[2]);
  C3 I129 (internal_0n[18], complete526_0n[3], complete526_0n[4], complete526_0n[5]);
  C3 I130 (internal_0n[19], complete526_0n[6], complete526_0n[7], complete526_0n[8]);
  C3 I131 (internal_0n[20], complete526_0n[9], complete526_0n[10], complete526_0n[11]);
  C3 I132 (internal_0n[21], complete526_0n[12], complete526_0n[13], complete526_0n[14]);
  C3 I133 (internal_0n[22], complete526_0n[15], complete526_0n[16], complete526_0n[17]);
  C3 I134 (internal_0n[23], complete526_0n[18], complete526_0n[19], complete526_0n[20]);
  C3 I135 (internal_0n[24], complete526_0n[21], complete526_0n[22], complete526_0n[23]);
  C3 I136 (internal_0n[25], complete526_0n[24], complete526_0n[25], complete526_0n[26]);
  C3 I137 (internal_0n[26], complete526_0n[27], complete526_0n[28], complete526_0n[29]);
  C3 I138 (internal_0n[27], complete526_0n[30], complete526_0n[31], complete526_0n[32]);
  C2 I139 (internal_0n[28], complete526_0n[33], complete526_0n[34]);
  C3 I140 (internal_0n[29], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I141 (internal_0n[30], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I142 (internal_0n[31], internal_0n[23], internal_0n[24], internal_0n[25]);
  C3 I143 (internal_0n[32], internal_0n[26], internal_0n[27], internal_0n[28]);
  C2 I144 (internal_0n[33], internal_0n[29], internal_0n[30]);
  C2 I145 (internal_0n[34], internal_0n[31], internal_0n[32]);
  C2 I146 (oaint_0n, internal_0n[33], internal_0n[34]);
  OR2 I147 (complete526_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I148 (complete526_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I149 (complete526_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I150 (complete526_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I151 (complete526_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I152 (complete526_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I153 (complete526_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I154 (complete526_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I155 (complete526_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I156 (complete526_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I157 (complete526_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I158 (complete526_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I159 (complete526_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I160 (complete526_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I161 (complete526_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I162 (complete526_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I163 (complete526_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I164 (complete526_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I165 (complete526_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I166 (complete526_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I167 (complete526_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I168 (complete526_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I169 (complete526_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I170 (complete526_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I171 (complete526_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I172 (complete526_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I173 (complete526_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I174 (complete526_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I175 (complete526_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I176 (complete526_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I177 (complete526_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I178 (complete526_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I179 (complete526_0n[32], o_0r0d[32], o_0r1d[32]);
  OR2 I180 (complete526_0n[33], o_0r0d[33], o_0r1d[33]);
  OR2 I181 (complete526_0n[34], o_0r0d[34], o_0r1d[34]);
  INV I182 (gate525_0n, o_0a);
  C2RI I183 (o_0r1d[0], otint_0n[0], gate525_0n, initialise);
  C2RI I184 (o_0r1d[1], otint_0n[1], gate525_0n, initialise);
  C2RI I185 (o_0r1d[2], otint_0n[2], gate525_0n, initialise);
  C2RI I186 (o_0r1d[3], otint_0n[3], gate525_0n, initialise);
  C2RI I187 (o_0r1d[4], otint_0n[4], gate525_0n, initialise);
  C2RI I188 (o_0r1d[5], otint_0n[5], gate525_0n, initialise);
  C2RI I189 (o_0r1d[6], otint_0n[6], gate525_0n, initialise);
  C2RI I190 (o_0r1d[7], otint_0n[7], gate525_0n, initialise);
  C2RI I191 (o_0r1d[8], otint_0n[8], gate525_0n, initialise);
  C2RI I192 (o_0r1d[9], otint_0n[9], gate525_0n, initialise);
  C2RI I193 (o_0r1d[10], otint_0n[10], gate525_0n, initialise);
  C2RI I194 (o_0r1d[11], otint_0n[11], gate525_0n, initialise);
  C2RI I195 (o_0r1d[12], otint_0n[12], gate525_0n, initialise);
  C2RI I196 (o_0r1d[13], otint_0n[13], gate525_0n, initialise);
  C2RI I197 (o_0r1d[14], otint_0n[14], gate525_0n, initialise);
  C2RI I198 (o_0r1d[15], otint_0n[15], gate525_0n, initialise);
  C2RI I199 (o_0r1d[16], otint_0n[16], gate525_0n, initialise);
  C2RI I200 (o_0r1d[17], otint_0n[17], gate525_0n, initialise);
  C2RI I201 (o_0r1d[18], otint_0n[18], gate525_0n, initialise);
  C2RI I202 (o_0r1d[19], otint_0n[19], gate525_0n, initialise);
  C2RI I203 (o_0r1d[20], otint_0n[20], gate525_0n, initialise);
  C2RI I204 (o_0r1d[21], otint_0n[21], gate525_0n, initialise);
  C2RI I205 (o_0r1d[22], otint_0n[22], gate525_0n, initialise);
  C2RI I206 (o_0r1d[23], otint_0n[23], gate525_0n, initialise);
  C2RI I207 (o_0r1d[24], otint_0n[24], gate525_0n, initialise);
  C2RI I208 (o_0r1d[25], otint_0n[25], gate525_0n, initialise);
  C2RI I209 (o_0r1d[26], otint_0n[26], gate525_0n, initialise);
  C2RI I210 (o_0r1d[27], otint_0n[27], gate525_0n, initialise);
  C2RI I211 (o_0r1d[28], otint_0n[28], gate525_0n, initialise);
  C2RI I212 (o_0r1d[29], otint_0n[29], gate525_0n, initialise);
  C2RI I213 (o_0r1d[30], otint_0n[30], gate525_0n, initialise);
  C2RI I214 (o_0r1d[31], otint_0n[31], gate525_0n, initialise);
  C2RI I215 (o_0r1d[32], otint_0n[32], gate525_0n, initialise);
  C2RI I216 (o_0r1d[33], otint_0n[33], gate525_0n, initialise);
  C2RI I217 (o_0r1d[34], otint_0n[34], gate525_0n, initialise);
  C2RI I218 (o_0r0d[0], ofint_0n[0], gate525_0n, initialise);
  C2RI I219 (o_0r0d[1], ofint_0n[1], gate525_0n, initialise);
  C2RI I220 (o_0r0d[2], ofint_0n[2], gate525_0n, initialise);
  C2RI I221 (o_0r0d[3], ofint_0n[3], gate525_0n, initialise);
  C2RI I222 (o_0r0d[4], ofint_0n[4], gate525_0n, initialise);
  C2RI I223 (o_0r0d[5], ofint_0n[5], gate525_0n, initialise);
  C2RI I224 (o_0r0d[6], ofint_0n[6], gate525_0n, initialise);
  C2RI I225 (o_0r0d[7], ofint_0n[7], gate525_0n, initialise);
  C2RI I226 (o_0r0d[8], ofint_0n[8], gate525_0n, initialise);
  C2RI I227 (o_0r0d[9], ofint_0n[9], gate525_0n, initialise);
  C2RI I228 (o_0r0d[10], ofint_0n[10], gate525_0n, initialise);
  C2RI I229 (o_0r0d[11], ofint_0n[11], gate525_0n, initialise);
  C2RI I230 (o_0r0d[12], ofint_0n[12], gate525_0n, initialise);
  C2RI I231 (o_0r0d[13], ofint_0n[13], gate525_0n, initialise);
  C2RI I232 (o_0r0d[14], ofint_0n[14], gate525_0n, initialise);
  C2RI I233 (o_0r0d[15], ofint_0n[15], gate525_0n, initialise);
  C2RI I234 (o_0r0d[16], ofint_0n[16], gate525_0n, initialise);
  C2RI I235 (o_0r0d[17], ofint_0n[17], gate525_0n, initialise);
  C2RI I236 (o_0r0d[18], ofint_0n[18], gate525_0n, initialise);
  C2RI I237 (o_0r0d[19], ofint_0n[19], gate525_0n, initialise);
  C2RI I238 (o_0r0d[20], ofint_0n[20], gate525_0n, initialise);
  C2RI I239 (o_0r0d[21], ofint_0n[21], gate525_0n, initialise);
  C2RI I240 (o_0r0d[22], ofint_0n[22], gate525_0n, initialise);
  C2RI I241 (o_0r0d[23], ofint_0n[23], gate525_0n, initialise);
  C2RI I242 (o_0r0d[24], ofint_0n[24], gate525_0n, initialise);
  C2RI I243 (o_0r0d[25], ofint_0n[25], gate525_0n, initialise);
  C2RI I244 (o_0r0d[26], ofint_0n[26], gate525_0n, initialise);
  C2RI I245 (o_0r0d[27], ofint_0n[27], gate525_0n, initialise);
  C2RI I246 (o_0r0d[28], ofint_0n[28], gate525_0n, initialise);
  C2RI I247 (o_0r0d[29], ofint_0n[29], gate525_0n, initialise);
  C2RI I248 (o_0r0d[30], ofint_0n[30], gate525_0n, initialise);
  C2RI I249 (o_0r0d[31], ofint_0n[31], gate525_0n, initialise);
  C2RI I250 (o_0r0d[32], ofint_0n[32], gate525_0n, initialise);
  C2RI I251 (o_0r0d[33], ofint_0n[33], gate525_0n, initialise);
  C2RI I252 (o_0r0d[34], ofint_0n[34], gate525_0n, initialise);
  assign otint_0n[0] = itint_0n[0];
  assign otint_0n[1] = itint_0n[1];
  assign otint_0n[2] = itint_1n[0];
  assign otint_0n[3] = itint_1n[1];
  assign otint_0n[4] = itint_1n[2];
  assign otint_0n[5] = itint_1n[3];
  assign otint_0n[6] = itint_1n[4];
  assign otint_0n[7] = itint_1n[5];
  assign otint_0n[8] = itint_1n[6];
  assign otint_0n[9] = itint_1n[7];
  assign otint_0n[10] = itint_1n[8];
  assign otint_0n[11] = itint_1n[9];
  assign otint_0n[12] = itint_1n[10];
  assign otint_0n[13] = itint_1n[11];
  assign otint_0n[14] = itint_1n[12];
  assign otint_0n[15] = itint_1n[13];
  assign otint_0n[16] = itint_1n[14];
  assign otint_0n[17] = itint_1n[15];
  assign otint_0n[18] = itint_1n[16];
  assign otint_0n[19] = itint_1n[17];
  assign otint_0n[20] = itint_1n[18];
  assign otint_0n[21] = itint_1n[19];
  assign otint_0n[22] = itint_1n[20];
  assign otint_0n[23] = itint_1n[21];
  assign otint_0n[24] = itint_1n[22];
  assign otint_0n[25] = itint_1n[23];
  assign otint_0n[26] = itint_1n[24];
  assign otint_0n[27] = itint_1n[25];
  assign otint_0n[28] = itint_1n[26];
  assign otint_0n[29] = itint_1n[27];
  assign otint_0n[30] = itint_1n[28];
  assign otint_0n[31] = itint_1n[29];
  assign otint_0n[32] = itint_1n[30];
  assign otint_0n[33] = itint_1n[31];
  assign otint_0n[34] = itint_1n[32];
  assign ofint_0n[0] = ifint_0n[0];
  assign ofint_0n[1] = ifint_0n[1];
  assign ofint_0n[2] = ifint_1n[0];
  assign ofint_0n[3] = ifint_1n[1];
  assign ofint_0n[4] = ifint_1n[2];
  assign ofint_0n[5] = ifint_1n[3];
  assign ofint_0n[6] = ifint_1n[4];
  assign ofint_0n[7] = ifint_1n[5];
  assign ofint_0n[8] = ifint_1n[6];
  assign ofint_0n[9] = ifint_1n[7];
  assign ofint_0n[10] = ifint_1n[8];
  assign ofint_0n[11] = ifint_1n[9];
  assign ofint_0n[12] = ifint_1n[10];
  assign ofint_0n[13] = ifint_1n[11];
  assign ofint_0n[14] = ifint_1n[12];
  assign ofint_0n[15] = ifint_1n[13];
  assign ofint_0n[16] = ifint_1n[14];
  assign ofint_0n[17] = ifint_1n[15];
  assign ofint_0n[18] = ifint_1n[16];
  assign ofint_0n[19] = ifint_1n[17];
  assign ofint_0n[20] = ifint_1n[18];
  assign ofint_0n[21] = ifint_1n[19];
  assign ofint_0n[22] = ifint_1n[20];
  assign ofint_0n[23] = ifint_1n[21];
  assign ofint_0n[24] = ifint_1n[22];
  assign ofint_0n[25] = ifint_1n[23];
  assign ofint_0n[26] = ifint_1n[24];
  assign ofint_0n[27] = ifint_1n[25];
  assign ofint_0n[28] = ifint_1n[26];
  assign ofint_0n[29] = ifint_1n[27];
  assign ofint_0n[30] = ifint_1n[28];
  assign ofint_0n[31] = ifint_1n[29];
  assign ofint_0n[32] = ifint_1n[30];
  assign ofint_0n[33] = ifint_1n[31];
  assign ofint_0n[34] = ifint_1n[32];
endmodule

module BrzJ_l11__283_200_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [2:0] i_0r0d;
  input [2:0] i_0r1d;
  output i_0a;
  input i_1r;
  output i_1a;
  output [2:0] o_0r0d;
  output [2:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [2:0] ofint_0n;
  wire [2:0] otint_0n;
  wire oaint_0n;
  wire [2:0] ifint_0n;
  wire ifint_1n;
  wire [2:0] itint_0n;
  wire iaint_0n;
  wire iaint_1n;
  wire gate545_0n;
  wire [2:0] complete542_0n;
  wire gate541_0n;
  wire [2:0] complete538_0n;
  wire gate537_0n;
  wire [2:0] joint_0n;
  wire [2:0] joinf_0n;
  wire icomplete_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign i_1a = ifint_1n;
  INV I3 (gate545_0n, iaint_1n);
  C2RI I4 (ifint_1n, i_1r, gate545_0n, initialise);
  C3 I5 (i_0a, complete542_0n[0], complete542_0n[1], complete542_0n[2]);
  OR2 I6 (complete542_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I7 (complete542_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I8 (complete542_0n[2], ifint_0n[2], itint_0n[2]);
  INV I9 (gate541_0n, iaint_0n);
  C2RI I10 (itint_0n[0], i_0r1d[0], gate541_0n, initialise);
  C2RI I11 (itint_0n[1], i_0r1d[1], gate541_0n, initialise);
  C2RI I12 (itint_0n[2], i_0r1d[2], gate541_0n, initialise);
  C2RI I13 (ifint_0n[0], i_0r0d[0], gate541_0n, initialise);
  C2RI I14 (ifint_0n[1], i_0r0d[1], gate541_0n, initialise);
  C2RI I15 (ifint_0n[2], i_0r0d[2], gate541_0n, initialise);
  C3 I16 (oaint_0n, complete538_0n[0], complete538_0n[1], complete538_0n[2]);
  OR2 I17 (complete538_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I18 (complete538_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I19 (complete538_0n[2], o_0r0d[2], o_0r1d[2]);
  INV I20 (gate537_0n, o_0a);
  C2RI I21 (o_0r1d[0], otint_0n[0], gate537_0n, initialise);
  C2RI I22 (o_0r1d[1], otint_0n[1], gate537_0n, initialise);
  C2RI I23 (o_0r1d[2], otint_0n[2], gate537_0n, initialise);
  C2RI I24 (o_0r0d[0], ofint_0n[0], gate537_0n, initialise);
  C2RI I25 (o_0r0d[1], ofint_0n[1], gate537_0n, initialise);
  C2RI I26 (o_0r0d[2], ofint_0n[2], gate537_0n, initialise);
  assign otint_0n[1] = joint_0n[1];
  assign otint_0n[2] = joint_0n[2];
  assign ofint_0n[1] = joinf_0n[1];
  assign ofint_0n[2] = joinf_0n[2];
  C2 I31 (otint_0n[0], joint_0n[0], icomplete_0n);
  C2 I32 (ofint_0n[0], joinf_0n[0], icomplete_0n);
  assign icomplete_0n = ifint_1n;
  assign joint_0n[0] = itint_0n[0];
  assign joint_0n[1] = itint_0n[1];
  assign joint_0n[2] = itint_0n[2];
  assign joinf_0n[0] = ifint_0n[0];
  assign joinf_0n[1] = ifint_0n[1];
  assign joinf_0n[2] = ifint_0n[2];
endmodule

module BrzJ_l12__2832_200_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [31:0] i_0r0d;
  input [31:0] i_0r1d;
  output i_0a;
  input i_1r;
  output i_1a;
  output [31:0] o_0r0d;
  output [31:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [33:0] internal_0n;
  wire [31:0] ofint_0n;
  wire [31:0] otint_0n;
  wire oaint_0n;
  wire [31:0] ifint_0n;
  wire ifint_1n;
  wire [31:0] itint_0n;
  wire iaint_0n;
  wire iaint_1n;
  wire gate556_0n;
  wire [31:0] complete553_0n;
  wire gate552_0n;
  wire [31:0] complete549_0n;
  wire gate548_0n;
  wire [31:0] joint_0n;
  wire [31:0] joinf_0n;
  wire icomplete_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign i_1a = ifint_1n;
  INV I3 (gate556_0n, iaint_1n);
  C2RI I4 (ifint_1n, i_1r, gate556_0n, initialise);
  C3 I5 (internal_0n[0], complete553_0n[0], complete553_0n[1], complete553_0n[2]);
  C3 I6 (internal_0n[1], complete553_0n[3], complete553_0n[4], complete553_0n[5]);
  C3 I7 (internal_0n[2], complete553_0n[6], complete553_0n[7], complete553_0n[8]);
  C3 I8 (internal_0n[3], complete553_0n[9], complete553_0n[10], complete553_0n[11]);
  C3 I9 (internal_0n[4], complete553_0n[12], complete553_0n[13], complete553_0n[14]);
  C3 I10 (internal_0n[5], complete553_0n[15], complete553_0n[16], complete553_0n[17]);
  C3 I11 (internal_0n[6], complete553_0n[18], complete553_0n[19], complete553_0n[20]);
  C3 I12 (internal_0n[7], complete553_0n[21], complete553_0n[22], complete553_0n[23]);
  C3 I13 (internal_0n[8], complete553_0n[24], complete553_0n[25], complete553_0n[26]);
  C3 I14 (internal_0n[9], complete553_0n[27], complete553_0n[28], complete553_0n[29]);
  C2 I15 (internal_0n[10], complete553_0n[30], complete553_0n[31]);
  C3 I16 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I17 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I18 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I19 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I20 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I21 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I22 (i_0a, internal_0n[15], internal_0n[16]);
  OR2 I23 (complete553_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I24 (complete553_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I25 (complete553_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I26 (complete553_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I27 (complete553_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I28 (complete553_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I29 (complete553_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I30 (complete553_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I31 (complete553_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I32 (complete553_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I33 (complete553_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I34 (complete553_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I35 (complete553_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I36 (complete553_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I37 (complete553_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I38 (complete553_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I39 (complete553_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I40 (complete553_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I41 (complete553_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I42 (complete553_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I43 (complete553_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I44 (complete553_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I45 (complete553_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I46 (complete553_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I47 (complete553_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I48 (complete553_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I49 (complete553_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I50 (complete553_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I51 (complete553_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I52 (complete553_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I53 (complete553_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I54 (complete553_0n[31], ifint_0n[31], itint_0n[31]);
  INV I55 (gate552_0n, iaint_0n);
  C2RI I56 (itint_0n[0], i_0r1d[0], gate552_0n, initialise);
  C2RI I57 (itint_0n[1], i_0r1d[1], gate552_0n, initialise);
  C2RI I58 (itint_0n[2], i_0r1d[2], gate552_0n, initialise);
  C2RI I59 (itint_0n[3], i_0r1d[3], gate552_0n, initialise);
  C2RI I60 (itint_0n[4], i_0r1d[4], gate552_0n, initialise);
  C2RI I61 (itint_0n[5], i_0r1d[5], gate552_0n, initialise);
  C2RI I62 (itint_0n[6], i_0r1d[6], gate552_0n, initialise);
  C2RI I63 (itint_0n[7], i_0r1d[7], gate552_0n, initialise);
  C2RI I64 (itint_0n[8], i_0r1d[8], gate552_0n, initialise);
  C2RI I65 (itint_0n[9], i_0r1d[9], gate552_0n, initialise);
  C2RI I66 (itint_0n[10], i_0r1d[10], gate552_0n, initialise);
  C2RI I67 (itint_0n[11], i_0r1d[11], gate552_0n, initialise);
  C2RI I68 (itint_0n[12], i_0r1d[12], gate552_0n, initialise);
  C2RI I69 (itint_0n[13], i_0r1d[13], gate552_0n, initialise);
  C2RI I70 (itint_0n[14], i_0r1d[14], gate552_0n, initialise);
  C2RI I71 (itint_0n[15], i_0r1d[15], gate552_0n, initialise);
  C2RI I72 (itint_0n[16], i_0r1d[16], gate552_0n, initialise);
  C2RI I73 (itint_0n[17], i_0r1d[17], gate552_0n, initialise);
  C2RI I74 (itint_0n[18], i_0r1d[18], gate552_0n, initialise);
  C2RI I75 (itint_0n[19], i_0r1d[19], gate552_0n, initialise);
  C2RI I76 (itint_0n[20], i_0r1d[20], gate552_0n, initialise);
  C2RI I77 (itint_0n[21], i_0r1d[21], gate552_0n, initialise);
  C2RI I78 (itint_0n[22], i_0r1d[22], gate552_0n, initialise);
  C2RI I79 (itint_0n[23], i_0r1d[23], gate552_0n, initialise);
  C2RI I80 (itint_0n[24], i_0r1d[24], gate552_0n, initialise);
  C2RI I81 (itint_0n[25], i_0r1d[25], gate552_0n, initialise);
  C2RI I82 (itint_0n[26], i_0r1d[26], gate552_0n, initialise);
  C2RI I83 (itint_0n[27], i_0r1d[27], gate552_0n, initialise);
  C2RI I84 (itint_0n[28], i_0r1d[28], gate552_0n, initialise);
  C2RI I85 (itint_0n[29], i_0r1d[29], gate552_0n, initialise);
  C2RI I86 (itint_0n[30], i_0r1d[30], gate552_0n, initialise);
  C2RI I87 (itint_0n[31], i_0r1d[31], gate552_0n, initialise);
  C2RI I88 (ifint_0n[0], i_0r0d[0], gate552_0n, initialise);
  C2RI I89 (ifint_0n[1], i_0r0d[1], gate552_0n, initialise);
  C2RI I90 (ifint_0n[2], i_0r0d[2], gate552_0n, initialise);
  C2RI I91 (ifint_0n[3], i_0r0d[3], gate552_0n, initialise);
  C2RI I92 (ifint_0n[4], i_0r0d[4], gate552_0n, initialise);
  C2RI I93 (ifint_0n[5], i_0r0d[5], gate552_0n, initialise);
  C2RI I94 (ifint_0n[6], i_0r0d[6], gate552_0n, initialise);
  C2RI I95 (ifint_0n[7], i_0r0d[7], gate552_0n, initialise);
  C2RI I96 (ifint_0n[8], i_0r0d[8], gate552_0n, initialise);
  C2RI I97 (ifint_0n[9], i_0r0d[9], gate552_0n, initialise);
  C2RI I98 (ifint_0n[10], i_0r0d[10], gate552_0n, initialise);
  C2RI I99 (ifint_0n[11], i_0r0d[11], gate552_0n, initialise);
  C2RI I100 (ifint_0n[12], i_0r0d[12], gate552_0n, initialise);
  C2RI I101 (ifint_0n[13], i_0r0d[13], gate552_0n, initialise);
  C2RI I102 (ifint_0n[14], i_0r0d[14], gate552_0n, initialise);
  C2RI I103 (ifint_0n[15], i_0r0d[15], gate552_0n, initialise);
  C2RI I104 (ifint_0n[16], i_0r0d[16], gate552_0n, initialise);
  C2RI I105 (ifint_0n[17], i_0r0d[17], gate552_0n, initialise);
  C2RI I106 (ifint_0n[18], i_0r0d[18], gate552_0n, initialise);
  C2RI I107 (ifint_0n[19], i_0r0d[19], gate552_0n, initialise);
  C2RI I108 (ifint_0n[20], i_0r0d[20], gate552_0n, initialise);
  C2RI I109 (ifint_0n[21], i_0r0d[21], gate552_0n, initialise);
  C2RI I110 (ifint_0n[22], i_0r0d[22], gate552_0n, initialise);
  C2RI I111 (ifint_0n[23], i_0r0d[23], gate552_0n, initialise);
  C2RI I112 (ifint_0n[24], i_0r0d[24], gate552_0n, initialise);
  C2RI I113 (ifint_0n[25], i_0r0d[25], gate552_0n, initialise);
  C2RI I114 (ifint_0n[26], i_0r0d[26], gate552_0n, initialise);
  C2RI I115 (ifint_0n[27], i_0r0d[27], gate552_0n, initialise);
  C2RI I116 (ifint_0n[28], i_0r0d[28], gate552_0n, initialise);
  C2RI I117 (ifint_0n[29], i_0r0d[29], gate552_0n, initialise);
  C2RI I118 (ifint_0n[30], i_0r0d[30], gate552_0n, initialise);
  C2RI I119 (ifint_0n[31], i_0r0d[31], gate552_0n, initialise);
  C3 I120 (internal_0n[17], complete549_0n[0], complete549_0n[1], complete549_0n[2]);
  C3 I121 (internal_0n[18], complete549_0n[3], complete549_0n[4], complete549_0n[5]);
  C3 I122 (internal_0n[19], complete549_0n[6], complete549_0n[7], complete549_0n[8]);
  C3 I123 (internal_0n[20], complete549_0n[9], complete549_0n[10], complete549_0n[11]);
  C3 I124 (internal_0n[21], complete549_0n[12], complete549_0n[13], complete549_0n[14]);
  C3 I125 (internal_0n[22], complete549_0n[15], complete549_0n[16], complete549_0n[17]);
  C3 I126 (internal_0n[23], complete549_0n[18], complete549_0n[19], complete549_0n[20]);
  C3 I127 (internal_0n[24], complete549_0n[21], complete549_0n[22], complete549_0n[23]);
  C3 I128 (internal_0n[25], complete549_0n[24], complete549_0n[25], complete549_0n[26]);
  C3 I129 (internal_0n[26], complete549_0n[27], complete549_0n[28], complete549_0n[29]);
  C2 I130 (internal_0n[27], complete549_0n[30], complete549_0n[31]);
  C3 I131 (internal_0n[28], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I132 (internal_0n[29], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I133 (internal_0n[30], internal_0n[23], internal_0n[24], internal_0n[25]);
  C2 I134 (internal_0n[31], internal_0n[26], internal_0n[27]);
  C2 I135 (internal_0n[32], internal_0n[28], internal_0n[29]);
  C2 I136 (internal_0n[33], internal_0n[30], internal_0n[31]);
  C2 I137 (oaint_0n, internal_0n[32], internal_0n[33]);
  OR2 I138 (complete549_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I139 (complete549_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I140 (complete549_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I141 (complete549_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I142 (complete549_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I143 (complete549_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I144 (complete549_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I145 (complete549_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I146 (complete549_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I147 (complete549_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I148 (complete549_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I149 (complete549_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I150 (complete549_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I151 (complete549_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I152 (complete549_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I153 (complete549_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I154 (complete549_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I155 (complete549_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I156 (complete549_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I157 (complete549_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I158 (complete549_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I159 (complete549_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I160 (complete549_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I161 (complete549_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I162 (complete549_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I163 (complete549_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I164 (complete549_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I165 (complete549_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I166 (complete549_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I167 (complete549_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I168 (complete549_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I169 (complete549_0n[31], o_0r0d[31], o_0r1d[31]);
  INV I170 (gate548_0n, o_0a);
  C2RI I171 (o_0r1d[0], otint_0n[0], gate548_0n, initialise);
  C2RI I172 (o_0r1d[1], otint_0n[1], gate548_0n, initialise);
  C2RI I173 (o_0r1d[2], otint_0n[2], gate548_0n, initialise);
  C2RI I174 (o_0r1d[3], otint_0n[3], gate548_0n, initialise);
  C2RI I175 (o_0r1d[4], otint_0n[4], gate548_0n, initialise);
  C2RI I176 (o_0r1d[5], otint_0n[5], gate548_0n, initialise);
  C2RI I177 (o_0r1d[6], otint_0n[6], gate548_0n, initialise);
  C2RI I178 (o_0r1d[7], otint_0n[7], gate548_0n, initialise);
  C2RI I179 (o_0r1d[8], otint_0n[8], gate548_0n, initialise);
  C2RI I180 (o_0r1d[9], otint_0n[9], gate548_0n, initialise);
  C2RI I181 (o_0r1d[10], otint_0n[10], gate548_0n, initialise);
  C2RI I182 (o_0r1d[11], otint_0n[11], gate548_0n, initialise);
  C2RI I183 (o_0r1d[12], otint_0n[12], gate548_0n, initialise);
  C2RI I184 (o_0r1d[13], otint_0n[13], gate548_0n, initialise);
  C2RI I185 (o_0r1d[14], otint_0n[14], gate548_0n, initialise);
  C2RI I186 (o_0r1d[15], otint_0n[15], gate548_0n, initialise);
  C2RI I187 (o_0r1d[16], otint_0n[16], gate548_0n, initialise);
  C2RI I188 (o_0r1d[17], otint_0n[17], gate548_0n, initialise);
  C2RI I189 (o_0r1d[18], otint_0n[18], gate548_0n, initialise);
  C2RI I190 (o_0r1d[19], otint_0n[19], gate548_0n, initialise);
  C2RI I191 (o_0r1d[20], otint_0n[20], gate548_0n, initialise);
  C2RI I192 (o_0r1d[21], otint_0n[21], gate548_0n, initialise);
  C2RI I193 (o_0r1d[22], otint_0n[22], gate548_0n, initialise);
  C2RI I194 (o_0r1d[23], otint_0n[23], gate548_0n, initialise);
  C2RI I195 (o_0r1d[24], otint_0n[24], gate548_0n, initialise);
  C2RI I196 (o_0r1d[25], otint_0n[25], gate548_0n, initialise);
  C2RI I197 (o_0r1d[26], otint_0n[26], gate548_0n, initialise);
  C2RI I198 (o_0r1d[27], otint_0n[27], gate548_0n, initialise);
  C2RI I199 (o_0r1d[28], otint_0n[28], gate548_0n, initialise);
  C2RI I200 (o_0r1d[29], otint_0n[29], gate548_0n, initialise);
  C2RI I201 (o_0r1d[30], otint_0n[30], gate548_0n, initialise);
  C2RI I202 (o_0r1d[31], otint_0n[31], gate548_0n, initialise);
  C2RI I203 (o_0r0d[0], ofint_0n[0], gate548_0n, initialise);
  C2RI I204 (o_0r0d[1], ofint_0n[1], gate548_0n, initialise);
  C2RI I205 (o_0r0d[2], ofint_0n[2], gate548_0n, initialise);
  C2RI I206 (o_0r0d[3], ofint_0n[3], gate548_0n, initialise);
  C2RI I207 (o_0r0d[4], ofint_0n[4], gate548_0n, initialise);
  C2RI I208 (o_0r0d[5], ofint_0n[5], gate548_0n, initialise);
  C2RI I209 (o_0r0d[6], ofint_0n[6], gate548_0n, initialise);
  C2RI I210 (o_0r0d[7], ofint_0n[7], gate548_0n, initialise);
  C2RI I211 (o_0r0d[8], ofint_0n[8], gate548_0n, initialise);
  C2RI I212 (o_0r0d[9], ofint_0n[9], gate548_0n, initialise);
  C2RI I213 (o_0r0d[10], ofint_0n[10], gate548_0n, initialise);
  C2RI I214 (o_0r0d[11], ofint_0n[11], gate548_0n, initialise);
  C2RI I215 (o_0r0d[12], ofint_0n[12], gate548_0n, initialise);
  C2RI I216 (o_0r0d[13], ofint_0n[13], gate548_0n, initialise);
  C2RI I217 (o_0r0d[14], ofint_0n[14], gate548_0n, initialise);
  C2RI I218 (o_0r0d[15], ofint_0n[15], gate548_0n, initialise);
  C2RI I219 (o_0r0d[16], ofint_0n[16], gate548_0n, initialise);
  C2RI I220 (o_0r0d[17], ofint_0n[17], gate548_0n, initialise);
  C2RI I221 (o_0r0d[18], ofint_0n[18], gate548_0n, initialise);
  C2RI I222 (o_0r0d[19], ofint_0n[19], gate548_0n, initialise);
  C2RI I223 (o_0r0d[20], ofint_0n[20], gate548_0n, initialise);
  C2RI I224 (o_0r0d[21], ofint_0n[21], gate548_0n, initialise);
  C2RI I225 (o_0r0d[22], ofint_0n[22], gate548_0n, initialise);
  C2RI I226 (o_0r0d[23], ofint_0n[23], gate548_0n, initialise);
  C2RI I227 (o_0r0d[24], ofint_0n[24], gate548_0n, initialise);
  C2RI I228 (o_0r0d[25], ofint_0n[25], gate548_0n, initialise);
  C2RI I229 (o_0r0d[26], ofint_0n[26], gate548_0n, initialise);
  C2RI I230 (o_0r0d[27], ofint_0n[27], gate548_0n, initialise);
  C2RI I231 (o_0r0d[28], ofint_0n[28], gate548_0n, initialise);
  C2RI I232 (o_0r0d[29], ofint_0n[29], gate548_0n, initialise);
  C2RI I233 (o_0r0d[30], ofint_0n[30], gate548_0n, initialise);
  C2RI I234 (o_0r0d[31], ofint_0n[31], gate548_0n, initialise);
  assign otint_0n[1] = joint_0n[1];
  assign otint_0n[2] = joint_0n[2];
  assign otint_0n[3] = joint_0n[3];
  assign otint_0n[4] = joint_0n[4];
  assign otint_0n[5] = joint_0n[5];
  assign otint_0n[6] = joint_0n[6];
  assign otint_0n[7] = joint_0n[7];
  assign otint_0n[8] = joint_0n[8];
  assign otint_0n[9] = joint_0n[9];
  assign otint_0n[10] = joint_0n[10];
  assign otint_0n[11] = joint_0n[11];
  assign otint_0n[12] = joint_0n[12];
  assign otint_0n[13] = joint_0n[13];
  assign otint_0n[14] = joint_0n[14];
  assign otint_0n[15] = joint_0n[15];
  assign otint_0n[16] = joint_0n[16];
  assign otint_0n[17] = joint_0n[17];
  assign otint_0n[18] = joint_0n[18];
  assign otint_0n[19] = joint_0n[19];
  assign otint_0n[20] = joint_0n[20];
  assign otint_0n[21] = joint_0n[21];
  assign otint_0n[22] = joint_0n[22];
  assign otint_0n[23] = joint_0n[23];
  assign otint_0n[24] = joint_0n[24];
  assign otint_0n[25] = joint_0n[25];
  assign otint_0n[26] = joint_0n[26];
  assign otint_0n[27] = joint_0n[27];
  assign otint_0n[28] = joint_0n[28];
  assign otint_0n[29] = joint_0n[29];
  assign otint_0n[30] = joint_0n[30];
  assign otint_0n[31] = joint_0n[31];
  assign ofint_0n[1] = joinf_0n[1];
  assign ofint_0n[2] = joinf_0n[2];
  assign ofint_0n[3] = joinf_0n[3];
  assign ofint_0n[4] = joinf_0n[4];
  assign ofint_0n[5] = joinf_0n[5];
  assign ofint_0n[6] = joinf_0n[6];
  assign ofint_0n[7] = joinf_0n[7];
  assign ofint_0n[8] = joinf_0n[8];
  assign ofint_0n[9] = joinf_0n[9];
  assign ofint_0n[10] = joinf_0n[10];
  assign ofint_0n[11] = joinf_0n[11];
  assign ofint_0n[12] = joinf_0n[12];
  assign ofint_0n[13] = joinf_0n[13];
  assign ofint_0n[14] = joinf_0n[14];
  assign ofint_0n[15] = joinf_0n[15];
  assign ofint_0n[16] = joinf_0n[16];
  assign ofint_0n[17] = joinf_0n[17];
  assign ofint_0n[18] = joinf_0n[18];
  assign ofint_0n[19] = joinf_0n[19];
  assign ofint_0n[20] = joinf_0n[20];
  assign ofint_0n[21] = joinf_0n[21];
  assign ofint_0n[22] = joinf_0n[22];
  assign ofint_0n[23] = joinf_0n[23];
  assign ofint_0n[24] = joinf_0n[24];
  assign ofint_0n[25] = joinf_0n[25];
  assign ofint_0n[26] = joinf_0n[26];
  assign ofint_0n[27] = joinf_0n[27];
  assign ofint_0n[28] = joinf_0n[28];
  assign ofint_0n[29] = joinf_0n[29];
  assign ofint_0n[30] = joinf_0n[30];
  assign ofint_0n[31] = joinf_0n[31];
  C2 I297 (otint_0n[0], joint_0n[0], icomplete_0n);
  C2 I298 (ofint_0n[0], joinf_0n[0], icomplete_0n);
  assign icomplete_0n = ifint_1n;
  assign joint_0n[0] = itint_0n[0];
  assign joint_0n[1] = itint_0n[1];
  assign joint_0n[2] = itint_0n[2];
  assign joint_0n[3] = itint_0n[3];
  assign joint_0n[4] = itint_0n[4];
  assign joint_0n[5] = itint_0n[5];
  assign joint_0n[6] = itint_0n[6];
  assign joint_0n[7] = itint_0n[7];
  assign joint_0n[8] = itint_0n[8];
  assign joint_0n[9] = itint_0n[9];
  assign joint_0n[10] = itint_0n[10];
  assign joint_0n[11] = itint_0n[11];
  assign joint_0n[12] = itint_0n[12];
  assign joint_0n[13] = itint_0n[13];
  assign joint_0n[14] = itint_0n[14];
  assign joint_0n[15] = itint_0n[15];
  assign joint_0n[16] = itint_0n[16];
  assign joint_0n[17] = itint_0n[17];
  assign joint_0n[18] = itint_0n[18];
  assign joint_0n[19] = itint_0n[19];
  assign joint_0n[20] = itint_0n[20];
  assign joint_0n[21] = itint_0n[21];
  assign joint_0n[22] = itint_0n[22];
  assign joint_0n[23] = itint_0n[23];
  assign joint_0n[24] = itint_0n[24];
  assign joint_0n[25] = itint_0n[25];
  assign joint_0n[26] = itint_0n[26];
  assign joint_0n[27] = itint_0n[27];
  assign joint_0n[28] = itint_0n[28];
  assign joint_0n[29] = itint_0n[29];
  assign joint_0n[30] = itint_0n[30];
  assign joint_0n[31] = itint_0n[31];
  assign joinf_0n[0] = ifint_0n[0];
  assign joinf_0n[1] = ifint_0n[1];
  assign joinf_0n[2] = ifint_0n[2];
  assign joinf_0n[3] = ifint_0n[3];
  assign joinf_0n[4] = ifint_0n[4];
  assign joinf_0n[5] = ifint_0n[5];
  assign joinf_0n[6] = ifint_0n[6];
  assign joinf_0n[7] = ifint_0n[7];
  assign joinf_0n[8] = ifint_0n[8];
  assign joinf_0n[9] = ifint_0n[9];
  assign joinf_0n[10] = ifint_0n[10];
  assign joinf_0n[11] = ifint_0n[11];
  assign joinf_0n[12] = ifint_0n[12];
  assign joinf_0n[13] = ifint_0n[13];
  assign joinf_0n[14] = ifint_0n[14];
  assign joinf_0n[15] = ifint_0n[15];
  assign joinf_0n[16] = ifint_0n[16];
  assign joinf_0n[17] = ifint_0n[17];
  assign joinf_0n[18] = ifint_0n[18];
  assign joinf_0n[19] = ifint_0n[19];
  assign joinf_0n[20] = ifint_0n[20];
  assign joinf_0n[21] = ifint_0n[21];
  assign joinf_0n[22] = ifint_0n[22];
  assign joinf_0n[23] = ifint_0n[23];
  assign joinf_0n[24] = ifint_0n[24];
  assign joinf_0n[25] = ifint_0n[25];
  assign joinf_0n[26] = ifint_0n[26];
  assign joinf_0n[27] = ifint_0n[27];
  assign joinf_0n[28] = ifint_0n[28];
  assign joinf_0n[29] = ifint_0n[29];
  assign joinf_0n[30] = ifint_0n[30];
  assign joinf_0n[31] = ifint_0n[31];
endmodule

module BrzJ_l12__2832_201_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [31:0] i_0r0d;
  input [31:0] i_0r1d;
  output i_0a;
  input i_1r0d;
  input i_1r1d;
  output i_1a;
  output [32:0] o_0r0d;
  output [32:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [33:0] internal_0n;
  wire [32:0] ofint_0n;
  wire [32:0] otint_0n;
  wire oaint_0n;
  wire [31:0] ifint_0n;
  wire ifint_1n;
  wire [31:0] itint_0n;
  wire itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire complete568_0n;
  wire gate567_0n;
  wire [31:0] complete564_0n;
  wire gate563_0n;
  wire [32:0] complete560_0n;
  wire gate559_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign i_1a = complete568_0n;
  OR2 I3 (complete568_0n, ifint_1n, itint_1n);
  INV I4 (gate567_0n, iaint_1n);
  C2RI I5 (itint_1n, i_1r1d, gate567_0n, initialise);
  C2RI I6 (ifint_1n, i_1r0d, gate567_0n, initialise);
  C3 I7 (internal_0n[0], complete564_0n[0], complete564_0n[1], complete564_0n[2]);
  C3 I8 (internal_0n[1], complete564_0n[3], complete564_0n[4], complete564_0n[5]);
  C3 I9 (internal_0n[2], complete564_0n[6], complete564_0n[7], complete564_0n[8]);
  C3 I10 (internal_0n[3], complete564_0n[9], complete564_0n[10], complete564_0n[11]);
  C3 I11 (internal_0n[4], complete564_0n[12], complete564_0n[13], complete564_0n[14]);
  C3 I12 (internal_0n[5], complete564_0n[15], complete564_0n[16], complete564_0n[17]);
  C3 I13 (internal_0n[6], complete564_0n[18], complete564_0n[19], complete564_0n[20]);
  C3 I14 (internal_0n[7], complete564_0n[21], complete564_0n[22], complete564_0n[23]);
  C3 I15 (internal_0n[8], complete564_0n[24], complete564_0n[25], complete564_0n[26]);
  C3 I16 (internal_0n[9], complete564_0n[27], complete564_0n[28], complete564_0n[29]);
  C2 I17 (internal_0n[10], complete564_0n[30], complete564_0n[31]);
  C3 I18 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I19 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I20 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I21 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I22 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I23 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I24 (i_0a, internal_0n[15], internal_0n[16]);
  OR2 I25 (complete564_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I26 (complete564_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I27 (complete564_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I28 (complete564_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I29 (complete564_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I30 (complete564_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I31 (complete564_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I32 (complete564_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I33 (complete564_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I34 (complete564_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I35 (complete564_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I36 (complete564_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I37 (complete564_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I38 (complete564_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I39 (complete564_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I40 (complete564_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I41 (complete564_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I42 (complete564_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I43 (complete564_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I44 (complete564_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I45 (complete564_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I46 (complete564_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I47 (complete564_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I48 (complete564_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I49 (complete564_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I50 (complete564_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I51 (complete564_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I52 (complete564_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I53 (complete564_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I54 (complete564_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I55 (complete564_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I56 (complete564_0n[31], ifint_0n[31], itint_0n[31]);
  INV I57 (gate563_0n, iaint_0n);
  C2RI I58 (itint_0n[0], i_0r1d[0], gate563_0n, initialise);
  C2RI I59 (itint_0n[1], i_0r1d[1], gate563_0n, initialise);
  C2RI I60 (itint_0n[2], i_0r1d[2], gate563_0n, initialise);
  C2RI I61 (itint_0n[3], i_0r1d[3], gate563_0n, initialise);
  C2RI I62 (itint_0n[4], i_0r1d[4], gate563_0n, initialise);
  C2RI I63 (itint_0n[5], i_0r1d[5], gate563_0n, initialise);
  C2RI I64 (itint_0n[6], i_0r1d[6], gate563_0n, initialise);
  C2RI I65 (itint_0n[7], i_0r1d[7], gate563_0n, initialise);
  C2RI I66 (itint_0n[8], i_0r1d[8], gate563_0n, initialise);
  C2RI I67 (itint_0n[9], i_0r1d[9], gate563_0n, initialise);
  C2RI I68 (itint_0n[10], i_0r1d[10], gate563_0n, initialise);
  C2RI I69 (itint_0n[11], i_0r1d[11], gate563_0n, initialise);
  C2RI I70 (itint_0n[12], i_0r1d[12], gate563_0n, initialise);
  C2RI I71 (itint_0n[13], i_0r1d[13], gate563_0n, initialise);
  C2RI I72 (itint_0n[14], i_0r1d[14], gate563_0n, initialise);
  C2RI I73 (itint_0n[15], i_0r1d[15], gate563_0n, initialise);
  C2RI I74 (itint_0n[16], i_0r1d[16], gate563_0n, initialise);
  C2RI I75 (itint_0n[17], i_0r1d[17], gate563_0n, initialise);
  C2RI I76 (itint_0n[18], i_0r1d[18], gate563_0n, initialise);
  C2RI I77 (itint_0n[19], i_0r1d[19], gate563_0n, initialise);
  C2RI I78 (itint_0n[20], i_0r1d[20], gate563_0n, initialise);
  C2RI I79 (itint_0n[21], i_0r1d[21], gate563_0n, initialise);
  C2RI I80 (itint_0n[22], i_0r1d[22], gate563_0n, initialise);
  C2RI I81 (itint_0n[23], i_0r1d[23], gate563_0n, initialise);
  C2RI I82 (itint_0n[24], i_0r1d[24], gate563_0n, initialise);
  C2RI I83 (itint_0n[25], i_0r1d[25], gate563_0n, initialise);
  C2RI I84 (itint_0n[26], i_0r1d[26], gate563_0n, initialise);
  C2RI I85 (itint_0n[27], i_0r1d[27], gate563_0n, initialise);
  C2RI I86 (itint_0n[28], i_0r1d[28], gate563_0n, initialise);
  C2RI I87 (itint_0n[29], i_0r1d[29], gate563_0n, initialise);
  C2RI I88 (itint_0n[30], i_0r1d[30], gate563_0n, initialise);
  C2RI I89 (itint_0n[31], i_0r1d[31], gate563_0n, initialise);
  C2RI I90 (ifint_0n[0], i_0r0d[0], gate563_0n, initialise);
  C2RI I91 (ifint_0n[1], i_0r0d[1], gate563_0n, initialise);
  C2RI I92 (ifint_0n[2], i_0r0d[2], gate563_0n, initialise);
  C2RI I93 (ifint_0n[3], i_0r0d[3], gate563_0n, initialise);
  C2RI I94 (ifint_0n[4], i_0r0d[4], gate563_0n, initialise);
  C2RI I95 (ifint_0n[5], i_0r0d[5], gate563_0n, initialise);
  C2RI I96 (ifint_0n[6], i_0r0d[6], gate563_0n, initialise);
  C2RI I97 (ifint_0n[7], i_0r0d[7], gate563_0n, initialise);
  C2RI I98 (ifint_0n[8], i_0r0d[8], gate563_0n, initialise);
  C2RI I99 (ifint_0n[9], i_0r0d[9], gate563_0n, initialise);
  C2RI I100 (ifint_0n[10], i_0r0d[10], gate563_0n, initialise);
  C2RI I101 (ifint_0n[11], i_0r0d[11], gate563_0n, initialise);
  C2RI I102 (ifint_0n[12], i_0r0d[12], gate563_0n, initialise);
  C2RI I103 (ifint_0n[13], i_0r0d[13], gate563_0n, initialise);
  C2RI I104 (ifint_0n[14], i_0r0d[14], gate563_0n, initialise);
  C2RI I105 (ifint_0n[15], i_0r0d[15], gate563_0n, initialise);
  C2RI I106 (ifint_0n[16], i_0r0d[16], gate563_0n, initialise);
  C2RI I107 (ifint_0n[17], i_0r0d[17], gate563_0n, initialise);
  C2RI I108 (ifint_0n[18], i_0r0d[18], gate563_0n, initialise);
  C2RI I109 (ifint_0n[19], i_0r0d[19], gate563_0n, initialise);
  C2RI I110 (ifint_0n[20], i_0r0d[20], gate563_0n, initialise);
  C2RI I111 (ifint_0n[21], i_0r0d[21], gate563_0n, initialise);
  C2RI I112 (ifint_0n[22], i_0r0d[22], gate563_0n, initialise);
  C2RI I113 (ifint_0n[23], i_0r0d[23], gate563_0n, initialise);
  C2RI I114 (ifint_0n[24], i_0r0d[24], gate563_0n, initialise);
  C2RI I115 (ifint_0n[25], i_0r0d[25], gate563_0n, initialise);
  C2RI I116 (ifint_0n[26], i_0r0d[26], gate563_0n, initialise);
  C2RI I117 (ifint_0n[27], i_0r0d[27], gate563_0n, initialise);
  C2RI I118 (ifint_0n[28], i_0r0d[28], gate563_0n, initialise);
  C2RI I119 (ifint_0n[29], i_0r0d[29], gate563_0n, initialise);
  C2RI I120 (ifint_0n[30], i_0r0d[30], gate563_0n, initialise);
  C2RI I121 (ifint_0n[31], i_0r0d[31], gate563_0n, initialise);
  C3 I122 (internal_0n[17], complete560_0n[0], complete560_0n[1], complete560_0n[2]);
  C3 I123 (internal_0n[18], complete560_0n[3], complete560_0n[4], complete560_0n[5]);
  C3 I124 (internal_0n[19], complete560_0n[6], complete560_0n[7], complete560_0n[8]);
  C3 I125 (internal_0n[20], complete560_0n[9], complete560_0n[10], complete560_0n[11]);
  C3 I126 (internal_0n[21], complete560_0n[12], complete560_0n[13], complete560_0n[14]);
  C3 I127 (internal_0n[22], complete560_0n[15], complete560_0n[16], complete560_0n[17]);
  C3 I128 (internal_0n[23], complete560_0n[18], complete560_0n[19], complete560_0n[20]);
  C3 I129 (internal_0n[24], complete560_0n[21], complete560_0n[22], complete560_0n[23]);
  C3 I130 (internal_0n[25], complete560_0n[24], complete560_0n[25], complete560_0n[26]);
  C3 I131 (internal_0n[26], complete560_0n[27], complete560_0n[28], complete560_0n[29]);
  C3 I132 (internal_0n[27], complete560_0n[30], complete560_0n[31], complete560_0n[32]);
  C3 I133 (internal_0n[28], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I134 (internal_0n[29], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I135 (internal_0n[30], internal_0n[23], internal_0n[24], internal_0n[25]);
  C2 I136 (internal_0n[31], internal_0n[26], internal_0n[27]);
  C2 I137 (internal_0n[32], internal_0n[28], internal_0n[29]);
  C2 I138 (internal_0n[33], internal_0n[30], internal_0n[31]);
  C2 I139 (oaint_0n, internal_0n[32], internal_0n[33]);
  OR2 I140 (complete560_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I141 (complete560_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I142 (complete560_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I143 (complete560_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I144 (complete560_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I145 (complete560_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I146 (complete560_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I147 (complete560_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I148 (complete560_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I149 (complete560_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I150 (complete560_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I151 (complete560_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I152 (complete560_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I153 (complete560_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I154 (complete560_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I155 (complete560_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I156 (complete560_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I157 (complete560_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I158 (complete560_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I159 (complete560_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I160 (complete560_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I161 (complete560_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I162 (complete560_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I163 (complete560_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I164 (complete560_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I165 (complete560_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I166 (complete560_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I167 (complete560_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I168 (complete560_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I169 (complete560_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I170 (complete560_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I171 (complete560_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I172 (complete560_0n[32], o_0r0d[32], o_0r1d[32]);
  INV I173 (gate559_0n, o_0a);
  C2RI I174 (o_0r1d[0], otint_0n[0], gate559_0n, initialise);
  C2RI I175 (o_0r1d[1], otint_0n[1], gate559_0n, initialise);
  C2RI I176 (o_0r1d[2], otint_0n[2], gate559_0n, initialise);
  C2RI I177 (o_0r1d[3], otint_0n[3], gate559_0n, initialise);
  C2RI I178 (o_0r1d[4], otint_0n[4], gate559_0n, initialise);
  C2RI I179 (o_0r1d[5], otint_0n[5], gate559_0n, initialise);
  C2RI I180 (o_0r1d[6], otint_0n[6], gate559_0n, initialise);
  C2RI I181 (o_0r1d[7], otint_0n[7], gate559_0n, initialise);
  C2RI I182 (o_0r1d[8], otint_0n[8], gate559_0n, initialise);
  C2RI I183 (o_0r1d[9], otint_0n[9], gate559_0n, initialise);
  C2RI I184 (o_0r1d[10], otint_0n[10], gate559_0n, initialise);
  C2RI I185 (o_0r1d[11], otint_0n[11], gate559_0n, initialise);
  C2RI I186 (o_0r1d[12], otint_0n[12], gate559_0n, initialise);
  C2RI I187 (o_0r1d[13], otint_0n[13], gate559_0n, initialise);
  C2RI I188 (o_0r1d[14], otint_0n[14], gate559_0n, initialise);
  C2RI I189 (o_0r1d[15], otint_0n[15], gate559_0n, initialise);
  C2RI I190 (o_0r1d[16], otint_0n[16], gate559_0n, initialise);
  C2RI I191 (o_0r1d[17], otint_0n[17], gate559_0n, initialise);
  C2RI I192 (o_0r1d[18], otint_0n[18], gate559_0n, initialise);
  C2RI I193 (o_0r1d[19], otint_0n[19], gate559_0n, initialise);
  C2RI I194 (o_0r1d[20], otint_0n[20], gate559_0n, initialise);
  C2RI I195 (o_0r1d[21], otint_0n[21], gate559_0n, initialise);
  C2RI I196 (o_0r1d[22], otint_0n[22], gate559_0n, initialise);
  C2RI I197 (o_0r1d[23], otint_0n[23], gate559_0n, initialise);
  C2RI I198 (o_0r1d[24], otint_0n[24], gate559_0n, initialise);
  C2RI I199 (o_0r1d[25], otint_0n[25], gate559_0n, initialise);
  C2RI I200 (o_0r1d[26], otint_0n[26], gate559_0n, initialise);
  C2RI I201 (o_0r1d[27], otint_0n[27], gate559_0n, initialise);
  C2RI I202 (o_0r1d[28], otint_0n[28], gate559_0n, initialise);
  C2RI I203 (o_0r1d[29], otint_0n[29], gate559_0n, initialise);
  C2RI I204 (o_0r1d[30], otint_0n[30], gate559_0n, initialise);
  C2RI I205 (o_0r1d[31], otint_0n[31], gate559_0n, initialise);
  C2RI I206 (o_0r1d[32], otint_0n[32], gate559_0n, initialise);
  C2RI I207 (o_0r0d[0], ofint_0n[0], gate559_0n, initialise);
  C2RI I208 (o_0r0d[1], ofint_0n[1], gate559_0n, initialise);
  C2RI I209 (o_0r0d[2], ofint_0n[2], gate559_0n, initialise);
  C2RI I210 (o_0r0d[3], ofint_0n[3], gate559_0n, initialise);
  C2RI I211 (o_0r0d[4], ofint_0n[4], gate559_0n, initialise);
  C2RI I212 (o_0r0d[5], ofint_0n[5], gate559_0n, initialise);
  C2RI I213 (o_0r0d[6], ofint_0n[6], gate559_0n, initialise);
  C2RI I214 (o_0r0d[7], ofint_0n[7], gate559_0n, initialise);
  C2RI I215 (o_0r0d[8], ofint_0n[8], gate559_0n, initialise);
  C2RI I216 (o_0r0d[9], ofint_0n[9], gate559_0n, initialise);
  C2RI I217 (o_0r0d[10], ofint_0n[10], gate559_0n, initialise);
  C2RI I218 (o_0r0d[11], ofint_0n[11], gate559_0n, initialise);
  C2RI I219 (o_0r0d[12], ofint_0n[12], gate559_0n, initialise);
  C2RI I220 (o_0r0d[13], ofint_0n[13], gate559_0n, initialise);
  C2RI I221 (o_0r0d[14], ofint_0n[14], gate559_0n, initialise);
  C2RI I222 (o_0r0d[15], ofint_0n[15], gate559_0n, initialise);
  C2RI I223 (o_0r0d[16], ofint_0n[16], gate559_0n, initialise);
  C2RI I224 (o_0r0d[17], ofint_0n[17], gate559_0n, initialise);
  C2RI I225 (o_0r0d[18], ofint_0n[18], gate559_0n, initialise);
  C2RI I226 (o_0r0d[19], ofint_0n[19], gate559_0n, initialise);
  C2RI I227 (o_0r0d[20], ofint_0n[20], gate559_0n, initialise);
  C2RI I228 (o_0r0d[21], ofint_0n[21], gate559_0n, initialise);
  C2RI I229 (o_0r0d[22], ofint_0n[22], gate559_0n, initialise);
  C2RI I230 (o_0r0d[23], ofint_0n[23], gate559_0n, initialise);
  C2RI I231 (o_0r0d[24], ofint_0n[24], gate559_0n, initialise);
  C2RI I232 (o_0r0d[25], ofint_0n[25], gate559_0n, initialise);
  C2RI I233 (o_0r0d[26], ofint_0n[26], gate559_0n, initialise);
  C2RI I234 (o_0r0d[27], ofint_0n[27], gate559_0n, initialise);
  C2RI I235 (o_0r0d[28], ofint_0n[28], gate559_0n, initialise);
  C2RI I236 (o_0r0d[29], ofint_0n[29], gate559_0n, initialise);
  C2RI I237 (o_0r0d[30], ofint_0n[30], gate559_0n, initialise);
  C2RI I238 (o_0r0d[31], ofint_0n[31], gate559_0n, initialise);
  C2RI I239 (o_0r0d[32], ofint_0n[32], gate559_0n, initialise);
  assign otint_0n[0] = itint_0n[0];
  assign otint_0n[1] = itint_0n[1];
  assign otint_0n[2] = itint_0n[2];
  assign otint_0n[3] = itint_0n[3];
  assign otint_0n[4] = itint_0n[4];
  assign otint_0n[5] = itint_0n[5];
  assign otint_0n[6] = itint_0n[6];
  assign otint_0n[7] = itint_0n[7];
  assign otint_0n[8] = itint_0n[8];
  assign otint_0n[9] = itint_0n[9];
  assign otint_0n[10] = itint_0n[10];
  assign otint_0n[11] = itint_0n[11];
  assign otint_0n[12] = itint_0n[12];
  assign otint_0n[13] = itint_0n[13];
  assign otint_0n[14] = itint_0n[14];
  assign otint_0n[15] = itint_0n[15];
  assign otint_0n[16] = itint_0n[16];
  assign otint_0n[17] = itint_0n[17];
  assign otint_0n[18] = itint_0n[18];
  assign otint_0n[19] = itint_0n[19];
  assign otint_0n[20] = itint_0n[20];
  assign otint_0n[21] = itint_0n[21];
  assign otint_0n[22] = itint_0n[22];
  assign otint_0n[23] = itint_0n[23];
  assign otint_0n[24] = itint_0n[24];
  assign otint_0n[25] = itint_0n[25];
  assign otint_0n[26] = itint_0n[26];
  assign otint_0n[27] = itint_0n[27];
  assign otint_0n[28] = itint_0n[28];
  assign otint_0n[29] = itint_0n[29];
  assign otint_0n[30] = itint_0n[30];
  assign otint_0n[31] = itint_0n[31];
  assign otint_0n[32] = itint_1n;
  assign ofint_0n[0] = ifint_0n[0];
  assign ofint_0n[1] = ifint_0n[1];
  assign ofint_0n[2] = ifint_0n[2];
  assign ofint_0n[3] = ifint_0n[3];
  assign ofint_0n[4] = ifint_0n[4];
  assign ofint_0n[5] = ifint_0n[5];
  assign ofint_0n[6] = ifint_0n[6];
  assign ofint_0n[7] = ifint_0n[7];
  assign ofint_0n[8] = ifint_0n[8];
  assign ofint_0n[9] = ifint_0n[9];
  assign ofint_0n[10] = ifint_0n[10];
  assign ofint_0n[11] = ifint_0n[11];
  assign ofint_0n[12] = ifint_0n[12];
  assign ofint_0n[13] = ifint_0n[13];
  assign ofint_0n[14] = ifint_0n[14];
  assign ofint_0n[15] = ifint_0n[15];
  assign ofint_0n[16] = ifint_0n[16];
  assign ofint_0n[17] = ifint_0n[17];
  assign ofint_0n[18] = ifint_0n[18];
  assign ofint_0n[19] = ifint_0n[19];
  assign ofint_0n[20] = ifint_0n[20];
  assign ofint_0n[21] = ifint_0n[21];
  assign ofint_0n[22] = ifint_0n[22];
  assign ofint_0n[23] = ifint_0n[23];
  assign ofint_0n[24] = ifint_0n[24];
  assign ofint_0n[25] = ifint_0n[25];
  assign ofint_0n[26] = ifint_0n[26];
  assign ofint_0n[27] = ifint_0n[27];
  assign ofint_0n[28] = ifint_0n[28];
  assign ofint_0n[29] = ifint_0n[29];
  assign ofint_0n[30] = ifint_0n[30];
  assign ofint_0n[31] = ifint_0n[31];
  assign ofint_0n[32] = ifint_1n;
endmodule

module BrzJ_l12__2832_202_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [31:0] i_0r0d;
  input [31:0] i_0r1d;
  output i_0a;
  input [1:0] i_1r0d;
  input [1:0] i_1r1d;
  output i_1a;
  output [33:0] o_0r0d;
  output [33:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [34:0] internal_0n;
  wire [33:0] ofint_0n;
  wire [33:0] otint_0n;
  wire oaint_0n;
  wire [31:0] ifint_0n;
  wire [1:0] ifint_1n;
  wire [31:0] itint_0n;
  wire [1:0] itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [1:0] complete580_0n;
  wire gate579_0n;
  wire [31:0] complete576_0n;
  wire gate575_0n;
  wire [33:0] complete572_0n;
  wire gate571_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  C2 I2 (i_1a, complete580_0n[0], complete580_0n[1]);
  OR2 I3 (complete580_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I4 (complete580_0n[1], ifint_1n[1], itint_1n[1]);
  INV I5 (gate579_0n, iaint_1n);
  C2RI I6 (itint_1n[0], i_1r1d[0], gate579_0n, initialise);
  C2RI I7 (itint_1n[1], i_1r1d[1], gate579_0n, initialise);
  C2RI I8 (ifint_1n[0], i_1r0d[0], gate579_0n, initialise);
  C2RI I9 (ifint_1n[1], i_1r0d[1], gate579_0n, initialise);
  C3 I10 (internal_0n[0], complete576_0n[0], complete576_0n[1], complete576_0n[2]);
  C3 I11 (internal_0n[1], complete576_0n[3], complete576_0n[4], complete576_0n[5]);
  C3 I12 (internal_0n[2], complete576_0n[6], complete576_0n[7], complete576_0n[8]);
  C3 I13 (internal_0n[3], complete576_0n[9], complete576_0n[10], complete576_0n[11]);
  C3 I14 (internal_0n[4], complete576_0n[12], complete576_0n[13], complete576_0n[14]);
  C3 I15 (internal_0n[5], complete576_0n[15], complete576_0n[16], complete576_0n[17]);
  C3 I16 (internal_0n[6], complete576_0n[18], complete576_0n[19], complete576_0n[20]);
  C3 I17 (internal_0n[7], complete576_0n[21], complete576_0n[22], complete576_0n[23]);
  C3 I18 (internal_0n[8], complete576_0n[24], complete576_0n[25], complete576_0n[26]);
  C3 I19 (internal_0n[9], complete576_0n[27], complete576_0n[28], complete576_0n[29]);
  C2 I20 (internal_0n[10], complete576_0n[30], complete576_0n[31]);
  C3 I21 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I22 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I23 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I24 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I25 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I26 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I27 (i_0a, internal_0n[15], internal_0n[16]);
  OR2 I28 (complete576_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I29 (complete576_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I30 (complete576_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I31 (complete576_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I32 (complete576_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I33 (complete576_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I34 (complete576_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I35 (complete576_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I36 (complete576_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I37 (complete576_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I38 (complete576_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I39 (complete576_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I40 (complete576_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I41 (complete576_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I42 (complete576_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I43 (complete576_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I44 (complete576_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I45 (complete576_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I46 (complete576_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I47 (complete576_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I48 (complete576_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I49 (complete576_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I50 (complete576_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I51 (complete576_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I52 (complete576_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I53 (complete576_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I54 (complete576_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I55 (complete576_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I56 (complete576_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I57 (complete576_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I58 (complete576_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I59 (complete576_0n[31], ifint_0n[31], itint_0n[31]);
  INV I60 (gate575_0n, iaint_0n);
  C2RI I61 (itint_0n[0], i_0r1d[0], gate575_0n, initialise);
  C2RI I62 (itint_0n[1], i_0r1d[1], gate575_0n, initialise);
  C2RI I63 (itint_0n[2], i_0r1d[2], gate575_0n, initialise);
  C2RI I64 (itint_0n[3], i_0r1d[3], gate575_0n, initialise);
  C2RI I65 (itint_0n[4], i_0r1d[4], gate575_0n, initialise);
  C2RI I66 (itint_0n[5], i_0r1d[5], gate575_0n, initialise);
  C2RI I67 (itint_0n[6], i_0r1d[6], gate575_0n, initialise);
  C2RI I68 (itint_0n[7], i_0r1d[7], gate575_0n, initialise);
  C2RI I69 (itint_0n[8], i_0r1d[8], gate575_0n, initialise);
  C2RI I70 (itint_0n[9], i_0r1d[9], gate575_0n, initialise);
  C2RI I71 (itint_0n[10], i_0r1d[10], gate575_0n, initialise);
  C2RI I72 (itint_0n[11], i_0r1d[11], gate575_0n, initialise);
  C2RI I73 (itint_0n[12], i_0r1d[12], gate575_0n, initialise);
  C2RI I74 (itint_0n[13], i_0r1d[13], gate575_0n, initialise);
  C2RI I75 (itint_0n[14], i_0r1d[14], gate575_0n, initialise);
  C2RI I76 (itint_0n[15], i_0r1d[15], gate575_0n, initialise);
  C2RI I77 (itint_0n[16], i_0r1d[16], gate575_0n, initialise);
  C2RI I78 (itint_0n[17], i_0r1d[17], gate575_0n, initialise);
  C2RI I79 (itint_0n[18], i_0r1d[18], gate575_0n, initialise);
  C2RI I80 (itint_0n[19], i_0r1d[19], gate575_0n, initialise);
  C2RI I81 (itint_0n[20], i_0r1d[20], gate575_0n, initialise);
  C2RI I82 (itint_0n[21], i_0r1d[21], gate575_0n, initialise);
  C2RI I83 (itint_0n[22], i_0r1d[22], gate575_0n, initialise);
  C2RI I84 (itint_0n[23], i_0r1d[23], gate575_0n, initialise);
  C2RI I85 (itint_0n[24], i_0r1d[24], gate575_0n, initialise);
  C2RI I86 (itint_0n[25], i_0r1d[25], gate575_0n, initialise);
  C2RI I87 (itint_0n[26], i_0r1d[26], gate575_0n, initialise);
  C2RI I88 (itint_0n[27], i_0r1d[27], gate575_0n, initialise);
  C2RI I89 (itint_0n[28], i_0r1d[28], gate575_0n, initialise);
  C2RI I90 (itint_0n[29], i_0r1d[29], gate575_0n, initialise);
  C2RI I91 (itint_0n[30], i_0r1d[30], gate575_0n, initialise);
  C2RI I92 (itint_0n[31], i_0r1d[31], gate575_0n, initialise);
  C2RI I93 (ifint_0n[0], i_0r0d[0], gate575_0n, initialise);
  C2RI I94 (ifint_0n[1], i_0r0d[1], gate575_0n, initialise);
  C2RI I95 (ifint_0n[2], i_0r0d[2], gate575_0n, initialise);
  C2RI I96 (ifint_0n[3], i_0r0d[3], gate575_0n, initialise);
  C2RI I97 (ifint_0n[4], i_0r0d[4], gate575_0n, initialise);
  C2RI I98 (ifint_0n[5], i_0r0d[5], gate575_0n, initialise);
  C2RI I99 (ifint_0n[6], i_0r0d[6], gate575_0n, initialise);
  C2RI I100 (ifint_0n[7], i_0r0d[7], gate575_0n, initialise);
  C2RI I101 (ifint_0n[8], i_0r0d[8], gate575_0n, initialise);
  C2RI I102 (ifint_0n[9], i_0r0d[9], gate575_0n, initialise);
  C2RI I103 (ifint_0n[10], i_0r0d[10], gate575_0n, initialise);
  C2RI I104 (ifint_0n[11], i_0r0d[11], gate575_0n, initialise);
  C2RI I105 (ifint_0n[12], i_0r0d[12], gate575_0n, initialise);
  C2RI I106 (ifint_0n[13], i_0r0d[13], gate575_0n, initialise);
  C2RI I107 (ifint_0n[14], i_0r0d[14], gate575_0n, initialise);
  C2RI I108 (ifint_0n[15], i_0r0d[15], gate575_0n, initialise);
  C2RI I109 (ifint_0n[16], i_0r0d[16], gate575_0n, initialise);
  C2RI I110 (ifint_0n[17], i_0r0d[17], gate575_0n, initialise);
  C2RI I111 (ifint_0n[18], i_0r0d[18], gate575_0n, initialise);
  C2RI I112 (ifint_0n[19], i_0r0d[19], gate575_0n, initialise);
  C2RI I113 (ifint_0n[20], i_0r0d[20], gate575_0n, initialise);
  C2RI I114 (ifint_0n[21], i_0r0d[21], gate575_0n, initialise);
  C2RI I115 (ifint_0n[22], i_0r0d[22], gate575_0n, initialise);
  C2RI I116 (ifint_0n[23], i_0r0d[23], gate575_0n, initialise);
  C2RI I117 (ifint_0n[24], i_0r0d[24], gate575_0n, initialise);
  C2RI I118 (ifint_0n[25], i_0r0d[25], gate575_0n, initialise);
  C2RI I119 (ifint_0n[26], i_0r0d[26], gate575_0n, initialise);
  C2RI I120 (ifint_0n[27], i_0r0d[27], gate575_0n, initialise);
  C2RI I121 (ifint_0n[28], i_0r0d[28], gate575_0n, initialise);
  C2RI I122 (ifint_0n[29], i_0r0d[29], gate575_0n, initialise);
  C2RI I123 (ifint_0n[30], i_0r0d[30], gate575_0n, initialise);
  C2RI I124 (ifint_0n[31], i_0r0d[31], gate575_0n, initialise);
  C3 I125 (internal_0n[17], complete572_0n[0], complete572_0n[1], complete572_0n[2]);
  C3 I126 (internal_0n[18], complete572_0n[3], complete572_0n[4], complete572_0n[5]);
  C3 I127 (internal_0n[19], complete572_0n[6], complete572_0n[7], complete572_0n[8]);
  C3 I128 (internal_0n[20], complete572_0n[9], complete572_0n[10], complete572_0n[11]);
  C3 I129 (internal_0n[21], complete572_0n[12], complete572_0n[13], complete572_0n[14]);
  C3 I130 (internal_0n[22], complete572_0n[15], complete572_0n[16], complete572_0n[17]);
  C3 I131 (internal_0n[23], complete572_0n[18], complete572_0n[19], complete572_0n[20]);
  C3 I132 (internal_0n[24], complete572_0n[21], complete572_0n[22], complete572_0n[23]);
  C3 I133 (internal_0n[25], complete572_0n[24], complete572_0n[25], complete572_0n[26]);
  C3 I134 (internal_0n[26], complete572_0n[27], complete572_0n[28], complete572_0n[29]);
  C2 I135 (internal_0n[27], complete572_0n[30], complete572_0n[31]);
  C2 I136 (internal_0n[28], complete572_0n[32], complete572_0n[33]);
  C3 I137 (internal_0n[29], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I138 (internal_0n[30], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I139 (internal_0n[31], internal_0n[23], internal_0n[24], internal_0n[25]);
  C3 I140 (internal_0n[32], internal_0n[26], internal_0n[27], internal_0n[28]);
  C2 I141 (internal_0n[33], internal_0n[29], internal_0n[30]);
  C2 I142 (internal_0n[34], internal_0n[31], internal_0n[32]);
  C2 I143 (oaint_0n, internal_0n[33], internal_0n[34]);
  OR2 I144 (complete572_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I145 (complete572_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I146 (complete572_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I147 (complete572_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I148 (complete572_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I149 (complete572_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I150 (complete572_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I151 (complete572_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I152 (complete572_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I153 (complete572_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I154 (complete572_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I155 (complete572_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I156 (complete572_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I157 (complete572_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I158 (complete572_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I159 (complete572_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I160 (complete572_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I161 (complete572_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I162 (complete572_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I163 (complete572_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I164 (complete572_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I165 (complete572_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I166 (complete572_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I167 (complete572_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I168 (complete572_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I169 (complete572_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I170 (complete572_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I171 (complete572_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I172 (complete572_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I173 (complete572_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I174 (complete572_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I175 (complete572_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I176 (complete572_0n[32], o_0r0d[32], o_0r1d[32]);
  OR2 I177 (complete572_0n[33], o_0r0d[33], o_0r1d[33]);
  INV I178 (gate571_0n, o_0a);
  C2RI I179 (o_0r1d[0], otint_0n[0], gate571_0n, initialise);
  C2RI I180 (o_0r1d[1], otint_0n[1], gate571_0n, initialise);
  C2RI I181 (o_0r1d[2], otint_0n[2], gate571_0n, initialise);
  C2RI I182 (o_0r1d[3], otint_0n[3], gate571_0n, initialise);
  C2RI I183 (o_0r1d[4], otint_0n[4], gate571_0n, initialise);
  C2RI I184 (o_0r1d[5], otint_0n[5], gate571_0n, initialise);
  C2RI I185 (o_0r1d[6], otint_0n[6], gate571_0n, initialise);
  C2RI I186 (o_0r1d[7], otint_0n[7], gate571_0n, initialise);
  C2RI I187 (o_0r1d[8], otint_0n[8], gate571_0n, initialise);
  C2RI I188 (o_0r1d[9], otint_0n[9], gate571_0n, initialise);
  C2RI I189 (o_0r1d[10], otint_0n[10], gate571_0n, initialise);
  C2RI I190 (o_0r1d[11], otint_0n[11], gate571_0n, initialise);
  C2RI I191 (o_0r1d[12], otint_0n[12], gate571_0n, initialise);
  C2RI I192 (o_0r1d[13], otint_0n[13], gate571_0n, initialise);
  C2RI I193 (o_0r1d[14], otint_0n[14], gate571_0n, initialise);
  C2RI I194 (o_0r1d[15], otint_0n[15], gate571_0n, initialise);
  C2RI I195 (o_0r1d[16], otint_0n[16], gate571_0n, initialise);
  C2RI I196 (o_0r1d[17], otint_0n[17], gate571_0n, initialise);
  C2RI I197 (o_0r1d[18], otint_0n[18], gate571_0n, initialise);
  C2RI I198 (o_0r1d[19], otint_0n[19], gate571_0n, initialise);
  C2RI I199 (o_0r1d[20], otint_0n[20], gate571_0n, initialise);
  C2RI I200 (o_0r1d[21], otint_0n[21], gate571_0n, initialise);
  C2RI I201 (o_0r1d[22], otint_0n[22], gate571_0n, initialise);
  C2RI I202 (o_0r1d[23], otint_0n[23], gate571_0n, initialise);
  C2RI I203 (o_0r1d[24], otint_0n[24], gate571_0n, initialise);
  C2RI I204 (o_0r1d[25], otint_0n[25], gate571_0n, initialise);
  C2RI I205 (o_0r1d[26], otint_0n[26], gate571_0n, initialise);
  C2RI I206 (o_0r1d[27], otint_0n[27], gate571_0n, initialise);
  C2RI I207 (o_0r1d[28], otint_0n[28], gate571_0n, initialise);
  C2RI I208 (o_0r1d[29], otint_0n[29], gate571_0n, initialise);
  C2RI I209 (o_0r1d[30], otint_0n[30], gate571_0n, initialise);
  C2RI I210 (o_0r1d[31], otint_0n[31], gate571_0n, initialise);
  C2RI I211 (o_0r1d[32], otint_0n[32], gate571_0n, initialise);
  C2RI I212 (o_0r1d[33], otint_0n[33], gate571_0n, initialise);
  C2RI I213 (o_0r0d[0], ofint_0n[0], gate571_0n, initialise);
  C2RI I214 (o_0r0d[1], ofint_0n[1], gate571_0n, initialise);
  C2RI I215 (o_0r0d[2], ofint_0n[2], gate571_0n, initialise);
  C2RI I216 (o_0r0d[3], ofint_0n[3], gate571_0n, initialise);
  C2RI I217 (o_0r0d[4], ofint_0n[4], gate571_0n, initialise);
  C2RI I218 (o_0r0d[5], ofint_0n[5], gate571_0n, initialise);
  C2RI I219 (o_0r0d[6], ofint_0n[6], gate571_0n, initialise);
  C2RI I220 (o_0r0d[7], ofint_0n[7], gate571_0n, initialise);
  C2RI I221 (o_0r0d[8], ofint_0n[8], gate571_0n, initialise);
  C2RI I222 (o_0r0d[9], ofint_0n[9], gate571_0n, initialise);
  C2RI I223 (o_0r0d[10], ofint_0n[10], gate571_0n, initialise);
  C2RI I224 (o_0r0d[11], ofint_0n[11], gate571_0n, initialise);
  C2RI I225 (o_0r0d[12], ofint_0n[12], gate571_0n, initialise);
  C2RI I226 (o_0r0d[13], ofint_0n[13], gate571_0n, initialise);
  C2RI I227 (o_0r0d[14], ofint_0n[14], gate571_0n, initialise);
  C2RI I228 (o_0r0d[15], ofint_0n[15], gate571_0n, initialise);
  C2RI I229 (o_0r0d[16], ofint_0n[16], gate571_0n, initialise);
  C2RI I230 (o_0r0d[17], ofint_0n[17], gate571_0n, initialise);
  C2RI I231 (o_0r0d[18], ofint_0n[18], gate571_0n, initialise);
  C2RI I232 (o_0r0d[19], ofint_0n[19], gate571_0n, initialise);
  C2RI I233 (o_0r0d[20], ofint_0n[20], gate571_0n, initialise);
  C2RI I234 (o_0r0d[21], ofint_0n[21], gate571_0n, initialise);
  C2RI I235 (o_0r0d[22], ofint_0n[22], gate571_0n, initialise);
  C2RI I236 (o_0r0d[23], ofint_0n[23], gate571_0n, initialise);
  C2RI I237 (o_0r0d[24], ofint_0n[24], gate571_0n, initialise);
  C2RI I238 (o_0r0d[25], ofint_0n[25], gate571_0n, initialise);
  C2RI I239 (o_0r0d[26], ofint_0n[26], gate571_0n, initialise);
  C2RI I240 (o_0r0d[27], ofint_0n[27], gate571_0n, initialise);
  C2RI I241 (o_0r0d[28], ofint_0n[28], gate571_0n, initialise);
  C2RI I242 (o_0r0d[29], ofint_0n[29], gate571_0n, initialise);
  C2RI I243 (o_0r0d[30], ofint_0n[30], gate571_0n, initialise);
  C2RI I244 (o_0r0d[31], ofint_0n[31], gate571_0n, initialise);
  C2RI I245 (o_0r0d[32], ofint_0n[32], gate571_0n, initialise);
  C2RI I246 (o_0r0d[33], ofint_0n[33], gate571_0n, initialise);
  assign otint_0n[0] = itint_0n[0];
  assign otint_0n[1] = itint_0n[1];
  assign otint_0n[2] = itint_0n[2];
  assign otint_0n[3] = itint_0n[3];
  assign otint_0n[4] = itint_0n[4];
  assign otint_0n[5] = itint_0n[5];
  assign otint_0n[6] = itint_0n[6];
  assign otint_0n[7] = itint_0n[7];
  assign otint_0n[8] = itint_0n[8];
  assign otint_0n[9] = itint_0n[9];
  assign otint_0n[10] = itint_0n[10];
  assign otint_0n[11] = itint_0n[11];
  assign otint_0n[12] = itint_0n[12];
  assign otint_0n[13] = itint_0n[13];
  assign otint_0n[14] = itint_0n[14];
  assign otint_0n[15] = itint_0n[15];
  assign otint_0n[16] = itint_0n[16];
  assign otint_0n[17] = itint_0n[17];
  assign otint_0n[18] = itint_0n[18];
  assign otint_0n[19] = itint_0n[19];
  assign otint_0n[20] = itint_0n[20];
  assign otint_0n[21] = itint_0n[21];
  assign otint_0n[22] = itint_0n[22];
  assign otint_0n[23] = itint_0n[23];
  assign otint_0n[24] = itint_0n[24];
  assign otint_0n[25] = itint_0n[25];
  assign otint_0n[26] = itint_0n[26];
  assign otint_0n[27] = itint_0n[27];
  assign otint_0n[28] = itint_0n[28];
  assign otint_0n[29] = itint_0n[29];
  assign otint_0n[30] = itint_0n[30];
  assign otint_0n[31] = itint_0n[31];
  assign otint_0n[32] = itint_1n[0];
  assign otint_0n[33] = itint_1n[1];
  assign ofint_0n[0] = ifint_0n[0];
  assign ofint_0n[1] = ifint_0n[1];
  assign ofint_0n[2] = ifint_0n[2];
  assign ofint_0n[3] = ifint_0n[3];
  assign ofint_0n[4] = ifint_0n[4];
  assign ofint_0n[5] = ifint_0n[5];
  assign ofint_0n[6] = ifint_0n[6];
  assign ofint_0n[7] = ifint_0n[7];
  assign ofint_0n[8] = ifint_0n[8];
  assign ofint_0n[9] = ifint_0n[9];
  assign ofint_0n[10] = ifint_0n[10];
  assign ofint_0n[11] = ifint_0n[11];
  assign ofint_0n[12] = ifint_0n[12];
  assign ofint_0n[13] = ifint_0n[13];
  assign ofint_0n[14] = ifint_0n[14];
  assign ofint_0n[15] = ifint_0n[15];
  assign ofint_0n[16] = ifint_0n[16];
  assign ofint_0n[17] = ifint_0n[17];
  assign ofint_0n[18] = ifint_0n[18];
  assign ofint_0n[19] = ifint_0n[19];
  assign ofint_0n[20] = ifint_0n[20];
  assign ofint_0n[21] = ifint_0n[21];
  assign ofint_0n[22] = ifint_0n[22];
  assign ofint_0n[23] = ifint_0n[23];
  assign ofint_0n[24] = ifint_0n[24];
  assign ofint_0n[25] = ifint_0n[25];
  assign ofint_0n[26] = ifint_0n[26];
  assign ofint_0n[27] = ifint_0n[27];
  assign ofint_0n[28] = ifint_0n[28];
  assign ofint_0n[29] = ifint_0n[29];
  assign ofint_0n[30] = ifint_0n[30];
  assign ofint_0n[31] = ifint_0n[31];
  assign ofint_0n[32] = ifint_1n[0];
  assign ofint_0n[33] = ifint_1n[1];
endmodule

module BrzJ_l12__2832_203_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [31:0] i_0r0d;
  input [31:0] i_0r1d;
  output i_0a;
  input [2:0] i_1r0d;
  input [2:0] i_1r1d;
  output i_1a;
  output [34:0] o_0r0d;
  output [34:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [34:0] internal_0n;
  wire [34:0] ofint_0n;
  wire [34:0] otint_0n;
  wire oaint_0n;
  wire [31:0] ifint_0n;
  wire [2:0] ifint_1n;
  wire [31:0] itint_0n;
  wire [2:0] itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [2:0] complete592_0n;
  wire gate591_0n;
  wire [31:0] complete588_0n;
  wire gate587_0n;
  wire [34:0] complete584_0n;
  wire gate583_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  C3 I2 (i_1a, complete592_0n[0], complete592_0n[1], complete592_0n[2]);
  OR2 I3 (complete592_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I4 (complete592_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I5 (complete592_0n[2], ifint_1n[2], itint_1n[2]);
  INV I6 (gate591_0n, iaint_1n);
  C2RI I7 (itint_1n[0], i_1r1d[0], gate591_0n, initialise);
  C2RI I8 (itint_1n[1], i_1r1d[1], gate591_0n, initialise);
  C2RI I9 (itint_1n[2], i_1r1d[2], gate591_0n, initialise);
  C2RI I10 (ifint_1n[0], i_1r0d[0], gate591_0n, initialise);
  C2RI I11 (ifint_1n[1], i_1r0d[1], gate591_0n, initialise);
  C2RI I12 (ifint_1n[2], i_1r0d[2], gate591_0n, initialise);
  C3 I13 (internal_0n[0], complete588_0n[0], complete588_0n[1], complete588_0n[2]);
  C3 I14 (internal_0n[1], complete588_0n[3], complete588_0n[4], complete588_0n[5]);
  C3 I15 (internal_0n[2], complete588_0n[6], complete588_0n[7], complete588_0n[8]);
  C3 I16 (internal_0n[3], complete588_0n[9], complete588_0n[10], complete588_0n[11]);
  C3 I17 (internal_0n[4], complete588_0n[12], complete588_0n[13], complete588_0n[14]);
  C3 I18 (internal_0n[5], complete588_0n[15], complete588_0n[16], complete588_0n[17]);
  C3 I19 (internal_0n[6], complete588_0n[18], complete588_0n[19], complete588_0n[20]);
  C3 I20 (internal_0n[7], complete588_0n[21], complete588_0n[22], complete588_0n[23]);
  C3 I21 (internal_0n[8], complete588_0n[24], complete588_0n[25], complete588_0n[26]);
  C3 I22 (internal_0n[9], complete588_0n[27], complete588_0n[28], complete588_0n[29]);
  C2 I23 (internal_0n[10], complete588_0n[30], complete588_0n[31]);
  C3 I24 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I25 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I26 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I27 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I28 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I29 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I30 (i_0a, internal_0n[15], internal_0n[16]);
  OR2 I31 (complete588_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I32 (complete588_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I33 (complete588_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I34 (complete588_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I35 (complete588_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I36 (complete588_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I37 (complete588_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I38 (complete588_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I39 (complete588_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I40 (complete588_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I41 (complete588_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I42 (complete588_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I43 (complete588_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I44 (complete588_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I45 (complete588_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I46 (complete588_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I47 (complete588_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I48 (complete588_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I49 (complete588_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I50 (complete588_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I51 (complete588_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I52 (complete588_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I53 (complete588_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I54 (complete588_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I55 (complete588_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I56 (complete588_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I57 (complete588_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I58 (complete588_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I59 (complete588_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I60 (complete588_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I61 (complete588_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I62 (complete588_0n[31], ifint_0n[31], itint_0n[31]);
  INV I63 (gate587_0n, iaint_0n);
  C2RI I64 (itint_0n[0], i_0r1d[0], gate587_0n, initialise);
  C2RI I65 (itint_0n[1], i_0r1d[1], gate587_0n, initialise);
  C2RI I66 (itint_0n[2], i_0r1d[2], gate587_0n, initialise);
  C2RI I67 (itint_0n[3], i_0r1d[3], gate587_0n, initialise);
  C2RI I68 (itint_0n[4], i_0r1d[4], gate587_0n, initialise);
  C2RI I69 (itint_0n[5], i_0r1d[5], gate587_0n, initialise);
  C2RI I70 (itint_0n[6], i_0r1d[6], gate587_0n, initialise);
  C2RI I71 (itint_0n[7], i_0r1d[7], gate587_0n, initialise);
  C2RI I72 (itint_0n[8], i_0r1d[8], gate587_0n, initialise);
  C2RI I73 (itint_0n[9], i_0r1d[9], gate587_0n, initialise);
  C2RI I74 (itint_0n[10], i_0r1d[10], gate587_0n, initialise);
  C2RI I75 (itint_0n[11], i_0r1d[11], gate587_0n, initialise);
  C2RI I76 (itint_0n[12], i_0r1d[12], gate587_0n, initialise);
  C2RI I77 (itint_0n[13], i_0r1d[13], gate587_0n, initialise);
  C2RI I78 (itint_0n[14], i_0r1d[14], gate587_0n, initialise);
  C2RI I79 (itint_0n[15], i_0r1d[15], gate587_0n, initialise);
  C2RI I80 (itint_0n[16], i_0r1d[16], gate587_0n, initialise);
  C2RI I81 (itint_0n[17], i_0r1d[17], gate587_0n, initialise);
  C2RI I82 (itint_0n[18], i_0r1d[18], gate587_0n, initialise);
  C2RI I83 (itint_0n[19], i_0r1d[19], gate587_0n, initialise);
  C2RI I84 (itint_0n[20], i_0r1d[20], gate587_0n, initialise);
  C2RI I85 (itint_0n[21], i_0r1d[21], gate587_0n, initialise);
  C2RI I86 (itint_0n[22], i_0r1d[22], gate587_0n, initialise);
  C2RI I87 (itint_0n[23], i_0r1d[23], gate587_0n, initialise);
  C2RI I88 (itint_0n[24], i_0r1d[24], gate587_0n, initialise);
  C2RI I89 (itint_0n[25], i_0r1d[25], gate587_0n, initialise);
  C2RI I90 (itint_0n[26], i_0r1d[26], gate587_0n, initialise);
  C2RI I91 (itint_0n[27], i_0r1d[27], gate587_0n, initialise);
  C2RI I92 (itint_0n[28], i_0r1d[28], gate587_0n, initialise);
  C2RI I93 (itint_0n[29], i_0r1d[29], gate587_0n, initialise);
  C2RI I94 (itint_0n[30], i_0r1d[30], gate587_0n, initialise);
  C2RI I95 (itint_0n[31], i_0r1d[31], gate587_0n, initialise);
  C2RI I96 (ifint_0n[0], i_0r0d[0], gate587_0n, initialise);
  C2RI I97 (ifint_0n[1], i_0r0d[1], gate587_0n, initialise);
  C2RI I98 (ifint_0n[2], i_0r0d[2], gate587_0n, initialise);
  C2RI I99 (ifint_0n[3], i_0r0d[3], gate587_0n, initialise);
  C2RI I100 (ifint_0n[4], i_0r0d[4], gate587_0n, initialise);
  C2RI I101 (ifint_0n[5], i_0r0d[5], gate587_0n, initialise);
  C2RI I102 (ifint_0n[6], i_0r0d[6], gate587_0n, initialise);
  C2RI I103 (ifint_0n[7], i_0r0d[7], gate587_0n, initialise);
  C2RI I104 (ifint_0n[8], i_0r0d[8], gate587_0n, initialise);
  C2RI I105 (ifint_0n[9], i_0r0d[9], gate587_0n, initialise);
  C2RI I106 (ifint_0n[10], i_0r0d[10], gate587_0n, initialise);
  C2RI I107 (ifint_0n[11], i_0r0d[11], gate587_0n, initialise);
  C2RI I108 (ifint_0n[12], i_0r0d[12], gate587_0n, initialise);
  C2RI I109 (ifint_0n[13], i_0r0d[13], gate587_0n, initialise);
  C2RI I110 (ifint_0n[14], i_0r0d[14], gate587_0n, initialise);
  C2RI I111 (ifint_0n[15], i_0r0d[15], gate587_0n, initialise);
  C2RI I112 (ifint_0n[16], i_0r0d[16], gate587_0n, initialise);
  C2RI I113 (ifint_0n[17], i_0r0d[17], gate587_0n, initialise);
  C2RI I114 (ifint_0n[18], i_0r0d[18], gate587_0n, initialise);
  C2RI I115 (ifint_0n[19], i_0r0d[19], gate587_0n, initialise);
  C2RI I116 (ifint_0n[20], i_0r0d[20], gate587_0n, initialise);
  C2RI I117 (ifint_0n[21], i_0r0d[21], gate587_0n, initialise);
  C2RI I118 (ifint_0n[22], i_0r0d[22], gate587_0n, initialise);
  C2RI I119 (ifint_0n[23], i_0r0d[23], gate587_0n, initialise);
  C2RI I120 (ifint_0n[24], i_0r0d[24], gate587_0n, initialise);
  C2RI I121 (ifint_0n[25], i_0r0d[25], gate587_0n, initialise);
  C2RI I122 (ifint_0n[26], i_0r0d[26], gate587_0n, initialise);
  C2RI I123 (ifint_0n[27], i_0r0d[27], gate587_0n, initialise);
  C2RI I124 (ifint_0n[28], i_0r0d[28], gate587_0n, initialise);
  C2RI I125 (ifint_0n[29], i_0r0d[29], gate587_0n, initialise);
  C2RI I126 (ifint_0n[30], i_0r0d[30], gate587_0n, initialise);
  C2RI I127 (ifint_0n[31], i_0r0d[31], gate587_0n, initialise);
  C3 I128 (internal_0n[17], complete584_0n[0], complete584_0n[1], complete584_0n[2]);
  C3 I129 (internal_0n[18], complete584_0n[3], complete584_0n[4], complete584_0n[5]);
  C3 I130 (internal_0n[19], complete584_0n[6], complete584_0n[7], complete584_0n[8]);
  C3 I131 (internal_0n[20], complete584_0n[9], complete584_0n[10], complete584_0n[11]);
  C3 I132 (internal_0n[21], complete584_0n[12], complete584_0n[13], complete584_0n[14]);
  C3 I133 (internal_0n[22], complete584_0n[15], complete584_0n[16], complete584_0n[17]);
  C3 I134 (internal_0n[23], complete584_0n[18], complete584_0n[19], complete584_0n[20]);
  C3 I135 (internal_0n[24], complete584_0n[21], complete584_0n[22], complete584_0n[23]);
  C3 I136 (internal_0n[25], complete584_0n[24], complete584_0n[25], complete584_0n[26]);
  C3 I137 (internal_0n[26], complete584_0n[27], complete584_0n[28], complete584_0n[29]);
  C3 I138 (internal_0n[27], complete584_0n[30], complete584_0n[31], complete584_0n[32]);
  C2 I139 (internal_0n[28], complete584_0n[33], complete584_0n[34]);
  C3 I140 (internal_0n[29], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I141 (internal_0n[30], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I142 (internal_0n[31], internal_0n[23], internal_0n[24], internal_0n[25]);
  C3 I143 (internal_0n[32], internal_0n[26], internal_0n[27], internal_0n[28]);
  C2 I144 (internal_0n[33], internal_0n[29], internal_0n[30]);
  C2 I145 (internal_0n[34], internal_0n[31], internal_0n[32]);
  C2 I146 (oaint_0n, internal_0n[33], internal_0n[34]);
  OR2 I147 (complete584_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I148 (complete584_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I149 (complete584_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I150 (complete584_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I151 (complete584_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I152 (complete584_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I153 (complete584_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I154 (complete584_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I155 (complete584_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I156 (complete584_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I157 (complete584_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I158 (complete584_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I159 (complete584_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I160 (complete584_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I161 (complete584_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I162 (complete584_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I163 (complete584_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I164 (complete584_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I165 (complete584_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I166 (complete584_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I167 (complete584_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I168 (complete584_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I169 (complete584_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I170 (complete584_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I171 (complete584_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I172 (complete584_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I173 (complete584_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I174 (complete584_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I175 (complete584_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I176 (complete584_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I177 (complete584_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I178 (complete584_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I179 (complete584_0n[32], o_0r0d[32], o_0r1d[32]);
  OR2 I180 (complete584_0n[33], o_0r0d[33], o_0r1d[33]);
  OR2 I181 (complete584_0n[34], o_0r0d[34], o_0r1d[34]);
  INV I182 (gate583_0n, o_0a);
  C2RI I183 (o_0r1d[0], otint_0n[0], gate583_0n, initialise);
  C2RI I184 (o_0r1d[1], otint_0n[1], gate583_0n, initialise);
  C2RI I185 (o_0r1d[2], otint_0n[2], gate583_0n, initialise);
  C2RI I186 (o_0r1d[3], otint_0n[3], gate583_0n, initialise);
  C2RI I187 (o_0r1d[4], otint_0n[4], gate583_0n, initialise);
  C2RI I188 (o_0r1d[5], otint_0n[5], gate583_0n, initialise);
  C2RI I189 (o_0r1d[6], otint_0n[6], gate583_0n, initialise);
  C2RI I190 (o_0r1d[7], otint_0n[7], gate583_0n, initialise);
  C2RI I191 (o_0r1d[8], otint_0n[8], gate583_0n, initialise);
  C2RI I192 (o_0r1d[9], otint_0n[9], gate583_0n, initialise);
  C2RI I193 (o_0r1d[10], otint_0n[10], gate583_0n, initialise);
  C2RI I194 (o_0r1d[11], otint_0n[11], gate583_0n, initialise);
  C2RI I195 (o_0r1d[12], otint_0n[12], gate583_0n, initialise);
  C2RI I196 (o_0r1d[13], otint_0n[13], gate583_0n, initialise);
  C2RI I197 (o_0r1d[14], otint_0n[14], gate583_0n, initialise);
  C2RI I198 (o_0r1d[15], otint_0n[15], gate583_0n, initialise);
  C2RI I199 (o_0r1d[16], otint_0n[16], gate583_0n, initialise);
  C2RI I200 (o_0r1d[17], otint_0n[17], gate583_0n, initialise);
  C2RI I201 (o_0r1d[18], otint_0n[18], gate583_0n, initialise);
  C2RI I202 (o_0r1d[19], otint_0n[19], gate583_0n, initialise);
  C2RI I203 (o_0r1d[20], otint_0n[20], gate583_0n, initialise);
  C2RI I204 (o_0r1d[21], otint_0n[21], gate583_0n, initialise);
  C2RI I205 (o_0r1d[22], otint_0n[22], gate583_0n, initialise);
  C2RI I206 (o_0r1d[23], otint_0n[23], gate583_0n, initialise);
  C2RI I207 (o_0r1d[24], otint_0n[24], gate583_0n, initialise);
  C2RI I208 (o_0r1d[25], otint_0n[25], gate583_0n, initialise);
  C2RI I209 (o_0r1d[26], otint_0n[26], gate583_0n, initialise);
  C2RI I210 (o_0r1d[27], otint_0n[27], gate583_0n, initialise);
  C2RI I211 (o_0r1d[28], otint_0n[28], gate583_0n, initialise);
  C2RI I212 (o_0r1d[29], otint_0n[29], gate583_0n, initialise);
  C2RI I213 (o_0r1d[30], otint_0n[30], gate583_0n, initialise);
  C2RI I214 (o_0r1d[31], otint_0n[31], gate583_0n, initialise);
  C2RI I215 (o_0r1d[32], otint_0n[32], gate583_0n, initialise);
  C2RI I216 (o_0r1d[33], otint_0n[33], gate583_0n, initialise);
  C2RI I217 (o_0r1d[34], otint_0n[34], gate583_0n, initialise);
  C2RI I218 (o_0r0d[0], ofint_0n[0], gate583_0n, initialise);
  C2RI I219 (o_0r0d[1], ofint_0n[1], gate583_0n, initialise);
  C2RI I220 (o_0r0d[2], ofint_0n[2], gate583_0n, initialise);
  C2RI I221 (o_0r0d[3], ofint_0n[3], gate583_0n, initialise);
  C2RI I222 (o_0r0d[4], ofint_0n[4], gate583_0n, initialise);
  C2RI I223 (o_0r0d[5], ofint_0n[5], gate583_0n, initialise);
  C2RI I224 (o_0r0d[6], ofint_0n[6], gate583_0n, initialise);
  C2RI I225 (o_0r0d[7], ofint_0n[7], gate583_0n, initialise);
  C2RI I226 (o_0r0d[8], ofint_0n[8], gate583_0n, initialise);
  C2RI I227 (o_0r0d[9], ofint_0n[9], gate583_0n, initialise);
  C2RI I228 (o_0r0d[10], ofint_0n[10], gate583_0n, initialise);
  C2RI I229 (o_0r0d[11], ofint_0n[11], gate583_0n, initialise);
  C2RI I230 (o_0r0d[12], ofint_0n[12], gate583_0n, initialise);
  C2RI I231 (o_0r0d[13], ofint_0n[13], gate583_0n, initialise);
  C2RI I232 (o_0r0d[14], ofint_0n[14], gate583_0n, initialise);
  C2RI I233 (o_0r0d[15], ofint_0n[15], gate583_0n, initialise);
  C2RI I234 (o_0r0d[16], ofint_0n[16], gate583_0n, initialise);
  C2RI I235 (o_0r0d[17], ofint_0n[17], gate583_0n, initialise);
  C2RI I236 (o_0r0d[18], ofint_0n[18], gate583_0n, initialise);
  C2RI I237 (o_0r0d[19], ofint_0n[19], gate583_0n, initialise);
  C2RI I238 (o_0r0d[20], ofint_0n[20], gate583_0n, initialise);
  C2RI I239 (o_0r0d[21], ofint_0n[21], gate583_0n, initialise);
  C2RI I240 (o_0r0d[22], ofint_0n[22], gate583_0n, initialise);
  C2RI I241 (o_0r0d[23], ofint_0n[23], gate583_0n, initialise);
  C2RI I242 (o_0r0d[24], ofint_0n[24], gate583_0n, initialise);
  C2RI I243 (o_0r0d[25], ofint_0n[25], gate583_0n, initialise);
  C2RI I244 (o_0r0d[26], ofint_0n[26], gate583_0n, initialise);
  C2RI I245 (o_0r0d[27], ofint_0n[27], gate583_0n, initialise);
  C2RI I246 (o_0r0d[28], ofint_0n[28], gate583_0n, initialise);
  C2RI I247 (o_0r0d[29], ofint_0n[29], gate583_0n, initialise);
  C2RI I248 (o_0r0d[30], ofint_0n[30], gate583_0n, initialise);
  C2RI I249 (o_0r0d[31], ofint_0n[31], gate583_0n, initialise);
  C2RI I250 (o_0r0d[32], ofint_0n[32], gate583_0n, initialise);
  C2RI I251 (o_0r0d[33], ofint_0n[33], gate583_0n, initialise);
  C2RI I252 (o_0r0d[34], ofint_0n[34], gate583_0n, initialise);
  assign otint_0n[0] = itint_0n[0];
  assign otint_0n[1] = itint_0n[1];
  assign otint_0n[2] = itint_0n[2];
  assign otint_0n[3] = itint_0n[3];
  assign otint_0n[4] = itint_0n[4];
  assign otint_0n[5] = itint_0n[5];
  assign otint_0n[6] = itint_0n[6];
  assign otint_0n[7] = itint_0n[7];
  assign otint_0n[8] = itint_0n[8];
  assign otint_0n[9] = itint_0n[9];
  assign otint_0n[10] = itint_0n[10];
  assign otint_0n[11] = itint_0n[11];
  assign otint_0n[12] = itint_0n[12];
  assign otint_0n[13] = itint_0n[13];
  assign otint_0n[14] = itint_0n[14];
  assign otint_0n[15] = itint_0n[15];
  assign otint_0n[16] = itint_0n[16];
  assign otint_0n[17] = itint_0n[17];
  assign otint_0n[18] = itint_0n[18];
  assign otint_0n[19] = itint_0n[19];
  assign otint_0n[20] = itint_0n[20];
  assign otint_0n[21] = itint_0n[21];
  assign otint_0n[22] = itint_0n[22];
  assign otint_0n[23] = itint_0n[23];
  assign otint_0n[24] = itint_0n[24];
  assign otint_0n[25] = itint_0n[25];
  assign otint_0n[26] = itint_0n[26];
  assign otint_0n[27] = itint_0n[27];
  assign otint_0n[28] = itint_0n[28];
  assign otint_0n[29] = itint_0n[29];
  assign otint_0n[30] = itint_0n[30];
  assign otint_0n[31] = itint_0n[31];
  assign otint_0n[32] = itint_1n[0];
  assign otint_0n[33] = itint_1n[1];
  assign otint_0n[34] = itint_1n[2];
  assign ofint_0n[0] = ifint_0n[0];
  assign ofint_0n[1] = ifint_0n[1];
  assign ofint_0n[2] = ifint_0n[2];
  assign ofint_0n[3] = ifint_0n[3];
  assign ofint_0n[4] = ifint_0n[4];
  assign ofint_0n[5] = ifint_0n[5];
  assign ofint_0n[6] = ifint_0n[6];
  assign ofint_0n[7] = ifint_0n[7];
  assign ofint_0n[8] = ifint_0n[8];
  assign ofint_0n[9] = ifint_0n[9];
  assign ofint_0n[10] = ifint_0n[10];
  assign ofint_0n[11] = ifint_0n[11];
  assign ofint_0n[12] = ifint_0n[12];
  assign ofint_0n[13] = ifint_0n[13];
  assign ofint_0n[14] = ifint_0n[14];
  assign ofint_0n[15] = ifint_0n[15];
  assign ofint_0n[16] = ifint_0n[16];
  assign ofint_0n[17] = ifint_0n[17];
  assign ofint_0n[18] = ifint_0n[18];
  assign ofint_0n[19] = ifint_0n[19];
  assign ofint_0n[20] = ifint_0n[20];
  assign ofint_0n[21] = ifint_0n[21];
  assign ofint_0n[22] = ifint_0n[22];
  assign ofint_0n[23] = ifint_0n[23];
  assign ofint_0n[24] = ifint_0n[24];
  assign ofint_0n[25] = ifint_0n[25];
  assign ofint_0n[26] = ifint_0n[26];
  assign ofint_0n[27] = ifint_0n[27];
  assign ofint_0n[28] = ifint_0n[28];
  assign ofint_0n[29] = ifint_0n[29];
  assign ofint_0n[30] = ifint_0n[30];
  assign ofint_0n[31] = ifint_0n[31];
  assign ofint_0n[32] = ifint_1n[0];
  assign ofint_0n[33] = ifint_1n[1];
  assign ofint_0n[34] = ifint_1n[2];
endmodule

module BrzJ_l12__2833_200_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [32:0] i_0r0d;
  input [32:0] i_0r1d;
  output i_0a;
  input i_1r;
  output i_1a;
  output [32:0] o_0r0d;
  output [32:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [33:0] internal_0n;
  wire [32:0] ofint_0n;
  wire [32:0] otint_0n;
  wire oaint_0n;
  wire [32:0] ifint_0n;
  wire ifint_1n;
  wire [32:0] itint_0n;
  wire iaint_0n;
  wire iaint_1n;
  wire gate603_0n;
  wire [32:0] complete600_0n;
  wire gate599_0n;
  wire [32:0] complete596_0n;
  wire gate595_0n;
  wire [32:0] joint_0n;
  wire [32:0] joinf_0n;
  wire icomplete_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign i_1a = ifint_1n;
  INV I3 (gate603_0n, iaint_1n);
  C2RI I4 (ifint_1n, i_1r, gate603_0n, initialise);
  C3 I5 (internal_0n[0], complete600_0n[0], complete600_0n[1], complete600_0n[2]);
  C3 I6 (internal_0n[1], complete600_0n[3], complete600_0n[4], complete600_0n[5]);
  C3 I7 (internal_0n[2], complete600_0n[6], complete600_0n[7], complete600_0n[8]);
  C3 I8 (internal_0n[3], complete600_0n[9], complete600_0n[10], complete600_0n[11]);
  C3 I9 (internal_0n[4], complete600_0n[12], complete600_0n[13], complete600_0n[14]);
  C3 I10 (internal_0n[5], complete600_0n[15], complete600_0n[16], complete600_0n[17]);
  C3 I11 (internal_0n[6], complete600_0n[18], complete600_0n[19], complete600_0n[20]);
  C3 I12 (internal_0n[7], complete600_0n[21], complete600_0n[22], complete600_0n[23]);
  C3 I13 (internal_0n[8], complete600_0n[24], complete600_0n[25], complete600_0n[26]);
  C3 I14 (internal_0n[9], complete600_0n[27], complete600_0n[28], complete600_0n[29]);
  C3 I15 (internal_0n[10], complete600_0n[30], complete600_0n[31], complete600_0n[32]);
  C3 I16 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I17 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I18 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I19 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I20 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I21 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I22 (i_0a, internal_0n[15], internal_0n[16]);
  OR2 I23 (complete600_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I24 (complete600_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I25 (complete600_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I26 (complete600_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I27 (complete600_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I28 (complete600_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I29 (complete600_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I30 (complete600_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I31 (complete600_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I32 (complete600_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I33 (complete600_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I34 (complete600_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I35 (complete600_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I36 (complete600_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I37 (complete600_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I38 (complete600_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I39 (complete600_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I40 (complete600_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I41 (complete600_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I42 (complete600_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I43 (complete600_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I44 (complete600_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I45 (complete600_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I46 (complete600_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I47 (complete600_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I48 (complete600_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I49 (complete600_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I50 (complete600_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I51 (complete600_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I52 (complete600_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I53 (complete600_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I54 (complete600_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I55 (complete600_0n[32], ifint_0n[32], itint_0n[32]);
  INV I56 (gate599_0n, iaint_0n);
  C2RI I57 (itint_0n[0], i_0r1d[0], gate599_0n, initialise);
  C2RI I58 (itint_0n[1], i_0r1d[1], gate599_0n, initialise);
  C2RI I59 (itint_0n[2], i_0r1d[2], gate599_0n, initialise);
  C2RI I60 (itint_0n[3], i_0r1d[3], gate599_0n, initialise);
  C2RI I61 (itint_0n[4], i_0r1d[4], gate599_0n, initialise);
  C2RI I62 (itint_0n[5], i_0r1d[5], gate599_0n, initialise);
  C2RI I63 (itint_0n[6], i_0r1d[6], gate599_0n, initialise);
  C2RI I64 (itint_0n[7], i_0r1d[7], gate599_0n, initialise);
  C2RI I65 (itint_0n[8], i_0r1d[8], gate599_0n, initialise);
  C2RI I66 (itint_0n[9], i_0r1d[9], gate599_0n, initialise);
  C2RI I67 (itint_0n[10], i_0r1d[10], gate599_0n, initialise);
  C2RI I68 (itint_0n[11], i_0r1d[11], gate599_0n, initialise);
  C2RI I69 (itint_0n[12], i_0r1d[12], gate599_0n, initialise);
  C2RI I70 (itint_0n[13], i_0r1d[13], gate599_0n, initialise);
  C2RI I71 (itint_0n[14], i_0r1d[14], gate599_0n, initialise);
  C2RI I72 (itint_0n[15], i_0r1d[15], gate599_0n, initialise);
  C2RI I73 (itint_0n[16], i_0r1d[16], gate599_0n, initialise);
  C2RI I74 (itint_0n[17], i_0r1d[17], gate599_0n, initialise);
  C2RI I75 (itint_0n[18], i_0r1d[18], gate599_0n, initialise);
  C2RI I76 (itint_0n[19], i_0r1d[19], gate599_0n, initialise);
  C2RI I77 (itint_0n[20], i_0r1d[20], gate599_0n, initialise);
  C2RI I78 (itint_0n[21], i_0r1d[21], gate599_0n, initialise);
  C2RI I79 (itint_0n[22], i_0r1d[22], gate599_0n, initialise);
  C2RI I80 (itint_0n[23], i_0r1d[23], gate599_0n, initialise);
  C2RI I81 (itint_0n[24], i_0r1d[24], gate599_0n, initialise);
  C2RI I82 (itint_0n[25], i_0r1d[25], gate599_0n, initialise);
  C2RI I83 (itint_0n[26], i_0r1d[26], gate599_0n, initialise);
  C2RI I84 (itint_0n[27], i_0r1d[27], gate599_0n, initialise);
  C2RI I85 (itint_0n[28], i_0r1d[28], gate599_0n, initialise);
  C2RI I86 (itint_0n[29], i_0r1d[29], gate599_0n, initialise);
  C2RI I87 (itint_0n[30], i_0r1d[30], gate599_0n, initialise);
  C2RI I88 (itint_0n[31], i_0r1d[31], gate599_0n, initialise);
  C2RI I89 (itint_0n[32], i_0r1d[32], gate599_0n, initialise);
  C2RI I90 (ifint_0n[0], i_0r0d[0], gate599_0n, initialise);
  C2RI I91 (ifint_0n[1], i_0r0d[1], gate599_0n, initialise);
  C2RI I92 (ifint_0n[2], i_0r0d[2], gate599_0n, initialise);
  C2RI I93 (ifint_0n[3], i_0r0d[3], gate599_0n, initialise);
  C2RI I94 (ifint_0n[4], i_0r0d[4], gate599_0n, initialise);
  C2RI I95 (ifint_0n[5], i_0r0d[5], gate599_0n, initialise);
  C2RI I96 (ifint_0n[6], i_0r0d[6], gate599_0n, initialise);
  C2RI I97 (ifint_0n[7], i_0r0d[7], gate599_0n, initialise);
  C2RI I98 (ifint_0n[8], i_0r0d[8], gate599_0n, initialise);
  C2RI I99 (ifint_0n[9], i_0r0d[9], gate599_0n, initialise);
  C2RI I100 (ifint_0n[10], i_0r0d[10], gate599_0n, initialise);
  C2RI I101 (ifint_0n[11], i_0r0d[11], gate599_0n, initialise);
  C2RI I102 (ifint_0n[12], i_0r0d[12], gate599_0n, initialise);
  C2RI I103 (ifint_0n[13], i_0r0d[13], gate599_0n, initialise);
  C2RI I104 (ifint_0n[14], i_0r0d[14], gate599_0n, initialise);
  C2RI I105 (ifint_0n[15], i_0r0d[15], gate599_0n, initialise);
  C2RI I106 (ifint_0n[16], i_0r0d[16], gate599_0n, initialise);
  C2RI I107 (ifint_0n[17], i_0r0d[17], gate599_0n, initialise);
  C2RI I108 (ifint_0n[18], i_0r0d[18], gate599_0n, initialise);
  C2RI I109 (ifint_0n[19], i_0r0d[19], gate599_0n, initialise);
  C2RI I110 (ifint_0n[20], i_0r0d[20], gate599_0n, initialise);
  C2RI I111 (ifint_0n[21], i_0r0d[21], gate599_0n, initialise);
  C2RI I112 (ifint_0n[22], i_0r0d[22], gate599_0n, initialise);
  C2RI I113 (ifint_0n[23], i_0r0d[23], gate599_0n, initialise);
  C2RI I114 (ifint_0n[24], i_0r0d[24], gate599_0n, initialise);
  C2RI I115 (ifint_0n[25], i_0r0d[25], gate599_0n, initialise);
  C2RI I116 (ifint_0n[26], i_0r0d[26], gate599_0n, initialise);
  C2RI I117 (ifint_0n[27], i_0r0d[27], gate599_0n, initialise);
  C2RI I118 (ifint_0n[28], i_0r0d[28], gate599_0n, initialise);
  C2RI I119 (ifint_0n[29], i_0r0d[29], gate599_0n, initialise);
  C2RI I120 (ifint_0n[30], i_0r0d[30], gate599_0n, initialise);
  C2RI I121 (ifint_0n[31], i_0r0d[31], gate599_0n, initialise);
  C2RI I122 (ifint_0n[32], i_0r0d[32], gate599_0n, initialise);
  C3 I123 (internal_0n[17], complete596_0n[0], complete596_0n[1], complete596_0n[2]);
  C3 I124 (internal_0n[18], complete596_0n[3], complete596_0n[4], complete596_0n[5]);
  C3 I125 (internal_0n[19], complete596_0n[6], complete596_0n[7], complete596_0n[8]);
  C3 I126 (internal_0n[20], complete596_0n[9], complete596_0n[10], complete596_0n[11]);
  C3 I127 (internal_0n[21], complete596_0n[12], complete596_0n[13], complete596_0n[14]);
  C3 I128 (internal_0n[22], complete596_0n[15], complete596_0n[16], complete596_0n[17]);
  C3 I129 (internal_0n[23], complete596_0n[18], complete596_0n[19], complete596_0n[20]);
  C3 I130 (internal_0n[24], complete596_0n[21], complete596_0n[22], complete596_0n[23]);
  C3 I131 (internal_0n[25], complete596_0n[24], complete596_0n[25], complete596_0n[26]);
  C3 I132 (internal_0n[26], complete596_0n[27], complete596_0n[28], complete596_0n[29]);
  C3 I133 (internal_0n[27], complete596_0n[30], complete596_0n[31], complete596_0n[32]);
  C3 I134 (internal_0n[28], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I135 (internal_0n[29], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I136 (internal_0n[30], internal_0n[23], internal_0n[24], internal_0n[25]);
  C2 I137 (internal_0n[31], internal_0n[26], internal_0n[27]);
  C2 I138 (internal_0n[32], internal_0n[28], internal_0n[29]);
  C2 I139 (internal_0n[33], internal_0n[30], internal_0n[31]);
  C2 I140 (oaint_0n, internal_0n[32], internal_0n[33]);
  OR2 I141 (complete596_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I142 (complete596_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I143 (complete596_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I144 (complete596_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I145 (complete596_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I146 (complete596_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I147 (complete596_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I148 (complete596_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I149 (complete596_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I150 (complete596_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I151 (complete596_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I152 (complete596_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I153 (complete596_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I154 (complete596_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I155 (complete596_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I156 (complete596_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I157 (complete596_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I158 (complete596_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I159 (complete596_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I160 (complete596_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I161 (complete596_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I162 (complete596_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I163 (complete596_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I164 (complete596_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I165 (complete596_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I166 (complete596_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I167 (complete596_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I168 (complete596_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I169 (complete596_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I170 (complete596_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I171 (complete596_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I172 (complete596_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I173 (complete596_0n[32], o_0r0d[32], o_0r1d[32]);
  INV I174 (gate595_0n, o_0a);
  C2RI I175 (o_0r1d[0], otint_0n[0], gate595_0n, initialise);
  C2RI I176 (o_0r1d[1], otint_0n[1], gate595_0n, initialise);
  C2RI I177 (o_0r1d[2], otint_0n[2], gate595_0n, initialise);
  C2RI I178 (o_0r1d[3], otint_0n[3], gate595_0n, initialise);
  C2RI I179 (o_0r1d[4], otint_0n[4], gate595_0n, initialise);
  C2RI I180 (o_0r1d[5], otint_0n[5], gate595_0n, initialise);
  C2RI I181 (o_0r1d[6], otint_0n[6], gate595_0n, initialise);
  C2RI I182 (o_0r1d[7], otint_0n[7], gate595_0n, initialise);
  C2RI I183 (o_0r1d[8], otint_0n[8], gate595_0n, initialise);
  C2RI I184 (o_0r1d[9], otint_0n[9], gate595_0n, initialise);
  C2RI I185 (o_0r1d[10], otint_0n[10], gate595_0n, initialise);
  C2RI I186 (o_0r1d[11], otint_0n[11], gate595_0n, initialise);
  C2RI I187 (o_0r1d[12], otint_0n[12], gate595_0n, initialise);
  C2RI I188 (o_0r1d[13], otint_0n[13], gate595_0n, initialise);
  C2RI I189 (o_0r1d[14], otint_0n[14], gate595_0n, initialise);
  C2RI I190 (o_0r1d[15], otint_0n[15], gate595_0n, initialise);
  C2RI I191 (o_0r1d[16], otint_0n[16], gate595_0n, initialise);
  C2RI I192 (o_0r1d[17], otint_0n[17], gate595_0n, initialise);
  C2RI I193 (o_0r1d[18], otint_0n[18], gate595_0n, initialise);
  C2RI I194 (o_0r1d[19], otint_0n[19], gate595_0n, initialise);
  C2RI I195 (o_0r1d[20], otint_0n[20], gate595_0n, initialise);
  C2RI I196 (o_0r1d[21], otint_0n[21], gate595_0n, initialise);
  C2RI I197 (o_0r1d[22], otint_0n[22], gate595_0n, initialise);
  C2RI I198 (o_0r1d[23], otint_0n[23], gate595_0n, initialise);
  C2RI I199 (o_0r1d[24], otint_0n[24], gate595_0n, initialise);
  C2RI I200 (o_0r1d[25], otint_0n[25], gate595_0n, initialise);
  C2RI I201 (o_0r1d[26], otint_0n[26], gate595_0n, initialise);
  C2RI I202 (o_0r1d[27], otint_0n[27], gate595_0n, initialise);
  C2RI I203 (o_0r1d[28], otint_0n[28], gate595_0n, initialise);
  C2RI I204 (o_0r1d[29], otint_0n[29], gate595_0n, initialise);
  C2RI I205 (o_0r1d[30], otint_0n[30], gate595_0n, initialise);
  C2RI I206 (o_0r1d[31], otint_0n[31], gate595_0n, initialise);
  C2RI I207 (o_0r1d[32], otint_0n[32], gate595_0n, initialise);
  C2RI I208 (o_0r0d[0], ofint_0n[0], gate595_0n, initialise);
  C2RI I209 (o_0r0d[1], ofint_0n[1], gate595_0n, initialise);
  C2RI I210 (o_0r0d[2], ofint_0n[2], gate595_0n, initialise);
  C2RI I211 (o_0r0d[3], ofint_0n[3], gate595_0n, initialise);
  C2RI I212 (o_0r0d[4], ofint_0n[4], gate595_0n, initialise);
  C2RI I213 (o_0r0d[5], ofint_0n[5], gate595_0n, initialise);
  C2RI I214 (o_0r0d[6], ofint_0n[6], gate595_0n, initialise);
  C2RI I215 (o_0r0d[7], ofint_0n[7], gate595_0n, initialise);
  C2RI I216 (o_0r0d[8], ofint_0n[8], gate595_0n, initialise);
  C2RI I217 (o_0r0d[9], ofint_0n[9], gate595_0n, initialise);
  C2RI I218 (o_0r0d[10], ofint_0n[10], gate595_0n, initialise);
  C2RI I219 (o_0r0d[11], ofint_0n[11], gate595_0n, initialise);
  C2RI I220 (o_0r0d[12], ofint_0n[12], gate595_0n, initialise);
  C2RI I221 (o_0r0d[13], ofint_0n[13], gate595_0n, initialise);
  C2RI I222 (o_0r0d[14], ofint_0n[14], gate595_0n, initialise);
  C2RI I223 (o_0r0d[15], ofint_0n[15], gate595_0n, initialise);
  C2RI I224 (o_0r0d[16], ofint_0n[16], gate595_0n, initialise);
  C2RI I225 (o_0r0d[17], ofint_0n[17], gate595_0n, initialise);
  C2RI I226 (o_0r0d[18], ofint_0n[18], gate595_0n, initialise);
  C2RI I227 (o_0r0d[19], ofint_0n[19], gate595_0n, initialise);
  C2RI I228 (o_0r0d[20], ofint_0n[20], gate595_0n, initialise);
  C2RI I229 (o_0r0d[21], ofint_0n[21], gate595_0n, initialise);
  C2RI I230 (o_0r0d[22], ofint_0n[22], gate595_0n, initialise);
  C2RI I231 (o_0r0d[23], ofint_0n[23], gate595_0n, initialise);
  C2RI I232 (o_0r0d[24], ofint_0n[24], gate595_0n, initialise);
  C2RI I233 (o_0r0d[25], ofint_0n[25], gate595_0n, initialise);
  C2RI I234 (o_0r0d[26], ofint_0n[26], gate595_0n, initialise);
  C2RI I235 (o_0r0d[27], ofint_0n[27], gate595_0n, initialise);
  C2RI I236 (o_0r0d[28], ofint_0n[28], gate595_0n, initialise);
  C2RI I237 (o_0r0d[29], ofint_0n[29], gate595_0n, initialise);
  C2RI I238 (o_0r0d[30], ofint_0n[30], gate595_0n, initialise);
  C2RI I239 (o_0r0d[31], ofint_0n[31], gate595_0n, initialise);
  C2RI I240 (o_0r0d[32], ofint_0n[32], gate595_0n, initialise);
  assign otint_0n[1] = joint_0n[1];
  assign otint_0n[2] = joint_0n[2];
  assign otint_0n[3] = joint_0n[3];
  assign otint_0n[4] = joint_0n[4];
  assign otint_0n[5] = joint_0n[5];
  assign otint_0n[6] = joint_0n[6];
  assign otint_0n[7] = joint_0n[7];
  assign otint_0n[8] = joint_0n[8];
  assign otint_0n[9] = joint_0n[9];
  assign otint_0n[10] = joint_0n[10];
  assign otint_0n[11] = joint_0n[11];
  assign otint_0n[12] = joint_0n[12];
  assign otint_0n[13] = joint_0n[13];
  assign otint_0n[14] = joint_0n[14];
  assign otint_0n[15] = joint_0n[15];
  assign otint_0n[16] = joint_0n[16];
  assign otint_0n[17] = joint_0n[17];
  assign otint_0n[18] = joint_0n[18];
  assign otint_0n[19] = joint_0n[19];
  assign otint_0n[20] = joint_0n[20];
  assign otint_0n[21] = joint_0n[21];
  assign otint_0n[22] = joint_0n[22];
  assign otint_0n[23] = joint_0n[23];
  assign otint_0n[24] = joint_0n[24];
  assign otint_0n[25] = joint_0n[25];
  assign otint_0n[26] = joint_0n[26];
  assign otint_0n[27] = joint_0n[27];
  assign otint_0n[28] = joint_0n[28];
  assign otint_0n[29] = joint_0n[29];
  assign otint_0n[30] = joint_0n[30];
  assign otint_0n[31] = joint_0n[31];
  assign otint_0n[32] = joint_0n[32];
  assign ofint_0n[1] = joinf_0n[1];
  assign ofint_0n[2] = joinf_0n[2];
  assign ofint_0n[3] = joinf_0n[3];
  assign ofint_0n[4] = joinf_0n[4];
  assign ofint_0n[5] = joinf_0n[5];
  assign ofint_0n[6] = joinf_0n[6];
  assign ofint_0n[7] = joinf_0n[7];
  assign ofint_0n[8] = joinf_0n[8];
  assign ofint_0n[9] = joinf_0n[9];
  assign ofint_0n[10] = joinf_0n[10];
  assign ofint_0n[11] = joinf_0n[11];
  assign ofint_0n[12] = joinf_0n[12];
  assign ofint_0n[13] = joinf_0n[13];
  assign ofint_0n[14] = joinf_0n[14];
  assign ofint_0n[15] = joinf_0n[15];
  assign ofint_0n[16] = joinf_0n[16];
  assign ofint_0n[17] = joinf_0n[17];
  assign ofint_0n[18] = joinf_0n[18];
  assign ofint_0n[19] = joinf_0n[19];
  assign ofint_0n[20] = joinf_0n[20];
  assign ofint_0n[21] = joinf_0n[21];
  assign ofint_0n[22] = joinf_0n[22];
  assign ofint_0n[23] = joinf_0n[23];
  assign ofint_0n[24] = joinf_0n[24];
  assign ofint_0n[25] = joinf_0n[25];
  assign ofint_0n[26] = joinf_0n[26];
  assign ofint_0n[27] = joinf_0n[27];
  assign ofint_0n[28] = joinf_0n[28];
  assign ofint_0n[29] = joinf_0n[29];
  assign ofint_0n[30] = joinf_0n[30];
  assign ofint_0n[31] = joinf_0n[31];
  assign ofint_0n[32] = joinf_0n[32];
  C2 I305 (otint_0n[0], joint_0n[0], icomplete_0n);
  C2 I306 (ofint_0n[0], joinf_0n[0], icomplete_0n);
  assign icomplete_0n = ifint_1n;
  assign joint_0n[0] = itint_0n[0];
  assign joint_0n[1] = itint_0n[1];
  assign joint_0n[2] = itint_0n[2];
  assign joint_0n[3] = itint_0n[3];
  assign joint_0n[4] = itint_0n[4];
  assign joint_0n[5] = itint_0n[5];
  assign joint_0n[6] = itint_0n[6];
  assign joint_0n[7] = itint_0n[7];
  assign joint_0n[8] = itint_0n[8];
  assign joint_0n[9] = itint_0n[9];
  assign joint_0n[10] = itint_0n[10];
  assign joint_0n[11] = itint_0n[11];
  assign joint_0n[12] = itint_0n[12];
  assign joint_0n[13] = itint_0n[13];
  assign joint_0n[14] = itint_0n[14];
  assign joint_0n[15] = itint_0n[15];
  assign joint_0n[16] = itint_0n[16];
  assign joint_0n[17] = itint_0n[17];
  assign joint_0n[18] = itint_0n[18];
  assign joint_0n[19] = itint_0n[19];
  assign joint_0n[20] = itint_0n[20];
  assign joint_0n[21] = itint_0n[21];
  assign joint_0n[22] = itint_0n[22];
  assign joint_0n[23] = itint_0n[23];
  assign joint_0n[24] = itint_0n[24];
  assign joint_0n[25] = itint_0n[25];
  assign joint_0n[26] = itint_0n[26];
  assign joint_0n[27] = itint_0n[27];
  assign joint_0n[28] = itint_0n[28];
  assign joint_0n[29] = itint_0n[29];
  assign joint_0n[30] = itint_0n[30];
  assign joint_0n[31] = itint_0n[31];
  assign joint_0n[32] = itint_0n[32];
  assign joinf_0n[0] = ifint_0n[0];
  assign joinf_0n[1] = ifint_0n[1];
  assign joinf_0n[2] = ifint_0n[2];
  assign joinf_0n[3] = ifint_0n[3];
  assign joinf_0n[4] = ifint_0n[4];
  assign joinf_0n[5] = ifint_0n[5];
  assign joinf_0n[6] = ifint_0n[6];
  assign joinf_0n[7] = ifint_0n[7];
  assign joinf_0n[8] = ifint_0n[8];
  assign joinf_0n[9] = ifint_0n[9];
  assign joinf_0n[10] = ifint_0n[10];
  assign joinf_0n[11] = ifint_0n[11];
  assign joinf_0n[12] = ifint_0n[12];
  assign joinf_0n[13] = ifint_0n[13];
  assign joinf_0n[14] = ifint_0n[14];
  assign joinf_0n[15] = ifint_0n[15];
  assign joinf_0n[16] = ifint_0n[16];
  assign joinf_0n[17] = ifint_0n[17];
  assign joinf_0n[18] = ifint_0n[18];
  assign joinf_0n[19] = ifint_0n[19];
  assign joinf_0n[20] = ifint_0n[20];
  assign joinf_0n[21] = ifint_0n[21];
  assign joinf_0n[22] = ifint_0n[22];
  assign joinf_0n[23] = ifint_0n[23];
  assign joinf_0n[24] = ifint_0n[24];
  assign joinf_0n[25] = ifint_0n[25];
  assign joinf_0n[26] = ifint_0n[26];
  assign joinf_0n[27] = ifint_0n[27];
  assign joinf_0n[28] = ifint_0n[28];
  assign joinf_0n[29] = ifint_0n[29];
  assign joinf_0n[30] = ifint_0n[30];
  assign joinf_0n[31] = ifint_0n[31];
  assign joinf_0n[32] = ifint_0n[32];
endmodule

module BrzJ_l12__2833_201_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [32:0] i_0r0d;
  input [32:0] i_0r1d;
  output i_0a;
  input i_1r0d;
  input i_1r1d;
  output i_1a;
  output [33:0] o_0r0d;
  output [33:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [34:0] internal_0n;
  wire [33:0] ofint_0n;
  wire [33:0] otint_0n;
  wire oaint_0n;
  wire [32:0] ifint_0n;
  wire ifint_1n;
  wire [32:0] itint_0n;
  wire itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire complete615_0n;
  wire gate614_0n;
  wire [32:0] complete611_0n;
  wire gate610_0n;
  wire [33:0] complete607_0n;
  wire gate606_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign i_1a = complete615_0n;
  OR2 I3 (complete615_0n, ifint_1n, itint_1n);
  INV I4 (gate614_0n, iaint_1n);
  C2RI I5 (itint_1n, i_1r1d, gate614_0n, initialise);
  C2RI I6 (ifint_1n, i_1r0d, gate614_0n, initialise);
  C3 I7 (internal_0n[0], complete611_0n[0], complete611_0n[1], complete611_0n[2]);
  C3 I8 (internal_0n[1], complete611_0n[3], complete611_0n[4], complete611_0n[5]);
  C3 I9 (internal_0n[2], complete611_0n[6], complete611_0n[7], complete611_0n[8]);
  C3 I10 (internal_0n[3], complete611_0n[9], complete611_0n[10], complete611_0n[11]);
  C3 I11 (internal_0n[4], complete611_0n[12], complete611_0n[13], complete611_0n[14]);
  C3 I12 (internal_0n[5], complete611_0n[15], complete611_0n[16], complete611_0n[17]);
  C3 I13 (internal_0n[6], complete611_0n[18], complete611_0n[19], complete611_0n[20]);
  C3 I14 (internal_0n[7], complete611_0n[21], complete611_0n[22], complete611_0n[23]);
  C3 I15 (internal_0n[8], complete611_0n[24], complete611_0n[25], complete611_0n[26]);
  C3 I16 (internal_0n[9], complete611_0n[27], complete611_0n[28], complete611_0n[29]);
  C3 I17 (internal_0n[10], complete611_0n[30], complete611_0n[31], complete611_0n[32]);
  C3 I18 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I19 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I20 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I21 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I22 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I23 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I24 (i_0a, internal_0n[15], internal_0n[16]);
  OR2 I25 (complete611_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I26 (complete611_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I27 (complete611_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I28 (complete611_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I29 (complete611_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I30 (complete611_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I31 (complete611_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I32 (complete611_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I33 (complete611_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I34 (complete611_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I35 (complete611_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I36 (complete611_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I37 (complete611_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I38 (complete611_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I39 (complete611_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I40 (complete611_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I41 (complete611_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I42 (complete611_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I43 (complete611_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I44 (complete611_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I45 (complete611_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I46 (complete611_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I47 (complete611_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I48 (complete611_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I49 (complete611_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I50 (complete611_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I51 (complete611_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I52 (complete611_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I53 (complete611_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I54 (complete611_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I55 (complete611_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I56 (complete611_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I57 (complete611_0n[32], ifint_0n[32], itint_0n[32]);
  INV I58 (gate610_0n, iaint_0n);
  C2RI I59 (itint_0n[0], i_0r1d[0], gate610_0n, initialise);
  C2RI I60 (itint_0n[1], i_0r1d[1], gate610_0n, initialise);
  C2RI I61 (itint_0n[2], i_0r1d[2], gate610_0n, initialise);
  C2RI I62 (itint_0n[3], i_0r1d[3], gate610_0n, initialise);
  C2RI I63 (itint_0n[4], i_0r1d[4], gate610_0n, initialise);
  C2RI I64 (itint_0n[5], i_0r1d[5], gate610_0n, initialise);
  C2RI I65 (itint_0n[6], i_0r1d[6], gate610_0n, initialise);
  C2RI I66 (itint_0n[7], i_0r1d[7], gate610_0n, initialise);
  C2RI I67 (itint_0n[8], i_0r1d[8], gate610_0n, initialise);
  C2RI I68 (itint_0n[9], i_0r1d[9], gate610_0n, initialise);
  C2RI I69 (itint_0n[10], i_0r1d[10], gate610_0n, initialise);
  C2RI I70 (itint_0n[11], i_0r1d[11], gate610_0n, initialise);
  C2RI I71 (itint_0n[12], i_0r1d[12], gate610_0n, initialise);
  C2RI I72 (itint_0n[13], i_0r1d[13], gate610_0n, initialise);
  C2RI I73 (itint_0n[14], i_0r1d[14], gate610_0n, initialise);
  C2RI I74 (itint_0n[15], i_0r1d[15], gate610_0n, initialise);
  C2RI I75 (itint_0n[16], i_0r1d[16], gate610_0n, initialise);
  C2RI I76 (itint_0n[17], i_0r1d[17], gate610_0n, initialise);
  C2RI I77 (itint_0n[18], i_0r1d[18], gate610_0n, initialise);
  C2RI I78 (itint_0n[19], i_0r1d[19], gate610_0n, initialise);
  C2RI I79 (itint_0n[20], i_0r1d[20], gate610_0n, initialise);
  C2RI I80 (itint_0n[21], i_0r1d[21], gate610_0n, initialise);
  C2RI I81 (itint_0n[22], i_0r1d[22], gate610_0n, initialise);
  C2RI I82 (itint_0n[23], i_0r1d[23], gate610_0n, initialise);
  C2RI I83 (itint_0n[24], i_0r1d[24], gate610_0n, initialise);
  C2RI I84 (itint_0n[25], i_0r1d[25], gate610_0n, initialise);
  C2RI I85 (itint_0n[26], i_0r1d[26], gate610_0n, initialise);
  C2RI I86 (itint_0n[27], i_0r1d[27], gate610_0n, initialise);
  C2RI I87 (itint_0n[28], i_0r1d[28], gate610_0n, initialise);
  C2RI I88 (itint_0n[29], i_0r1d[29], gate610_0n, initialise);
  C2RI I89 (itint_0n[30], i_0r1d[30], gate610_0n, initialise);
  C2RI I90 (itint_0n[31], i_0r1d[31], gate610_0n, initialise);
  C2RI I91 (itint_0n[32], i_0r1d[32], gate610_0n, initialise);
  C2RI I92 (ifint_0n[0], i_0r0d[0], gate610_0n, initialise);
  C2RI I93 (ifint_0n[1], i_0r0d[1], gate610_0n, initialise);
  C2RI I94 (ifint_0n[2], i_0r0d[2], gate610_0n, initialise);
  C2RI I95 (ifint_0n[3], i_0r0d[3], gate610_0n, initialise);
  C2RI I96 (ifint_0n[4], i_0r0d[4], gate610_0n, initialise);
  C2RI I97 (ifint_0n[5], i_0r0d[5], gate610_0n, initialise);
  C2RI I98 (ifint_0n[6], i_0r0d[6], gate610_0n, initialise);
  C2RI I99 (ifint_0n[7], i_0r0d[7], gate610_0n, initialise);
  C2RI I100 (ifint_0n[8], i_0r0d[8], gate610_0n, initialise);
  C2RI I101 (ifint_0n[9], i_0r0d[9], gate610_0n, initialise);
  C2RI I102 (ifint_0n[10], i_0r0d[10], gate610_0n, initialise);
  C2RI I103 (ifint_0n[11], i_0r0d[11], gate610_0n, initialise);
  C2RI I104 (ifint_0n[12], i_0r0d[12], gate610_0n, initialise);
  C2RI I105 (ifint_0n[13], i_0r0d[13], gate610_0n, initialise);
  C2RI I106 (ifint_0n[14], i_0r0d[14], gate610_0n, initialise);
  C2RI I107 (ifint_0n[15], i_0r0d[15], gate610_0n, initialise);
  C2RI I108 (ifint_0n[16], i_0r0d[16], gate610_0n, initialise);
  C2RI I109 (ifint_0n[17], i_0r0d[17], gate610_0n, initialise);
  C2RI I110 (ifint_0n[18], i_0r0d[18], gate610_0n, initialise);
  C2RI I111 (ifint_0n[19], i_0r0d[19], gate610_0n, initialise);
  C2RI I112 (ifint_0n[20], i_0r0d[20], gate610_0n, initialise);
  C2RI I113 (ifint_0n[21], i_0r0d[21], gate610_0n, initialise);
  C2RI I114 (ifint_0n[22], i_0r0d[22], gate610_0n, initialise);
  C2RI I115 (ifint_0n[23], i_0r0d[23], gate610_0n, initialise);
  C2RI I116 (ifint_0n[24], i_0r0d[24], gate610_0n, initialise);
  C2RI I117 (ifint_0n[25], i_0r0d[25], gate610_0n, initialise);
  C2RI I118 (ifint_0n[26], i_0r0d[26], gate610_0n, initialise);
  C2RI I119 (ifint_0n[27], i_0r0d[27], gate610_0n, initialise);
  C2RI I120 (ifint_0n[28], i_0r0d[28], gate610_0n, initialise);
  C2RI I121 (ifint_0n[29], i_0r0d[29], gate610_0n, initialise);
  C2RI I122 (ifint_0n[30], i_0r0d[30], gate610_0n, initialise);
  C2RI I123 (ifint_0n[31], i_0r0d[31], gate610_0n, initialise);
  C2RI I124 (ifint_0n[32], i_0r0d[32], gate610_0n, initialise);
  C3 I125 (internal_0n[17], complete607_0n[0], complete607_0n[1], complete607_0n[2]);
  C3 I126 (internal_0n[18], complete607_0n[3], complete607_0n[4], complete607_0n[5]);
  C3 I127 (internal_0n[19], complete607_0n[6], complete607_0n[7], complete607_0n[8]);
  C3 I128 (internal_0n[20], complete607_0n[9], complete607_0n[10], complete607_0n[11]);
  C3 I129 (internal_0n[21], complete607_0n[12], complete607_0n[13], complete607_0n[14]);
  C3 I130 (internal_0n[22], complete607_0n[15], complete607_0n[16], complete607_0n[17]);
  C3 I131 (internal_0n[23], complete607_0n[18], complete607_0n[19], complete607_0n[20]);
  C3 I132 (internal_0n[24], complete607_0n[21], complete607_0n[22], complete607_0n[23]);
  C3 I133 (internal_0n[25], complete607_0n[24], complete607_0n[25], complete607_0n[26]);
  C3 I134 (internal_0n[26], complete607_0n[27], complete607_0n[28], complete607_0n[29]);
  C2 I135 (internal_0n[27], complete607_0n[30], complete607_0n[31]);
  C2 I136 (internal_0n[28], complete607_0n[32], complete607_0n[33]);
  C3 I137 (internal_0n[29], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I138 (internal_0n[30], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I139 (internal_0n[31], internal_0n[23], internal_0n[24], internal_0n[25]);
  C3 I140 (internal_0n[32], internal_0n[26], internal_0n[27], internal_0n[28]);
  C2 I141 (internal_0n[33], internal_0n[29], internal_0n[30]);
  C2 I142 (internal_0n[34], internal_0n[31], internal_0n[32]);
  C2 I143 (oaint_0n, internal_0n[33], internal_0n[34]);
  OR2 I144 (complete607_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I145 (complete607_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I146 (complete607_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I147 (complete607_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I148 (complete607_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I149 (complete607_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I150 (complete607_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I151 (complete607_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I152 (complete607_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I153 (complete607_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I154 (complete607_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I155 (complete607_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I156 (complete607_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I157 (complete607_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I158 (complete607_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I159 (complete607_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I160 (complete607_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I161 (complete607_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I162 (complete607_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I163 (complete607_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I164 (complete607_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I165 (complete607_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I166 (complete607_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I167 (complete607_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I168 (complete607_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I169 (complete607_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I170 (complete607_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I171 (complete607_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I172 (complete607_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I173 (complete607_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I174 (complete607_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I175 (complete607_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I176 (complete607_0n[32], o_0r0d[32], o_0r1d[32]);
  OR2 I177 (complete607_0n[33], o_0r0d[33], o_0r1d[33]);
  INV I178 (gate606_0n, o_0a);
  C2RI I179 (o_0r1d[0], otint_0n[0], gate606_0n, initialise);
  C2RI I180 (o_0r1d[1], otint_0n[1], gate606_0n, initialise);
  C2RI I181 (o_0r1d[2], otint_0n[2], gate606_0n, initialise);
  C2RI I182 (o_0r1d[3], otint_0n[3], gate606_0n, initialise);
  C2RI I183 (o_0r1d[4], otint_0n[4], gate606_0n, initialise);
  C2RI I184 (o_0r1d[5], otint_0n[5], gate606_0n, initialise);
  C2RI I185 (o_0r1d[6], otint_0n[6], gate606_0n, initialise);
  C2RI I186 (o_0r1d[7], otint_0n[7], gate606_0n, initialise);
  C2RI I187 (o_0r1d[8], otint_0n[8], gate606_0n, initialise);
  C2RI I188 (o_0r1d[9], otint_0n[9], gate606_0n, initialise);
  C2RI I189 (o_0r1d[10], otint_0n[10], gate606_0n, initialise);
  C2RI I190 (o_0r1d[11], otint_0n[11], gate606_0n, initialise);
  C2RI I191 (o_0r1d[12], otint_0n[12], gate606_0n, initialise);
  C2RI I192 (o_0r1d[13], otint_0n[13], gate606_0n, initialise);
  C2RI I193 (o_0r1d[14], otint_0n[14], gate606_0n, initialise);
  C2RI I194 (o_0r1d[15], otint_0n[15], gate606_0n, initialise);
  C2RI I195 (o_0r1d[16], otint_0n[16], gate606_0n, initialise);
  C2RI I196 (o_0r1d[17], otint_0n[17], gate606_0n, initialise);
  C2RI I197 (o_0r1d[18], otint_0n[18], gate606_0n, initialise);
  C2RI I198 (o_0r1d[19], otint_0n[19], gate606_0n, initialise);
  C2RI I199 (o_0r1d[20], otint_0n[20], gate606_0n, initialise);
  C2RI I200 (o_0r1d[21], otint_0n[21], gate606_0n, initialise);
  C2RI I201 (o_0r1d[22], otint_0n[22], gate606_0n, initialise);
  C2RI I202 (o_0r1d[23], otint_0n[23], gate606_0n, initialise);
  C2RI I203 (o_0r1d[24], otint_0n[24], gate606_0n, initialise);
  C2RI I204 (o_0r1d[25], otint_0n[25], gate606_0n, initialise);
  C2RI I205 (o_0r1d[26], otint_0n[26], gate606_0n, initialise);
  C2RI I206 (o_0r1d[27], otint_0n[27], gate606_0n, initialise);
  C2RI I207 (o_0r1d[28], otint_0n[28], gate606_0n, initialise);
  C2RI I208 (o_0r1d[29], otint_0n[29], gate606_0n, initialise);
  C2RI I209 (o_0r1d[30], otint_0n[30], gate606_0n, initialise);
  C2RI I210 (o_0r1d[31], otint_0n[31], gate606_0n, initialise);
  C2RI I211 (o_0r1d[32], otint_0n[32], gate606_0n, initialise);
  C2RI I212 (o_0r1d[33], otint_0n[33], gate606_0n, initialise);
  C2RI I213 (o_0r0d[0], ofint_0n[0], gate606_0n, initialise);
  C2RI I214 (o_0r0d[1], ofint_0n[1], gate606_0n, initialise);
  C2RI I215 (o_0r0d[2], ofint_0n[2], gate606_0n, initialise);
  C2RI I216 (o_0r0d[3], ofint_0n[3], gate606_0n, initialise);
  C2RI I217 (o_0r0d[4], ofint_0n[4], gate606_0n, initialise);
  C2RI I218 (o_0r0d[5], ofint_0n[5], gate606_0n, initialise);
  C2RI I219 (o_0r0d[6], ofint_0n[6], gate606_0n, initialise);
  C2RI I220 (o_0r0d[7], ofint_0n[7], gate606_0n, initialise);
  C2RI I221 (o_0r0d[8], ofint_0n[8], gate606_0n, initialise);
  C2RI I222 (o_0r0d[9], ofint_0n[9], gate606_0n, initialise);
  C2RI I223 (o_0r0d[10], ofint_0n[10], gate606_0n, initialise);
  C2RI I224 (o_0r0d[11], ofint_0n[11], gate606_0n, initialise);
  C2RI I225 (o_0r0d[12], ofint_0n[12], gate606_0n, initialise);
  C2RI I226 (o_0r0d[13], ofint_0n[13], gate606_0n, initialise);
  C2RI I227 (o_0r0d[14], ofint_0n[14], gate606_0n, initialise);
  C2RI I228 (o_0r0d[15], ofint_0n[15], gate606_0n, initialise);
  C2RI I229 (o_0r0d[16], ofint_0n[16], gate606_0n, initialise);
  C2RI I230 (o_0r0d[17], ofint_0n[17], gate606_0n, initialise);
  C2RI I231 (o_0r0d[18], ofint_0n[18], gate606_0n, initialise);
  C2RI I232 (o_0r0d[19], ofint_0n[19], gate606_0n, initialise);
  C2RI I233 (o_0r0d[20], ofint_0n[20], gate606_0n, initialise);
  C2RI I234 (o_0r0d[21], ofint_0n[21], gate606_0n, initialise);
  C2RI I235 (o_0r0d[22], ofint_0n[22], gate606_0n, initialise);
  C2RI I236 (o_0r0d[23], ofint_0n[23], gate606_0n, initialise);
  C2RI I237 (o_0r0d[24], ofint_0n[24], gate606_0n, initialise);
  C2RI I238 (o_0r0d[25], ofint_0n[25], gate606_0n, initialise);
  C2RI I239 (o_0r0d[26], ofint_0n[26], gate606_0n, initialise);
  C2RI I240 (o_0r0d[27], ofint_0n[27], gate606_0n, initialise);
  C2RI I241 (o_0r0d[28], ofint_0n[28], gate606_0n, initialise);
  C2RI I242 (o_0r0d[29], ofint_0n[29], gate606_0n, initialise);
  C2RI I243 (o_0r0d[30], ofint_0n[30], gate606_0n, initialise);
  C2RI I244 (o_0r0d[31], ofint_0n[31], gate606_0n, initialise);
  C2RI I245 (o_0r0d[32], ofint_0n[32], gate606_0n, initialise);
  C2RI I246 (o_0r0d[33], ofint_0n[33], gate606_0n, initialise);
  assign otint_0n[0] = itint_0n[0];
  assign otint_0n[1] = itint_0n[1];
  assign otint_0n[2] = itint_0n[2];
  assign otint_0n[3] = itint_0n[3];
  assign otint_0n[4] = itint_0n[4];
  assign otint_0n[5] = itint_0n[5];
  assign otint_0n[6] = itint_0n[6];
  assign otint_0n[7] = itint_0n[7];
  assign otint_0n[8] = itint_0n[8];
  assign otint_0n[9] = itint_0n[9];
  assign otint_0n[10] = itint_0n[10];
  assign otint_0n[11] = itint_0n[11];
  assign otint_0n[12] = itint_0n[12];
  assign otint_0n[13] = itint_0n[13];
  assign otint_0n[14] = itint_0n[14];
  assign otint_0n[15] = itint_0n[15];
  assign otint_0n[16] = itint_0n[16];
  assign otint_0n[17] = itint_0n[17];
  assign otint_0n[18] = itint_0n[18];
  assign otint_0n[19] = itint_0n[19];
  assign otint_0n[20] = itint_0n[20];
  assign otint_0n[21] = itint_0n[21];
  assign otint_0n[22] = itint_0n[22];
  assign otint_0n[23] = itint_0n[23];
  assign otint_0n[24] = itint_0n[24];
  assign otint_0n[25] = itint_0n[25];
  assign otint_0n[26] = itint_0n[26];
  assign otint_0n[27] = itint_0n[27];
  assign otint_0n[28] = itint_0n[28];
  assign otint_0n[29] = itint_0n[29];
  assign otint_0n[30] = itint_0n[30];
  assign otint_0n[31] = itint_0n[31];
  assign otint_0n[32] = itint_0n[32];
  assign otint_0n[33] = itint_1n;
  assign ofint_0n[0] = ifint_0n[0];
  assign ofint_0n[1] = ifint_0n[1];
  assign ofint_0n[2] = ifint_0n[2];
  assign ofint_0n[3] = ifint_0n[3];
  assign ofint_0n[4] = ifint_0n[4];
  assign ofint_0n[5] = ifint_0n[5];
  assign ofint_0n[6] = ifint_0n[6];
  assign ofint_0n[7] = ifint_0n[7];
  assign ofint_0n[8] = ifint_0n[8];
  assign ofint_0n[9] = ifint_0n[9];
  assign ofint_0n[10] = ifint_0n[10];
  assign ofint_0n[11] = ifint_0n[11];
  assign ofint_0n[12] = ifint_0n[12];
  assign ofint_0n[13] = ifint_0n[13];
  assign ofint_0n[14] = ifint_0n[14];
  assign ofint_0n[15] = ifint_0n[15];
  assign ofint_0n[16] = ifint_0n[16];
  assign ofint_0n[17] = ifint_0n[17];
  assign ofint_0n[18] = ifint_0n[18];
  assign ofint_0n[19] = ifint_0n[19];
  assign ofint_0n[20] = ifint_0n[20];
  assign ofint_0n[21] = ifint_0n[21];
  assign ofint_0n[22] = ifint_0n[22];
  assign ofint_0n[23] = ifint_0n[23];
  assign ofint_0n[24] = ifint_0n[24];
  assign ofint_0n[25] = ifint_0n[25];
  assign ofint_0n[26] = ifint_0n[26];
  assign ofint_0n[27] = ifint_0n[27];
  assign ofint_0n[28] = ifint_0n[28];
  assign ofint_0n[29] = ifint_0n[29];
  assign ofint_0n[30] = ifint_0n[30];
  assign ofint_0n[31] = ifint_0n[31];
  assign ofint_0n[32] = ifint_0n[32];
  assign ofint_0n[33] = ifint_1n;
endmodule

module BrzJ_l12__2833_202_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [32:0] i_0r0d;
  input [32:0] i_0r1d;
  output i_0a;
  input [1:0] i_1r0d;
  input [1:0] i_1r1d;
  output i_1a;
  output [34:0] o_0r0d;
  output [34:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [34:0] internal_0n;
  wire [34:0] ofint_0n;
  wire [34:0] otint_0n;
  wire oaint_0n;
  wire [32:0] ifint_0n;
  wire [1:0] ifint_1n;
  wire [32:0] itint_0n;
  wire [1:0] itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [1:0] complete627_0n;
  wire gate626_0n;
  wire [32:0] complete623_0n;
  wire gate622_0n;
  wire [34:0] complete619_0n;
  wire gate618_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  C2 I2 (i_1a, complete627_0n[0], complete627_0n[1]);
  OR2 I3 (complete627_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I4 (complete627_0n[1], ifint_1n[1], itint_1n[1]);
  INV I5 (gate626_0n, iaint_1n);
  C2RI I6 (itint_1n[0], i_1r1d[0], gate626_0n, initialise);
  C2RI I7 (itint_1n[1], i_1r1d[1], gate626_0n, initialise);
  C2RI I8 (ifint_1n[0], i_1r0d[0], gate626_0n, initialise);
  C2RI I9 (ifint_1n[1], i_1r0d[1], gate626_0n, initialise);
  C3 I10 (internal_0n[0], complete623_0n[0], complete623_0n[1], complete623_0n[2]);
  C3 I11 (internal_0n[1], complete623_0n[3], complete623_0n[4], complete623_0n[5]);
  C3 I12 (internal_0n[2], complete623_0n[6], complete623_0n[7], complete623_0n[8]);
  C3 I13 (internal_0n[3], complete623_0n[9], complete623_0n[10], complete623_0n[11]);
  C3 I14 (internal_0n[4], complete623_0n[12], complete623_0n[13], complete623_0n[14]);
  C3 I15 (internal_0n[5], complete623_0n[15], complete623_0n[16], complete623_0n[17]);
  C3 I16 (internal_0n[6], complete623_0n[18], complete623_0n[19], complete623_0n[20]);
  C3 I17 (internal_0n[7], complete623_0n[21], complete623_0n[22], complete623_0n[23]);
  C3 I18 (internal_0n[8], complete623_0n[24], complete623_0n[25], complete623_0n[26]);
  C3 I19 (internal_0n[9], complete623_0n[27], complete623_0n[28], complete623_0n[29]);
  C3 I20 (internal_0n[10], complete623_0n[30], complete623_0n[31], complete623_0n[32]);
  C3 I21 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I22 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I23 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I24 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I25 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I26 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I27 (i_0a, internal_0n[15], internal_0n[16]);
  OR2 I28 (complete623_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I29 (complete623_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I30 (complete623_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I31 (complete623_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I32 (complete623_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I33 (complete623_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I34 (complete623_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I35 (complete623_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I36 (complete623_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I37 (complete623_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I38 (complete623_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I39 (complete623_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I40 (complete623_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I41 (complete623_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I42 (complete623_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I43 (complete623_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I44 (complete623_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I45 (complete623_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I46 (complete623_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I47 (complete623_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I48 (complete623_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I49 (complete623_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I50 (complete623_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I51 (complete623_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I52 (complete623_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I53 (complete623_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I54 (complete623_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I55 (complete623_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I56 (complete623_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I57 (complete623_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I58 (complete623_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I59 (complete623_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I60 (complete623_0n[32], ifint_0n[32], itint_0n[32]);
  INV I61 (gate622_0n, iaint_0n);
  C2RI I62 (itint_0n[0], i_0r1d[0], gate622_0n, initialise);
  C2RI I63 (itint_0n[1], i_0r1d[1], gate622_0n, initialise);
  C2RI I64 (itint_0n[2], i_0r1d[2], gate622_0n, initialise);
  C2RI I65 (itint_0n[3], i_0r1d[3], gate622_0n, initialise);
  C2RI I66 (itint_0n[4], i_0r1d[4], gate622_0n, initialise);
  C2RI I67 (itint_0n[5], i_0r1d[5], gate622_0n, initialise);
  C2RI I68 (itint_0n[6], i_0r1d[6], gate622_0n, initialise);
  C2RI I69 (itint_0n[7], i_0r1d[7], gate622_0n, initialise);
  C2RI I70 (itint_0n[8], i_0r1d[8], gate622_0n, initialise);
  C2RI I71 (itint_0n[9], i_0r1d[9], gate622_0n, initialise);
  C2RI I72 (itint_0n[10], i_0r1d[10], gate622_0n, initialise);
  C2RI I73 (itint_0n[11], i_0r1d[11], gate622_0n, initialise);
  C2RI I74 (itint_0n[12], i_0r1d[12], gate622_0n, initialise);
  C2RI I75 (itint_0n[13], i_0r1d[13], gate622_0n, initialise);
  C2RI I76 (itint_0n[14], i_0r1d[14], gate622_0n, initialise);
  C2RI I77 (itint_0n[15], i_0r1d[15], gate622_0n, initialise);
  C2RI I78 (itint_0n[16], i_0r1d[16], gate622_0n, initialise);
  C2RI I79 (itint_0n[17], i_0r1d[17], gate622_0n, initialise);
  C2RI I80 (itint_0n[18], i_0r1d[18], gate622_0n, initialise);
  C2RI I81 (itint_0n[19], i_0r1d[19], gate622_0n, initialise);
  C2RI I82 (itint_0n[20], i_0r1d[20], gate622_0n, initialise);
  C2RI I83 (itint_0n[21], i_0r1d[21], gate622_0n, initialise);
  C2RI I84 (itint_0n[22], i_0r1d[22], gate622_0n, initialise);
  C2RI I85 (itint_0n[23], i_0r1d[23], gate622_0n, initialise);
  C2RI I86 (itint_0n[24], i_0r1d[24], gate622_0n, initialise);
  C2RI I87 (itint_0n[25], i_0r1d[25], gate622_0n, initialise);
  C2RI I88 (itint_0n[26], i_0r1d[26], gate622_0n, initialise);
  C2RI I89 (itint_0n[27], i_0r1d[27], gate622_0n, initialise);
  C2RI I90 (itint_0n[28], i_0r1d[28], gate622_0n, initialise);
  C2RI I91 (itint_0n[29], i_0r1d[29], gate622_0n, initialise);
  C2RI I92 (itint_0n[30], i_0r1d[30], gate622_0n, initialise);
  C2RI I93 (itint_0n[31], i_0r1d[31], gate622_0n, initialise);
  C2RI I94 (itint_0n[32], i_0r1d[32], gate622_0n, initialise);
  C2RI I95 (ifint_0n[0], i_0r0d[0], gate622_0n, initialise);
  C2RI I96 (ifint_0n[1], i_0r0d[1], gate622_0n, initialise);
  C2RI I97 (ifint_0n[2], i_0r0d[2], gate622_0n, initialise);
  C2RI I98 (ifint_0n[3], i_0r0d[3], gate622_0n, initialise);
  C2RI I99 (ifint_0n[4], i_0r0d[4], gate622_0n, initialise);
  C2RI I100 (ifint_0n[5], i_0r0d[5], gate622_0n, initialise);
  C2RI I101 (ifint_0n[6], i_0r0d[6], gate622_0n, initialise);
  C2RI I102 (ifint_0n[7], i_0r0d[7], gate622_0n, initialise);
  C2RI I103 (ifint_0n[8], i_0r0d[8], gate622_0n, initialise);
  C2RI I104 (ifint_0n[9], i_0r0d[9], gate622_0n, initialise);
  C2RI I105 (ifint_0n[10], i_0r0d[10], gate622_0n, initialise);
  C2RI I106 (ifint_0n[11], i_0r0d[11], gate622_0n, initialise);
  C2RI I107 (ifint_0n[12], i_0r0d[12], gate622_0n, initialise);
  C2RI I108 (ifint_0n[13], i_0r0d[13], gate622_0n, initialise);
  C2RI I109 (ifint_0n[14], i_0r0d[14], gate622_0n, initialise);
  C2RI I110 (ifint_0n[15], i_0r0d[15], gate622_0n, initialise);
  C2RI I111 (ifint_0n[16], i_0r0d[16], gate622_0n, initialise);
  C2RI I112 (ifint_0n[17], i_0r0d[17], gate622_0n, initialise);
  C2RI I113 (ifint_0n[18], i_0r0d[18], gate622_0n, initialise);
  C2RI I114 (ifint_0n[19], i_0r0d[19], gate622_0n, initialise);
  C2RI I115 (ifint_0n[20], i_0r0d[20], gate622_0n, initialise);
  C2RI I116 (ifint_0n[21], i_0r0d[21], gate622_0n, initialise);
  C2RI I117 (ifint_0n[22], i_0r0d[22], gate622_0n, initialise);
  C2RI I118 (ifint_0n[23], i_0r0d[23], gate622_0n, initialise);
  C2RI I119 (ifint_0n[24], i_0r0d[24], gate622_0n, initialise);
  C2RI I120 (ifint_0n[25], i_0r0d[25], gate622_0n, initialise);
  C2RI I121 (ifint_0n[26], i_0r0d[26], gate622_0n, initialise);
  C2RI I122 (ifint_0n[27], i_0r0d[27], gate622_0n, initialise);
  C2RI I123 (ifint_0n[28], i_0r0d[28], gate622_0n, initialise);
  C2RI I124 (ifint_0n[29], i_0r0d[29], gate622_0n, initialise);
  C2RI I125 (ifint_0n[30], i_0r0d[30], gate622_0n, initialise);
  C2RI I126 (ifint_0n[31], i_0r0d[31], gate622_0n, initialise);
  C2RI I127 (ifint_0n[32], i_0r0d[32], gate622_0n, initialise);
  C3 I128 (internal_0n[17], complete619_0n[0], complete619_0n[1], complete619_0n[2]);
  C3 I129 (internal_0n[18], complete619_0n[3], complete619_0n[4], complete619_0n[5]);
  C3 I130 (internal_0n[19], complete619_0n[6], complete619_0n[7], complete619_0n[8]);
  C3 I131 (internal_0n[20], complete619_0n[9], complete619_0n[10], complete619_0n[11]);
  C3 I132 (internal_0n[21], complete619_0n[12], complete619_0n[13], complete619_0n[14]);
  C3 I133 (internal_0n[22], complete619_0n[15], complete619_0n[16], complete619_0n[17]);
  C3 I134 (internal_0n[23], complete619_0n[18], complete619_0n[19], complete619_0n[20]);
  C3 I135 (internal_0n[24], complete619_0n[21], complete619_0n[22], complete619_0n[23]);
  C3 I136 (internal_0n[25], complete619_0n[24], complete619_0n[25], complete619_0n[26]);
  C3 I137 (internal_0n[26], complete619_0n[27], complete619_0n[28], complete619_0n[29]);
  C3 I138 (internal_0n[27], complete619_0n[30], complete619_0n[31], complete619_0n[32]);
  C2 I139 (internal_0n[28], complete619_0n[33], complete619_0n[34]);
  C3 I140 (internal_0n[29], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I141 (internal_0n[30], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I142 (internal_0n[31], internal_0n[23], internal_0n[24], internal_0n[25]);
  C3 I143 (internal_0n[32], internal_0n[26], internal_0n[27], internal_0n[28]);
  C2 I144 (internal_0n[33], internal_0n[29], internal_0n[30]);
  C2 I145 (internal_0n[34], internal_0n[31], internal_0n[32]);
  C2 I146 (oaint_0n, internal_0n[33], internal_0n[34]);
  OR2 I147 (complete619_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I148 (complete619_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I149 (complete619_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I150 (complete619_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I151 (complete619_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I152 (complete619_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I153 (complete619_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I154 (complete619_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I155 (complete619_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I156 (complete619_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I157 (complete619_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I158 (complete619_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I159 (complete619_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I160 (complete619_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I161 (complete619_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I162 (complete619_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I163 (complete619_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I164 (complete619_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I165 (complete619_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I166 (complete619_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I167 (complete619_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I168 (complete619_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I169 (complete619_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I170 (complete619_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I171 (complete619_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I172 (complete619_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I173 (complete619_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I174 (complete619_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I175 (complete619_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I176 (complete619_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I177 (complete619_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I178 (complete619_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I179 (complete619_0n[32], o_0r0d[32], o_0r1d[32]);
  OR2 I180 (complete619_0n[33], o_0r0d[33], o_0r1d[33]);
  OR2 I181 (complete619_0n[34], o_0r0d[34], o_0r1d[34]);
  INV I182 (gate618_0n, o_0a);
  C2RI I183 (o_0r1d[0], otint_0n[0], gate618_0n, initialise);
  C2RI I184 (o_0r1d[1], otint_0n[1], gate618_0n, initialise);
  C2RI I185 (o_0r1d[2], otint_0n[2], gate618_0n, initialise);
  C2RI I186 (o_0r1d[3], otint_0n[3], gate618_0n, initialise);
  C2RI I187 (o_0r1d[4], otint_0n[4], gate618_0n, initialise);
  C2RI I188 (o_0r1d[5], otint_0n[5], gate618_0n, initialise);
  C2RI I189 (o_0r1d[6], otint_0n[6], gate618_0n, initialise);
  C2RI I190 (o_0r1d[7], otint_0n[7], gate618_0n, initialise);
  C2RI I191 (o_0r1d[8], otint_0n[8], gate618_0n, initialise);
  C2RI I192 (o_0r1d[9], otint_0n[9], gate618_0n, initialise);
  C2RI I193 (o_0r1d[10], otint_0n[10], gate618_0n, initialise);
  C2RI I194 (o_0r1d[11], otint_0n[11], gate618_0n, initialise);
  C2RI I195 (o_0r1d[12], otint_0n[12], gate618_0n, initialise);
  C2RI I196 (o_0r1d[13], otint_0n[13], gate618_0n, initialise);
  C2RI I197 (o_0r1d[14], otint_0n[14], gate618_0n, initialise);
  C2RI I198 (o_0r1d[15], otint_0n[15], gate618_0n, initialise);
  C2RI I199 (o_0r1d[16], otint_0n[16], gate618_0n, initialise);
  C2RI I200 (o_0r1d[17], otint_0n[17], gate618_0n, initialise);
  C2RI I201 (o_0r1d[18], otint_0n[18], gate618_0n, initialise);
  C2RI I202 (o_0r1d[19], otint_0n[19], gate618_0n, initialise);
  C2RI I203 (o_0r1d[20], otint_0n[20], gate618_0n, initialise);
  C2RI I204 (o_0r1d[21], otint_0n[21], gate618_0n, initialise);
  C2RI I205 (o_0r1d[22], otint_0n[22], gate618_0n, initialise);
  C2RI I206 (o_0r1d[23], otint_0n[23], gate618_0n, initialise);
  C2RI I207 (o_0r1d[24], otint_0n[24], gate618_0n, initialise);
  C2RI I208 (o_0r1d[25], otint_0n[25], gate618_0n, initialise);
  C2RI I209 (o_0r1d[26], otint_0n[26], gate618_0n, initialise);
  C2RI I210 (o_0r1d[27], otint_0n[27], gate618_0n, initialise);
  C2RI I211 (o_0r1d[28], otint_0n[28], gate618_0n, initialise);
  C2RI I212 (o_0r1d[29], otint_0n[29], gate618_0n, initialise);
  C2RI I213 (o_0r1d[30], otint_0n[30], gate618_0n, initialise);
  C2RI I214 (o_0r1d[31], otint_0n[31], gate618_0n, initialise);
  C2RI I215 (o_0r1d[32], otint_0n[32], gate618_0n, initialise);
  C2RI I216 (o_0r1d[33], otint_0n[33], gate618_0n, initialise);
  C2RI I217 (o_0r1d[34], otint_0n[34], gate618_0n, initialise);
  C2RI I218 (o_0r0d[0], ofint_0n[0], gate618_0n, initialise);
  C2RI I219 (o_0r0d[1], ofint_0n[1], gate618_0n, initialise);
  C2RI I220 (o_0r0d[2], ofint_0n[2], gate618_0n, initialise);
  C2RI I221 (o_0r0d[3], ofint_0n[3], gate618_0n, initialise);
  C2RI I222 (o_0r0d[4], ofint_0n[4], gate618_0n, initialise);
  C2RI I223 (o_0r0d[5], ofint_0n[5], gate618_0n, initialise);
  C2RI I224 (o_0r0d[6], ofint_0n[6], gate618_0n, initialise);
  C2RI I225 (o_0r0d[7], ofint_0n[7], gate618_0n, initialise);
  C2RI I226 (o_0r0d[8], ofint_0n[8], gate618_0n, initialise);
  C2RI I227 (o_0r0d[9], ofint_0n[9], gate618_0n, initialise);
  C2RI I228 (o_0r0d[10], ofint_0n[10], gate618_0n, initialise);
  C2RI I229 (o_0r0d[11], ofint_0n[11], gate618_0n, initialise);
  C2RI I230 (o_0r0d[12], ofint_0n[12], gate618_0n, initialise);
  C2RI I231 (o_0r0d[13], ofint_0n[13], gate618_0n, initialise);
  C2RI I232 (o_0r0d[14], ofint_0n[14], gate618_0n, initialise);
  C2RI I233 (o_0r0d[15], ofint_0n[15], gate618_0n, initialise);
  C2RI I234 (o_0r0d[16], ofint_0n[16], gate618_0n, initialise);
  C2RI I235 (o_0r0d[17], ofint_0n[17], gate618_0n, initialise);
  C2RI I236 (o_0r0d[18], ofint_0n[18], gate618_0n, initialise);
  C2RI I237 (o_0r0d[19], ofint_0n[19], gate618_0n, initialise);
  C2RI I238 (o_0r0d[20], ofint_0n[20], gate618_0n, initialise);
  C2RI I239 (o_0r0d[21], ofint_0n[21], gate618_0n, initialise);
  C2RI I240 (o_0r0d[22], ofint_0n[22], gate618_0n, initialise);
  C2RI I241 (o_0r0d[23], ofint_0n[23], gate618_0n, initialise);
  C2RI I242 (o_0r0d[24], ofint_0n[24], gate618_0n, initialise);
  C2RI I243 (o_0r0d[25], ofint_0n[25], gate618_0n, initialise);
  C2RI I244 (o_0r0d[26], ofint_0n[26], gate618_0n, initialise);
  C2RI I245 (o_0r0d[27], ofint_0n[27], gate618_0n, initialise);
  C2RI I246 (o_0r0d[28], ofint_0n[28], gate618_0n, initialise);
  C2RI I247 (o_0r0d[29], ofint_0n[29], gate618_0n, initialise);
  C2RI I248 (o_0r0d[30], ofint_0n[30], gate618_0n, initialise);
  C2RI I249 (o_0r0d[31], ofint_0n[31], gate618_0n, initialise);
  C2RI I250 (o_0r0d[32], ofint_0n[32], gate618_0n, initialise);
  C2RI I251 (o_0r0d[33], ofint_0n[33], gate618_0n, initialise);
  C2RI I252 (o_0r0d[34], ofint_0n[34], gate618_0n, initialise);
  assign otint_0n[0] = itint_0n[0];
  assign otint_0n[1] = itint_0n[1];
  assign otint_0n[2] = itint_0n[2];
  assign otint_0n[3] = itint_0n[3];
  assign otint_0n[4] = itint_0n[4];
  assign otint_0n[5] = itint_0n[5];
  assign otint_0n[6] = itint_0n[6];
  assign otint_0n[7] = itint_0n[7];
  assign otint_0n[8] = itint_0n[8];
  assign otint_0n[9] = itint_0n[9];
  assign otint_0n[10] = itint_0n[10];
  assign otint_0n[11] = itint_0n[11];
  assign otint_0n[12] = itint_0n[12];
  assign otint_0n[13] = itint_0n[13];
  assign otint_0n[14] = itint_0n[14];
  assign otint_0n[15] = itint_0n[15];
  assign otint_0n[16] = itint_0n[16];
  assign otint_0n[17] = itint_0n[17];
  assign otint_0n[18] = itint_0n[18];
  assign otint_0n[19] = itint_0n[19];
  assign otint_0n[20] = itint_0n[20];
  assign otint_0n[21] = itint_0n[21];
  assign otint_0n[22] = itint_0n[22];
  assign otint_0n[23] = itint_0n[23];
  assign otint_0n[24] = itint_0n[24];
  assign otint_0n[25] = itint_0n[25];
  assign otint_0n[26] = itint_0n[26];
  assign otint_0n[27] = itint_0n[27];
  assign otint_0n[28] = itint_0n[28];
  assign otint_0n[29] = itint_0n[29];
  assign otint_0n[30] = itint_0n[30];
  assign otint_0n[31] = itint_0n[31];
  assign otint_0n[32] = itint_0n[32];
  assign otint_0n[33] = itint_1n[0];
  assign otint_0n[34] = itint_1n[1];
  assign ofint_0n[0] = ifint_0n[0];
  assign ofint_0n[1] = ifint_0n[1];
  assign ofint_0n[2] = ifint_0n[2];
  assign ofint_0n[3] = ifint_0n[3];
  assign ofint_0n[4] = ifint_0n[4];
  assign ofint_0n[5] = ifint_0n[5];
  assign ofint_0n[6] = ifint_0n[6];
  assign ofint_0n[7] = ifint_0n[7];
  assign ofint_0n[8] = ifint_0n[8];
  assign ofint_0n[9] = ifint_0n[9];
  assign ofint_0n[10] = ifint_0n[10];
  assign ofint_0n[11] = ifint_0n[11];
  assign ofint_0n[12] = ifint_0n[12];
  assign ofint_0n[13] = ifint_0n[13];
  assign ofint_0n[14] = ifint_0n[14];
  assign ofint_0n[15] = ifint_0n[15];
  assign ofint_0n[16] = ifint_0n[16];
  assign ofint_0n[17] = ifint_0n[17];
  assign ofint_0n[18] = ifint_0n[18];
  assign ofint_0n[19] = ifint_0n[19];
  assign ofint_0n[20] = ifint_0n[20];
  assign ofint_0n[21] = ifint_0n[21];
  assign ofint_0n[22] = ifint_0n[22];
  assign ofint_0n[23] = ifint_0n[23];
  assign ofint_0n[24] = ifint_0n[24];
  assign ofint_0n[25] = ifint_0n[25];
  assign ofint_0n[26] = ifint_0n[26];
  assign ofint_0n[27] = ifint_0n[27];
  assign ofint_0n[28] = ifint_0n[28];
  assign ofint_0n[29] = ifint_0n[29];
  assign ofint_0n[30] = ifint_0n[30];
  assign ofint_0n[31] = ifint_0n[31];
  assign ofint_0n[32] = ifint_0n[32];
  assign ofint_0n[33] = ifint_1n[0];
  assign ofint_0n[34] = ifint_1n[1];
endmodule

module BrzJ_l13__2833_2033_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [32:0] i_0r0d;
  input [32:0] i_0r1d;
  output i_0a;
  input [32:0] i_1r0d;
  input [32:0] i_1r1d;
  output i_1a;
  output [65:0] o_0r0d;
  output [65:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [66:0] internal_0n;
  wire [65:0] ofint_0n;
  wire [65:0] otint_0n;
  wire oaint_0n;
  wire [32:0] ifint_0n;
  wire [32:0] ifint_1n;
  wire [32:0] itint_0n;
  wire [32:0] itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [32:0] complete639_0n;
  wire gate638_0n;
  wire [32:0] complete635_0n;
  wire gate634_0n;
  wire [65:0] complete631_0n;
  wire gate630_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  C3 I2 (internal_0n[0], complete639_0n[0], complete639_0n[1], complete639_0n[2]);
  C3 I3 (internal_0n[1], complete639_0n[3], complete639_0n[4], complete639_0n[5]);
  C3 I4 (internal_0n[2], complete639_0n[6], complete639_0n[7], complete639_0n[8]);
  C3 I5 (internal_0n[3], complete639_0n[9], complete639_0n[10], complete639_0n[11]);
  C3 I6 (internal_0n[4], complete639_0n[12], complete639_0n[13], complete639_0n[14]);
  C3 I7 (internal_0n[5], complete639_0n[15], complete639_0n[16], complete639_0n[17]);
  C3 I8 (internal_0n[6], complete639_0n[18], complete639_0n[19], complete639_0n[20]);
  C3 I9 (internal_0n[7], complete639_0n[21], complete639_0n[22], complete639_0n[23]);
  C3 I10 (internal_0n[8], complete639_0n[24], complete639_0n[25], complete639_0n[26]);
  C3 I11 (internal_0n[9], complete639_0n[27], complete639_0n[28], complete639_0n[29]);
  C3 I12 (internal_0n[10], complete639_0n[30], complete639_0n[31], complete639_0n[32]);
  C3 I13 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I14 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I15 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I16 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I17 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I18 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I19 (i_1a, internal_0n[15], internal_0n[16]);
  OR2 I20 (complete639_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I21 (complete639_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I22 (complete639_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I23 (complete639_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I24 (complete639_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I25 (complete639_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I26 (complete639_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I27 (complete639_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I28 (complete639_0n[8], ifint_1n[8], itint_1n[8]);
  OR2 I29 (complete639_0n[9], ifint_1n[9], itint_1n[9]);
  OR2 I30 (complete639_0n[10], ifint_1n[10], itint_1n[10]);
  OR2 I31 (complete639_0n[11], ifint_1n[11], itint_1n[11]);
  OR2 I32 (complete639_0n[12], ifint_1n[12], itint_1n[12]);
  OR2 I33 (complete639_0n[13], ifint_1n[13], itint_1n[13]);
  OR2 I34 (complete639_0n[14], ifint_1n[14], itint_1n[14]);
  OR2 I35 (complete639_0n[15], ifint_1n[15], itint_1n[15]);
  OR2 I36 (complete639_0n[16], ifint_1n[16], itint_1n[16]);
  OR2 I37 (complete639_0n[17], ifint_1n[17], itint_1n[17]);
  OR2 I38 (complete639_0n[18], ifint_1n[18], itint_1n[18]);
  OR2 I39 (complete639_0n[19], ifint_1n[19], itint_1n[19]);
  OR2 I40 (complete639_0n[20], ifint_1n[20], itint_1n[20]);
  OR2 I41 (complete639_0n[21], ifint_1n[21], itint_1n[21]);
  OR2 I42 (complete639_0n[22], ifint_1n[22], itint_1n[22]);
  OR2 I43 (complete639_0n[23], ifint_1n[23], itint_1n[23]);
  OR2 I44 (complete639_0n[24], ifint_1n[24], itint_1n[24]);
  OR2 I45 (complete639_0n[25], ifint_1n[25], itint_1n[25]);
  OR2 I46 (complete639_0n[26], ifint_1n[26], itint_1n[26]);
  OR2 I47 (complete639_0n[27], ifint_1n[27], itint_1n[27]);
  OR2 I48 (complete639_0n[28], ifint_1n[28], itint_1n[28]);
  OR2 I49 (complete639_0n[29], ifint_1n[29], itint_1n[29]);
  OR2 I50 (complete639_0n[30], ifint_1n[30], itint_1n[30]);
  OR2 I51 (complete639_0n[31], ifint_1n[31], itint_1n[31]);
  OR2 I52 (complete639_0n[32], ifint_1n[32], itint_1n[32]);
  INV I53 (gate638_0n, iaint_1n);
  C2RI I54 (itint_1n[0], i_1r1d[0], gate638_0n, initialise);
  C2RI I55 (itint_1n[1], i_1r1d[1], gate638_0n, initialise);
  C2RI I56 (itint_1n[2], i_1r1d[2], gate638_0n, initialise);
  C2RI I57 (itint_1n[3], i_1r1d[3], gate638_0n, initialise);
  C2RI I58 (itint_1n[4], i_1r1d[4], gate638_0n, initialise);
  C2RI I59 (itint_1n[5], i_1r1d[5], gate638_0n, initialise);
  C2RI I60 (itint_1n[6], i_1r1d[6], gate638_0n, initialise);
  C2RI I61 (itint_1n[7], i_1r1d[7], gate638_0n, initialise);
  C2RI I62 (itint_1n[8], i_1r1d[8], gate638_0n, initialise);
  C2RI I63 (itint_1n[9], i_1r1d[9], gate638_0n, initialise);
  C2RI I64 (itint_1n[10], i_1r1d[10], gate638_0n, initialise);
  C2RI I65 (itint_1n[11], i_1r1d[11], gate638_0n, initialise);
  C2RI I66 (itint_1n[12], i_1r1d[12], gate638_0n, initialise);
  C2RI I67 (itint_1n[13], i_1r1d[13], gate638_0n, initialise);
  C2RI I68 (itint_1n[14], i_1r1d[14], gate638_0n, initialise);
  C2RI I69 (itint_1n[15], i_1r1d[15], gate638_0n, initialise);
  C2RI I70 (itint_1n[16], i_1r1d[16], gate638_0n, initialise);
  C2RI I71 (itint_1n[17], i_1r1d[17], gate638_0n, initialise);
  C2RI I72 (itint_1n[18], i_1r1d[18], gate638_0n, initialise);
  C2RI I73 (itint_1n[19], i_1r1d[19], gate638_0n, initialise);
  C2RI I74 (itint_1n[20], i_1r1d[20], gate638_0n, initialise);
  C2RI I75 (itint_1n[21], i_1r1d[21], gate638_0n, initialise);
  C2RI I76 (itint_1n[22], i_1r1d[22], gate638_0n, initialise);
  C2RI I77 (itint_1n[23], i_1r1d[23], gate638_0n, initialise);
  C2RI I78 (itint_1n[24], i_1r1d[24], gate638_0n, initialise);
  C2RI I79 (itint_1n[25], i_1r1d[25], gate638_0n, initialise);
  C2RI I80 (itint_1n[26], i_1r1d[26], gate638_0n, initialise);
  C2RI I81 (itint_1n[27], i_1r1d[27], gate638_0n, initialise);
  C2RI I82 (itint_1n[28], i_1r1d[28], gate638_0n, initialise);
  C2RI I83 (itint_1n[29], i_1r1d[29], gate638_0n, initialise);
  C2RI I84 (itint_1n[30], i_1r1d[30], gate638_0n, initialise);
  C2RI I85 (itint_1n[31], i_1r1d[31], gate638_0n, initialise);
  C2RI I86 (itint_1n[32], i_1r1d[32], gate638_0n, initialise);
  C2RI I87 (ifint_1n[0], i_1r0d[0], gate638_0n, initialise);
  C2RI I88 (ifint_1n[1], i_1r0d[1], gate638_0n, initialise);
  C2RI I89 (ifint_1n[2], i_1r0d[2], gate638_0n, initialise);
  C2RI I90 (ifint_1n[3], i_1r0d[3], gate638_0n, initialise);
  C2RI I91 (ifint_1n[4], i_1r0d[4], gate638_0n, initialise);
  C2RI I92 (ifint_1n[5], i_1r0d[5], gate638_0n, initialise);
  C2RI I93 (ifint_1n[6], i_1r0d[6], gate638_0n, initialise);
  C2RI I94 (ifint_1n[7], i_1r0d[7], gate638_0n, initialise);
  C2RI I95 (ifint_1n[8], i_1r0d[8], gate638_0n, initialise);
  C2RI I96 (ifint_1n[9], i_1r0d[9], gate638_0n, initialise);
  C2RI I97 (ifint_1n[10], i_1r0d[10], gate638_0n, initialise);
  C2RI I98 (ifint_1n[11], i_1r0d[11], gate638_0n, initialise);
  C2RI I99 (ifint_1n[12], i_1r0d[12], gate638_0n, initialise);
  C2RI I100 (ifint_1n[13], i_1r0d[13], gate638_0n, initialise);
  C2RI I101 (ifint_1n[14], i_1r0d[14], gate638_0n, initialise);
  C2RI I102 (ifint_1n[15], i_1r0d[15], gate638_0n, initialise);
  C2RI I103 (ifint_1n[16], i_1r0d[16], gate638_0n, initialise);
  C2RI I104 (ifint_1n[17], i_1r0d[17], gate638_0n, initialise);
  C2RI I105 (ifint_1n[18], i_1r0d[18], gate638_0n, initialise);
  C2RI I106 (ifint_1n[19], i_1r0d[19], gate638_0n, initialise);
  C2RI I107 (ifint_1n[20], i_1r0d[20], gate638_0n, initialise);
  C2RI I108 (ifint_1n[21], i_1r0d[21], gate638_0n, initialise);
  C2RI I109 (ifint_1n[22], i_1r0d[22], gate638_0n, initialise);
  C2RI I110 (ifint_1n[23], i_1r0d[23], gate638_0n, initialise);
  C2RI I111 (ifint_1n[24], i_1r0d[24], gate638_0n, initialise);
  C2RI I112 (ifint_1n[25], i_1r0d[25], gate638_0n, initialise);
  C2RI I113 (ifint_1n[26], i_1r0d[26], gate638_0n, initialise);
  C2RI I114 (ifint_1n[27], i_1r0d[27], gate638_0n, initialise);
  C2RI I115 (ifint_1n[28], i_1r0d[28], gate638_0n, initialise);
  C2RI I116 (ifint_1n[29], i_1r0d[29], gate638_0n, initialise);
  C2RI I117 (ifint_1n[30], i_1r0d[30], gate638_0n, initialise);
  C2RI I118 (ifint_1n[31], i_1r0d[31], gate638_0n, initialise);
  C2RI I119 (ifint_1n[32], i_1r0d[32], gate638_0n, initialise);
  C3 I120 (internal_0n[17], complete635_0n[0], complete635_0n[1], complete635_0n[2]);
  C3 I121 (internal_0n[18], complete635_0n[3], complete635_0n[4], complete635_0n[5]);
  C3 I122 (internal_0n[19], complete635_0n[6], complete635_0n[7], complete635_0n[8]);
  C3 I123 (internal_0n[20], complete635_0n[9], complete635_0n[10], complete635_0n[11]);
  C3 I124 (internal_0n[21], complete635_0n[12], complete635_0n[13], complete635_0n[14]);
  C3 I125 (internal_0n[22], complete635_0n[15], complete635_0n[16], complete635_0n[17]);
  C3 I126 (internal_0n[23], complete635_0n[18], complete635_0n[19], complete635_0n[20]);
  C3 I127 (internal_0n[24], complete635_0n[21], complete635_0n[22], complete635_0n[23]);
  C3 I128 (internal_0n[25], complete635_0n[24], complete635_0n[25], complete635_0n[26]);
  C3 I129 (internal_0n[26], complete635_0n[27], complete635_0n[28], complete635_0n[29]);
  C3 I130 (internal_0n[27], complete635_0n[30], complete635_0n[31], complete635_0n[32]);
  C3 I131 (internal_0n[28], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I132 (internal_0n[29], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I133 (internal_0n[30], internal_0n[23], internal_0n[24], internal_0n[25]);
  C2 I134 (internal_0n[31], internal_0n[26], internal_0n[27]);
  C2 I135 (internal_0n[32], internal_0n[28], internal_0n[29]);
  C2 I136 (internal_0n[33], internal_0n[30], internal_0n[31]);
  C2 I137 (i_0a, internal_0n[32], internal_0n[33]);
  OR2 I138 (complete635_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I139 (complete635_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I140 (complete635_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I141 (complete635_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I142 (complete635_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I143 (complete635_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I144 (complete635_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I145 (complete635_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I146 (complete635_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I147 (complete635_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I148 (complete635_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I149 (complete635_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I150 (complete635_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I151 (complete635_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I152 (complete635_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I153 (complete635_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I154 (complete635_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I155 (complete635_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I156 (complete635_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I157 (complete635_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I158 (complete635_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I159 (complete635_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I160 (complete635_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I161 (complete635_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I162 (complete635_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I163 (complete635_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I164 (complete635_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I165 (complete635_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I166 (complete635_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I167 (complete635_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I168 (complete635_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I169 (complete635_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I170 (complete635_0n[32], ifint_0n[32], itint_0n[32]);
  INV I171 (gate634_0n, iaint_0n);
  C2RI I172 (itint_0n[0], i_0r1d[0], gate634_0n, initialise);
  C2RI I173 (itint_0n[1], i_0r1d[1], gate634_0n, initialise);
  C2RI I174 (itint_0n[2], i_0r1d[2], gate634_0n, initialise);
  C2RI I175 (itint_0n[3], i_0r1d[3], gate634_0n, initialise);
  C2RI I176 (itint_0n[4], i_0r1d[4], gate634_0n, initialise);
  C2RI I177 (itint_0n[5], i_0r1d[5], gate634_0n, initialise);
  C2RI I178 (itint_0n[6], i_0r1d[6], gate634_0n, initialise);
  C2RI I179 (itint_0n[7], i_0r1d[7], gate634_0n, initialise);
  C2RI I180 (itint_0n[8], i_0r1d[8], gate634_0n, initialise);
  C2RI I181 (itint_0n[9], i_0r1d[9], gate634_0n, initialise);
  C2RI I182 (itint_0n[10], i_0r1d[10], gate634_0n, initialise);
  C2RI I183 (itint_0n[11], i_0r1d[11], gate634_0n, initialise);
  C2RI I184 (itint_0n[12], i_0r1d[12], gate634_0n, initialise);
  C2RI I185 (itint_0n[13], i_0r1d[13], gate634_0n, initialise);
  C2RI I186 (itint_0n[14], i_0r1d[14], gate634_0n, initialise);
  C2RI I187 (itint_0n[15], i_0r1d[15], gate634_0n, initialise);
  C2RI I188 (itint_0n[16], i_0r1d[16], gate634_0n, initialise);
  C2RI I189 (itint_0n[17], i_0r1d[17], gate634_0n, initialise);
  C2RI I190 (itint_0n[18], i_0r1d[18], gate634_0n, initialise);
  C2RI I191 (itint_0n[19], i_0r1d[19], gate634_0n, initialise);
  C2RI I192 (itint_0n[20], i_0r1d[20], gate634_0n, initialise);
  C2RI I193 (itint_0n[21], i_0r1d[21], gate634_0n, initialise);
  C2RI I194 (itint_0n[22], i_0r1d[22], gate634_0n, initialise);
  C2RI I195 (itint_0n[23], i_0r1d[23], gate634_0n, initialise);
  C2RI I196 (itint_0n[24], i_0r1d[24], gate634_0n, initialise);
  C2RI I197 (itint_0n[25], i_0r1d[25], gate634_0n, initialise);
  C2RI I198 (itint_0n[26], i_0r1d[26], gate634_0n, initialise);
  C2RI I199 (itint_0n[27], i_0r1d[27], gate634_0n, initialise);
  C2RI I200 (itint_0n[28], i_0r1d[28], gate634_0n, initialise);
  C2RI I201 (itint_0n[29], i_0r1d[29], gate634_0n, initialise);
  C2RI I202 (itint_0n[30], i_0r1d[30], gate634_0n, initialise);
  C2RI I203 (itint_0n[31], i_0r1d[31], gate634_0n, initialise);
  C2RI I204 (itint_0n[32], i_0r1d[32], gate634_0n, initialise);
  C2RI I205 (ifint_0n[0], i_0r0d[0], gate634_0n, initialise);
  C2RI I206 (ifint_0n[1], i_0r0d[1], gate634_0n, initialise);
  C2RI I207 (ifint_0n[2], i_0r0d[2], gate634_0n, initialise);
  C2RI I208 (ifint_0n[3], i_0r0d[3], gate634_0n, initialise);
  C2RI I209 (ifint_0n[4], i_0r0d[4], gate634_0n, initialise);
  C2RI I210 (ifint_0n[5], i_0r0d[5], gate634_0n, initialise);
  C2RI I211 (ifint_0n[6], i_0r0d[6], gate634_0n, initialise);
  C2RI I212 (ifint_0n[7], i_0r0d[7], gate634_0n, initialise);
  C2RI I213 (ifint_0n[8], i_0r0d[8], gate634_0n, initialise);
  C2RI I214 (ifint_0n[9], i_0r0d[9], gate634_0n, initialise);
  C2RI I215 (ifint_0n[10], i_0r0d[10], gate634_0n, initialise);
  C2RI I216 (ifint_0n[11], i_0r0d[11], gate634_0n, initialise);
  C2RI I217 (ifint_0n[12], i_0r0d[12], gate634_0n, initialise);
  C2RI I218 (ifint_0n[13], i_0r0d[13], gate634_0n, initialise);
  C2RI I219 (ifint_0n[14], i_0r0d[14], gate634_0n, initialise);
  C2RI I220 (ifint_0n[15], i_0r0d[15], gate634_0n, initialise);
  C2RI I221 (ifint_0n[16], i_0r0d[16], gate634_0n, initialise);
  C2RI I222 (ifint_0n[17], i_0r0d[17], gate634_0n, initialise);
  C2RI I223 (ifint_0n[18], i_0r0d[18], gate634_0n, initialise);
  C2RI I224 (ifint_0n[19], i_0r0d[19], gate634_0n, initialise);
  C2RI I225 (ifint_0n[20], i_0r0d[20], gate634_0n, initialise);
  C2RI I226 (ifint_0n[21], i_0r0d[21], gate634_0n, initialise);
  C2RI I227 (ifint_0n[22], i_0r0d[22], gate634_0n, initialise);
  C2RI I228 (ifint_0n[23], i_0r0d[23], gate634_0n, initialise);
  C2RI I229 (ifint_0n[24], i_0r0d[24], gate634_0n, initialise);
  C2RI I230 (ifint_0n[25], i_0r0d[25], gate634_0n, initialise);
  C2RI I231 (ifint_0n[26], i_0r0d[26], gate634_0n, initialise);
  C2RI I232 (ifint_0n[27], i_0r0d[27], gate634_0n, initialise);
  C2RI I233 (ifint_0n[28], i_0r0d[28], gate634_0n, initialise);
  C2RI I234 (ifint_0n[29], i_0r0d[29], gate634_0n, initialise);
  C2RI I235 (ifint_0n[30], i_0r0d[30], gate634_0n, initialise);
  C2RI I236 (ifint_0n[31], i_0r0d[31], gate634_0n, initialise);
  C2RI I237 (ifint_0n[32], i_0r0d[32], gate634_0n, initialise);
  C3 I238 (internal_0n[34], complete631_0n[0], complete631_0n[1], complete631_0n[2]);
  C3 I239 (internal_0n[35], complete631_0n[3], complete631_0n[4], complete631_0n[5]);
  C3 I240 (internal_0n[36], complete631_0n[6], complete631_0n[7], complete631_0n[8]);
  C3 I241 (internal_0n[37], complete631_0n[9], complete631_0n[10], complete631_0n[11]);
  C3 I242 (internal_0n[38], complete631_0n[12], complete631_0n[13], complete631_0n[14]);
  C3 I243 (internal_0n[39], complete631_0n[15], complete631_0n[16], complete631_0n[17]);
  C3 I244 (internal_0n[40], complete631_0n[18], complete631_0n[19], complete631_0n[20]);
  C3 I245 (internal_0n[41], complete631_0n[21], complete631_0n[22], complete631_0n[23]);
  C3 I246 (internal_0n[42], complete631_0n[24], complete631_0n[25], complete631_0n[26]);
  C3 I247 (internal_0n[43], complete631_0n[27], complete631_0n[28], complete631_0n[29]);
  C3 I248 (internal_0n[44], complete631_0n[30], complete631_0n[31], complete631_0n[32]);
  C3 I249 (internal_0n[45], complete631_0n[33], complete631_0n[34], complete631_0n[35]);
  C3 I250 (internal_0n[46], complete631_0n[36], complete631_0n[37], complete631_0n[38]);
  C3 I251 (internal_0n[47], complete631_0n[39], complete631_0n[40], complete631_0n[41]);
  C3 I252 (internal_0n[48], complete631_0n[42], complete631_0n[43], complete631_0n[44]);
  C3 I253 (internal_0n[49], complete631_0n[45], complete631_0n[46], complete631_0n[47]);
  C3 I254 (internal_0n[50], complete631_0n[48], complete631_0n[49], complete631_0n[50]);
  C3 I255 (internal_0n[51], complete631_0n[51], complete631_0n[52], complete631_0n[53]);
  C3 I256 (internal_0n[52], complete631_0n[54], complete631_0n[55], complete631_0n[56]);
  C3 I257 (internal_0n[53], complete631_0n[57], complete631_0n[58], complete631_0n[59]);
  C3 I258 (internal_0n[54], complete631_0n[60], complete631_0n[61], complete631_0n[62]);
  C3 I259 (internal_0n[55], complete631_0n[63], complete631_0n[64], complete631_0n[65]);
  C3 I260 (internal_0n[56], internal_0n[34], internal_0n[35], internal_0n[36]);
  C3 I261 (internal_0n[57], internal_0n[37], internal_0n[38], internal_0n[39]);
  C3 I262 (internal_0n[58], internal_0n[40], internal_0n[41], internal_0n[42]);
  C3 I263 (internal_0n[59], internal_0n[43], internal_0n[44], internal_0n[45]);
  C3 I264 (internal_0n[60], internal_0n[46], internal_0n[47], internal_0n[48]);
  C3 I265 (internal_0n[61], internal_0n[49], internal_0n[50], internal_0n[51]);
  C2 I266 (internal_0n[62], internal_0n[52], internal_0n[53]);
  C2 I267 (internal_0n[63], internal_0n[54], internal_0n[55]);
  C3 I268 (internal_0n[64], internal_0n[56], internal_0n[57], internal_0n[58]);
  C3 I269 (internal_0n[65], internal_0n[59], internal_0n[60], internal_0n[61]);
  C2 I270 (internal_0n[66], internal_0n[62], internal_0n[63]);
  C3 I271 (oaint_0n, internal_0n[64], internal_0n[65], internal_0n[66]);
  OR2 I272 (complete631_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I273 (complete631_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I274 (complete631_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I275 (complete631_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I276 (complete631_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I277 (complete631_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I278 (complete631_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I279 (complete631_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I280 (complete631_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I281 (complete631_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I282 (complete631_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I283 (complete631_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I284 (complete631_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I285 (complete631_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I286 (complete631_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I287 (complete631_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I288 (complete631_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I289 (complete631_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I290 (complete631_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I291 (complete631_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I292 (complete631_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I293 (complete631_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I294 (complete631_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I295 (complete631_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I296 (complete631_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I297 (complete631_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I298 (complete631_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I299 (complete631_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I300 (complete631_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I301 (complete631_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I302 (complete631_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I303 (complete631_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I304 (complete631_0n[32], o_0r0d[32], o_0r1d[32]);
  OR2 I305 (complete631_0n[33], o_0r0d[33], o_0r1d[33]);
  OR2 I306 (complete631_0n[34], o_0r0d[34], o_0r1d[34]);
  OR2 I307 (complete631_0n[35], o_0r0d[35], o_0r1d[35]);
  OR2 I308 (complete631_0n[36], o_0r0d[36], o_0r1d[36]);
  OR2 I309 (complete631_0n[37], o_0r0d[37], o_0r1d[37]);
  OR2 I310 (complete631_0n[38], o_0r0d[38], o_0r1d[38]);
  OR2 I311 (complete631_0n[39], o_0r0d[39], o_0r1d[39]);
  OR2 I312 (complete631_0n[40], o_0r0d[40], o_0r1d[40]);
  OR2 I313 (complete631_0n[41], o_0r0d[41], o_0r1d[41]);
  OR2 I314 (complete631_0n[42], o_0r0d[42], o_0r1d[42]);
  OR2 I315 (complete631_0n[43], o_0r0d[43], o_0r1d[43]);
  OR2 I316 (complete631_0n[44], o_0r0d[44], o_0r1d[44]);
  OR2 I317 (complete631_0n[45], o_0r0d[45], o_0r1d[45]);
  OR2 I318 (complete631_0n[46], o_0r0d[46], o_0r1d[46]);
  OR2 I319 (complete631_0n[47], o_0r0d[47], o_0r1d[47]);
  OR2 I320 (complete631_0n[48], o_0r0d[48], o_0r1d[48]);
  OR2 I321 (complete631_0n[49], o_0r0d[49], o_0r1d[49]);
  OR2 I322 (complete631_0n[50], o_0r0d[50], o_0r1d[50]);
  OR2 I323 (complete631_0n[51], o_0r0d[51], o_0r1d[51]);
  OR2 I324 (complete631_0n[52], o_0r0d[52], o_0r1d[52]);
  OR2 I325 (complete631_0n[53], o_0r0d[53], o_0r1d[53]);
  OR2 I326 (complete631_0n[54], o_0r0d[54], o_0r1d[54]);
  OR2 I327 (complete631_0n[55], o_0r0d[55], o_0r1d[55]);
  OR2 I328 (complete631_0n[56], o_0r0d[56], o_0r1d[56]);
  OR2 I329 (complete631_0n[57], o_0r0d[57], o_0r1d[57]);
  OR2 I330 (complete631_0n[58], o_0r0d[58], o_0r1d[58]);
  OR2 I331 (complete631_0n[59], o_0r0d[59], o_0r1d[59]);
  OR2 I332 (complete631_0n[60], o_0r0d[60], o_0r1d[60]);
  OR2 I333 (complete631_0n[61], o_0r0d[61], o_0r1d[61]);
  OR2 I334 (complete631_0n[62], o_0r0d[62], o_0r1d[62]);
  OR2 I335 (complete631_0n[63], o_0r0d[63], o_0r1d[63]);
  OR2 I336 (complete631_0n[64], o_0r0d[64], o_0r1d[64]);
  OR2 I337 (complete631_0n[65], o_0r0d[65], o_0r1d[65]);
  INV I338 (gate630_0n, o_0a);
  C2RI I339 (o_0r1d[0], otint_0n[0], gate630_0n, initialise);
  C2RI I340 (o_0r1d[1], otint_0n[1], gate630_0n, initialise);
  C2RI I341 (o_0r1d[2], otint_0n[2], gate630_0n, initialise);
  C2RI I342 (o_0r1d[3], otint_0n[3], gate630_0n, initialise);
  C2RI I343 (o_0r1d[4], otint_0n[4], gate630_0n, initialise);
  C2RI I344 (o_0r1d[5], otint_0n[5], gate630_0n, initialise);
  C2RI I345 (o_0r1d[6], otint_0n[6], gate630_0n, initialise);
  C2RI I346 (o_0r1d[7], otint_0n[7], gate630_0n, initialise);
  C2RI I347 (o_0r1d[8], otint_0n[8], gate630_0n, initialise);
  C2RI I348 (o_0r1d[9], otint_0n[9], gate630_0n, initialise);
  C2RI I349 (o_0r1d[10], otint_0n[10], gate630_0n, initialise);
  C2RI I350 (o_0r1d[11], otint_0n[11], gate630_0n, initialise);
  C2RI I351 (o_0r1d[12], otint_0n[12], gate630_0n, initialise);
  C2RI I352 (o_0r1d[13], otint_0n[13], gate630_0n, initialise);
  C2RI I353 (o_0r1d[14], otint_0n[14], gate630_0n, initialise);
  C2RI I354 (o_0r1d[15], otint_0n[15], gate630_0n, initialise);
  C2RI I355 (o_0r1d[16], otint_0n[16], gate630_0n, initialise);
  C2RI I356 (o_0r1d[17], otint_0n[17], gate630_0n, initialise);
  C2RI I357 (o_0r1d[18], otint_0n[18], gate630_0n, initialise);
  C2RI I358 (o_0r1d[19], otint_0n[19], gate630_0n, initialise);
  C2RI I359 (o_0r1d[20], otint_0n[20], gate630_0n, initialise);
  C2RI I360 (o_0r1d[21], otint_0n[21], gate630_0n, initialise);
  C2RI I361 (o_0r1d[22], otint_0n[22], gate630_0n, initialise);
  C2RI I362 (o_0r1d[23], otint_0n[23], gate630_0n, initialise);
  C2RI I363 (o_0r1d[24], otint_0n[24], gate630_0n, initialise);
  C2RI I364 (o_0r1d[25], otint_0n[25], gate630_0n, initialise);
  C2RI I365 (o_0r1d[26], otint_0n[26], gate630_0n, initialise);
  C2RI I366 (o_0r1d[27], otint_0n[27], gate630_0n, initialise);
  C2RI I367 (o_0r1d[28], otint_0n[28], gate630_0n, initialise);
  C2RI I368 (o_0r1d[29], otint_0n[29], gate630_0n, initialise);
  C2RI I369 (o_0r1d[30], otint_0n[30], gate630_0n, initialise);
  C2RI I370 (o_0r1d[31], otint_0n[31], gate630_0n, initialise);
  C2RI I371 (o_0r1d[32], otint_0n[32], gate630_0n, initialise);
  C2RI I372 (o_0r1d[33], otint_0n[33], gate630_0n, initialise);
  C2RI I373 (o_0r1d[34], otint_0n[34], gate630_0n, initialise);
  C2RI I374 (o_0r1d[35], otint_0n[35], gate630_0n, initialise);
  C2RI I375 (o_0r1d[36], otint_0n[36], gate630_0n, initialise);
  C2RI I376 (o_0r1d[37], otint_0n[37], gate630_0n, initialise);
  C2RI I377 (o_0r1d[38], otint_0n[38], gate630_0n, initialise);
  C2RI I378 (o_0r1d[39], otint_0n[39], gate630_0n, initialise);
  C2RI I379 (o_0r1d[40], otint_0n[40], gate630_0n, initialise);
  C2RI I380 (o_0r1d[41], otint_0n[41], gate630_0n, initialise);
  C2RI I381 (o_0r1d[42], otint_0n[42], gate630_0n, initialise);
  C2RI I382 (o_0r1d[43], otint_0n[43], gate630_0n, initialise);
  C2RI I383 (o_0r1d[44], otint_0n[44], gate630_0n, initialise);
  C2RI I384 (o_0r1d[45], otint_0n[45], gate630_0n, initialise);
  C2RI I385 (o_0r1d[46], otint_0n[46], gate630_0n, initialise);
  C2RI I386 (o_0r1d[47], otint_0n[47], gate630_0n, initialise);
  C2RI I387 (o_0r1d[48], otint_0n[48], gate630_0n, initialise);
  C2RI I388 (o_0r1d[49], otint_0n[49], gate630_0n, initialise);
  C2RI I389 (o_0r1d[50], otint_0n[50], gate630_0n, initialise);
  C2RI I390 (o_0r1d[51], otint_0n[51], gate630_0n, initialise);
  C2RI I391 (o_0r1d[52], otint_0n[52], gate630_0n, initialise);
  C2RI I392 (o_0r1d[53], otint_0n[53], gate630_0n, initialise);
  C2RI I393 (o_0r1d[54], otint_0n[54], gate630_0n, initialise);
  C2RI I394 (o_0r1d[55], otint_0n[55], gate630_0n, initialise);
  C2RI I395 (o_0r1d[56], otint_0n[56], gate630_0n, initialise);
  C2RI I396 (o_0r1d[57], otint_0n[57], gate630_0n, initialise);
  C2RI I397 (o_0r1d[58], otint_0n[58], gate630_0n, initialise);
  C2RI I398 (o_0r1d[59], otint_0n[59], gate630_0n, initialise);
  C2RI I399 (o_0r1d[60], otint_0n[60], gate630_0n, initialise);
  C2RI I400 (o_0r1d[61], otint_0n[61], gate630_0n, initialise);
  C2RI I401 (o_0r1d[62], otint_0n[62], gate630_0n, initialise);
  C2RI I402 (o_0r1d[63], otint_0n[63], gate630_0n, initialise);
  C2RI I403 (o_0r1d[64], otint_0n[64], gate630_0n, initialise);
  C2RI I404 (o_0r1d[65], otint_0n[65], gate630_0n, initialise);
  C2RI I405 (o_0r0d[0], ofint_0n[0], gate630_0n, initialise);
  C2RI I406 (o_0r0d[1], ofint_0n[1], gate630_0n, initialise);
  C2RI I407 (o_0r0d[2], ofint_0n[2], gate630_0n, initialise);
  C2RI I408 (o_0r0d[3], ofint_0n[3], gate630_0n, initialise);
  C2RI I409 (o_0r0d[4], ofint_0n[4], gate630_0n, initialise);
  C2RI I410 (o_0r0d[5], ofint_0n[5], gate630_0n, initialise);
  C2RI I411 (o_0r0d[6], ofint_0n[6], gate630_0n, initialise);
  C2RI I412 (o_0r0d[7], ofint_0n[7], gate630_0n, initialise);
  C2RI I413 (o_0r0d[8], ofint_0n[8], gate630_0n, initialise);
  C2RI I414 (o_0r0d[9], ofint_0n[9], gate630_0n, initialise);
  C2RI I415 (o_0r0d[10], ofint_0n[10], gate630_0n, initialise);
  C2RI I416 (o_0r0d[11], ofint_0n[11], gate630_0n, initialise);
  C2RI I417 (o_0r0d[12], ofint_0n[12], gate630_0n, initialise);
  C2RI I418 (o_0r0d[13], ofint_0n[13], gate630_0n, initialise);
  C2RI I419 (o_0r0d[14], ofint_0n[14], gate630_0n, initialise);
  C2RI I420 (o_0r0d[15], ofint_0n[15], gate630_0n, initialise);
  C2RI I421 (o_0r0d[16], ofint_0n[16], gate630_0n, initialise);
  C2RI I422 (o_0r0d[17], ofint_0n[17], gate630_0n, initialise);
  C2RI I423 (o_0r0d[18], ofint_0n[18], gate630_0n, initialise);
  C2RI I424 (o_0r0d[19], ofint_0n[19], gate630_0n, initialise);
  C2RI I425 (o_0r0d[20], ofint_0n[20], gate630_0n, initialise);
  C2RI I426 (o_0r0d[21], ofint_0n[21], gate630_0n, initialise);
  C2RI I427 (o_0r0d[22], ofint_0n[22], gate630_0n, initialise);
  C2RI I428 (o_0r0d[23], ofint_0n[23], gate630_0n, initialise);
  C2RI I429 (o_0r0d[24], ofint_0n[24], gate630_0n, initialise);
  C2RI I430 (o_0r0d[25], ofint_0n[25], gate630_0n, initialise);
  C2RI I431 (o_0r0d[26], ofint_0n[26], gate630_0n, initialise);
  C2RI I432 (o_0r0d[27], ofint_0n[27], gate630_0n, initialise);
  C2RI I433 (o_0r0d[28], ofint_0n[28], gate630_0n, initialise);
  C2RI I434 (o_0r0d[29], ofint_0n[29], gate630_0n, initialise);
  C2RI I435 (o_0r0d[30], ofint_0n[30], gate630_0n, initialise);
  C2RI I436 (o_0r0d[31], ofint_0n[31], gate630_0n, initialise);
  C2RI I437 (o_0r0d[32], ofint_0n[32], gate630_0n, initialise);
  C2RI I438 (o_0r0d[33], ofint_0n[33], gate630_0n, initialise);
  C2RI I439 (o_0r0d[34], ofint_0n[34], gate630_0n, initialise);
  C2RI I440 (o_0r0d[35], ofint_0n[35], gate630_0n, initialise);
  C2RI I441 (o_0r0d[36], ofint_0n[36], gate630_0n, initialise);
  C2RI I442 (o_0r0d[37], ofint_0n[37], gate630_0n, initialise);
  C2RI I443 (o_0r0d[38], ofint_0n[38], gate630_0n, initialise);
  C2RI I444 (o_0r0d[39], ofint_0n[39], gate630_0n, initialise);
  C2RI I445 (o_0r0d[40], ofint_0n[40], gate630_0n, initialise);
  C2RI I446 (o_0r0d[41], ofint_0n[41], gate630_0n, initialise);
  C2RI I447 (o_0r0d[42], ofint_0n[42], gate630_0n, initialise);
  C2RI I448 (o_0r0d[43], ofint_0n[43], gate630_0n, initialise);
  C2RI I449 (o_0r0d[44], ofint_0n[44], gate630_0n, initialise);
  C2RI I450 (o_0r0d[45], ofint_0n[45], gate630_0n, initialise);
  C2RI I451 (o_0r0d[46], ofint_0n[46], gate630_0n, initialise);
  C2RI I452 (o_0r0d[47], ofint_0n[47], gate630_0n, initialise);
  C2RI I453 (o_0r0d[48], ofint_0n[48], gate630_0n, initialise);
  C2RI I454 (o_0r0d[49], ofint_0n[49], gate630_0n, initialise);
  C2RI I455 (o_0r0d[50], ofint_0n[50], gate630_0n, initialise);
  C2RI I456 (o_0r0d[51], ofint_0n[51], gate630_0n, initialise);
  C2RI I457 (o_0r0d[52], ofint_0n[52], gate630_0n, initialise);
  C2RI I458 (o_0r0d[53], ofint_0n[53], gate630_0n, initialise);
  C2RI I459 (o_0r0d[54], ofint_0n[54], gate630_0n, initialise);
  C2RI I460 (o_0r0d[55], ofint_0n[55], gate630_0n, initialise);
  C2RI I461 (o_0r0d[56], ofint_0n[56], gate630_0n, initialise);
  C2RI I462 (o_0r0d[57], ofint_0n[57], gate630_0n, initialise);
  C2RI I463 (o_0r0d[58], ofint_0n[58], gate630_0n, initialise);
  C2RI I464 (o_0r0d[59], ofint_0n[59], gate630_0n, initialise);
  C2RI I465 (o_0r0d[60], ofint_0n[60], gate630_0n, initialise);
  C2RI I466 (o_0r0d[61], ofint_0n[61], gate630_0n, initialise);
  C2RI I467 (o_0r0d[62], ofint_0n[62], gate630_0n, initialise);
  C2RI I468 (o_0r0d[63], ofint_0n[63], gate630_0n, initialise);
  C2RI I469 (o_0r0d[64], ofint_0n[64], gate630_0n, initialise);
  C2RI I470 (o_0r0d[65], ofint_0n[65], gate630_0n, initialise);
  assign otint_0n[0] = itint_0n[0];
  assign otint_0n[1] = itint_0n[1];
  assign otint_0n[2] = itint_0n[2];
  assign otint_0n[3] = itint_0n[3];
  assign otint_0n[4] = itint_0n[4];
  assign otint_0n[5] = itint_0n[5];
  assign otint_0n[6] = itint_0n[6];
  assign otint_0n[7] = itint_0n[7];
  assign otint_0n[8] = itint_0n[8];
  assign otint_0n[9] = itint_0n[9];
  assign otint_0n[10] = itint_0n[10];
  assign otint_0n[11] = itint_0n[11];
  assign otint_0n[12] = itint_0n[12];
  assign otint_0n[13] = itint_0n[13];
  assign otint_0n[14] = itint_0n[14];
  assign otint_0n[15] = itint_0n[15];
  assign otint_0n[16] = itint_0n[16];
  assign otint_0n[17] = itint_0n[17];
  assign otint_0n[18] = itint_0n[18];
  assign otint_0n[19] = itint_0n[19];
  assign otint_0n[20] = itint_0n[20];
  assign otint_0n[21] = itint_0n[21];
  assign otint_0n[22] = itint_0n[22];
  assign otint_0n[23] = itint_0n[23];
  assign otint_0n[24] = itint_0n[24];
  assign otint_0n[25] = itint_0n[25];
  assign otint_0n[26] = itint_0n[26];
  assign otint_0n[27] = itint_0n[27];
  assign otint_0n[28] = itint_0n[28];
  assign otint_0n[29] = itint_0n[29];
  assign otint_0n[30] = itint_0n[30];
  assign otint_0n[31] = itint_0n[31];
  assign otint_0n[32] = itint_0n[32];
  assign otint_0n[33] = itint_1n[0];
  assign otint_0n[34] = itint_1n[1];
  assign otint_0n[35] = itint_1n[2];
  assign otint_0n[36] = itint_1n[3];
  assign otint_0n[37] = itint_1n[4];
  assign otint_0n[38] = itint_1n[5];
  assign otint_0n[39] = itint_1n[6];
  assign otint_0n[40] = itint_1n[7];
  assign otint_0n[41] = itint_1n[8];
  assign otint_0n[42] = itint_1n[9];
  assign otint_0n[43] = itint_1n[10];
  assign otint_0n[44] = itint_1n[11];
  assign otint_0n[45] = itint_1n[12];
  assign otint_0n[46] = itint_1n[13];
  assign otint_0n[47] = itint_1n[14];
  assign otint_0n[48] = itint_1n[15];
  assign otint_0n[49] = itint_1n[16];
  assign otint_0n[50] = itint_1n[17];
  assign otint_0n[51] = itint_1n[18];
  assign otint_0n[52] = itint_1n[19];
  assign otint_0n[53] = itint_1n[20];
  assign otint_0n[54] = itint_1n[21];
  assign otint_0n[55] = itint_1n[22];
  assign otint_0n[56] = itint_1n[23];
  assign otint_0n[57] = itint_1n[24];
  assign otint_0n[58] = itint_1n[25];
  assign otint_0n[59] = itint_1n[26];
  assign otint_0n[60] = itint_1n[27];
  assign otint_0n[61] = itint_1n[28];
  assign otint_0n[62] = itint_1n[29];
  assign otint_0n[63] = itint_1n[30];
  assign otint_0n[64] = itint_1n[31];
  assign otint_0n[65] = itint_1n[32];
  assign ofint_0n[0] = ifint_0n[0];
  assign ofint_0n[1] = ifint_0n[1];
  assign ofint_0n[2] = ifint_0n[2];
  assign ofint_0n[3] = ifint_0n[3];
  assign ofint_0n[4] = ifint_0n[4];
  assign ofint_0n[5] = ifint_0n[5];
  assign ofint_0n[6] = ifint_0n[6];
  assign ofint_0n[7] = ifint_0n[7];
  assign ofint_0n[8] = ifint_0n[8];
  assign ofint_0n[9] = ifint_0n[9];
  assign ofint_0n[10] = ifint_0n[10];
  assign ofint_0n[11] = ifint_0n[11];
  assign ofint_0n[12] = ifint_0n[12];
  assign ofint_0n[13] = ifint_0n[13];
  assign ofint_0n[14] = ifint_0n[14];
  assign ofint_0n[15] = ifint_0n[15];
  assign ofint_0n[16] = ifint_0n[16];
  assign ofint_0n[17] = ifint_0n[17];
  assign ofint_0n[18] = ifint_0n[18];
  assign ofint_0n[19] = ifint_0n[19];
  assign ofint_0n[20] = ifint_0n[20];
  assign ofint_0n[21] = ifint_0n[21];
  assign ofint_0n[22] = ifint_0n[22];
  assign ofint_0n[23] = ifint_0n[23];
  assign ofint_0n[24] = ifint_0n[24];
  assign ofint_0n[25] = ifint_0n[25];
  assign ofint_0n[26] = ifint_0n[26];
  assign ofint_0n[27] = ifint_0n[27];
  assign ofint_0n[28] = ifint_0n[28];
  assign ofint_0n[29] = ifint_0n[29];
  assign ofint_0n[30] = ifint_0n[30];
  assign ofint_0n[31] = ifint_0n[31];
  assign ofint_0n[32] = ifint_0n[32];
  assign ofint_0n[33] = ifint_1n[0];
  assign ofint_0n[34] = ifint_1n[1];
  assign ofint_0n[35] = ifint_1n[2];
  assign ofint_0n[36] = ifint_1n[3];
  assign ofint_0n[37] = ifint_1n[4];
  assign ofint_0n[38] = ifint_1n[5];
  assign ofint_0n[39] = ifint_1n[6];
  assign ofint_0n[40] = ifint_1n[7];
  assign ofint_0n[41] = ifint_1n[8];
  assign ofint_0n[42] = ifint_1n[9];
  assign ofint_0n[43] = ifint_1n[10];
  assign ofint_0n[44] = ifint_1n[11];
  assign ofint_0n[45] = ifint_1n[12];
  assign ofint_0n[46] = ifint_1n[13];
  assign ofint_0n[47] = ifint_1n[14];
  assign ofint_0n[48] = ifint_1n[15];
  assign ofint_0n[49] = ifint_1n[16];
  assign ofint_0n[50] = ifint_1n[17];
  assign ofint_0n[51] = ifint_1n[18];
  assign ofint_0n[52] = ifint_1n[19];
  assign ofint_0n[53] = ifint_1n[20];
  assign ofint_0n[54] = ifint_1n[21];
  assign ofint_0n[55] = ifint_1n[22];
  assign ofint_0n[56] = ifint_1n[23];
  assign ofint_0n[57] = ifint_1n[24];
  assign ofint_0n[58] = ifint_1n[25];
  assign ofint_0n[59] = ifint_1n[26];
  assign ofint_0n[60] = ifint_1n[27];
  assign ofint_0n[61] = ifint_1n[28];
  assign ofint_0n[62] = ifint_1n[29];
  assign ofint_0n[63] = ifint_1n[30];
  assign ofint_0n[64] = ifint_1n[31];
  assign ofint_0n[65] = ifint_1n[32];
endmodule

module BrzJ_l12__2834_200_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [33:0] i_0r0d;
  input [33:0] i_0r1d;
  output i_0a;
  input i_1r;
  output i_1a;
  output [33:0] o_0r0d;
  output [33:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [35:0] internal_0n;
  wire [33:0] ofint_0n;
  wire [33:0] otint_0n;
  wire oaint_0n;
  wire [33:0] ifint_0n;
  wire ifint_1n;
  wire [33:0] itint_0n;
  wire iaint_0n;
  wire iaint_1n;
  wire gate650_0n;
  wire [33:0] complete647_0n;
  wire gate646_0n;
  wire [33:0] complete643_0n;
  wire gate642_0n;
  wire [33:0] joint_0n;
  wire [33:0] joinf_0n;
  wire icomplete_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign i_1a = ifint_1n;
  INV I3 (gate650_0n, iaint_1n);
  C2RI I4 (ifint_1n, i_1r, gate650_0n, initialise);
  C3 I5 (internal_0n[0], complete647_0n[0], complete647_0n[1], complete647_0n[2]);
  C3 I6 (internal_0n[1], complete647_0n[3], complete647_0n[4], complete647_0n[5]);
  C3 I7 (internal_0n[2], complete647_0n[6], complete647_0n[7], complete647_0n[8]);
  C3 I8 (internal_0n[3], complete647_0n[9], complete647_0n[10], complete647_0n[11]);
  C3 I9 (internal_0n[4], complete647_0n[12], complete647_0n[13], complete647_0n[14]);
  C3 I10 (internal_0n[5], complete647_0n[15], complete647_0n[16], complete647_0n[17]);
  C3 I11 (internal_0n[6], complete647_0n[18], complete647_0n[19], complete647_0n[20]);
  C3 I12 (internal_0n[7], complete647_0n[21], complete647_0n[22], complete647_0n[23]);
  C3 I13 (internal_0n[8], complete647_0n[24], complete647_0n[25], complete647_0n[26]);
  C3 I14 (internal_0n[9], complete647_0n[27], complete647_0n[28], complete647_0n[29]);
  C2 I15 (internal_0n[10], complete647_0n[30], complete647_0n[31]);
  C2 I16 (internal_0n[11], complete647_0n[32], complete647_0n[33]);
  C3 I17 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I18 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I19 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I20 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I21 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I22 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I23 (i_0a, internal_0n[16], internal_0n[17]);
  OR2 I24 (complete647_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I25 (complete647_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I26 (complete647_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I27 (complete647_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I28 (complete647_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I29 (complete647_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I30 (complete647_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I31 (complete647_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I32 (complete647_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I33 (complete647_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I34 (complete647_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I35 (complete647_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I36 (complete647_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I37 (complete647_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I38 (complete647_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I39 (complete647_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I40 (complete647_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I41 (complete647_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I42 (complete647_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I43 (complete647_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I44 (complete647_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I45 (complete647_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I46 (complete647_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I47 (complete647_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I48 (complete647_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I49 (complete647_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I50 (complete647_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I51 (complete647_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I52 (complete647_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I53 (complete647_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I54 (complete647_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I55 (complete647_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I56 (complete647_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I57 (complete647_0n[33], ifint_0n[33], itint_0n[33]);
  INV I58 (gate646_0n, iaint_0n);
  C2RI I59 (itint_0n[0], i_0r1d[0], gate646_0n, initialise);
  C2RI I60 (itint_0n[1], i_0r1d[1], gate646_0n, initialise);
  C2RI I61 (itint_0n[2], i_0r1d[2], gate646_0n, initialise);
  C2RI I62 (itint_0n[3], i_0r1d[3], gate646_0n, initialise);
  C2RI I63 (itint_0n[4], i_0r1d[4], gate646_0n, initialise);
  C2RI I64 (itint_0n[5], i_0r1d[5], gate646_0n, initialise);
  C2RI I65 (itint_0n[6], i_0r1d[6], gate646_0n, initialise);
  C2RI I66 (itint_0n[7], i_0r1d[7], gate646_0n, initialise);
  C2RI I67 (itint_0n[8], i_0r1d[8], gate646_0n, initialise);
  C2RI I68 (itint_0n[9], i_0r1d[9], gate646_0n, initialise);
  C2RI I69 (itint_0n[10], i_0r1d[10], gate646_0n, initialise);
  C2RI I70 (itint_0n[11], i_0r1d[11], gate646_0n, initialise);
  C2RI I71 (itint_0n[12], i_0r1d[12], gate646_0n, initialise);
  C2RI I72 (itint_0n[13], i_0r1d[13], gate646_0n, initialise);
  C2RI I73 (itint_0n[14], i_0r1d[14], gate646_0n, initialise);
  C2RI I74 (itint_0n[15], i_0r1d[15], gate646_0n, initialise);
  C2RI I75 (itint_0n[16], i_0r1d[16], gate646_0n, initialise);
  C2RI I76 (itint_0n[17], i_0r1d[17], gate646_0n, initialise);
  C2RI I77 (itint_0n[18], i_0r1d[18], gate646_0n, initialise);
  C2RI I78 (itint_0n[19], i_0r1d[19], gate646_0n, initialise);
  C2RI I79 (itint_0n[20], i_0r1d[20], gate646_0n, initialise);
  C2RI I80 (itint_0n[21], i_0r1d[21], gate646_0n, initialise);
  C2RI I81 (itint_0n[22], i_0r1d[22], gate646_0n, initialise);
  C2RI I82 (itint_0n[23], i_0r1d[23], gate646_0n, initialise);
  C2RI I83 (itint_0n[24], i_0r1d[24], gate646_0n, initialise);
  C2RI I84 (itint_0n[25], i_0r1d[25], gate646_0n, initialise);
  C2RI I85 (itint_0n[26], i_0r1d[26], gate646_0n, initialise);
  C2RI I86 (itint_0n[27], i_0r1d[27], gate646_0n, initialise);
  C2RI I87 (itint_0n[28], i_0r1d[28], gate646_0n, initialise);
  C2RI I88 (itint_0n[29], i_0r1d[29], gate646_0n, initialise);
  C2RI I89 (itint_0n[30], i_0r1d[30], gate646_0n, initialise);
  C2RI I90 (itint_0n[31], i_0r1d[31], gate646_0n, initialise);
  C2RI I91 (itint_0n[32], i_0r1d[32], gate646_0n, initialise);
  C2RI I92 (itint_0n[33], i_0r1d[33], gate646_0n, initialise);
  C2RI I93 (ifint_0n[0], i_0r0d[0], gate646_0n, initialise);
  C2RI I94 (ifint_0n[1], i_0r0d[1], gate646_0n, initialise);
  C2RI I95 (ifint_0n[2], i_0r0d[2], gate646_0n, initialise);
  C2RI I96 (ifint_0n[3], i_0r0d[3], gate646_0n, initialise);
  C2RI I97 (ifint_0n[4], i_0r0d[4], gate646_0n, initialise);
  C2RI I98 (ifint_0n[5], i_0r0d[5], gate646_0n, initialise);
  C2RI I99 (ifint_0n[6], i_0r0d[6], gate646_0n, initialise);
  C2RI I100 (ifint_0n[7], i_0r0d[7], gate646_0n, initialise);
  C2RI I101 (ifint_0n[8], i_0r0d[8], gate646_0n, initialise);
  C2RI I102 (ifint_0n[9], i_0r0d[9], gate646_0n, initialise);
  C2RI I103 (ifint_0n[10], i_0r0d[10], gate646_0n, initialise);
  C2RI I104 (ifint_0n[11], i_0r0d[11], gate646_0n, initialise);
  C2RI I105 (ifint_0n[12], i_0r0d[12], gate646_0n, initialise);
  C2RI I106 (ifint_0n[13], i_0r0d[13], gate646_0n, initialise);
  C2RI I107 (ifint_0n[14], i_0r0d[14], gate646_0n, initialise);
  C2RI I108 (ifint_0n[15], i_0r0d[15], gate646_0n, initialise);
  C2RI I109 (ifint_0n[16], i_0r0d[16], gate646_0n, initialise);
  C2RI I110 (ifint_0n[17], i_0r0d[17], gate646_0n, initialise);
  C2RI I111 (ifint_0n[18], i_0r0d[18], gate646_0n, initialise);
  C2RI I112 (ifint_0n[19], i_0r0d[19], gate646_0n, initialise);
  C2RI I113 (ifint_0n[20], i_0r0d[20], gate646_0n, initialise);
  C2RI I114 (ifint_0n[21], i_0r0d[21], gate646_0n, initialise);
  C2RI I115 (ifint_0n[22], i_0r0d[22], gate646_0n, initialise);
  C2RI I116 (ifint_0n[23], i_0r0d[23], gate646_0n, initialise);
  C2RI I117 (ifint_0n[24], i_0r0d[24], gate646_0n, initialise);
  C2RI I118 (ifint_0n[25], i_0r0d[25], gate646_0n, initialise);
  C2RI I119 (ifint_0n[26], i_0r0d[26], gate646_0n, initialise);
  C2RI I120 (ifint_0n[27], i_0r0d[27], gate646_0n, initialise);
  C2RI I121 (ifint_0n[28], i_0r0d[28], gate646_0n, initialise);
  C2RI I122 (ifint_0n[29], i_0r0d[29], gate646_0n, initialise);
  C2RI I123 (ifint_0n[30], i_0r0d[30], gate646_0n, initialise);
  C2RI I124 (ifint_0n[31], i_0r0d[31], gate646_0n, initialise);
  C2RI I125 (ifint_0n[32], i_0r0d[32], gate646_0n, initialise);
  C2RI I126 (ifint_0n[33], i_0r0d[33], gate646_0n, initialise);
  C3 I127 (internal_0n[18], complete643_0n[0], complete643_0n[1], complete643_0n[2]);
  C3 I128 (internal_0n[19], complete643_0n[3], complete643_0n[4], complete643_0n[5]);
  C3 I129 (internal_0n[20], complete643_0n[6], complete643_0n[7], complete643_0n[8]);
  C3 I130 (internal_0n[21], complete643_0n[9], complete643_0n[10], complete643_0n[11]);
  C3 I131 (internal_0n[22], complete643_0n[12], complete643_0n[13], complete643_0n[14]);
  C3 I132 (internal_0n[23], complete643_0n[15], complete643_0n[16], complete643_0n[17]);
  C3 I133 (internal_0n[24], complete643_0n[18], complete643_0n[19], complete643_0n[20]);
  C3 I134 (internal_0n[25], complete643_0n[21], complete643_0n[22], complete643_0n[23]);
  C3 I135 (internal_0n[26], complete643_0n[24], complete643_0n[25], complete643_0n[26]);
  C3 I136 (internal_0n[27], complete643_0n[27], complete643_0n[28], complete643_0n[29]);
  C2 I137 (internal_0n[28], complete643_0n[30], complete643_0n[31]);
  C2 I138 (internal_0n[29], complete643_0n[32], complete643_0n[33]);
  C3 I139 (internal_0n[30], internal_0n[18], internal_0n[19], internal_0n[20]);
  C3 I140 (internal_0n[31], internal_0n[21], internal_0n[22], internal_0n[23]);
  C3 I141 (internal_0n[32], internal_0n[24], internal_0n[25], internal_0n[26]);
  C3 I142 (internal_0n[33], internal_0n[27], internal_0n[28], internal_0n[29]);
  C2 I143 (internal_0n[34], internal_0n[30], internal_0n[31]);
  C2 I144 (internal_0n[35], internal_0n[32], internal_0n[33]);
  C2 I145 (oaint_0n, internal_0n[34], internal_0n[35]);
  OR2 I146 (complete643_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I147 (complete643_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I148 (complete643_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I149 (complete643_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I150 (complete643_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I151 (complete643_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I152 (complete643_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I153 (complete643_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I154 (complete643_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I155 (complete643_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I156 (complete643_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I157 (complete643_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I158 (complete643_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I159 (complete643_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I160 (complete643_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I161 (complete643_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I162 (complete643_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I163 (complete643_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I164 (complete643_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I165 (complete643_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I166 (complete643_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I167 (complete643_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I168 (complete643_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I169 (complete643_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I170 (complete643_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I171 (complete643_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I172 (complete643_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I173 (complete643_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I174 (complete643_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I175 (complete643_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I176 (complete643_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I177 (complete643_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I178 (complete643_0n[32], o_0r0d[32], o_0r1d[32]);
  OR2 I179 (complete643_0n[33], o_0r0d[33], o_0r1d[33]);
  INV I180 (gate642_0n, o_0a);
  C2RI I181 (o_0r1d[0], otint_0n[0], gate642_0n, initialise);
  C2RI I182 (o_0r1d[1], otint_0n[1], gate642_0n, initialise);
  C2RI I183 (o_0r1d[2], otint_0n[2], gate642_0n, initialise);
  C2RI I184 (o_0r1d[3], otint_0n[3], gate642_0n, initialise);
  C2RI I185 (o_0r1d[4], otint_0n[4], gate642_0n, initialise);
  C2RI I186 (o_0r1d[5], otint_0n[5], gate642_0n, initialise);
  C2RI I187 (o_0r1d[6], otint_0n[6], gate642_0n, initialise);
  C2RI I188 (o_0r1d[7], otint_0n[7], gate642_0n, initialise);
  C2RI I189 (o_0r1d[8], otint_0n[8], gate642_0n, initialise);
  C2RI I190 (o_0r1d[9], otint_0n[9], gate642_0n, initialise);
  C2RI I191 (o_0r1d[10], otint_0n[10], gate642_0n, initialise);
  C2RI I192 (o_0r1d[11], otint_0n[11], gate642_0n, initialise);
  C2RI I193 (o_0r1d[12], otint_0n[12], gate642_0n, initialise);
  C2RI I194 (o_0r1d[13], otint_0n[13], gate642_0n, initialise);
  C2RI I195 (o_0r1d[14], otint_0n[14], gate642_0n, initialise);
  C2RI I196 (o_0r1d[15], otint_0n[15], gate642_0n, initialise);
  C2RI I197 (o_0r1d[16], otint_0n[16], gate642_0n, initialise);
  C2RI I198 (o_0r1d[17], otint_0n[17], gate642_0n, initialise);
  C2RI I199 (o_0r1d[18], otint_0n[18], gate642_0n, initialise);
  C2RI I200 (o_0r1d[19], otint_0n[19], gate642_0n, initialise);
  C2RI I201 (o_0r1d[20], otint_0n[20], gate642_0n, initialise);
  C2RI I202 (o_0r1d[21], otint_0n[21], gate642_0n, initialise);
  C2RI I203 (o_0r1d[22], otint_0n[22], gate642_0n, initialise);
  C2RI I204 (o_0r1d[23], otint_0n[23], gate642_0n, initialise);
  C2RI I205 (o_0r1d[24], otint_0n[24], gate642_0n, initialise);
  C2RI I206 (o_0r1d[25], otint_0n[25], gate642_0n, initialise);
  C2RI I207 (o_0r1d[26], otint_0n[26], gate642_0n, initialise);
  C2RI I208 (o_0r1d[27], otint_0n[27], gate642_0n, initialise);
  C2RI I209 (o_0r1d[28], otint_0n[28], gate642_0n, initialise);
  C2RI I210 (o_0r1d[29], otint_0n[29], gate642_0n, initialise);
  C2RI I211 (o_0r1d[30], otint_0n[30], gate642_0n, initialise);
  C2RI I212 (o_0r1d[31], otint_0n[31], gate642_0n, initialise);
  C2RI I213 (o_0r1d[32], otint_0n[32], gate642_0n, initialise);
  C2RI I214 (o_0r1d[33], otint_0n[33], gate642_0n, initialise);
  C2RI I215 (o_0r0d[0], ofint_0n[0], gate642_0n, initialise);
  C2RI I216 (o_0r0d[1], ofint_0n[1], gate642_0n, initialise);
  C2RI I217 (o_0r0d[2], ofint_0n[2], gate642_0n, initialise);
  C2RI I218 (o_0r0d[3], ofint_0n[3], gate642_0n, initialise);
  C2RI I219 (o_0r0d[4], ofint_0n[4], gate642_0n, initialise);
  C2RI I220 (o_0r0d[5], ofint_0n[5], gate642_0n, initialise);
  C2RI I221 (o_0r0d[6], ofint_0n[6], gate642_0n, initialise);
  C2RI I222 (o_0r0d[7], ofint_0n[7], gate642_0n, initialise);
  C2RI I223 (o_0r0d[8], ofint_0n[8], gate642_0n, initialise);
  C2RI I224 (o_0r0d[9], ofint_0n[9], gate642_0n, initialise);
  C2RI I225 (o_0r0d[10], ofint_0n[10], gate642_0n, initialise);
  C2RI I226 (o_0r0d[11], ofint_0n[11], gate642_0n, initialise);
  C2RI I227 (o_0r0d[12], ofint_0n[12], gate642_0n, initialise);
  C2RI I228 (o_0r0d[13], ofint_0n[13], gate642_0n, initialise);
  C2RI I229 (o_0r0d[14], ofint_0n[14], gate642_0n, initialise);
  C2RI I230 (o_0r0d[15], ofint_0n[15], gate642_0n, initialise);
  C2RI I231 (o_0r0d[16], ofint_0n[16], gate642_0n, initialise);
  C2RI I232 (o_0r0d[17], ofint_0n[17], gate642_0n, initialise);
  C2RI I233 (o_0r0d[18], ofint_0n[18], gate642_0n, initialise);
  C2RI I234 (o_0r0d[19], ofint_0n[19], gate642_0n, initialise);
  C2RI I235 (o_0r0d[20], ofint_0n[20], gate642_0n, initialise);
  C2RI I236 (o_0r0d[21], ofint_0n[21], gate642_0n, initialise);
  C2RI I237 (o_0r0d[22], ofint_0n[22], gate642_0n, initialise);
  C2RI I238 (o_0r0d[23], ofint_0n[23], gate642_0n, initialise);
  C2RI I239 (o_0r0d[24], ofint_0n[24], gate642_0n, initialise);
  C2RI I240 (o_0r0d[25], ofint_0n[25], gate642_0n, initialise);
  C2RI I241 (o_0r0d[26], ofint_0n[26], gate642_0n, initialise);
  C2RI I242 (o_0r0d[27], ofint_0n[27], gate642_0n, initialise);
  C2RI I243 (o_0r0d[28], ofint_0n[28], gate642_0n, initialise);
  C2RI I244 (o_0r0d[29], ofint_0n[29], gate642_0n, initialise);
  C2RI I245 (o_0r0d[30], ofint_0n[30], gate642_0n, initialise);
  C2RI I246 (o_0r0d[31], ofint_0n[31], gate642_0n, initialise);
  C2RI I247 (o_0r0d[32], ofint_0n[32], gate642_0n, initialise);
  C2RI I248 (o_0r0d[33], ofint_0n[33], gate642_0n, initialise);
  assign otint_0n[1] = joint_0n[1];
  assign otint_0n[2] = joint_0n[2];
  assign otint_0n[3] = joint_0n[3];
  assign otint_0n[4] = joint_0n[4];
  assign otint_0n[5] = joint_0n[5];
  assign otint_0n[6] = joint_0n[6];
  assign otint_0n[7] = joint_0n[7];
  assign otint_0n[8] = joint_0n[8];
  assign otint_0n[9] = joint_0n[9];
  assign otint_0n[10] = joint_0n[10];
  assign otint_0n[11] = joint_0n[11];
  assign otint_0n[12] = joint_0n[12];
  assign otint_0n[13] = joint_0n[13];
  assign otint_0n[14] = joint_0n[14];
  assign otint_0n[15] = joint_0n[15];
  assign otint_0n[16] = joint_0n[16];
  assign otint_0n[17] = joint_0n[17];
  assign otint_0n[18] = joint_0n[18];
  assign otint_0n[19] = joint_0n[19];
  assign otint_0n[20] = joint_0n[20];
  assign otint_0n[21] = joint_0n[21];
  assign otint_0n[22] = joint_0n[22];
  assign otint_0n[23] = joint_0n[23];
  assign otint_0n[24] = joint_0n[24];
  assign otint_0n[25] = joint_0n[25];
  assign otint_0n[26] = joint_0n[26];
  assign otint_0n[27] = joint_0n[27];
  assign otint_0n[28] = joint_0n[28];
  assign otint_0n[29] = joint_0n[29];
  assign otint_0n[30] = joint_0n[30];
  assign otint_0n[31] = joint_0n[31];
  assign otint_0n[32] = joint_0n[32];
  assign otint_0n[33] = joint_0n[33];
  assign ofint_0n[1] = joinf_0n[1];
  assign ofint_0n[2] = joinf_0n[2];
  assign ofint_0n[3] = joinf_0n[3];
  assign ofint_0n[4] = joinf_0n[4];
  assign ofint_0n[5] = joinf_0n[5];
  assign ofint_0n[6] = joinf_0n[6];
  assign ofint_0n[7] = joinf_0n[7];
  assign ofint_0n[8] = joinf_0n[8];
  assign ofint_0n[9] = joinf_0n[9];
  assign ofint_0n[10] = joinf_0n[10];
  assign ofint_0n[11] = joinf_0n[11];
  assign ofint_0n[12] = joinf_0n[12];
  assign ofint_0n[13] = joinf_0n[13];
  assign ofint_0n[14] = joinf_0n[14];
  assign ofint_0n[15] = joinf_0n[15];
  assign ofint_0n[16] = joinf_0n[16];
  assign ofint_0n[17] = joinf_0n[17];
  assign ofint_0n[18] = joinf_0n[18];
  assign ofint_0n[19] = joinf_0n[19];
  assign ofint_0n[20] = joinf_0n[20];
  assign ofint_0n[21] = joinf_0n[21];
  assign ofint_0n[22] = joinf_0n[22];
  assign ofint_0n[23] = joinf_0n[23];
  assign ofint_0n[24] = joinf_0n[24];
  assign ofint_0n[25] = joinf_0n[25];
  assign ofint_0n[26] = joinf_0n[26];
  assign ofint_0n[27] = joinf_0n[27];
  assign ofint_0n[28] = joinf_0n[28];
  assign ofint_0n[29] = joinf_0n[29];
  assign ofint_0n[30] = joinf_0n[30];
  assign ofint_0n[31] = joinf_0n[31];
  assign ofint_0n[32] = joinf_0n[32];
  assign ofint_0n[33] = joinf_0n[33];
  C2 I315 (otint_0n[0], joint_0n[0], icomplete_0n);
  C2 I316 (ofint_0n[0], joinf_0n[0], icomplete_0n);
  assign icomplete_0n = ifint_1n;
  assign joint_0n[0] = itint_0n[0];
  assign joint_0n[1] = itint_0n[1];
  assign joint_0n[2] = itint_0n[2];
  assign joint_0n[3] = itint_0n[3];
  assign joint_0n[4] = itint_0n[4];
  assign joint_0n[5] = itint_0n[5];
  assign joint_0n[6] = itint_0n[6];
  assign joint_0n[7] = itint_0n[7];
  assign joint_0n[8] = itint_0n[8];
  assign joint_0n[9] = itint_0n[9];
  assign joint_0n[10] = itint_0n[10];
  assign joint_0n[11] = itint_0n[11];
  assign joint_0n[12] = itint_0n[12];
  assign joint_0n[13] = itint_0n[13];
  assign joint_0n[14] = itint_0n[14];
  assign joint_0n[15] = itint_0n[15];
  assign joint_0n[16] = itint_0n[16];
  assign joint_0n[17] = itint_0n[17];
  assign joint_0n[18] = itint_0n[18];
  assign joint_0n[19] = itint_0n[19];
  assign joint_0n[20] = itint_0n[20];
  assign joint_0n[21] = itint_0n[21];
  assign joint_0n[22] = itint_0n[22];
  assign joint_0n[23] = itint_0n[23];
  assign joint_0n[24] = itint_0n[24];
  assign joint_0n[25] = itint_0n[25];
  assign joint_0n[26] = itint_0n[26];
  assign joint_0n[27] = itint_0n[27];
  assign joint_0n[28] = itint_0n[28];
  assign joint_0n[29] = itint_0n[29];
  assign joint_0n[30] = itint_0n[30];
  assign joint_0n[31] = itint_0n[31];
  assign joint_0n[32] = itint_0n[32];
  assign joint_0n[33] = itint_0n[33];
  assign joinf_0n[0] = ifint_0n[0];
  assign joinf_0n[1] = ifint_0n[1];
  assign joinf_0n[2] = ifint_0n[2];
  assign joinf_0n[3] = ifint_0n[3];
  assign joinf_0n[4] = ifint_0n[4];
  assign joinf_0n[5] = ifint_0n[5];
  assign joinf_0n[6] = ifint_0n[6];
  assign joinf_0n[7] = ifint_0n[7];
  assign joinf_0n[8] = ifint_0n[8];
  assign joinf_0n[9] = ifint_0n[9];
  assign joinf_0n[10] = ifint_0n[10];
  assign joinf_0n[11] = ifint_0n[11];
  assign joinf_0n[12] = ifint_0n[12];
  assign joinf_0n[13] = ifint_0n[13];
  assign joinf_0n[14] = ifint_0n[14];
  assign joinf_0n[15] = ifint_0n[15];
  assign joinf_0n[16] = ifint_0n[16];
  assign joinf_0n[17] = ifint_0n[17];
  assign joinf_0n[18] = ifint_0n[18];
  assign joinf_0n[19] = ifint_0n[19];
  assign joinf_0n[20] = ifint_0n[20];
  assign joinf_0n[21] = ifint_0n[21];
  assign joinf_0n[22] = ifint_0n[22];
  assign joinf_0n[23] = ifint_0n[23];
  assign joinf_0n[24] = ifint_0n[24];
  assign joinf_0n[25] = ifint_0n[25];
  assign joinf_0n[26] = ifint_0n[26];
  assign joinf_0n[27] = ifint_0n[27];
  assign joinf_0n[28] = ifint_0n[28];
  assign joinf_0n[29] = ifint_0n[29];
  assign joinf_0n[30] = ifint_0n[30];
  assign joinf_0n[31] = ifint_0n[31];
  assign joinf_0n[32] = ifint_0n[32];
  assign joinf_0n[33] = ifint_0n[33];
endmodule

module BrzJ_l12__2834_201_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [33:0] i_0r0d;
  input [33:0] i_0r1d;
  output i_0a;
  input i_1r0d;
  input i_1r1d;
  output i_1a;
  output [34:0] o_0r0d;
  output [34:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [35:0] internal_0n;
  wire [34:0] ofint_0n;
  wire [34:0] otint_0n;
  wire oaint_0n;
  wire [33:0] ifint_0n;
  wire ifint_1n;
  wire [33:0] itint_0n;
  wire itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire complete662_0n;
  wire gate661_0n;
  wire [33:0] complete658_0n;
  wire gate657_0n;
  wire [34:0] complete654_0n;
  wire gate653_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign i_1a = complete662_0n;
  OR2 I3 (complete662_0n, ifint_1n, itint_1n);
  INV I4 (gate661_0n, iaint_1n);
  C2RI I5 (itint_1n, i_1r1d, gate661_0n, initialise);
  C2RI I6 (ifint_1n, i_1r0d, gate661_0n, initialise);
  C3 I7 (internal_0n[0], complete658_0n[0], complete658_0n[1], complete658_0n[2]);
  C3 I8 (internal_0n[1], complete658_0n[3], complete658_0n[4], complete658_0n[5]);
  C3 I9 (internal_0n[2], complete658_0n[6], complete658_0n[7], complete658_0n[8]);
  C3 I10 (internal_0n[3], complete658_0n[9], complete658_0n[10], complete658_0n[11]);
  C3 I11 (internal_0n[4], complete658_0n[12], complete658_0n[13], complete658_0n[14]);
  C3 I12 (internal_0n[5], complete658_0n[15], complete658_0n[16], complete658_0n[17]);
  C3 I13 (internal_0n[6], complete658_0n[18], complete658_0n[19], complete658_0n[20]);
  C3 I14 (internal_0n[7], complete658_0n[21], complete658_0n[22], complete658_0n[23]);
  C3 I15 (internal_0n[8], complete658_0n[24], complete658_0n[25], complete658_0n[26]);
  C3 I16 (internal_0n[9], complete658_0n[27], complete658_0n[28], complete658_0n[29]);
  C2 I17 (internal_0n[10], complete658_0n[30], complete658_0n[31]);
  C2 I18 (internal_0n[11], complete658_0n[32], complete658_0n[33]);
  C3 I19 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I20 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I21 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I22 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I23 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I24 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I25 (i_0a, internal_0n[16], internal_0n[17]);
  OR2 I26 (complete658_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I27 (complete658_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I28 (complete658_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I29 (complete658_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I30 (complete658_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I31 (complete658_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I32 (complete658_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I33 (complete658_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I34 (complete658_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I35 (complete658_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I36 (complete658_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I37 (complete658_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I38 (complete658_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I39 (complete658_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I40 (complete658_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I41 (complete658_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I42 (complete658_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I43 (complete658_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I44 (complete658_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I45 (complete658_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I46 (complete658_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I47 (complete658_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I48 (complete658_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I49 (complete658_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I50 (complete658_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I51 (complete658_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I52 (complete658_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I53 (complete658_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I54 (complete658_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I55 (complete658_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I56 (complete658_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I57 (complete658_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I58 (complete658_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I59 (complete658_0n[33], ifint_0n[33], itint_0n[33]);
  INV I60 (gate657_0n, iaint_0n);
  C2RI I61 (itint_0n[0], i_0r1d[0], gate657_0n, initialise);
  C2RI I62 (itint_0n[1], i_0r1d[1], gate657_0n, initialise);
  C2RI I63 (itint_0n[2], i_0r1d[2], gate657_0n, initialise);
  C2RI I64 (itint_0n[3], i_0r1d[3], gate657_0n, initialise);
  C2RI I65 (itint_0n[4], i_0r1d[4], gate657_0n, initialise);
  C2RI I66 (itint_0n[5], i_0r1d[5], gate657_0n, initialise);
  C2RI I67 (itint_0n[6], i_0r1d[6], gate657_0n, initialise);
  C2RI I68 (itint_0n[7], i_0r1d[7], gate657_0n, initialise);
  C2RI I69 (itint_0n[8], i_0r1d[8], gate657_0n, initialise);
  C2RI I70 (itint_0n[9], i_0r1d[9], gate657_0n, initialise);
  C2RI I71 (itint_0n[10], i_0r1d[10], gate657_0n, initialise);
  C2RI I72 (itint_0n[11], i_0r1d[11], gate657_0n, initialise);
  C2RI I73 (itint_0n[12], i_0r1d[12], gate657_0n, initialise);
  C2RI I74 (itint_0n[13], i_0r1d[13], gate657_0n, initialise);
  C2RI I75 (itint_0n[14], i_0r1d[14], gate657_0n, initialise);
  C2RI I76 (itint_0n[15], i_0r1d[15], gate657_0n, initialise);
  C2RI I77 (itint_0n[16], i_0r1d[16], gate657_0n, initialise);
  C2RI I78 (itint_0n[17], i_0r1d[17], gate657_0n, initialise);
  C2RI I79 (itint_0n[18], i_0r1d[18], gate657_0n, initialise);
  C2RI I80 (itint_0n[19], i_0r1d[19], gate657_0n, initialise);
  C2RI I81 (itint_0n[20], i_0r1d[20], gate657_0n, initialise);
  C2RI I82 (itint_0n[21], i_0r1d[21], gate657_0n, initialise);
  C2RI I83 (itint_0n[22], i_0r1d[22], gate657_0n, initialise);
  C2RI I84 (itint_0n[23], i_0r1d[23], gate657_0n, initialise);
  C2RI I85 (itint_0n[24], i_0r1d[24], gate657_0n, initialise);
  C2RI I86 (itint_0n[25], i_0r1d[25], gate657_0n, initialise);
  C2RI I87 (itint_0n[26], i_0r1d[26], gate657_0n, initialise);
  C2RI I88 (itint_0n[27], i_0r1d[27], gate657_0n, initialise);
  C2RI I89 (itint_0n[28], i_0r1d[28], gate657_0n, initialise);
  C2RI I90 (itint_0n[29], i_0r1d[29], gate657_0n, initialise);
  C2RI I91 (itint_0n[30], i_0r1d[30], gate657_0n, initialise);
  C2RI I92 (itint_0n[31], i_0r1d[31], gate657_0n, initialise);
  C2RI I93 (itint_0n[32], i_0r1d[32], gate657_0n, initialise);
  C2RI I94 (itint_0n[33], i_0r1d[33], gate657_0n, initialise);
  C2RI I95 (ifint_0n[0], i_0r0d[0], gate657_0n, initialise);
  C2RI I96 (ifint_0n[1], i_0r0d[1], gate657_0n, initialise);
  C2RI I97 (ifint_0n[2], i_0r0d[2], gate657_0n, initialise);
  C2RI I98 (ifint_0n[3], i_0r0d[3], gate657_0n, initialise);
  C2RI I99 (ifint_0n[4], i_0r0d[4], gate657_0n, initialise);
  C2RI I100 (ifint_0n[5], i_0r0d[5], gate657_0n, initialise);
  C2RI I101 (ifint_0n[6], i_0r0d[6], gate657_0n, initialise);
  C2RI I102 (ifint_0n[7], i_0r0d[7], gate657_0n, initialise);
  C2RI I103 (ifint_0n[8], i_0r0d[8], gate657_0n, initialise);
  C2RI I104 (ifint_0n[9], i_0r0d[9], gate657_0n, initialise);
  C2RI I105 (ifint_0n[10], i_0r0d[10], gate657_0n, initialise);
  C2RI I106 (ifint_0n[11], i_0r0d[11], gate657_0n, initialise);
  C2RI I107 (ifint_0n[12], i_0r0d[12], gate657_0n, initialise);
  C2RI I108 (ifint_0n[13], i_0r0d[13], gate657_0n, initialise);
  C2RI I109 (ifint_0n[14], i_0r0d[14], gate657_0n, initialise);
  C2RI I110 (ifint_0n[15], i_0r0d[15], gate657_0n, initialise);
  C2RI I111 (ifint_0n[16], i_0r0d[16], gate657_0n, initialise);
  C2RI I112 (ifint_0n[17], i_0r0d[17], gate657_0n, initialise);
  C2RI I113 (ifint_0n[18], i_0r0d[18], gate657_0n, initialise);
  C2RI I114 (ifint_0n[19], i_0r0d[19], gate657_0n, initialise);
  C2RI I115 (ifint_0n[20], i_0r0d[20], gate657_0n, initialise);
  C2RI I116 (ifint_0n[21], i_0r0d[21], gate657_0n, initialise);
  C2RI I117 (ifint_0n[22], i_0r0d[22], gate657_0n, initialise);
  C2RI I118 (ifint_0n[23], i_0r0d[23], gate657_0n, initialise);
  C2RI I119 (ifint_0n[24], i_0r0d[24], gate657_0n, initialise);
  C2RI I120 (ifint_0n[25], i_0r0d[25], gate657_0n, initialise);
  C2RI I121 (ifint_0n[26], i_0r0d[26], gate657_0n, initialise);
  C2RI I122 (ifint_0n[27], i_0r0d[27], gate657_0n, initialise);
  C2RI I123 (ifint_0n[28], i_0r0d[28], gate657_0n, initialise);
  C2RI I124 (ifint_0n[29], i_0r0d[29], gate657_0n, initialise);
  C2RI I125 (ifint_0n[30], i_0r0d[30], gate657_0n, initialise);
  C2RI I126 (ifint_0n[31], i_0r0d[31], gate657_0n, initialise);
  C2RI I127 (ifint_0n[32], i_0r0d[32], gate657_0n, initialise);
  C2RI I128 (ifint_0n[33], i_0r0d[33], gate657_0n, initialise);
  C3 I129 (internal_0n[18], complete654_0n[0], complete654_0n[1], complete654_0n[2]);
  C3 I130 (internal_0n[19], complete654_0n[3], complete654_0n[4], complete654_0n[5]);
  C3 I131 (internal_0n[20], complete654_0n[6], complete654_0n[7], complete654_0n[8]);
  C3 I132 (internal_0n[21], complete654_0n[9], complete654_0n[10], complete654_0n[11]);
  C3 I133 (internal_0n[22], complete654_0n[12], complete654_0n[13], complete654_0n[14]);
  C3 I134 (internal_0n[23], complete654_0n[15], complete654_0n[16], complete654_0n[17]);
  C3 I135 (internal_0n[24], complete654_0n[18], complete654_0n[19], complete654_0n[20]);
  C3 I136 (internal_0n[25], complete654_0n[21], complete654_0n[22], complete654_0n[23]);
  C3 I137 (internal_0n[26], complete654_0n[24], complete654_0n[25], complete654_0n[26]);
  C3 I138 (internal_0n[27], complete654_0n[27], complete654_0n[28], complete654_0n[29]);
  C3 I139 (internal_0n[28], complete654_0n[30], complete654_0n[31], complete654_0n[32]);
  C2 I140 (internal_0n[29], complete654_0n[33], complete654_0n[34]);
  C3 I141 (internal_0n[30], internal_0n[18], internal_0n[19], internal_0n[20]);
  C3 I142 (internal_0n[31], internal_0n[21], internal_0n[22], internal_0n[23]);
  C3 I143 (internal_0n[32], internal_0n[24], internal_0n[25], internal_0n[26]);
  C3 I144 (internal_0n[33], internal_0n[27], internal_0n[28], internal_0n[29]);
  C2 I145 (internal_0n[34], internal_0n[30], internal_0n[31]);
  C2 I146 (internal_0n[35], internal_0n[32], internal_0n[33]);
  C2 I147 (oaint_0n, internal_0n[34], internal_0n[35]);
  OR2 I148 (complete654_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I149 (complete654_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I150 (complete654_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I151 (complete654_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I152 (complete654_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I153 (complete654_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I154 (complete654_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I155 (complete654_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I156 (complete654_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I157 (complete654_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I158 (complete654_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I159 (complete654_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I160 (complete654_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I161 (complete654_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I162 (complete654_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I163 (complete654_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I164 (complete654_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I165 (complete654_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I166 (complete654_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I167 (complete654_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I168 (complete654_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I169 (complete654_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I170 (complete654_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I171 (complete654_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I172 (complete654_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I173 (complete654_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I174 (complete654_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I175 (complete654_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I176 (complete654_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I177 (complete654_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I178 (complete654_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I179 (complete654_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I180 (complete654_0n[32], o_0r0d[32], o_0r1d[32]);
  OR2 I181 (complete654_0n[33], o_0r0d[33], o_0r1d[33]);
  OR2 I182 (complete654_0n[34], o_0r0d[34], o_0r1d[34]);
  INV I183 (gate653_0n, o_0a);
  C2RI I184 (o_0r1d[0], otint_0n[0], gate653_0n, initialise);
  C2RI I185 (o_0r1d[1], otint_0n[1], gate653_0n, initialise);
  C2RI I186 (o_0r1d[2], otint_0n[2], gate653_0n, initialise);
  C2RI I187 (o_0r1d[3], otint_0n[3], gate653_0n, initialise);
  C2RI I188 (o_0r1d[4], otint_0n[4], gate653_0n, initialise);
  C2RI I189 (o_0r1d[5], otint_0n[5], gate653_0n, initialise);
  C2RI I190 (o_0r1d[6], otint_0n[6], gate653_0n, initialise);
  C2RI I191 (o_0r1d[7], otint_0n[7], gate653_0n, initialise);
  C2RI I192 (o_0r1d[8], otint_0n[8], gate653_0n, initialise);
  C2RI I193 (o_0r1d[9], otint_0n[9], gate653_0n, initialise);
  C2RI I194 (o_0r1d[10], otint_0n[10], gate653_0n, initialise);
  C2RI I195 (o_0r1d[11], otint_0n[11], gate653_0n, initialise);
  C2RI I196 (o_0r1d[12], otint_0n[12], gate653_0n, initialise);
  C2RI I197 (o_0r1d[13], otint_0n[13], gate653_0n, initialise);
  C2RI I198 (o_0r1d[14], otint_0n[14], gate653_0n, initialise);
  C2RI I199 (o_0r1d[15], otint_0n[15], gate653_0n, initialise);
  C2RI I200 (o_0r1d[16], otint_0n[16], gate653_0n, initialise);
  C2RI I201 (o_0r1d[17], otint_0n[17], gate653_0n, initialise);
  C2RI I202 (o_0r1d[18], otint_0n[18], gate653_0n, initialise);
  C2RI I203 (o_0r1d[19], otint_0n[19], gate653_0n, initialise);
  C2RI I204 (o_0r1d[20], otint_0n[20], gate653_0n, initialise);
  C2RI I205 (o_0r1d[21], otint_0n[21], gate653_0n, initialise);
  C2RI I206 (o_0r1d[22], otint_0n[22], gate653_0n, initialise);
  C2RI I207 (o_0r1d[23], otint_0n[23], gate653_0n, initialise);
  C2RI I208 (o_0r1d[24], otint_0n[24], gate653_0n, initialise);
  C2RI I209 (o_0r1d[25], otint_0n[25], gate653_0n, initialise);
  C2RI I210 (o_0r1d[26], otint_0n[26], gate653_0n, initialise);
  C2RI I211 (o_0r1d[27], otint_0n[27], gate653_0n, initialise);
  C2RI I212 (o_0r1d[28], otint_0n[28], gate653_0n, initialise);
  C2RI I213 (o_0r1d[29], otint_0n[29], gate653_0n, initialise);
  C2RI I214 (o_0r1d[30], otint_0n[30], gate653_0n, initialise);
  C2RI I215 (o_0r1d[31], otint_0n[31], gate653_0n, initialise);
  C2RI I216 (o_0r1d[32], otint_0n[32], gate653_0n, initialise);
  C2RI I217 (o_0r1d[33], otint_0n[33], gate653_0n, initialise);
  C2RI I218 (o_0r1d[34], otint_0n[34], gate653_0n, initialise);
  C2RI I219 (o_0r0d[0], ofint_0n[0], gate653_0n, initialise);
  C2RI I220 (o_0r0d[1], ofint_0n[1], gate653_0n, initialise);
  C2RI I221 (o_0r0d[2], ofint_0n[2], gate653_0n, initialise);
  C2RI I222 (o_0r0d[3], ofint_0n[3], gate653_0n, initialise);
  C2RI I223 (o_0r0d[4], ofint_0n[4], gate653_0n, initialise);
  C2RI I224 (o_0r0d[5], ofint_0n[5], gate653_0n, initialise);
  C2RI I225 (o_0r0d[6], ofint_0n[6], gate653_0n, initialise);
  C2RI I226 (o_0r0d[7], ofint_0n[7], gate653_0n, initialise);
  C2RI I227 (o_0r0d[8], ofint_0n[8], gate653_0n, initialise);
  C2RI I228 (o_0r0d[9], ofint_0n[9], gate653_0n, initialise);
  C2RI I229 (o_0r0d[10], ofint_0n[10], gate653_0n, initialise);
  C2RI I230 (o_0r0d[11], ofint_0n[11], gate653_0n, initialise);
  C2RI I231 (o_0r0d[12], ofint_0n[12], gate653_0n, initialise);
  C2RI I232 (o_0r0d[13], ofint_0n[13], gate653_0n, initialise);
  C2RI I233 (o_0r0d[14], ofint_0n[14], gate653_0n, initialise);
  C2RI I234 (o_0r0d[15], ofint_0n[15], gate653_0n, initialise);
  C2RI I235 (o_0r0d[16], ofint_0n[16], gate653_0n, initialise);
  C2RI I236 (o_0r0d[17], ofint_0n[17], gate653_0n, initialise);
  C2RI I237 (o_0r0d[18], ofint_0n[18], gate653_0n, initialise);
  C2RI I238 (o_0r0d[19], ofint_0n[19], gate653_0n, initialise);
  C2RI I239 (o_0r0d[20], ofint_0n[20], gate653_0n, initialise);
  C2RI I240 (o_0r0d[21], ofint_0n[21], gate653_0n, initialise);
  C2RI I241 (o_0r0d[22], ofint_0n[22], gate653_0n, initialise);
  C2RI I242 (o_0r0d[23], ofint_0n[23], gate653_0n, initialise);
  C2RI I243 (o_0r0d[24], ofint_0n[24], gate653_0n, initialise);
  C2RI I244 (o_0r0d[25], ofint_0n[25], gate653_0n, initialise);
  C2RI I245 (o_0r0d[26], ofint_0n[26], gate653_0n, initialise);
  C2RI I246 (o_0r0d[27], ofint_0n[27], gate653_0n, initialise);
  C2RI I247 (o_0r0d[28], ofint_0n[28], gate653_0n, initialise);
  C2RI I248 (o_0r0d[29], ofint_0n[29], gate653_0n, initialise);
  C2RI I249 (o_0r0d[30], ofint_0n[30], gate653_0n, initialise);
  C2RI I250 (o_0r0d[31], ofint_0n[31], gate653_0n, initialise);
  C2RI I251 (o_0r0d[32], ofint_0n[32], gate653_0n, initialise);
  C2RI I252 (o_0r0d[33], ofint_0n[33], gate653_0n, initialise);
  C2RI I253 (o_0r0d[34], ofint_0n[34], gate653_0n, initialise);
  assign otint_0n[0] = itint_0n[0];
  assign otint_0n[1] = itint_0n[1];
  assign otint_0n[2] = itint_0n[2];
  assign otint_0n[3] = itint_0n[3];
  assign otint_0n[4] = itint_0n[4];
  assign otint_0n[5] = itint_0n[5];
  assign otint_0n[6] = itint_0n[6];
  assign otint_0n[7] = itint_0n[7];
  assign otint_0n[8] = itint_0n[8];
  assign otint_0n[9] = itint_0n[9];
  assign otint_0n[10] = itint_0n[10];
  assign otint_0n[11] = itint_0n[11];
  assign otint_0n[12] = itint_0n[12];
  assign otint_0n[13] = itint_0n[13];
  assign otint_0n[14] = itint_0n[14];
  assign otint_0n[15] = itint_0n[15];
  assign otint_0n[16] = itint_0n[16];
  assign otint_0n[17] = itint_0n[17];
  assign otint_0n[18] = itint_0n[18];
  assign otint_0n[19] = itint_0n[19];
  assign otint_0n[20] = itint_0n[20];
  assign otint_0n[21] = itint_0n[21];
  assign otint_0n[22] = itint_0n[22];
  assign otint_0n[23] = itint_0n[23];
  assign otint_0n[24] = itint_0n[24];
  assign otint_0n[25] = itint_0n[25];
  assign otint_0n[26] = itint_0n[26];
  assign otint_0n[27] = itint_0n[27];
  assign otint_0n[28] = itint_0n[28];
  assign otint_0n[29] = itint_0n[29];
  assign otint_0n[30] = itint_0n[30];
  assign otint_0n[31] = itint_0n[31];
  assign otint_0n[32] = itint_0n[32];
  assign otint_0n[33] = itint_0n[33];
  assign otint_0n[34] = itint_1n;
  assign ofint_0n[0] = ifint_0n[0];
  assign ofint_0n[1] = ifint_0n[1];
  assign ofint_0n[2] = ifint_0n[2];
  assign ofint_0n[3] = ifint_0n[3];
  assign ofint_0n[4] = ifint_0n[4];
  assign ofint_0n[5] = ifint_0n[5];
  assign ofint_0n[6] = ifint_0n[6];
  assign ofint_0n[7] = ifint_0n[7];
  assign ofint_0n[8] = ifint_0n[8];
  assign ofint_0n[9] = ifint_0n[9];
  assign ofint_0n[10] = ifint_0n[10];
  assign ofint_0n[11] = ifint_0n[11];
  assign ofint_0n[12] = ifint_0n[12];
  assign ofint_0n[13] = ifint_0n[13];
  assign ofint_0n[14] = ifint_0n[14];
  assign ofint_0n[15] = ifint_0n[15];
  assign ofint_0n[16] = ifint_0n[16];
  assign ofint_0n[17] = ifint_0n[17];
  assign ofint_0n[18] = ifint_0n[18];
  assign ofint_0n[19] = ifint_0n[19];
  assign ofint_0n[20] = ifint_0n[20];
  assign ofint_0n[21] = ifint_0n[21];
  assign ofint_0n[22] = ifint_0n[22];
  assign ofint_0n[23] = ifint_0n[23];
  assign ofint_0n[24] = ifint_0n[24];
  assign ofint_0n[25] = ifint_0n[25];
  assign ofint_0n[26] = ifint_0n[26];
  assign ofint_0n[27] = ifint_0n[27];
  assign ofint_0n[28] = ifint_0n[28];
  assign ofint_0n[29] = ifint_0n[29];
  assign ofint_0n[30] = ifint_0n[30];
  assign ofint_0n[31] = ifint_0n[31];
  assign ofint_0n[32] = ifint_0n[32];
  assign ofint_0n[33] = ifint_0n[33];
  assign ofint_0n[34] = ifint_1n;
endmodule

module BrzJ_l12__2835_200_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [34:0] i_0r0d;
  input [34:0] i_0r1d;
  output i_0a;
  input i_1r;
  output i_1a;
  output [34:0] o_0r0d;
  output [34:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [35:0] internal_0n;
  wire [34:0] ofint_0n;
  wire [34:0] otint_0n;
  wire oaint_0n;
  wire [34:0] ifint_0n;
  wire ifint_1n;
  wire [34:0] itint_0n;
  wire iaint_0n;
  wire iaint_1n;
  wire gate673_0n;
  wire [34:0] complete670_0n;
  wire gate669_0n;
  wire [34:0] complete666_0n;
  wire gate665_0n;
  wire [34:0] joint_0n;
  wire [34:0] joinf_0n;
  wire icomplete_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign i_1a = ifint_1n;
  INV I3 (gate673_0n, iaint_1n);
  C2RI I4 (ifint_1n, i_1r, gate673_0n, initialise);
  C3 I5 (internal_0n[0], complete670_0n[0], complete670_0n[1], complete670_0n[2]);
  C3 I6 (internal_0n[1], complete670_0n[3], complete670_0n[4], complete670_0n[5]);
  C3 I7 (internal_0n[2], complete670_0n[6], complete670_0n[7], complete670_0n[8]);
  C3 I8 (internal_0n[3], complete670_0n[9], complete670_0n[10], complete670_0n[11]);
  C3 I9 (internal_0n[4], complete670_0n[12], complete670_0n[13], complete670_0n[14]);
  C3 I10 (internal_0n[5], complete670_0n[15], complete670_0n[16], complete670_0n[17]);
  C3 I11 (internal_0n[6], complete670_0n[18], complete670_0n[19], complete670_0n[20]);
  C3 I12 (internal_0n[7], complete670_0n[21], complete670_0n[22], complete670_0n[23]);
  C3 I13 (internal_0n[8], complete670_0n[24], complete670_0n[25], complete670_0n[26]);
  C3 I14 (internal_0n[9], complete670_0n[27], complete670_0n[28], complete670_0n[29]);
  C3 I15 (internal_0n[10], complete670_0n[30], complete670_0n[31], complete670_0n[32]);
  C2 I16 (internal_0n[11], complete670_0n[33], complete670_0n[34]);
  C3 I17 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I18 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I19 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I20 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I21 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I22 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I23 (i_0a, internal_0n[16], internal_0n[17]);
  OR2 I24 (complete670_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I25 (complete670_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I26 (complete670_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I27 (complete670_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I28 (complete670_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I29 (complete670_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I30 (complete670_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I31 (complete670_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I32 (complete670_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I33 (complete670_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I34 (complete670_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I35 (complete670_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I36 (complete670_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I37 (complete670_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I38 (complete670_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I39 (complete670_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I40 (complete670_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I41 (complete670_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I42 (complete670_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I43 (complete670_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I44 (complete670_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I45 (complete670_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I46 (complete670_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I47 (complete670_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I48 (complete670_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I49 (complete670_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I50 (complete670_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I51 (complete670_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I52 (complete670_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I53 (complete670_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I54 (complete670_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I55 (complete670_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I56 (complete670_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I57 (complete670_0n[33], ifint_0n[33], itint_0n[33]);
  OR2 I58 (complete670_0n[34], ifint_0n[34], itint_0n[34]);
  INV I59 (gate669_0n, iaint_0n);
  C2RI I60 (itint_0n[0], i_0r1d[0], gate669_0n, initialise);
  C2RI I61 (itint_0n[1], i_0r1d[1], gate669_0n, initialise);
  C2RI I62 (itint_0n[2], i_0r1d[2], gate669_0n, initialise);
  C2RI I63 (itint_0n[3], i_0r1d[3], gate669_0n, initialise);
  C2RI I64 (itint_0n[4], i_0r1d[4], gate669_0n, initialise);
  C2RI I65 (itint_0n[5], i_0r1d[5], gate669_0n, initialise);
  C2RI I66 (itint_0n[6], i_0r1d[6], gate669_0n, initialise);
  C2RI I67 (itint_0n[7], i_0r1d[7], gate669_0n, initialise);
  C2RI I68 (itint_0n[8], i_0r1d[8], gate669_0n, initialise);
  C2RI I69 (itint_0n[9], i_0r1d[9], gate669_0n, initialise);
  C2RI I70 (itint_0n[10], i_0r1d[10], gate669_0n, initialise);
  C2RI I71 (itint_0n[11], i_0r1d[11], gate669_0n, initialise);
  C2RI I72 (itint_0n[12], i_0r1d[12], gate669_0n, initialise);
  C2RI I73 (itint_0n[13], i_0r1d[13], gate669_0n, initialise);
  C2RI I74 (itint_0n[14], i_0r1d[14], gate669_0n, initialise);
  C2RI I75 (itint_0n[15], i_0r1d[15], gate669_0n, initialise);
  C2RI I76 (itint_0n[16], i_0r1d[16], gate669_0n, initialise);
  C2RI I77 (itint_0n[17], i_0r1d[17], gate669_0n, initialise);
  C2RI I78 (itint_0n[18], i_0r1d[18], gate669_0n, initialise);
  C2RI I79 (itint_0n[19], i_0r1d[19], gate669_0n, initialise);
  C2RI I80 (itint_0n[20], i_0r1d[20], gate669_0n, initialise);
  C2RI I81 (itint_0n[21], i_0r1d[21], gate669_0n, initialise);
  C2RI I82 (itint_0n[22], i_0r1d[22], gate669_0n, initialise);
  C2RI I83 (itint_0n[23], i_0r1d[23], gate669_0n, initialise);
  C2RI I84 (itint_0n[24], i_0r1d[24], gate669_0n, initialise);
  C2RI I85 (itint_0n[25], i_0r1d[25], gate669_0n, initialise);
  C2RI I86 (itint_0n[26], i_0r1d[26], gate669_0n, initialise);
  C2RI I87 (itint_0n[27], i_0r1d[27], gate669_0n, initialise);
  C2RI I88 (itint_0n[28], i_0r1d[28], gate669_0n, initialise);
  C2RI I89 (itint_0n[29], i_0r1d[29], gate669_0n, initialise);
  C2RI I90 (itint_0n[30], i_0r1d[30], gate669_0n, initialise);
  C2RI I91 (itint_0n[31], i_0r1d[31], gate669_0n, initialise);
  C2RI I92 (itint_0n[32], i_0r1d[32], gate669_0n, initialise);
  C2RI I93 (itint_0n[33], i_0r1d[33], gate669_0n, initialise);
  C2RI I94 (itint_0n[34], i_0r1d[34], gate669_0n, initialise);
  C2RI I95 (ifint_0n[0], i_0r0d[0], gate669_0n, initialise);
  C2RI I96 (ifint_0n[1], i_0r0d[1], gate669_0n, initialise);
  C2RI I97 (ifint_0n[2], i_0r0d[2], gate669_0n, initialise);
  C2RI I98 (ifint_0n[3], i_0r0d[3], gate669_0n, initialise);
  C2RI I99 (ifint_0n[4], i_0r0d[4], gate669_0n, initialise);
  C2RI I100 (ifint_0n[5], i_0r0d[5], gate669_0n, initialise);
  C2RI I101 (ifint_0n[6], i_0r0d[6], gate669_0n, initialise);
  C2RI I102 (ifint_0n[7], i_0r0d[7], gate669_0n, initialise);
  C2RI I103 (ifint_0n[8], i_0r0d[8], gate669_0n, initialise);
  C2RI I104 (ifint_0n[9], i_0r0d[9], gate669_0n, initialise);
  C2RI I105 (ifint_0n[10], i_0r0d[10], gate669_0n, initialise);
  C2RI I106 (ifint_0n[11], i_0r0d[11], gate669_0n, initialise);
  C2RI I107 (ifint_0n[12], i_0r0d[12], gate669_0n, initialise);
  C2RI I108 (ifint_0n[13], i_0r0d[13], gate669_0n, initialise);
  C2RI I109 (ifint_0n[14], i_0r0d[14], gate669_0n, initialise);
  C2RI I110 (ifint_0n[15], i_0r0d[15], gate669_0n, initialise);
  C2RI I111 (ifint_0n[16], i_0r0d[16], gate669_0n, initialise);
  C2RI I112 (ifint_0n[17], i_0r0d[17], gate669_0n, initialise);
  C2RI I113 (ifint_0n[18], i_0r0d[18], gate669_0n, initialise);
  C2RI I114 (ifint_0n[19], i_0r0d[19], gate669_0n, initialise);
  C2RI I115 (ifint_0n[20], i_0r0d[20], gate669_0n, initialise);
  C2RI I116 (ifint_0n[21], i_0r0d[21], gate669_0n, initialise);
  C2RI I117 (ifint_0n[22], i_0r0d[22], gate669_0n, initialise);
  C2RI I118 (ifint_0n[23], i_0r0d[23], gate669_0n, initialise);
  C2RI I119 (ifint_0n[24], i_0r0d[24], gate669_0n, initialise);
  C2RI I120 (ifint_0n[25], i_0r0d[25], gate669_0n, initialise);
  C2RI I121 (ifint_0n[26], i_0r0d[26], gate669_0n, initialise);
  C2RI I122 (ifint_0n[27], i_0r0d[27], gate669_0n, initialise);
  C2RI I123 (ifint_0n[28], i_0r0d[28], gate669_0n, initialise);
  C2RI I124 (ifint_0n[29], i_0r0d[29], gate669_0n, initialise);
  C2RI I125 (ifint_0n[30], i_0r0d[30], gate669_0n, initialise);
  C2RI I126 (ifint_0n[31], i_0r0d[31], gate669_0n, initialise);
  C2RI I127 (ifint_0n[32], i_0r0d[32], gate669_0n, initialise);
  C2RI I128 (ifint_0n[33], i_0r0d[33], gate669_0n, initialise);
  C2RI I129 (ifint_0n[34], i_0r0d[34], gate669_0n, initialise);
  C3 I130 (internal_0n[18], complete666_0n[0], complete666_0n[1], complete666_0n[2]);
  C3 I131 (internal_0n[19], complete666_0n[3], complete666_0n[4], complete666_0n[5]);
  C3 I132 (internal_0n[20], complete666_0n[6], complete666_0n[7], complete666_0n[8]);
  C3 I133 (internal_0n[21], complete666_0n[9], complete666_0n[10], complete666_0n[11]);
  C3 I134 (internal_0n[22], complete666_0n[12], complete666_0n[13], complete666_0n[14]);
  C3 I135 (internal_0n[23], complete666_0n[15], complete666_0n[16], complete666_0n[17]);
  C3 I136 (internal_0n[24], complete666_0n[18], complete666_0n[19], complete666_0n[20]);
  C3 I137 (internal_0n[25], complete666_0n[21], complete666_0n[22], complete666_0n[23]);
  C3 I138 (internal_0n[26], complete666_0n[24], complete666_0n[25], complete666_0n[26]);
  C3 I139 (internal_0n[27], complete666_0n[27], complete666_0n[28], complete666_0n[29]);
  C3 I140 (internal_0n[28], complete666_0n[30], complete666_0n[31], complete666_0n[32]);
  C2 I141 (internal_0n[29], complete666_0n[33], complete666_0n[34]);
  C3 I142 (internal_0n[30], internal_0n[18], internal_0n[19], internal_0n[20]);
  C3 I143 (internal_0n[31], internal_0n[21], internal_0n[22], internal_0n[23]);
  C3 I144 (internal_0n[32], internal_0n[24], internal_0n[25], internal_0n[26]);
  C3 I145 (internal_0n[33], internal_0n[27], internal_0n[28], internal_0n[29]);
  C2 I146 (internal_0n[34], internal_0n[30], internal_0n[31]);
  C2 I147 (internal_0n[35], internal_0n[32], internal_0n[33]);
  C2 I148 (oaint_0n, internal_0n[34], internal_0n[35]);
  OR2 I149 (complete666_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I150 (complete666_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I151 (complete666_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I152 (complete666_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I153 (complete666_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I154 (complete666_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I155 (complete666_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I156 (complete666_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I157 (complete666_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I158 (complete666_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I159 (complete666_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I160 (complete666_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I161 (complete666_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I162 (complete666_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I163 (complete666_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I164 (complete666_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I165 (complete666_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I166 (complete666_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I167 (complete666_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I168 (complete666_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I169 (complete666_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I170 (complete666_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I171 (complete666_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I172 (complete666_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I173 (complete666_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I174 (complete666_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I175 (complete666_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I176 (complete666_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I177 (complete666_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I178 (complete666_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I179 (complete666_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I180 (complete666_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I181 (complete666_0n[32], o_0r0d[32], o_0r1d[32]);
  OR2 I182 (complete666_0n[33], o_0r0d[33], o_0r1d[33]);
  OR2 I183 (complete666_0n[34], o_0r0d[34], o_0r1d[34]);
  INV I184 (gate665_0n, o_0a);
  C2RI I185 (o_0r1d[0], otint_0n[0], gate665_0n, initialise);
  C2RI I186 (o_0r1d[1], otint_0n[1], gate665_0n, initialise);
  C2RI I187 (o_0r1d[2], otint_0n[2], gate665_0n, initialise);
  C2RI I188 (o_0r1d[3], otint_0n[3], gate665_0n, initialise);
  C2RI I189 (o_0r1d[4], otint_0n[4], gate665_0n, initialise);
  C2RI I190 (o_0r1d[5], otint_0n[5], gate665_0n, initialise);
  C2RI I191 (o_0r1d[6], otint_0n[6], gate665_0n, initialise);
  C2RI I192 (o_0r1d[7], otint_0n[7], gate665_0n, initialise);
  C2RI I193 (o_0r1d[8], otint_0n[8], gate665_0n, initialise);
  C2RI I194 (o_0r1d[9], otint_0n[9], gate665_0n, initialise);
  C2RI I195 (o_0r1d[10], otint_0n[10], gate665_0n, initialise);
  C2RI I196 (o_0r1d[11], otint_0n[11], gate665_0n, initialise);
  C2RI I197 (o_0r1d[12], otint_0n[12], gate665_0n, initialise);
  C2RI I198 (o_0r1d[13], otint_0n[13], gate665_0n, initialise);
  C2RI I199 (o_0r1d[14], otint_0n[14], gate665_0n, initialise);
  C2RI I200 (o_0r1d[15], otint_0n[15], gate665_0n, initialise);
  C2RI I201 (o_0r1d[16], otint_0n[16], gate665_0n, initialise);
  C2RI I202 (o_0r1d[17], otint_0n[17], gate665_0n, initialise);
  C2RI I203 (o_0r1d[18], otint_0n[18], gate665_0n, initialise);
  C2RI I204 (o_0r1d[19], otint_0n[19], gate665_0n, initialise);
  C2RI I205 (o_0r1d[20], otint_0n[20], gate665_0n, initialise);
  C2RI I206 (o_0r1d[21], otint_0n[21], gate665_0n, initialise);
  C2RI I207 (o_0r1d[22], otint_0n[22], gate665_0n, initialise);
  C2RI I208 (o_0r1d[23], otint_0n[23], gate665_0n, initialise);
  C2RI I209 (o_0r1d[24], otint_0n[24], gate665_0n, initialise);
  C2RI I210 (o_0r1d[25], otint_0n[25], gate665_0n, initialise);
  C2RI I211 (o_0r1d[26], otint_0n[26], gate665_0n, initialise);
  C2RI I212 (o_0r1d[27], otint_0n[27], gate665_0n, initialise);
  C2RI I213 (o_0r1d[28], otint_0n[28], gate665_0n, initialise);
  C2RI I214 (o_0r1d[29], otint_0n[29], gate665_0n, initialise);
  C2RI I215 (o_0r1d[30], otint_0n[30], gate665_0n, initialise);
  C2RI I216 (o_0r1d[31], otint_0n[31], gate665_0n, initialise);
  C2RI I217 (o_0r1d[32], otint_0n[32], gate665_0n, initialise);
  C2RI I218 (o_0r1d[33], otint_0n[33], gate665_0n, initialise);
  C2RI I219 (o_0r1d[34], otint_0n[34], gate665_0n, initialise);
  C2RI I220 (o_0r0d[0], ofint_0n[0], gate665_0n, initialise);
  C2RI I221 (o_0r0d[1], ofint_0n[1], gate665_0n, initialise);
  C2RI I222 (o_0r0d[2], ofint_0n[2], gate665_0n, initialise);
  C2RI I223 (o_0r0d[3], ofint_0n[3], gate665_0n, initialise);
  C2RI I224 (o_0r0d[4], ofint_0n[4], gate665_0n, initialise);
  C2RI I225 (o_0r0d[5], ofint_0n[5], gate665_0n, initialise);
  C2RI I226 (o_0r0d[6], ofint_0n[6], gate665_0n, initialise);
  C2RI I227 (o_0r0d[7], ofint_0n[7], gate665_0n, initialise);
  C2RI I228 (o_0r0d[8], ofint_0n[8], gate665_0n, initialise);
  C2RI I229 (o_0r0d[9], ofint_0n[9], gate665_0n, initialise);
  C2RI I230 (o_0r0d[10], ofint_0n[10], gate665_0n, initialise);
  C2RI I231 (o_0r0d[11], ofint_0n[11], gate665_0n, initialise);
  C2RI I232 (o_0r0d[12], ofint_0n[12], gate665_0n, initialise);
  C2RI I233 (o_0r0d[13], ofint_0n[13], gate665_0n, initialise);
  C2RI I234 (o_0r0d[14], ofint_0n[14], gate665_0n, initialise);
  C2RI I235 (o_0r0d[15], ofint_0n[15], gate665_0n, initialise);
  C2RI I236 (o_0r0d[16], ofint_0n[16], gate665_0n, initialise);
  C2RI I237 (o_0r0d[17], ofint_0n[17], gate665_0n, initialise);
  C2RI I238 (o_0r0d[18], ofint_0n[18], gate665_0n, initialise);
  C2RI I239 (o_0r0d[19], ofint_0n[19], gate665_0n, initialise);
  C2RI I240 (o_0r0d[20], ofint_0n[20], gate665_0n, initialise);
  C2RI I241 (o_0r0d[21], ofint_0n[21], gate665_0n, initialise);
  C2RI I242 (o_0r0d[22], ofint_0n[22], gate665_0n, initialise);
  C2RI I243 (o_0r0d[23], ofint_0n[23], gate665_0n, initialise);
  C2RI I244 (o_0r0d[24], ofint_0n[24], gate665_0n, initialise);
  C2RI I245 (o_0r0d[25], ofint_0n[25], gate665_0n, initialise);
  C2RI I246 (o_0r0d[26], ofint_0n[26], gate665_0n, initialise);
  C2RI I247 (o_0r0d[27], ofint_0n[27], gate665_0n, initialise);
  C2RI I248 (o_0r0d[28], ofint_0n[28], gate665_0n, initialise);
  C2RI I249 (o_0r0d[29], ofint_0n[29], gate665_0n, initialise);
  C2RI I250 (o_0r0d[30], ofint_0n[30], gate665_0n, initialise);
  C2RI I251 (o_0r0d[31], ofint_0n[31], gate665_0n, initialise);
  C2RI I252 (o_0r0d[32], ofint_0n[32], gate665_0n, initialise);
  C2RI I253 (o_0r0d[33], ofint_0n[33], gate665_0n, initialise);
  C2RI I254 (o_0r0d[34], ofint_0n[34], gate665_0n, initialise);
  assign otint_0n[1] = joint_0n[1];
  assign otint_0n[2] = joint_0n[2];
  assign otint_0n[3] = joint_0n[3];
  assign otint_0n[4] = joint_0n[4];
  assign otint_0n[5] = joint_0n[5];
  assign otint_0n[6] = joint_0n[6];
  assign otint_0n[7] = joint_0n[7];
  assign otint_0n[8] = joint_0n[8];
  assign otint_0n[9] = joint_0n[9];
  assign otint_0n[10] = joint_0n[10];
  assign otint_0n[11] = joint_0n[11];
  assign otint_0n[12] = joint_0n[12];
  assign otint_0n[13] = joint_0n[13];
  assign otint_0n[14] = joint_0n[14];
  assign otint_0n[15] = joint_0n[15];
  assign otint_0n[16] = joint_0n[16];
  assign otint_0n[17] = joint_0n[17];
  assign otint_0n[18] = joint_0n[18];
  assign otint_0n[19] = joint_0n[19];
  assign otint_0n[20] = joint_0n[20];
  assign otint_0n[21] = joint_0n[21];
  assign otint_0n[22] = joint_0n[22];
  assign otint_0n[23] = joint_0n[23];
  assign otint_0n[24] = joint_0n[24];
  assign otint_0n[25] = joint_0n[25];
  assign otint_0n[26] = joint_0n[26];
  assign otint_0n[27] = joint_0n[27];
  assign otint_0n[28] = joint_0n[28];
  assign otint_0n[29] = joint_0n[29];
  assign otint_0n[30] = joint_0n[30];
  assign otint_0n[31] = joint_0n[31];
  assign otint_0n[32] = joint_0n[32];
  assign otint_0n[33] = joint_0n[33];
  assign otint_0n[34] = joint_0n[34];
  assign ofint_0n[1] = joinf_0n[1];
  assign ofint_0n[2] = joinf_0n[2];
  assign ofint_0n[3] = joinf_0n[3];
  assign ofint_0n[4] = joinf_0n[4];
  assign ofint_0n[5] = joinf_0n[5];
  assign ofint_0n[6] = joinf_0n[6];
  assign ofint_0n[7] = joinf_0n[7];
  assign ofint_0n[8] = joinf_0n[8];
  assign ofint_0n[9] = joinf_0n[9];
  assign ofint_0n[10] = joinf_0n[10];
  assign ofint_0n[11] = joinf_0n[11];
  assign ofint_0n[12] = joinf_0n[12];
  assign ofint_0n[13] = joinf_0n[13];
  assign ofint_0n[14] = joinf_0n[14];
  assign ofint_0n[15] = joinf_0n[15];
  assign ofint_0n[16] = joinf_0n[16];
  assign ofint_0n[17] = joinf_0n[17];
  assign ofint_0n[18] = joinf_0n[18];
  assign ofint_0n[19] = joinf_0n[19];
  assign ofint_0n[20] = joinf_0n[20];
  assign ofint_0n[21] = joinf_0n[21];
  assign ofint_0n[22] = joinf_0n[22];
  assign ofint_0n[23] = joinf_0n[23];
  assign ofint_0n[24] = joinf_0n[24];
  assign ofint_0n[25] = joinf_0n[25];
  assign ofint_0n[26] = joinf_0n[26];
  assign ofint_0n[27] = joinf_0n[27];
  assign ofint_0n[28] = joinf_0n[28];
  assign ofint_0n[29] = joinf_0n[29];
  assign ofint_0n[30] = joinf_0n[30];
  assign ofint_0n[31] = joinf_0n[31];
  assign ofint_0n[32] = joinf_0n[32];
  assign ofint_0n[33] = joinf_0n[33];
  assign ofint_0n[34] = joinf_0n[34];
  C2 I323 (otint_0n[0], joint_0n[0], icomplete_0n);
  C2 I324 (ofint_0n[0], joinf_0n[0], icomplete_0n);
  assign icomplete_0n = ifint_1n;
  assign joint_0n[0] = itint_0n[0];
  assign joint_0n[1] = itint_0n[1];
  assign joint_0n[2] = itint_0n[2];
  assign joint_0n[3] = itint_0n[3];
  assign joint_0n[4] = itint_0n[4];
  assign joint_0n[5] = itint_0n[5];
  assign joint_0n[6] = itint_0n[6];
  assign joint_0n[7] = itint_0n[7];
  assign joint_0n[8] = itint_0n[8];
  assign joint_0n[9] = itint_0n[9];
  assign joint_0n[10] = itint_0n[10];
  assign joint_0n[11] = itint_0n[11];
  assign joint_0n[12] = itint_0n[12];
  assign joint_0n[13] = itint_0n[13];
  assign joint_0n[14] = itint_0n[14];
  assign joint_0n[15] = itint_0n[15];
  assign joint_0n[16] = itint_0n[16];
  assign joint_0n[17] = itint_0n[17];
  assign joint_0n[18] = itint_0n[18];
  assign joint_0n[19] = itint_0n[19];
  assign joint_0n[20] = itint_0n[20];
  assign joint_0n[21] = itint_0n[21];
  assign joint_0n[22] = itint_0n[22];
  assign joint_0n[23] = itint_0n[23];
  assign joint_0n[24] = itint_0n[24];
  assign joint_0n[25] = itint_0n[25];
  assign joint_0n[26] = itint_0n[26];
  assign joint_0n[27] = itint_0n[27];
  assign joint_0n[28] = itint_0n[28];
  assign joint_0n[29] = itint_0n[29];
  assign joint_0n[30] = itint_0n[30];
  assign joint_0n[31] = itint_0n[31];
  assign joint_0n[32] = itint_0n[32];
  assign joint_0n[33] = itint_0n[33];
  assign joint_0n[34] = itint_0n[34];
  assign joinf_0n[0] = ifint_0n[0];
  assign joinf_0n[1] = ifint_0n[1];
  assign joinf_0n[2] = ifint_0n[2];
  assign joinf_0n[3] = ifint_0n[3];
  assign joinf_0n[4] = ifint_0n[4];
  assign joinf_0n[5] = ifint_0n[5];
  assign joinf_0n[6] = ifint_0n[6];
  assign joinf_0n[7] = ifint_0n[7];
  assign joinf_0n[8] = ifint_0n[8];
  assign joinf_0n[9] = ifint_0n[9];
  assign joinf_0n[10] = ifint_0n[10];
  assign joinf_0n[11] = ifint_0n[11];
  assign joinf_0n[12] = ifint_0n[12];
  assign joinf_0n[13] = ifint_0n[13];
  assign joinf_0n[14] = ifint_0n[14];
  assign joinf_0n[15] = ifint_0n[15];
  assign joinf_0n[16] = ifint_0n[16];
  assign joinf_0n[17] = ifint_0n[17];
  assign joinf_0n[18] = ifint_0n[18];
  assign joinf_0n[19] = ifint_0n[19];
  assign joinf_0n[20] = ifint_0n[20];
  assign joinf_0n[21] = ifint_0n[21];
  assign joinf_0n[22] = ifint_0n[22];
  assign joinf_0n[23] = ifint_0n[23];
  assign joinf_0n[24] = ifint_0n[24];
  assign joinf_0n[25] = ifint_0n[25];
  assign joinf_0n[26] = ifint_0n[26];
  assign joinf_0n[27] = ifint_0n[27];
  assign joinf_0n[28] = ifint_0n[28];
  assign joinf_0n[29] = ifint_0n[29];
  assign joinf_0n[30] = ifint_0n[30];
  assign joinf_0n[31] = ifint_0n[31];
  assign joinf_0n[32] = ifint_0n[32];
  assign joinf_0n[33] = ifint_0n[33];
  assign joinf_0n[34] = ifint_0n[34];
endmodule

module BrzJ_l13__2835_2035_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [34:0] i_0r0d;
  input [34:0] i_0r1d;
  output i_0a;
  input [34:0] i_1r0d;
  input [34:0] i_1r1d;
  output i_1a;
  output [69:0] o_0r0d;
  output [69:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [70:0] internal_0n;
  wire [69:0] ofint_0n;
  wire [69:0] otint_0n;
  wire oaint_0n;
  wire [34:0] ifint_0n;
  wire [34:0] ifint_1n;
  wire [34:0] itint_0n;
  wire [34:0] itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [34:0] complete685_0n;
  wire gate684_0n;
  wire [34:0] complete681_0n;
  wire gate680_0n;
  wire [69:0] complete677_0n;
  wire gate676_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  C3 I2 (internal_0n[0], complete685_0n[0], complete685_0n[1], complete685_0n[2]);
  C3 I3 (internal_0n[1], complete685_0n[3], complete685_0n[4], complete685_0n[5]);
  C3 I4 (internal_0n[2], complete685_0n[6], complete685_0n[7], complete685_0n[8]);
  C3 I5 (internal_0n[3], complete685_0n[9], complete685_0n[10], complete685_0n[11]);
  C3 I6 (internal_0n[4], complete685_0n[12], complete685_0n[13], complete685_0n[14]);
  C3 I7 (internal_0n[5], complete685_0n[15], complete685_0n[16], complete685_0n[17]);
  C3 I8 (internal_0n[6], complete685_0n[18], complete685_0n[19], complete685_0n[20]);
  C3 I9 (internal_0n[7], complete685_0n[21], complete685_0n[22], complete685_0n[23]);
  C3 I10 (internal_0n[8], complete685_0n[24], complete685_0n[25], complete685_0n[26]);
  C3 I11 (internal_0n[9], complete685_0n[27], complete685_0n[28], complete685_0n[29]);
  C3 I12 (internal_0n[10], complete685_0n[30], complete685_0n[31], complete685_0n[32]);
  C2 I13 (internal_0n[11], complete685_0n[33], complete685_0n[34]);
  C3 I14 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I15 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I16 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I17 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I18 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I19 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I20 (i_1a, internal_0n[16], internal_0n[17]);
  OR2 I21 (complete685_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I22 (complete685_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I23 (complete685_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I24 (complete685_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I25 (complete685_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I26 (complete685_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I27 (complete685_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I28 (complete685_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I29 (complete685_0n[8], ifint_1n[8], itint_1n[8]);
  OR2 I30 (complete685_0n[9], ifint_1n[9], itint_1n[9]);
  OR2 I31 (complete685_0n[10], ifint_1n[10], itint_1n[10]);
  OR2 I32 (complete685_0n[11], ifint_1n[11], itint_1n[11]);
  OR2 I33 (complete685_0n[12], ifint_1n[12], itint_1n[12]);
  OR2 I34 (complete685_0n[13], ifint_1n[13], itint_1n[13]);
  OR2 I35 (complete685_0n[14], ifint_1n[14], itint_1n[14]);
  OR2 I36 (complete685_0n[15], ifint_1n[15], itint_1n[15]);
  OR2 I37 (complete685_0n[16], ifint_1n[16], itint_1n[16]);
  OR2 I38 (complete685_0n[17], ifint_1n[17], itint_1n[17]);
  OR2 I39 (complete685_0n[18], ifint_1n[18], itint_1n[18]);
  OR2 I40 (complete685_0n[19], ifint_1n[19], itint_1n[19]);
  OR2 I41 (complete685_0n[20], ifint_1n[20], itint_1n[20]);
  OR2 I42 (complete685_0n[21], ifint_1n[21], itint_1n[21]);
  OR2 I43 (complete685_0n[22], ifint_1n[22], itint_1n[22]);
  OR2 I44 (complete685_0n[23], ifint_1n[23], itint_1n[23]);
  OR2 I45 (complete685_0n[24], ifint_1n[24], itint_1n[24]);
  OR2 I46 (complete685_0n[25], ifint_1n[25], itint_1n[25]);
  OR2 I47 (complete685_0n[26], ifint_1n[26], itint_1n[26]);
  OR2 I48 (complete685_0n[27], ifint_1n[27], itint_1n[27]);
  OR2 I49 (complete685_0n[28], ifint_1n[28], itint_1n[28]);
  OR2 I50 (complete685_0n[29], ifint_1n[29], itint_1n[29]);
  OR2 I51 (complete685_0n[30], ifint_1n[30], itint_1n[30]);
  OR2 I52 (complete685_0n[31], ifint_1n[31], itint_1n[31]);
  OR2 I53 (complete685_0n[32], ifint_1n[32], itint_1n[32]);
  OR2 I54 (complete685_0n[33], ifint_1n[33], itint_1n[33]);
  OR2 I55 (complete685_0n[34], ifint_1n[34], itint_1n[34]);
  INV I56 (gate684_0n, iaint_1n);
  C2RI I57 (itint_1n[0], i_1r1d[0], gate684_0n, initialise);
  C2RI I58 (itint_1n[1], i_1r1d[1], gate684_0n, initialise);
  C2RI I59 (itint_1n[2], i_1r1d[2], gate684_0n, initialise);
  C2RI I60 (itint_1n[3], i_1r1d[3], gate684_0n, initialise);
  C2RI I61 (itint_1n[4], i_1r1d[4], gate684_0n, initialise);
  C2RI I62 (itint_1n[5], i_1r1d[5], gate684_0n, initialise);
  C2RI I63 (itint_1n[6], i_1r1d[6], gate684_0n, initialise);
  C2RI I64 (itint_1n[7], i_1r1d[7], gate684_0n, initialise);
  C2RI I65 (itint_1n[8], i_1r1d[8], gate684_0n, initialise);
  C2RI I66 (itint_1n[9], i_1r1d[9], gate684_0n, initialise);
  C2RI I67 (itint_1n[10], i_1r1d[10], gate684_0n, initialise);
  C2RI I68 (itint_1n[11], i_1r1d[11], gate684_0n, initialise);
  C2RI I69 (itint_1n[12], i_1r1d[12], gate684_0n, initialise);
  C2RI I70 (itint_1n[13], i_1r1d[13], gate684_0n, initialise);
  C2RI I71 (itint_1n[14], i_1r1d[14], gate684_0n, initialise);
  C2RI I72 (itint_1n[15], i_1r1d[15], gate684_0n, initialise);
  C2RI I73 (itint_1n[16], i_1r1d[16], gate684_0n, initialise);
  C2RI I74 (itint_1n[17], i_1r1d[17], gate684_0n, initialise);
  C2RI I75 (itint_1n[18], i_1r1d[18], gate684_0n, initialise);
  C2RI I76 (itint_1n[19], i_1r1d[19], gate684_0n, initialise);
  C2RI I77 (itint_1n[20], i_1r1d[20], gate684_0n, initialise);
  C2RI I78 (itint_1n[21], i_1r1d[21], gate684_0n, initialise);
  C2RI I79 (itint_1n[22], i_1r1d[22], gate684_0n, initialise);
  C2RI I80 (itint_1n[23], i_1r1d[23], gate684_0n, initialise);
  C2RI I81 (itint_1n[24], i_1r1d[24], gate684_0n, initialise);
  C2RI I82 (itint_1n[25], i_1r1d[25], gate684_0n, initialise);
  C2RI I83 (itint_1n[26], i_1r1d[26], gate684_0n, initialise);
  C2RI I84 (itint_1n[27], i_1r1d[27], gate684_0n, initialise);
  C2RI I85 (itint_1n[28], i_1r1d[28], gate684_0n, initialise);
  C2RI I86 (itint_1n[29], i_1r1d[29], gate684_0n, initialise);
  C2RI I87 (itint_1n[30], i_1r1d[30], gate684_0n, initialise);
  C2RI I88 (itint_1n[31], i_1r1d[31], gate684_0n, initialise);
  C2RI I89 (itint_1n[32], i_1r1d[32], gate684_0n, initialise);
  C2RI I90 (itint_1n[33], i_1r1d[33], gate684_0n, initialise);
  C2RI I91 (itint_1n[34], i_1r1d[34], gate684_0n, initialise);
  C2RI I92 (ifint_1n[0], i_1r0d[0], gate684_0n, initialise);
  C2RI I93 (ifint_1n[1], i_1r0d[1], gate684_0n, initialise);
  C2RI I94 (ifint_1n[2], i_1r0d[2], gate684_0n, initialise);
  C2RI I95 (ifint_1n[3], i_1r0d[3], gate684_0n, initialise);
  C2RI I96 (ifint_1n[4], i_1r0d[4], gate684_0n, initialise);
  C2RI I97 (ifint_1n[5], i_1r0d[5], gate684_0n, initialise);
  C2RI I98 (ifint_1n[6], i_1r0d[6], gate684_0n, initialise);
  C2RI I99 (ifint_1n[7], i_1r0d[7], gate684_0n, initialise);
  C2RI I100 (ifint_1n[8], i_1r0d[8], gate684_0n, initialise);
  C2RI I101 (ifint_1n[9], i_1r0d[9], gate684_0n, initialise);
  C2RI I102 (ifint_1n[10], i_1r0d[10], gate684_0n, initialise);
  C2RI I103 (ifint_1n[11], i_1r0d[11], gate684_0n, initialise);
  C2RI I104 (ifint_1n[12], i_1r0d[12], gate684_0n, initialise);
  C2RI I105 (ifint_1n[13], i_1r0d[13], gate684_0n, initialise);
  C2RI I106 (ifint_1n[14], i_1r0d[14], gate684_0n, initialise);
  C2RI I107 (ifint_1n[15], i_1r0d[15], gate684_0n, initialise);
  C2RI I108 (ifint_1n[16], i_1r0d[16], gate684_0n, initialise);
  C2RI I109 (ifint_1n[17], i_1r0d[17], gate684_0n, initialise);
  C2RI I110 (ifint_1n[18], i_1r0d[18], gate684_0n, initialise);
  C2RI I111 (ifint_1n[19], i_1r0d[19], gate684_0n, initialise);
  C2RI I112 (ifint_1n[20], i_1r0d[20], gate684_0n, initialise);
  C2RI I113 (ifint_1n[21], i_1r0d[21], gate684_0n, initialise);
  C2RI I114 (ifint_1n[22], i_1r0d[22], gate684_0n, initialise);
  C2RI I115 (ifint_1n[23], i_1r0d[23], gate684_0n, initialise);
  C2RI I116 (ifint_1n[24], i_1r0d[24], gate684_0n, initialise);
  C2RI I117 (ifint_1n[25], i_1r0d[25], gate684_0n, initialise);
  C2RI I118 (ifint_1n[26], i_1r0d[26], gate684_0n, initialise);
  C2RI I119 (ifint_1n[27], i_1r0d[27], gate684_0n, initialise);
  C2RI I120 (ifint_1n[28], i_1r0d[28], gate684_0n, initialise);
  C2RI I121 (ifint_1n[29], i_1r0d[29], gate684_0n, initialise);
  C2RI I122 (ifint_1n[30], i_1r0d[30], gate684_0n, initialise);
  C2RI I123 (ifint_1n[31], i_1r0d[31], gate684_0n, initialise);
  C2RI I124 (ifint_1n[32], i_1r0d[32], gate684_0n, initialise);
  C2RI I125 (ifint_1n[33], i_1r0d[33], gate684_0n, initialise);
  C2RI I126 (ifint_1n[34], i_1r0d[34], gate684_0n, initialise);
  C3 I127 (internal_0n[18], complete681_0n[0], complete681_0n[1], complete681_0n[2]);
  C3 I128 (internal_0n[19], complete681_0n[3], complete681_0n[4], complete681_0n[5]);
  C3 I129 (internal_0n[20], complete681_0n[6], complete681_0n[7], complete681_0n[8]);
  C3 I130 (internal_0n[21], complete681_0n[9], complete681_0n[10], complete681_0n[11]);
  C3 I131 (internal_0n[22], complete681_0n[12], complete681_0n[13], complete681_0n[14]);
  C3 I132 (internal_0n[23], complete681_0n[15], complete681_0n[16], complete681_0n[17]);
  C3 I133 (internal_0n[24], complete681_0n[18], complete681_0n[19], complete681_0n[20]);
  C3 I134 (internal_0n[25], complete681_0n[21], complete681_0n[22], complete681_0n[23]);
  C3 I135 (internal_0n[26], complete681_0n[24], complete681_0n[25], complete681_0n[26]);
  C3 I136 (internal_0n[27], complete681_0n[27], complete681_0n[28], complete681_0n[29]);
  C3 I137 (internal_0n[28], complete681_0n[30], complete681_0n[31], complete681_0n[32]);
  C2 I138 (internal_0n[29], complete681_0n[33], complete681_0n[34]);
  C3 I139 (internal_0n[30], internal_0n[18], internal_0n[19], internal_0n[20]);
  C3 I140 (internal_0n[31], internal_0n[21], internal_0n[22], internal_0n[23]);
  C3 I141 (internal_0n[32], internal_0n[24], internal_0n[25], internal_0n[26]);
  C3 I142 (internal_0n[33], internal_0n[27], internal_0n[28], internal_0n[29]);
  C2 I143 (internal_0n[34], internal_0n[30], internal_0n[31]);
  C2 I144 (internal_0n[35], internal_0n[32], internal_0n[33]);
  C2 I145 (i_0a, internal_0n[34], internal_0n[35]);
  OR2 I146 (complete681_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I147 (complete681_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I148 (complete681_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I149 (complete681_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I150 (complete681_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I151 (complete681_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I152 (complete681_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I153 (complete681_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I154 (complete681_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I155 (complete681_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I156 (complete681_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I157 (complete681_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I158 (complete681_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I159 (complete681_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I160 (complete681_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I161 (complete681_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I162 (complete681_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I163 (complete681_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I164 (complete681_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I165 (complete681_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I166 (complete681_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I167 (complete681_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I168 (complete681_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I169 (complete681_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I170 (complete681_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I171 (complete681_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I172 (complete681_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I173 (complete681_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I174 (complete681_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I175 (complete681_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I176 (complete681_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I177 (complete681_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I178 (complete681_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I179 (complete681_0n[33], ifint_0n[33], itint_0n[33]);
  OR2 I180 (complete681_0n[34], ifint_0n[34], itint_0n[34]);
  INV I181 (gate680_0n, iaint_0n);
  C2RI I182 (itint_0n[0], i_0r1d[0], gate680_0n, initialise);
  C2RI I183 (itint_0n[1], i_0r1d[1], gate680_0n, initialise);
  C2RI I184 (itint_0n[2], i_0r1d[2], gate680_0n, initialise);
  C2RI I185 (itint_0n[3], i_0r1d[3], gate680_0n, initialise);
  C2RI I186 (itint_0n[4], i_0r1d[4], gate680_0n, initialise);
  C2RI I187 (itint_0n[5], i_0r1d[5], gate680_0n, initialise);
  C2RI I188 (itint_0n[6], i_0r1d[6], gate680_0n, initialise);
  C2RI I189 (itint_0n[7], i_0r1d[7], gate680_0n, initialise);
  C2RI I190 (itint_0n[8], i_0r1d[8], gate680_0n, initialise);
  C2RI I191 (itint_0n[9], i_0r1d[9], gate680_0n, initialise);
  C2RI I192 (itint_0n[10], i_0r1d[10], gate680_0n, initialise);
  C2RI I193 (itint_0n[11], i_0r1d[11], gate680_0n, initialise);
  C2RI I194 (itint_0n[12], i_0r1d[12], gate680_0n, initialise);
  C2RI I195 (itint_0n[13], i_0r1d[13], gate680_0n, initialise);
  C2RI I196 (itint_0n[14], i_0r1d[14], gate680_0n, initialise);
  C2RI I197 (itint_0n[15], i_0r1d[15], gate680_0n, initialise);
  C2RI I198 (itint_0n[16], i_0r1d[16], gate680_0n, initialise);
  C2RI I199 (itint_0n[17], i_0r1d[17], gate680_0n, initialise);
  C2RI I200 (itint_0n[18], i_0r1d[18], gate680_0n, initialise);
  C2RI I201 (itint_0n[19], i_0r1d[19], gate680_0n, initialise);
  C2RI I202 (itint_0n[20], i_0r1d[20], gate680_0n, initialise);
  C2RI I203 (itint_0n[21], i_0r1d[21], gate680_0n, initialise);
  C2RI I204 (itint_0n[22], i_0r1d[22], gate680_0n, initialise);
  C2RI I205 (itint_0n[23], i_0r1d[23], gate680_0n, initialise);
  C2RI I206 (itint_0n[24], i_0r1d[24], gate680_0n, initialise);
  C2RI I207 (itint_0n[25], i_0r1d[25], gate680_0n, initialise);
  C2RI I208 (itint_0n[26], i_0r1d[26], gate680_0n, initialise);
  C2RI I209 (itint_0n[27], i_0r1d[27], gate680_0n, initialise);
  C2RI I210 (itint_0n[28], i_0r1d[28], gate680_0n, initialise);
  C2RI I211 (itint_0n[29], i_0r1d[29], gate680_0n, initialise);
  C2RI I212 (itint_0n[30], i_0r1d[30], gate680_0n, initialise);
  C2RI I213 (itint_0n[31], i_0r1d[31], gate680_0n, initialise);
  C2RI I214 (itint_0n[32], i_0r1d[32], gate680_0n, initialise);
  C2RI I215 (itint_0n[33], i_0r1d[33], gate680_0n, initialise);
  C2RI I216 (itint_0n[34], i_0r1d[34], gate680_0n, initialise);
  C2RI I217 (ifint_0n[0], i_0r0d[0], gate680_0n, initialise);
  C2RI I218 (ifint_0n[1], i_0r0d[1], gate680_0n, initialise);
  C2RI I219 (ifint_0n[2], i_0r0d[2], gate680_0n, initialise);
  C2RI I220 (ifint_0n[3], i_0r0d[3], gate680_0n, initialise);
  C2RI I221 (ifint_0n[4], i_0r0d[4], gate680_0n, initialise);
  C2RI I222 (ifint_0n[5], i_0r0d[5], gate680_0n, initialise);
  C2RI I223 (ifint_0n[6], i_0r0d[6], gate680_0n, initialise);
  C2RI I224 (ifint_0n[7], i_0r0d[7], gate680_0n, initialise);
  C2RI I225 (ifint_0n[8], i_0r0d[8], gate680_0n, initialise);
  C2RI I226 (ifint_0n[9], i_0r0d[9], gate680_0n, initialise);
  C2RI I227 (ifint_0n[10], i_0r0d[10], gate680_0n, initialise);
  C2RI I228 (ifint_0n[11], i_0r0d[11], gate680_0n, initialise);
  C2RI I229 (ifint_0n[12], i_0r0d[12], gate680_0n, initialise);
  C2RI I230 (ifint_0n[13], i_0r0d[13], gate680_0n, initialise);
  C2RI I231 (ifint_0n[14], i_0r0d[14], gate680_0n, initialise);
  C2RI I232 (ifint_0n[15], i_0r0d[15], gate680_0n, initialise);
  C2RI I233 (ifint_0n[16], i_0r0d[16], gate680_0n, initialise);
  C2RI I234 (ifint_0n[17], i_0r0d[17], gate680_0n, initialise);
  C2RI I235 (ifint_0n[18], i_0r0d[18], gate680_0n, initialise);
  C2RI I236 (ifint_0n[19], i_0r0d[19], gate680_0n, initialise);
  C2RI I237 (ifint_0n[20], i_0r0d[20], gate680_0n, initialise);
  C2RI I238 (ifint_0n[21], i_0r0d[21], gate680_0n, initialise);
  C2RI I239 (ifint_0n[22], i_0r0d[22], gate680_0n, initialise);
  C2RI I240 (ifint_0n[23], i_0r0d[23], gate680_0n, initialise);
  C2RI I241 (ifint_0n[24], i_0r0d[24], gate680_0n, initialise);
  C2RI I242 (ifint_0n[25], i_0r0d[25], gate680_0n, initialise);
  C2RI I243 (ifint_0n[26], i_0r0d[26], gate680_0n, initialise);
  C2RI I244 (ifint_0n[27], i_0r0d[27], gate680_0n, initialise);
  C2RI I245 (ifint_0n[28], i_0r0d[28], gate680_0n, initialise);
  C2RI I246 (ifint_0n[29], i_0r0d[29], gate680_0n, initialise);
  C2RI I247 (ifint_0n[30], i_0r0d[30], gate680_0n, initialise);
  C2RI I248 (ifint_0n[31], i_0r0d[31], gate680_0n, initialise);
  C2RI I249 (ifint_0n[32], i_0r0d[32], gate680_0n, initialise);
  C2RI I250 (ifint_0n[33], i_0r0d[33], gate680_0n, initialise);
  C2RI I251 (ifint_0n[34], i_0r0d[34], gate680_0n, initialise);
  C3 I252 (internal_0n[36], complete677_0n[0], complete677_0n[1], complete677_0n[2]);
  C3 I253 (internal_0n[37], complete677_0n[3], complete677_0n[4], complete677_0n[5]);
  C3 I254 (internal_0n[38], complete677_0n[6], complete677_0n[7], complete677_0n[8]);
  C3 I255 (internal_0n[39], complete677_0n[9], complete677_0n[10], complete677_0n[11]);
  C3 I256 (internal_0n[40], complete677_0n[12], complete677_0n[13], complete677_0n[14]);
  C3 I257 (internal_0n[41], complete677_0n[15], complete677_0n[16], complete677_0n[17]);
  C3 I258 (internal_0n[42], complete677_0n[18], complete677_0n[19], complete677_0n[20]);
  C3 I259 (internal_0n[43], complete677_0n[21], complete677_0n[22], complete677_0n[23]);
  C3 I260 (internal_0n[44], complete677_0n[24], complete677_0n[25], complete677_0n[26]);
  C3 I261 (internal_0n[45], complete677_0n[27], complete677_0n[28], complete677_0n[29]);
  C3 I262 (internal_0n[46], complete677_0n[30], complete677_0n[31], complete677_0n[32]);
  C3 I263 (internal_0n[47], complete677_0n[33], complete677_0n[34], complete677_0n[35]);
  C3 I264 (internal_0n[48], complete677_0n[36], complete677_0n[37], complete677_0n[38]);
  C3 I265 (internal_0n[49], complete677_0n[39], complete677_0n[40], complete677_0n[41]);
  C3 I266 (internal_0n[50], complete677_0n[42], complete677_0n[43], complete677_0n[44]);
  C3 I267 (internal_0n[51], complete677_0n[45], complete677_0n[46], complete677_0n[47]);
  C3 I268 (internal_0n[52], complete677_0n[48], complete677_0n[49], complete677_0n[50]);
  C3 I269 (internal_0n[53], complete677_0n[51], complete677_0n[52], complete677_0n[53]);
  C3 I270 (internal_0n[54], complete677_0n[54], complete677_0n[55], complete677_0n[56]);
  C3 I271 (internal_0n[55], complete677_0n[57], complete677_0n[58], complete677_0n[59]);
  C3 I272 (internal_0n[56], complete677_0n[60], complete677_0n[61], complete677_0n[62]);
  C3 I273 (internal_0n[57], complete677_0n[63], complete677_0n[64], complete677_0n[65]);
  C2 I274 (internal_0n[58], complete677_0n[66], complete677_0n[67]);
  C2 I275 (internal_0n[59], complete677_0n[68], complete677_0n[69]);
  C3 I276 (internal_0n[60], internal_0n[36], internal_0n[37], internal_0n[38]);
  C3 I277 (internal_0n[61], internal_0n[39], internal_0n[40], internal_0n[41]);
  C3 I278 (internal_0n[62], internal_0n[42], internal_0n[43], internal_0n[44]);
  C3 I279 (internal_0n[63], internal_0n[45], internal_0n[46], internal_0n[47]);
  C3 I280 (internal_0n[64], internal_0n[48], internal_0n[49], internal_0n[50]);
  C3 I281 (internal_0n[65], internal_0n[51], internal_0n[52], internal_0n[53]);
  C3 I282 (internal_0n[66], internal_0n[54], internal_0n[55], internal_0n[56]);
  C3 I283 (internal_0n[67], internal_0n[57], internal_0n[58], internal_0n[59]);
  C3 I284 (internal_0n[68], internal_0n[60], internal_0n[61], internal_0n[62]);
  C3 I285 (internal_0n[69], internal_0n[63], internal_0n[64], internal_0n[65]);
  C2 I286 (internal_0n[70], internal_0n[66], internal_0n[67]);
  C3 I287 (oaint_0n, internal_0n[68], internal_0n[69], internal_0n[70]);
  OR2 I288 (complete677_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I289 (complete677_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I290 (complete677_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I291 (complete677_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I292 (complete677_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I293 (complete677_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I294 (complete677_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I295 (complete677_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I296 (complete677_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I297 (complete677_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I298 (complete677_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I299 (complete677_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I300 (complete677_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I301 (complete677_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I302 (complete677_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I303 (complete677_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I304 (complete677_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I305 (complete677_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I306 (complete677_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I307 (complete677_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I308 (complete677_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I309 (complete677_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I310 (complete677_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I311 (complete677_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I312 (complete677_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I313 (complete677_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I314 (complete677_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I315 (complete677_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I316 (complete677_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I317 (complete677_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I318 (complete677_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I319 (complete677_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I320 (complete677_0n[32], o_0r0d[32], o_0r1d[32]);
  OR2 I321 (complete677_0n[33], o_0r0d[33], o_0r1d[33]);
  OR2 I322 (complete677_0n[34], o_0r0d[34], o_0r1d[34]);
  OR2 I323 (complete677_0n[35], o_0r0d[35], o_0r1d[35]);
  OR2 I324 (complete677_0n[36], o_0r0d[36], o_0r1d[36]);
  OR2 I325 (complete677_0n[37], o_0r0d[37], o_0r1d[37]);
  OR2 I326 (complete677_0n[38], o_0r0d[38], o_0r1d[38]);
  OR2 I327 (complete677_0n[39], o_0r0d[39], o_0r1d[39]);
  OR2 I328 (complete677_0n[40], o_0r0d[40], o_0r1d[40]);
  OR2 I329 (complete677_0n[41], o_0r0d[41], o_0r1d[41]);
  OR2 I330 (complete677_0n[42], o_0r0d[42], o_0r1d[42]);
  OR2 I331 (complete677_0n[43], o_0r0d[43], o_0r1d[43]);
  OR2 I332 (complete677_0n[44], o_0r0d[44], o_0r1d[44]);
  OR2 I333 (complete677_0n[45], o_0r0d[45], o_0r1d[45]);
  OR2 I334 (complete677_0n[46], o_0r0d[46], o_0r1d[46]);
  OR2 I335 (complete677_0n[47], o_0r0d[47], o_0r1d[47]);
  OR2 I336 (complete677_0n[48], o_0r0d[48], o_0r1d[48]);
  OR2 I337 (complete677_0n[49], o_0r0d[49], o_0r1d[49]);
  OR2 I338 (complete677_0n[50], o_0r0d[50], o_0r1d[50]);
  OR2 I339 (complete677_0n[51], o_0r0d[51], o_0r1d[51]);
  OR2 I340 (complete677_0n[52], o_0r0d[52], o_0r1d[52]);
  OR2 I341 (complete677_0n[53], o_0r0d[53], o_0r1d[53]);
  OR2 I342 (complete677_0n[54], o_0r0d[54], o_0r1d[54]);
  OR2 I343 (complete677_0n[55], o_0r0d[55], o_0r1d[55]);
  OR2 I344 (complete677_0n[56], o_0r0d[56], o_0r1d[56]);
  OR2 I345 (complete677_0n[57], o_0r0d[57], o_0r1d[57]);
  OR2 I346 (complete677_0n[58], o_0r0d[58], o_0r1d[58]);
  OR2 I347 (complete677_0n[59], o_0r0d[59], o_0r1d[59]);
  OR2 I348 (complete677_0n[60], o_0r0d[60], o_0r1d[60]);
  OR2 I349 (complete677_0n[61], o_0r0d[61], o_0r1d[61]);
  OR2 I350 (complete677_0n[62], o_0r0d[62], o_0r1d[62]);
  OR2 I351 (complete677_0n[63], o_0r0d[63], o_0r1d[63]);
  OR2 I352 (complete677_0n[64], o_0r0d[64], o_0r1d[64]);
  OR2 I353 (complete677_0n[65], o_0r0d[65], o_0r1d[65]);
  OR2 I354 (complete677_0n[66], o_0r0d[66], o_0r1d[66]);
  OR2 I355 (complete677_0n[67], o_0r0d[67], o_0r1d[67]);
  OR2 I356 (complete677_0n[68], o_0r0d[68], o_0r1d[68]);
  OR2 I357 (complete677_0n[69], o_0r0d[69], o_0r1d[69]);
  INV I358 (gate676_0n, o_0a);
  C2RI I359 (o_0r1d[0], otint_0n[0], gate676_0n, initialise);
  C2RI I360 (o_0r1d[1], otint_0n[1], gate676_0n, initialise);
  C2RI I361 (o_0r1d[2], otint_0n[2], gate676_0n, initialise);
  C2RI I362 (o_0r1d[3], otint_0n[3], gate676_0n, initialise);
  C2RI I363 (o_0r1d[4], otint_0n[4], gate676_0n, initialise);
  C2RI I364 (o_0r1d[5], otint_0n[5], gate676_0n, initialise);
  C2RI I365 (o_0r1d[6], otint_0n[6], gate676_0n, initialise);
  C2RI I366 (o_0r1d[7], otint_0n[7], gate676_0n, initialise);
  C2RI I367 (o_0r1d[8], otint_0n[8], gate676_0n, initialise);
  C2RI I368 (o_0r1d[9], otint_0n[9], gate676_0n, initialise);
  C2RI I369 (o_0r1d[10], otint_0n[10], gate676_0n, initialise);
  C2RI I370 (o_0r1d[11], otint_0n[11], gate676_0n, initialise);
  C2RI I371 (o_0r1d[12], otint_0n[12], gate676_0n, initialise);
  C2RI I372 (o_0r1d[13], otint_0n[13], gate676_0n, initialise);
  C2RI I373 (o_0r1d[14], otint_0n[14], gate676_0n, initialise);
  C2RI I374 (o_0r1d[15], otint_0n[15], gate676_0n, initialise);
  C2RI I375 (o_0r1d[16], otint_0n[16], gate676_0n, initialise);
  C2RI I376 (o_0r1d[17], otint_0n[17], gate676_0n, initialise);
  C2RI I377 (o_0r1d[18], otint_0n[18], gate676_0n, initialise);
  C2RI I378 (o_0r1d[19], otint_0n[19], gate676_0n, initialise);
  C2RI I379 (o_0r1d[20], otint_0n[20], gate676_0n, initialise);
  C2RI I380 (o_0r1d[21], otint_0n[21], gate676_0n, initialise);
  C2RI I381 (o_0r1d[22], otint_0n[22], gate676_0n, initialise);
  C2RI I382 (o_0r1d[23], otint_0n[23], gate676_0n, initialise);
  C2RI I383 (o_0r1d[24], otint_0n[24], gate676_0n, initialise);
  C2RI I384 (o_0r1d[25], otint_0n[25], gate676_0n, initialise);
  C2RI I385 (o_0r1d[26], otint_0n[26], gate676_0n, initialise);
  C2RI I386 (o_0r1d[27], otint_0n[27], gate676_0n, initialise);
  C2RI I387 (o_0r1d[28], otint_0n[28], gate676_0n, initialise);
  C2RI I388 (o_0r1d[29], otint_0n[29], gate676_0n, initialise);
  C2RI I389 (o_0r1d[30], otint_0n[30], gate676_0n, initialise);
  C2RI I390 (o_0r1d[31], otint_0n[31], gate676_0n, initialise);
  C2RI I391 (o_0r1d[32], otint_0n[32], gate676_0n, initialise);
  C2RI I392 (o_0r1d[33], otint_0n[33], gate676_0n, initialise);
  C2RI I393 (o_0r1d[34], otint_0n[34], gate676_0n, initialise);
  C2RI I394 (o_0r1d[35], otint_0n[35], gate676_0n, initialise);
  C2RI I395 (o_0r1d[36], otint_0n[36], gate676_0n, initialise);
  C2RI I396 (o_0r1d[37], otint_0n[37], gate676_0n, initialise);
  C2RI I397 (o_0r1d[38], otint_0n[38], gate676_0n, initialise);
  C2RI I398 (o_0r1d[39], otint_0n[39], gate676_0n, initialise);
  C2RI I399 (o_0r1d[40], otint_0n[40], gate676_0n, initialise);
  C2RI I400 (o_0r1d[41], otint_0n[41], gate676_0n, initialise);
  C2RI I401 (o_0r1d[42], otint_0n[42], gate676_0n, initialise);
  C2RI I402 (o_0r1d[43], otint_0n[43], gate676_0n, initialise);
  C2RI I403 (o_0r1d[44], otint_0n[44], gate676_0n, initialise);
  C2RI I404 (o_0r1d[45], otint_0n[45], gate676_0n, initialise);
  C2RI I405 (o_0r1d[46], otint_0n[46], gate676_0n, initialise);
  C2RI I406 (o_0r1d[47], otint_0n[47], gate676_0n, initialise);
  C2RI I407 (o_0r1d[48], otint_0n[48], gate676_0n, initialise);
  C2RI I408 (o_0r1d[49], otint_0n[49], gate676_0n, initialise);
  C2RI I409 (o_0r1d[50], otint_0n[50], gate676_0n, initialise);
  C2RI I410 (o_0r1d[51], otint_0n[51], gate676_0n, initialise);
  C2RI I411 (o_0r1d[52], otint_0n[52], gate676_0n, initialise);
  C2RI I412 (o_0r1d[53], otint_0n[53], gate676_0n, initialise);
  C2RI I413 (o_0r1d[54], otint_0n[54], gate676_0n, initialise);
  C2RI I414 (o_0r1d[55], otint_0n[55], gate676_0n, initialise);
  C2RI I415 (o_0r1d[56], otint_0n[56], gate676_0n, initialise);
  C2RI I416 (o_0r1d[57], otint_0n[57], gate676_0n, initialise);
  C2RI I417 (o_0r1d[58], otint_0n[58], gate676_0n, initialise);
  C2RI I418 (o_0r1d[59], otint_0n[59], gate676_0n, initialise);
  C2RI I419 (o_0r1d[60], otint_0n[60], gate676_0n, initialise);
  C2RI I420 (o_0r1d[61], otint_0n[61], gate676_0n, initialise);
  C2RI I421 (o_0r1d[62], otint_0n[62], gate676_0n, initialise);
  C2RI I422 (o_0r1d[63], otint_0n[63], gate676_0n, initialise);
  C2RI I423 (o_0r1d[64], otint_0n[64], gate676_0n, initialise);
  C2RI I424 (o_0r1d[65], otint_0n[65], gate676_0n, initialise);
  C2RI I425 (o_0r1d[66], otint_0n[66], gate676_0n, initialise);
  C2RI I426 (o_0r1d[67], otint_0n[67], gate676_0n, initialise);
  C2RI I427 (o_0r1d[68], otint_0n[68], gate676_0n, initialise);
  C2RI I428 (o_0r1d[69], otint_0n[69], gate676_0n, initialise);
  C2RI I429 (o_0r0d[0], ofint_0n[0], gate676_0n, initialise);
  C2RI I430 (o_0r0d[1], ofint_0n[1], gate676_0n, initialise);
  C2RI I431 (o_0r0d[2], ofint_0n[2], gate676_0n, initialise);
  C2RI I432 (o_0r0d[3], ofint_0n[3], gate676_0n, initialise);
  C2RI I433 (o_0r0d[4], ofint_0n[4], gate676_0n, initialise);
  C2RI I434 (o_0r0d[5], ofint_0n[5], gate676_0n, initialise);
  C2RI I435 (o_0r0d[6], ofint_0n[6], gate676_0n, initialise);
  C2RI I436 (o_0r0d[7], ofint_0n[7], gate676_0n, initialise);
  C2RI I437 (o_0r0d[8], ofint_0n[8], gate676_0n, initialise);
  C2RI I438 (o_0r0d[9], ofint_0n[9], gate676_0n, initialise);
  C2RI I439 (o_0r0d[10], ofint_0n[10], gate676_0n, initialise);
  C2RI I440 (o_0r0d[11], ofint_0n[11], gate676_0n, initialise);
  C2RI I441 (o_0r0d[12], ofint_0n[12], gate676_0n, initialise);
  C2RI I442 (o_0r0d[13], ofint_0n[13], gate676_0n, initialise);
  C2RI I443 (o_0r0d[14], ofint_0n[14], gate676_0n, initialise);
  C2RI I444 (o_0r0d[15], ofint_0n[15], gate676_0n, initialise);
  C2RI I445 (o_0r0d[16], ofint_0n[16], gate676_0n, initialise);
  C2RI I446 (o_0r0d[17], ofint_0n[17], gate676_0n, initialise);
  C2RI I447 (o_0r0d[18], ofint_0n[18], gate676_0n, initialise);
  C2RI I448 (o_0r0d[19], ofint_0n[19], gate676_0n, initialise);
  C2RI I449 (o_0r0d[20], ofint_0n[20], gate676_0n, initialise);
  C2RI I450 (o_0r0d[21], ofint_0n[21], gate676_0n, initialise);
  C2RI I451 (o_0r0d[22], ofint_0n[22], gate676_0n, initialise);
  C2RI I452 (o_0r0d[23], ofint_0n[23], gate676_0n, initialise);
  C2RI I453 (o_0r0d[24], ofint_0n[24], gate676_0n, initialise);
  C2RI I454 (o_0r0d[25], ofint_0n[25], gate676_0n, initialise);
  C2RI I455 (o_0r0d[26], ofint_0n[26], gate676_0n, initialise);
  C2RI I456 (o_0r0d[27], ofint_0n[27], gate676_0n, initialise);
  C2RI I457 (o_0r0d[28], ofint_0n[28], gate676_0n, initialise);
  C2RI I458 (o_0r0d[29], ofint_0n[29], gate676_0n, initialise);
  C2RI I459 (o_0r0d[30], ofint_0n[30], gate676_0n, initialise);
  C2RI I460 (o_0r0d[31], ofint_0n[31], gate676_0n, initialise);
  C2RI I461 (o_0r0d[32], ofint_0n[32], gate676_0n, initialise);
  C2RI I462 (o_0r0d[33], ofint_0n[33], gate676_0n, initialise);
  C2RI I463 (o_0r0d[34], ofint_0n[34], gate676_0n, initialise);
  C2RI I464 (o_0r0d[35], ofint_0n[35], gate676_0n, initialise);
  C2RI I465 (o_0r0d[36], ofint_0n[36], gate676_0n, initialise);
  C2RI I466 (o_0r0d[37], ofint_0n[37], gate676_0n, initialise);
  C2RI I467 (o_0r0d[38], ofint_0n[38], gate676_0n, initialise);
  C2RI I468 (o_0r0d[39], ofint_0n[39], gate676_0n, initialise);
  C2RI I469 (o_0r0d[40], ofint_0n[40], gate676_0n, initialise);
  C2RI I470 (o_0r0d[41], ofint_0n[41], gate676_0n, initialise);
  C2RI I471 (o_0r0d[42], ofint_0n[42], gate676_0n, initialise);
  C2RI I472 (o_0r0d[43], ofint_0n[43], gate676_0n, initialise);
  C2RI I473 (o_0r0d[44], ofint_0n[44], gate676_0n, initialise);
  C2RI I474 (o_0r0d[45], ofint_0n[45], gate676_0n, initialise);
  C2RI I475 (o_0r0d[46], ofint_0n[46], gate676_0n, initialise);
  C2RI I476 (o_0r0d[47], ofint_0n[47], gate676_0n, initialise);
  C2RI I477 (o_0r0d[48], ofint_0n[48], gate676_0n, initialise);
  C2RI I478 (o_0r0d[49], ofint_0n[49], gate676_0n, initialise);
  C2RI I479 (o_0r0d[50], ofint_0n[50], gate676_0n, initialise);
  C2RI I480 (o_0r0d[51], ofint_0n[51], gate676_0n, initialise);
  C2RI I481 (o_0r0d[52], ofint_0n[52], gate676_0n, initialise);
  C2RI I482 (o_0r0d[53], ofint_0n[53], gate676_0n, initialise);
  C2RI I483 (o_0r0d[54], ofint_0n[54], gate676_0n, initialise);
  C2RI I484 (o_0r0d[55], ofint_0n[55], gate676_0n, initialise);
  C2RI I485 (o_0r0d[56], ofint_0n[56], gate676_0n, initialise);
  C2RI I486 (o_0r0d[57], ofint_0n[57], gate676_0n, initialise);
  C2RI I487 (o_0r0d[58], ofint_0n[58], gate676_0n, initialise);
  C2RI I488 (o_0r0d[59], ofint_0n[59], gate676_0n, initialise);
  C2RI I489 (o_0r0d[60], ofint_0n[60], gate676_0n, initialise);
  C2RI I490 (o_0r0d[61], ofint_0n[61], gate676_0n, initialise);
  C2RI I491 (o_0r0d[62], ofint_0n[62], gate676_0n, initialise);
  C2RI I492 (o_0r0d[63], ofint_0n[63], gate676_0n, initialise);
  C2RI I493 (o_0r0d[64], ofint_0n[64], gate676_0n, initialise);
  C2RI I494 (o_0r0d[65], ofint_0n[65], gate676_0n, initialise);
  C2RI I495 (o_0r0d[66], ofint_0n[66], gate676_0n, initialise);
  C2RI I496 (o_0r0d[67], ofint_0n[67], gate676_0n, initialise);
  C2RI I497 (o_0r0d[68], ofint_0n[68], gate676_0n, initialise);
  C2RI I498 (o_0r0d[69], ofint_0n[69], gate676_0n, initialise);
  assign otint_0n[0] = itint_0n[0];
  assign otint_0n[1] = itint_0n[1];
  assign otint_0n[2] = itint_0n[2];
  assign otint_0n[3] = itint_0n[3];
  assign otint_0n[4] = itint_0n[4];
  assign otint_0n[5] = itint_0n[5];
  assign otint_0n[6] = itint_0n[6];
  assign otint_0n[7] = itint_0n[7];
  assign otint_0n[8] = itint_0n[8];
  assign otint_0n[9] = itint_0n[9];
  assign otint_0n[10] = itint_0n[10];
  assign otint_0n[11] = itint_0n[11];
  assign otint_0n[12] = itint_0n[12];
  assign otint_0n[13] = itint_0n[13];
  assign otint_0n[14] = itint_0n[14];
  assign otint_0n[15] = itint_0n[15];
  assign otint_0n[16] = itint_0n[16];
  assign otint_0n[17] = itint_0n[17];
  assign otint_0n[18] = itint_0n[18];
  assign otint_0n[19] = itint_0n[19];
  assign otint_0n[20] = itint_0n[20];
  assign otint_0n[21] = itint_0n[21];
  assign otint_0n[22] = itint_0n[22];
  assign otint_0n[23] = itint_0n[23];
  assign otint_0n[24] = itint_0n[24];
  assign otint_0n[25] = itint_0n[25];
  assign otint_0n[26] = itint_0n[26];
  assign otint_0n[27] = itint_0n[27];
  assign otint_0n[28] = itint_0n[28];
  assign otint_0n[29] = itint_0n[29];
  assign otint_0n[30] = itint_0n[30];
  assign otint_0n[31] = itint_0n[31];
  assign otint_0n[32] = itint_0n[32];
  assign otint_0n[33] = itint_0n[33];
  assign otint_0n[34] = itint_0n[34];
  assign otint_0n[35] = itint_1n[0];
  assign otint_0n[36] = itint_1n[1];
  assign otint_0n[37] = itint_1n[2];
  assign otint_0n[38] = itint_1n[3];
  assign otint_0n[39] = itint_1n[4];
  assign otint_0n[40] = itint_1n[5];
  assign otint_0n[41] = itint_1n[6];
  assign otint_0n[42] = itint_1n[7];
  assign otint_0n[43] = itint_1n[8];
  assign otint_0n[44] = itint_1n[9];
  assign otint_0n[45] = itint_1n[10];
  assign otint_0n[46] = itint_1n[11];
  assign otint_0n[47] = itint_1n[12];
  assign otint_0n[48] = itint_1n[13];
  assign otint_0n[49] = itint_1n[14];
  assign otint_0n[50] = itint_1n[15];
  assign otint_0n[51] = itint_1n[16];
  assign otint_0n[52] = itint_1n[17];
  assign otint_0n[53] = itint_1n[18];
  assign otint_0n[54] = itint_1n[19];
  assign otint_0n[55] = itint_1n[20];
  assign otint_0n[56] = itint_1n[21];
  assign otint_0n[57] = itint_1n[22];
  assign otint_0n[58] = itint_1n[23];
  assign otint_0n[59] = itint_1n[24];
  assign otint_0n[60] = itint_1n[25];
  assign otint_0n[61] = itint_1n[26];
  assign otint_0n[62] = itint_1n[27];
  assign otint_0n[63] = itint_1n[28];
  assign otint_0n[64] = itint_1n[29];
  assign otint_0n[65] = itint_1n[30];
  assign otint_0n[66] = itint_1n[31];
  assign otint_0n[67] = itint_1n[32];
  assign otint_0n[68] = itint_1n[33];
  assign otint_0n[69] = itint_1n[34];
  assign ofint_0n[0] = ifint_0n[0];
  assign ofint_0n[1] = ifint_0n[1];
  assign ofint_0n[2] = ifint_0n[2];
  assign ofint_0n[3] = ifint_0n[3];
  assign ofint_0n[4] = ifint_0n[4];
  assign ofint_0n[5] = ifint_0n[5];
  assign ofint_0n[6] = ifint_0n[6];
  assign ofint_0n[7] = ifint_0n[7];
  assign ofint_0n[8] = ifint_0n[8];
  assign ofint_0n[9] = ifint_0n[9];
  assign ofint_0n[10] = ifint_0n[10];
  assign ofint_0n[11] = ifint_0n[11];
  assign ofint_0n[12] = ifint_0n[12];
  assign ofint_0n[13] = ifint_0n[13];
  assign ofint_0n[14] = ifint_0n[14];
  assign ofint_0n[15] = ifint_0n[15];
  assign ofint_0n[16] = ifint_0n[16];
  assign ofint_0n[17] = ifint_0n[17];
  assign ofint_0n[18] = ifint_0n[18];
  assign ofint_0n[19] = ifint_0n[19];
  assign ofint_0n[20] = ifint_0n[20];
  assign ofint_0n[21] = ifint_0n[21];
  assign ofint_0n[22] = ifint_0n[22];
  assign ofint_0n[23] = ifint_0n[23];
  assign ofint_0n[24] = ifint_0n[24];
  assign ofint_0n[25] = ifint_0n[25];
  assign ofint_0n[26] = ifint_0n[26];
  assign ofint_0n[27] = ifint_0n[27];
  assign ofint_0n[28] = ifint_0n[28];
  assign ofint_0n[29] = ifint_0n[29];
  assign ofint_0n[30] = ifint_0n[30];
  assign ofint_0n[31] = ifint_0n[31];
  assign ofint_0n[32] = ifint_0n[32];
  assign ofint_0n[33] = ifint_0n[33];
  assign ofint_0n[34] = ifint_0n[34];
  assign ofint_0n[35] = ifint_1n[0];
  assign ofint_0n[36] = ifint_1n[1];
  assign ofint_0n[37] = ifint_1n[2];
  assign ofint_0n[38] = ifint_1n[3];
  assign ofint_0n[39] = ifint_1n[4];
  assign ofint_0n[40] = ifint_1n[5];
  assign ofint_0n[41] = ifint_1n[6];
  assign ofint_0n[42] = ifint_1n[7];
  assign ofint_0n[43] = ifint_1n[8];
  assign ofint_0n[44] = ifint_1n[9];
  assign ofint_0n[45] = ifint_1n[10];
  assign ofint_0n[46] = ifint_1n[11];
  assign ofint_0n[47] = ifint_1n[12];
  assign ofint_0n[48] = ifint_1n[13];
  assign ofint_0n[49] = ifint_1n[14];
  assign ofint_0n[50] = ifint_1n[15];
  assign ofint_0n[51] = ifint_1n[16];
  assign ofint_0n[52] = ifint_1n[17];
  assign ofint_0n[53] = ifint_1n[18];
  assign ofint_0n[54] = ifint_1n[19];
  assign ofint_0n[55] = ifint_1n[20];
  assign ofint_0n[56] = ifint_1n[21];
  assign ofint_0n[57] = ifint_1n[22];
  assign ofint_0n[58] = ifint_1n[23];
  assign ofint_0n[59] = ifint_1n[24];
  assign ofint_0n[60] = ifint_1n[25];
  assign ofint_0n[61] = ifint_1n[26];
  assign ofint_0n[62] = ifint_1n[27];
  assign ofint_0n[63] = ifint_1n[28];
  assign ofint_0n[64] = ifint_1n[29];
  assign ofint_0n[65] = ifint_1n[30];
  assign ofint_0n[66] = ifint_1n[31];
  assign ofint_0n[67] = ifint_1n[32];
  assign ofint_0n[68] = ifint_1n[33];
  assign ofint_0n[69] = ifint_1n[34];
endmodule

module BrzJ_l12__2836_200_29 (
  i_0r0d, i_0r1d, i_0a,
  i_1r, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [35:0] i_0r0d;
  input [35:0] i_0r1d;
  output i_0a;
  input i_1r;
  output i_1a;
  output [35:0] o_0r0d;
  output [35:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [35:0] internal_0n;
  wire [35:0] ofint_0n;
  wire [35:0] otint_0n;
  wire oaint_0n;
  wire [35:0] ifint_0n;
  wire ifint_1n;
  wire [35:0] itint_0n;
  wire iaint_0n;
  wire iaint_1n;
  wire gate696_0n;
  wire [35:0] complete693_0n;
  wire gate692_0n;
  wire [35:0] complete689_0n;
  wire gate688_0n;
  wire [35:0] joint_0n;
  wire [35:0] joinf_0n;
  wire icomplete_0n;
  assign iaint_0n = oaint_0n;
  assign iaint_1n = oaint_0n;
  assign i_1a = ifint_1n;
  INV I3 (gate696_0n, iaint_1n);
  C2RI I4 (ifint_1n, i_1r, gate696_0n, initialise);
  C3 I5 (internal_0n[0], complete693_0n[0], complete693_0n[1], complete693_0n[2]);
  C3 I6 (internal_0n[1], complete693_0n[3], complete693_0n[4], complete693_0n[5]);
  C3 I7 (internal_0n[2], complete693_0n[6], complete693_0n[7], complete693_0n[8]);
  C3 I8 (internal_0n[3], complete693_0n[9], complete693_0n[10], complete693_0n[11]);
  C3 I9 (internal_0n[4], complete693_0n[12], complete693_0n[13], complete693_0n[14]);
  C3 I10 (internal_0n[5], complete693_0n[15], complete693_0n[16], complete693_0n[17]);
  C3 I11 (internal_0n[6], complete693_0n[18], complete693_0n[19], complete693_0n[20]);
  C3 I12 (internal_0n[7], complete693_0n[21], complete693_0n[22], complete693_0n[23]);
  C3 I13 (internal_0n[8], complete693_0n[24], complete693_0n[25], complete693_0n[26]);
  C3 I14 (internal_0n[9], complete693_0n[27], complete693_0n[28], complete693_0n[29]);
  C3 I15 (internal_0n[10], complete693_0n[30], complete693_0n[31], complete693_0n[32]);
  C3 I16 (internal_0n[11], complete693_0n[33], complete693_0n[34], complete693_0n[35]);
  C3 I17 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I18 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I19 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I20 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I21 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I22 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I23 (i_0a, internal_0n[16], internal_0n[17]);
  OR2 I24 (complete693_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I25 (complete693_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I26 (complete693_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I27 (complete693_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I28 (complete693_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I29 (complete693_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I30 (complete693_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I31 (complete693_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I32 (complete693_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I33 (complete693_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I34 (complete693_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I35 (complete693_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I36 (complete693_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I37 (complete693_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I38 (complete693_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I39 (complete693_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I40 (complete693_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I41 (complete693_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I42 (complete693_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I43 (complete693_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I44 (complete693_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I45 (complete693_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I46 (complete693_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I47 (complete693_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I48 (complete693_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I49 (complete693_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I50 (complete693_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I51 (complete693_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I52 (complete693_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I53 (complete693_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I54 (complete693_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I55 (complete693_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I56 (complete693_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I57 (complete693_0n[33], ifint_0n[33], itint_0n[33]);
  OR2 I58 (complete693_0n[34], ifint_0n[34], itint_0n[34]);
  OR2 I59 (complete693_0n[35], ifint_0n[35], itint_0n[35]);
  INV I60 (gate692_0n, iaint_0n);
  C2RI I61 (itint_0n[0], i_0r1d[0], gate692_0n, initialise);
  C2RI I62 (itint_0n[1], i_0r1d[1], gate692_0n, initialise);
  C2RI I63 (itint_0n[2], i_0r1d[2], gate692_0n, initialise);
  C2RI I64 (itint_0n[3], i_0r1d[3], gate692_0n, initialise);
  C2RI I65 (itint_0n[4], i_0r1d[4], gate692_0n, initialise);
  C2RI I66 (itint_0n[5], i_0r1d[5], gate692_0n, initialise);
  C2RI I67 (itint_0n[6], i_0r1d[6], gate692_0n, initialise);
  C2RI I68 (itint_0n[7], i_0r1d[7], gate692_0n, initialise);
  C2RI I69 (itint_0n[8], i_0r1d[8], gate692_0n, initialise);
  C2RI I70 (itint_0n[9], i_0r1d[9], gate692_0n, initialise);
  C2RI I71 (itint_0n[10], i_0r1d[10], gate692_0n, initialise);
  C2RI I72 (itint_0n[11], i_0r1d[11], gate692_0n, initialise);
  C2RI I73 (itint_0n[12], i_0r1d[12], gate692_0n, initialise);
  C2RI I74 (itint_0n[13], i_0r1d[13], gate692_0n, initialise);
  C2RI I75 (itint_0n[14], i_0r1d[14], gate692_0n, initialise);
  C2RI I76 (itint_0n[15], i_0r1d[15], gate692_0n, initialise);
  C2RI I77 (itint_0n[16], i_0r1d[16], gate692_0n, initialise);
  C2RI I78 (itint_0n[17], i_0r1d[17], gate692_0n, initialise);
  C2RI I79 (itint_0n[18], i_0r1d[18], gate692_0n, initialise);
  C2RI I80 (itint_0n[19], i_0r1d[19], gate692_0n, initialise);
  C2RI I81 (itint_0n[20], i_0r1d[20], gate692_0n, initialise);
  C2RI I82 (itint_0n[21], i_0r1d[21], gate692_0n, initialise);
  C2RI I83 (itint_0n[22], i_0r1d[22], gate692_0n, initialise);
  C2RI I84 (itint_0n[23], i_0r1d[23], gate692_0n, initialise);
  C2RI I85 (itint_0n[24], i_0r1d[24], gate692_0n, initialise);
  C2RI I86 (itint_0n[25], i_0r1d[25], gate692_0n, initialise);
  C2RI I87 (itint_0n[26], i_0r1d[26], gate692_0n, initialise);
  C2RI I88 (itint_0n[27], i_0r1d[27], gate692_0n, initialise);
  C2RI I89 (itint_0n[28], i_0r1d[28], gate692_0n, initialise);
  C2RI I90 (itint_0n[29], i_0r1d[29], gate692_0n, initialise);
  C2RI I91 (itint_0n[30], i_0r1d[30], gate692_0n, initialise);
  C2RI I92 (itint_0n[31], i_0r1d[31], gate692_0n, initialise);
  C2RI I93 (itint_0n[32], i_0r1d[32], gate692_0n, initialise);
  C2RI I94 (itint_0n[33], i_0r1d[33], gate692_0n, initialise);
  C2RI I95 (itint_0n[34], i_0r1d[34], gate692_0n, initialise);
  C2RI I96 (itint_0n[35], i_0r1d[35], gate692_0n, initialise);
  C2RI I97 (ifint_0n[0], i_0r0d[0], gate692_0n, initialise);
  C2RI I98 (ifint_0n[1], i_0r0d[1], gate692_0n, initialise);
  C2RI I99 (ifint_0n[2], i_0r0d[2], gate692_0n, initialise);
  C2RI I100 (ifint_0n[3], i_0r0d[3], gate692_0n, initialise);
  C2RI I101 (ifint_0n[4], i_0r0d[4], gate692_0n, initialise);
  C2RI I102 (ifint_0n[5], i_0r0d[5], gate692_0n, initialise);
  C2RI I103 (ifint_0n[6], i_0r0d[6], gate692_0n, initialise);
  C2RI I104 (ifint_0n[7], i_0r0d[7], gate692_0n, initialise);
  C2RI I105 (ifint_0n[8], i_0r0d[8], gate692_0n, initialise);
  C2RI I106 (ifint_0n[9], i_0r0d[9], gate692_0n, initialise);
  C2RI I107 (ifint_0n[10], i_0r0d[10], gate692_0n, initialise);
  C2RI I108 (ifint_0n[11], i_0r0d[11], gate692_0n, initialise);
  C2RI I109 (ifint_0n[12], i_0r0d[12], gate692_0n, initialise);
  C2RI I110 (ifint_0n[13], i_0r0d[13], gate692_0n, initialise);
  C2RI I111 (ifint_0n[14], i_0r0d[14], gate692_0n, initialise);
  C2RI I112 (ifint_0n[15], i_0r0d[15], gate692_0n, initialise);
  C2RI I113 (ifint_0n[16], i_0r0d[16], gate692_0n, initialise);
  C2RI I114 (ifint_0n[17], i_0r0d[17], gate692_0n, initialise);
  C2RI I115 (ifint_0n[18], i_0r0d[18], gate692_0n, initialise);
  C2RI I116 (ifint_0n[19], i_0r0d[19], gate692_0n, initialise);
  C2RI I117 (ifint_0n[20], i_0r0d[20], gate692_0n, initialise);
  C2RI I118 (ifint_0n[21], i_0r0d[21], gate692_0n, initialise);
  C2RI I119 (ifint_0n[22], i_0r0d[22], gate692_0n, initialise);
  C2RI I120 (ifint_0n[23], i_0r0d[23], gate692_0n, initialise);
  C2RI I121 (ifint_0n[24], i_0r0d[24], gate692_0n, initialise);
  C2RI I122 (ifint_0n[25], i_0r0d[25], gate692_0n, initialise);
  C2RI I123 (ifint_0n[26], i_0r0d[26], gate692_0n, initialise);
  C2RI I124 (ifint_0n[27], i_0r0d[27], gate692_0n, initialise);
  C2RI I125 (ifint_0n[28], i_0r0d[28], gate692_0n, initialise);
  C2RI I126 (ifint_0n[29], i_0r0d[29], gate692_0n, initialise);
  C2RI I127 (ifint_0n[30], i_0r0d[30], gate692_0n, initialise);
  C2RI I128 (ifint_0n[31], i_0r0d[31], gate692_0n, initialise);
  C2RI I129 (ifint_0n[32], i_0r0d[32], gate692_0n, initialise);
  C2RI I130 (ifint_0n[33], i_0r0d[33], gate692_0n, initialise);
  C2RI I131 (ifint_0n[34], i_0r0d[34], gate692_0n, initialise);
  C2RI I132 (ifint_0n[35], i_0r0d[35], gate692_0n, initialise);
  C3 I133 (internal_0n[18], complete689_0n[0], complete689_0n[1], complete689_0n[2]);
  C3 I134 (internal_0n[19], complete689_0n[3], complete689_0n[4], complete689_0n[5]);
  C3 I135 (internal_0n[20], complete689_0n[6], complete689_0n[7], complete689_0n[8]);
  C3 I136 (internal_0n[21], complete689_0n[9], complete689_0n[10], complete689_0n[11]);
  C3 I137 (internal_0n[22], complete689_0n[12], complete689_0n[13], complete689_0n[14]);
  C3 I138 (internal_0n[23], complete689_0n[15], complete689_0n[16], complete689_0n[17]);
  C3 I139 (internal_0n[24], complete689_0n[18], complete689_0n[19], complete689_0n[20]);
  C3 I140 (internal_0n[25], complete689_0n[21], complete689_0n[22], complete689_0n[23]);
  C3 I141 (internal_0n[26], complete689_0n[24], complete689_0n[25], complete689_0n[26]);
  C3 I142 (internal_0n[27], complete689_0n[27], complete689_0n[28], complete689_0n[29]);
  C3 I143 (internal_0n[28], complete689_0n[30], complete689_0n[31], complete689_0n[32]);
  C3 I144 (internal_0n[29], complete689_0n[33], complete689_0n[34], complete689_0n[35]);
  C3 I145 (internal_0n[30], internal_0n[18], internal_0n[19], internal_0n[20]);
  C3 I146 (internal_0n[31], internal_0n[21], internal_0n[22], internal_0n[23]);
  C3 I147 (internal_0n[32], internal_0n[24], internal_0n[25], internal_0n[26]);
  C3 I148 (internal_0n[33], internal_0n[27], internal_0n[28], internal_0n[29]);
  C2 I149 (internal_0n[34], internal_0n[30], internal_0n[31]);
  C2 I150 (internal_0n[35], internal_0n[32], internal_0n[33]);
  C2 I151 (oaint_0n, internal_0n[34], internal_0n[35]);
  OR2 I152 (complete689_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I153 (complete689_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I154 (complete689_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I155 (complete689_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I156 (complete689_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I157 (complete689_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I158 (complete689_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I159 (complete689_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I160 (complete689_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I161 (complete689_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I162 (complete689_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I163 (complete689_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I164 (complete689_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I165 (complete689_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I166 (complete689_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I167 (complete689_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I168 (complete689_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I169 (complete689_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I170 (complete689_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I171 (complete689_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I172 (complete689_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I173 (complete689_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I174 (complete689_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I175 (complete689_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I176 (complete689_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I177 (complete689_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I178 (complete689_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I179 (complete689_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I180 (complete689_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I181 (complete689_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I182 (complete689_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I183 (complete689_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I184 (complete689_0n[32], o_0r0d[32], o_0r1d[32]);
  OR2 I185 (complete689_0n[33], o_0r0d[33], o_0r1d[33]);
  OR2 I186 (complete689_0n[34], o_0r0d[34], o_0r1d[34]);
  OR2 I187 (complete689_0n[35], o_0r0d[35], o_0r1d[35]);
  INV I188 (gate688_0n, o_0a);
  C2RI I189 (o_0r1d[0], otint_0n[0], gate688_0n, initialise);
  C2RI I190 (o_0r1d[1], otint_0n[1], gate688_0n, initialise);
  C2RI I191 (o_0r1d[2], otint_0n[2], gate688_0n, initialise);
  C2RI I192 (o_0r1d[3], otint_0n[3], gate688_0n, initialise);
  C2RI I193 (o_0r1d[4], otint_0n[4], gate688_0n, initialise);
  C2RI I194 (o_0r1d[5], otint_0n[5], gate688_0n, initialise);
  C2RI I195 (o_0r1d[6], otint_0n[6], gate688_0n, initialise);
  C2RI I196 (o_0r1d[7], otint_0n[7], gate688_0n, initialise);
  C2RI I197 (o_0r1d[8], otint_0n[8], gate688_0n, initialise);
  C2RI I198 (o_0r1d[9], otint_0n[9], gate688_0n, initialise);
  C2RI I199 (o_0r1d[10], otint_0n[10], gate688_0n, initialise);
  C2RI I200 (o_0r1d[11], otint_0n[11], gate688_0n, initialise);
  C2RI I201 (o_0r1d[12], otint_0n[12], gate688_0n, initialise);
  C2RI I202 (o_0r1d[13], otint_0n[13], gate688_0n, initialise);
  C2RI I203 (o_0r1d[14], otint_0n[14], gate688_0n, initialise);
  C2RI I204 (o_0r1d[15], otint_0n[15], gate688_0n, initialise);
  C2RI I205 (o_0r1d[16], otint_0n[16], gate688_0n, initialise);
  C2RI I206 (o_0r1d[17], otint_0n[17], gate688_0n, initialise);
  C2RI I207 (o_0r1d[18], otint_0n[18], gate688_0n, initialise);
  C2RI I208 (o_0r1d[19], otint_0n[19], gate688_0n, initialise);
  C2RI I209 (o_0r1d[20], otint_0n[20], gate688_0n, initialise);
  C2RI I210 (o_0r1d[21], otint_0n[21], gate688_0n, initialise);
  C2RI I211 (o_0r1d[22], otint_0n[22], gate688_0n, initialise);
  C2RI I212 (o_0r1d[23], otint_0n[23], gate688_0n, initialise);
  C2RI I213 (o_0r1d[24], otint_0n[24], gate688_0n, initialise);
  C2RI I214 (o_0r1d[25], otint_0n[25], gate688_0n, initialise);
  C2RI I215 (o_0r1d[26], otint_0n[26], gate688_0n, initialise);
  C2RI I216 (o_0r1d[27], otint_0n[27], gate688_0n, initialise);
  C2RI I217 (o_0r1d[28], otint_0n[28], gate688_0n, initialise);
  C2RI I218 (o_0r1d[29], otint_0n[29], gate688_0n, initialise);
  C2RI I219 (o_0r1d[30], otint_0n[30], gate688_0n, initialise);
  C2RI I220 (o_0r1d[31], otint_0n[31], gate688_0n, initialise);
  C2RI I221 (o_0r1d[32], otint_0n[32], gate688_0n, initialise);
  C2RI I222 (o_0r1d[33], otint_0n[33], gate688_0n, initialise);
  C2RI I223 (o_0r1d[34], otint_0n[34], gate688_0n, initialise);
  C2RI I224 (o_0r1d[35], otint_0n[35], gate688_0n, initialise);
  C2RI I225 (o_0r0d[0], ofint_0n[0], gate688_0n, initialise);
  C2RI I226 (o_0r0d[1], ofint_0n[1], gate688_0n, initialise);
  C2RI I227 (o_0r0d[2], ofint_0n[2], gate688_0n, initialise);
  C2RI I228 (o_0r0d[3], ofint_0n[3], gate688_0n, initialise);
  C2RI I229 (o_0r0d[4], ofint_0n[4], gate688_0n, initialise);
  C2RI I230 (o_0r0d[5], ofint_0n[5], gate688_0n, initialise);
  C2RI I231 (o_0r0d[6], ofint_0n[6], gate688_0n, initialise);
  C2RI I232 (o_0r0d[7], ofint_0n[7], gate688_0n, initialise);
  C2RI I233 (o_0r0d[8], ofint_0n[8], gate688_0n, initialise);
  C2RI I234 (o_0r0d[9], ofint_0n[9], gate688_0n, initialise);
  C2RI I235 (o_0r0d[10], ofint_0n[10], gate688_0n, initialise);
  C2RI I236 (o_0r0d[11], ofint_0n[11], gate688_0n, initialise);
  C2RI I237 (o_0r0d[12], ofint_0n[12], gate688_0n, initialise);
  C2RI I238 (o_0r0d[13], ofint_0n[13], gate688_0n, initialise);
  C2RI I239 (o_0r0d[14], ofint_0n[14], gate688_0n, initialise);
  C2RI I240 (o_0r0d[15], ofint_0n[15], gate688_0n, initialise);
  C2RI I241 (o_0r0d[16], ofint_0n[16], gate688_0n, initialise);
  C2RI I242 (o_0r0d[17], ofint_0n[17], gate688_0n, initialise);
  C2RI I243 (o_0r0d[18], ofint_0n[18], gate688_0n, initialise);
  C2RI I244 (o_0r0d[19], ofint_0n[19], gate688_0n, initialise);
  C2RI I245 (o_0r0d[20], ofint_0n[20], gate688_0n, initialise);
  C2RI I246 (o_0r0d[21], ofint_0n[21], gate688_0n, initialise);
  C2RI I247 (o_0r0d[22], ofint_0n[22], gate688_0n, initialise);
  C2RI I248 (o_0r0d[23], ofint_0n[23], gate688_0n, initialise);
  C2RI I249 (o_0r0d[24], ofint_0n[24], gate688_0n, initialise);
  C2RI I250 (o_0r0d[25], ofint_0n[25], gate688_0n, initialise);
  C2RI I251 (o_0r0d[26], ofint_0n[26], gate688_0n, initialise);
  C2RI I252 (o_0r0d[27], ofint_0n[27], gate688_0n, initialise);
  C2RI I253 (o_0r0d[28], ofint_0n[28], gate688_0n, initialise);
  C2RI I254 (o_0r0d[29], ofint_0n[29], gate688_0n, initialise);
  C2RI I255 (o_0r0d[30], ofint_0n[30], gate688_0n, initialise);
  C2RI I256 (o_0r0d[31], ofint_0n[31], gate688_0n, initialise);
  C2RI I257 (o_0r0d[32], ofint_0n[32], gate688_0n, initialise);
  C2RI I258 (o_0r0d[33], ofint_0n[33], gate688_0n, initialise);
  C2RI I259 (o_0r0d[34], ofint_0n[34], gate688_0n, initialise);
  C2RI I260 (o_0r0d[35], ofint_0n[35], gate688_0n, initialise);
  assign otint_0n[1] = joint_0n[1];
  assign otint_0n[2] = joint_0n[2];
  assign otint_0n[3] = joint_0n[3];
  assign otint_0n[4] = joint_0n[4];
  assign otint_0n[5] = joint_0n[5];
  assign otint_0n[6] = joint_0n[6];
  assign otint_0n[7] = joint_0n[7];
  assign otint_0n[8] = joint_0n[8];
  assign otint_0n[9] = joint_0n[9];
  assign otint_0n[10] = joint_0n[10];
  assign otint_0n[11] = joint_0n[11];
  assign otint_0n[12] = joint_0n[12];
  assign otint_0n[13] = joint_0n[13];
  assign otint_0n[14] = joint_0n[14];
  assign otint_0n[15] = joint_0n[15];
  assign otint_0n[16] = joint_0n[16];
  assign otint_0n[17] = joint_0n[17];
  assign otint_0n[18] = joint_0n[18];
  assign otint_0n[19] = joint_0n[19];
  assign otint_0n[20] = joint_0n[20];
  assign otint_0n[21] = joint_0n[21];
  assign otint_0n[22] = joint_0n[22];
  assign otint_0n[23] = joint_0n[23];
  assign otint_0n[24] = joint_0n[24];
  assign otint_0n[25] = joint_0n[25];
  assign otint_0n[26] = joint_0n[26];
  assign otint_0n[27] = joint_0n[27];
  assign otint_0n[28] = joint_0n[28];
  assign otint_0n[29] = joint_0n[29];
  assign otint_0n[30] = joint_0n[30];
  assign otint_0n[31] = joint_0n[31];
  assign otint_0n[32] = joint_0n[32];
  assign otint_0n[33] = joint_0n[33];
  assign otint_0n[34] = joint_0n[34];
  assign otint_0n[35] = joint_0n[35];
  assign ofint_0n[1] = joinf_0n[1];
  assign ofint_0n[2] = joinf_0n[2];
  assign ofint_0n[3] = joinf_0n[3];
  assign ofint_0n[4] = joinf_0n[4];
  assign ofint_0n[5] = joinf_0n[5];
  assign ofint_0n[6] = joinf_0n[6];
  assign ofint_0n[7] = joinf_0n[7];
  assign ofint_0n[8] = joinf_0n[8];
  assign ofint_0n[9] = joinf_0n[9];
  assign ofint_0n[10] = joinf_0n[10];
  assign ofint_0n[11] = joinf_0n[11];
  assign ofint_0n[12] = joinf_0n[12];
  assign ofint_0n[13] = joinf_0n[13];
  assign ofint_0n[14] = joinf_0n[14];
  assign ofint_0n[15] = joinf_0n[15];
  assign ofint_0n[16] = joinf_0n[16];
  assign ofint_0n[17] = joinf_0n[17];
  assign ofint_0n[18] = joinf_0n[18];
  assign ofint_0n[19] = joinf_0n[19];
  assign ofint_0n[20] = joinf_0n[20];
  assign ofint_0n[21] = joinf_0n[21];
  assign ofint_0n[22] = joinf_0n[22];
  assign ofint_0n[23] = joinf_0n[23];
  assign ofint_0n[24] = joinf_0n[24];
  assign ofint_0n[25] = joinf_0n[25];
  assign ofint_0n[26] = joinf_0n[26];
  assign ofint_0n[27] = joinf_0n[27];
  assign ofint_0n[28] = joinf_0n[28];
  assign ofint_0n[29] = joinf_0n[29];
  assign ofint_0n[30] = joinf_0n[30];
  assign ofint_0n[31] = joinf_0n[31];
  assign ofint_0n[32] = joinf_0n[32];
  assign ofint_0n[33] = joinf_0n[33];
  assign ofint_0n[34] = joinf_0n[34];
  assign ofint_0n[35] = joinf_0n[35];
  C2 I331 (otint_0n[0], joint_0n[0], icomplete_0n);
  C2 I332 (ofint_0n[0], joinf_0n[0], icomplete_0n);
  assign icomplete_0n = ifint_1n;
  assign joint_0n[0] = itint_0n[0];
  assign joint_0n[1] = itint_0n[1];
  assign joint_0n[2] = itint_0n[2];
  assign joint_0n[3] = itint_0n[3];
  assign joint_0n[4] = itint_0n[4];
  assign joint_0n[5] = itint_0n[5];
  assign joint_0n[6] = itint_0n[6];
  assign joint_0n[7] = itint_0n[7];
  assign joint_0n[8] = itint_0n[8];
  assign joint_0n[9] = itint_0n[9];
  assign joint_0n[10] = itint_0n[10];
  assign joint_0n[11] = itint_0n[11];
  assign joint_0n[12] = itint_0n[12];
  assign joint_0n[13] = itint_0n[13];
  assign joint_0n[14] = itint_0n[14];
  assign joint_0n[15] = itint_0n[15];
  assign joint_0n[16] = itint_0n[16];
  assign joint_0n[17] = itint_0n[17];
  assign joint_0n[18] = itint_0n[18];
  assign joint_0n[19] = itint_0n[19];
  assign joint_0n[20] = itint_0n[20];
  assign joint_0n[21] = itint_0n[21];
  assign joint_0n[22] = itint_0n[22];
  assign joint_0n[23] = itint_0n[23];
  assign joint_0n[24] = itint_0n[24];
  assign joint_0n[25] = itint_0n[25];
  assign joint_0n[26] = itint_0n[26];
  assign joint_0n[27] = itint_0n[27];
  assign joint_0n[28] = itint_0n[28];
  assign joint_0n[29] = itint_0n[29];
  assign joint_0n[30] = itint_0n[30];
  assign joint_0n[31] = itint_0n[31];
  assign joint_0n[32] = itint_0n[32];
  assign joint_0n[33] = itint_0n[33];
  assign joint_0n[34] = itint_0n[34];
  assign joint_0n[35] = itint_0n[35];
  assign joinf_0n[0] = ifint_0n[0];
  assign joinf_0n[1] = ifint_0n[1];
  assign joinf_0n[2] = ifint_0n[2];
  assign joinf_0n[3] = ifint_0n[3];
  assign joinf_0n[4] = ifint_0n[4];
  assign joinf_0n[5] = ifint_0n[5];
  assign joinf_0n[6] = ifint_0n[6];
  assign joinf_0n[7] = ifint_0n[7];
  assign joinf_0n[8] = ifint_0n[8];
  assign joinf_0n[9] = ifint_0n[9];
  assign joinf_0n[10] = ifint_0n[10];
  assign joinf_0n[11] = ifint_0n[11];
  assign joinf_0n[12] = ifint_0n[12];
  assign joinf_0n[13] = ifint_0n[13];
  assign joinf_0n[14] = ifint_0n[14];
  assign joinf_0n[15] = ifint_0n[15];
  assign joinf_0n[16] = ifint_0n[16];
  assign joinf_0n[17] = ifint_0n[17];
  assign joinf_0n[18] = ifint_0n[18];
  assign joinf_0n[19] = ifint_0n[19];
  assign joinf_0n[20] = ifint_0n[20];
  assign joinf_0n[21] = ifint_0n[21];
  assign joinf_0n[22] = ifint_0n[22];
  assign joinf_0n[23] = ifint_0n[23];
  assign joinf_0n[24] = ifint_0n[24];
  assign joinf_0n[25] = ifint_0n[25];
  assign joinf_0n[26] = ifint_0n[26];
  assign joinf_0n[27] = ifint_0n[27];
  assign joinf_0n[28] = ifint_0n[28];
  assign joinf_0n[29] = ifint_0n[29];
  assign joinf_0n[30] = ifint_0n[30];
  assign joinf_0n[31] = ifint_0n[31];
  assign joinf_0n[32] = ifint_0n[32];
  assign joinf_0n[33] = ifint_0n[33];
  assign joinf_0n[34] = ifint_0n[34];
  assign joinf_0n[35] = ifint_0n[35];
endmodule

module BrzM_0_2 (
  i_0r, i_0a,
  i_1r, i_1a,
  o_0r, o_0a,
  initialise
);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  output o_0r;
  input o_0a;
  input initialise;
  wire [1:0] sel_0n;
  wire ofint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire ifint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [1:0] gate_0n;
  wire gfint_0n;
  wire gfint_1n;
  wire gate705_0n;
  wire gate702_0n;
  wire gate699_0n;
  assign i_1a = ifint_1n;
  INV I1 (gate705_0n, iaint_1n);
  C2RI I2 (ifint_1n, i_1r, gate705_0n, initialise);
  assign i_0a = ifint_0n;
  INV I4 (gate702_0n, iaint_0n);
  C2RI I5 (ifint_0n, i_0r, gate702_0n, initialise);
  assign oaint_0n = o_0r;
  INV I7 (gate699_0n, o_0a);
  C2RI I8 (o_0r, ofint_0n, gate699_0n, initialise);
  C2RI I9 (iaint_0n, sel_0n[0], oaint_0n, initialise);
  C2RI I10 (iaint_1n, sel_0n[1], oaint_0n, initialise);
  assign gfint_0n = ifint_0n;
  assign gfint_1n = ifint_1n;
  assign sel_0n[0] = gfint_0n;
  assign sel_0n[1] = gfint_1n;
  OR2 I15 (ofint_0n, gfint_0n, gfint_1n);
endmodule

module BrzM_0_9 (
  i_0r, i_0a,
  i_1r, i_1a,
  i_2r, i_2a,
  i_3r, i_3a,
  i_4r, i_4a,
  i_5r, i_5a,
  i_6r, i_6a,
  i_7r, i_7a,
  i_8r, i_8a,
  o_0r, o_0a,
  initialise
);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  input i_4r;
  output i_4a;
  input i_5r;
  output i_5a;
  input i_6r;
  output i_6a;
  input i_7r;
  output i_7a;
  input i_8r;
  output i_8a;
  output o_0r;
  input o_0a;
  input initialise;
  wire [2:0] internal_0n;
  wire [8:0] sel_0n;
  wire ofint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire ifint_1n;
  wire ifint_2n;
  wire ifint_3n;
  wire ifint_4n;
  wire ifint_5n;
  wire ifint_6n;
  wire ifint_7n;
  wire ifint_8n;
  wire iaint_0n;
  wire iaint_1n;
  wire iaint_2n;
  wire iaint_3n;
  wire iaint_4n;
  wire iaint_5n;
  wire iaint_6n;
  wire iaint_7n;
  wire iaint_8n;
  wire [8:0] gate_0n;
  wire gfint_0n;
  wire gfint_1n;
  wire gfint_2n;
  wire gfint_3n;
  wire gfint_4n;
  wire gfint_5n;
  wire gfint_6n;
  wire gfint_7n;
  wire gfint_8n;
  wire gate735_0n;
  wire gate732_0n;
  wire gate729_0n;
  wire gate726_0n;
  wire gate723_0n;
  wire gate720_0n;
  wire gate717_0n;
  wire gate714_0n;
  wire gate711_0n;
  wire gate708_0n;
  assign i_8a = ifint_8n;
  INV I1 (gate735_0n, iaint_8n);
  C2RI I2 (ifint_8n, i_8r, gate735_0n, initialise);
  assign i_7a = ifint_7n;
  INV I4 (gate732_0n, iaint_7n);
  C2RI I5 (ifint_7n, i_7r, gate732_0n, initialise);
  assign i_6a = ifint_6n;
  INV I7 (gate729_0n, iaint_6n);
  C2RI I8 (ifint_6n, i_6r, gate729_0n, initialise);
  assign i_5a = ifint_5n;
  INV I10 (gate726_0n, iaint_5n);
  C2RI I11 (ifint_5n, i_5r, gate726_0n, initialise);
  assign i_4a = ifint_4n;
  INV I13 (gate723_0n, iaint_4n);
  C2RI I14 (ifint_4n, i_4r, gate723_0n, initialise);
  assign i_3a = ifint_3n;
  INV I16 (gate720_0n, iaint_3n);
  C2RI I17 (ifint_3n, i_3r, gate720_0n, initialise);
  assign i_2a = ifint_2n;
  INV I19 (gate717_0n, iaint_2n);
  C2RI I20 (ifint_2n, i_2r, gate717_0n, initialise);
  assign i_1a = ifint_1n;
  INV I22 (gate714_0n, iaint_1n);
  C2RI I23 (ifint_1n, i_1r, gate714_0n, initialise);
  assign i_0a = ifint_0n;
  INV I25 (gate711_0n, iaint_0n);
  C2RI I26 (ifint_0n, i_0r, gate711_0n, initialise);
  assign oaint_0n = o_0r;
  INV I28 (gate708_0n, o_0a);
  C2RI I29 (o_0r, ofint_0n, gate708_0n, initialise);
  C2RI I30 (iaint_0n, sel_0n[0], oaint_0n, initialise);
  C2RI I31 (iaint_1n, sel_0n[1], oaint_0n, initialise);
  C2RI I32 (iaint_2n, sel_0n[2], oaint_0n, initialise);
  C2RI I33 (iaint_3n, sel_0n[3], oaint_0n, initialise);
  C2RI I34 (iaint_4n, sel_0n[4], oaint_0n, initialise);
  C2RI I35 (iaint_5n, sel_0n[5], oaint_0n, initialise);
  C2RI I36 (iaint_6n, sel_0n[6], oaint_0n, initialise);
  C2RI I37 (iaint_7n, sel_0n[7], oaint_0n, initialise);
  C2RI I38 (iaint_8n, sel_0n[8], oaint_0n, initialise);
  assign gfint_0n = ifint_0n;
  assign gfint_1n = ifint_1n;
  assign gfint_2n = ifint_2n;
  assign gfint_3n = ifint_3n;
  assign gfint_4n = ifint_4n;
  assign gfint_5n = ifint_5n;
  assign gfint_6n = ifint_6n;
  assign gfint_7n = ifint_7n;
  assign gfint_8n = ifint_8n;
  assign sel_0n[0] = gfint_0n;
  assign sel_0n[1] = gfint_1n;
  assign sel_0n[2] = gfint_2n;
  assign sel_0n[3] = gfint_3n;
  assign sel_0n[4] = gfint_4n;
  assign sel_0n[5] = gfint_5n;
  assign sel_0n[6] = gfint_6n;
  assign sel_0n[7] = gfint_7n;
  assign sel_0n[8] = gfint_8n;
  NOR3 I57 (internal_0n[0], gfint_0n, gfint_1n, gfint_2n);
  NOR3 I58 (internal_0n[1], gfint_3n, gfint_4n, gfint_5n);
  NOR3 I59 (internal_0n[2], gfint_6n, gfint_7n, gfint_8n);
  NAND3 I60 (ofint_0n, internal_0n[0], internal_0n[1], internal_0n[2]);
endmodule

module BrzM_1_2 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input i_0r0d;
  input i_0r1d;
  output i_0a;
  input i_1r0d;
  input i_1r1d;
  output i_1a;
  output o_0r0d;
  output o_0r1d;
  input o_0a;
  input initialise;
  wire [1:0] sel_0n;
  wire ofint_0n;
  wire otint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire ifint_1n;
  wire itint_0n;
  wire itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [1:0] gate_0n;
  wire gfint_0n;
  wire gfint_1n;
  wire gtint_0n;
  wire gtint_1n;
  wire complete749_0n;
  wire gate748_0n;
  wire complete745_0n;
  wire gate744_0n;
  wire complete741_0n;
  wire gate740_0n;
  wire complete737_0n;
  wire complete736_0n;
  wire selcomp_0n;
  wire selcomp_1n;
  assign i_1a = complete749_0n;
  OR2 I1 (complete749_0n, ifint_1n, itint_1n);
  INV I2 (gate748_0n, iaint_1n);
  C2RI I3 (itint_1n, i_1r1d, gate748_0n, initialise);
  C2RI I4 (ifint_1n, i_1r0d, gate748_0n, initialise);
  assign i_0a = complete745_0n;
  OR2 I6 (complete745_0n, ifint_0n, itint_0n);
  INV I7 (gate744_0n, iaint_0n);
  C2RI I8 (itint_0n, i_0r1d, gate744_0n, initialise);
  C2RI I9 (ifint_0n, i_0r0d, gate744_0n, initialise);
  assign oaint_0n = complete741_0n;
  OR2 I11 (complete741_0n, o_0r0d, o_0r1d);
  INV I12 (gate740_0n, o_0a);
  C2RI I13 (o_0r1d, otint_0n, gate740_0n, initialise);
  C2RI I14 (o_0r0d, ofint_0n, gate740_0n, initialise);
  C2RI I15 (iaint_0n, sel_0n[0], oaint_0n, initialise);
  C2RI I16 (iaint_1n, sel_0n[1], oaint_0n, initialise);
  assign gate_0n[0] = sel_0n[0];
  assign gate_0n[1] = sel_0n[1];
  assign sel_0n[0] = selcomp_0n;
  assign sel_0n[1] = selcomp_1n;
  assign selcomp_1n = complete737_0n;
  OR2 I22 (complete737_0n, ifint_1n, itint_1n);
  assign selcomp_0n = complete736_0n;
  OR2 I24 (complete736_0n, ifint_0n, itint_0n);
  AND2 I25 (gfint_0n, gate_0n[0], ifint_0n);
  AND2 I26 (gfint_1n, gate_0n[1], ifint_1n);
  AND2 I27 (gtint_0n, gate_0n[0], itint_0n);
  AND2 I28 (gtint_1n, gate_0n[1], itint_1n);
  OR2 I29 (otint_0n, gtint_0n, gtint_1n);
  OR2 I30 (ofint_0n, gfint_0n, gfint_1n);
endmodule

module BrzM_1_3 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  i_2r0d, i_2r1d, i_2a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input i_0r0d;
  input i_0r1d;
  output i_0a;
  input i_1r0d;
  input i_1r1d;
  output i_1a;
  input i_2r0d;
  input i_2r1d;
  output i_2a;
  output o_0r0d;
  output o_0r1d;
  input o_0a;
  input initialise;
  wire [2:0] sel_0n;
  wire ofint_0n;
  wire otint_0n;
  wire oaint_0n;
  wire ifint_0n;
  wire ifint_1n;
  wire ifint_2n;
  wire itint_0n;
  wire itint_1n;
  wire itint_2n;
  wire iaint_0n;
  wire iaint_1n;
  wire iaint_2n;
  wire [2:0] gate_0n;
  wire gfint_0n;
  wire gfint_1n;
  wire gfint_2n;
  wire gtint_0n;
  wire gtint_1n;
  wire gtint_2n;
  wire complete768_0n;
  wire gate767_0n;
  wire complete764_0n;
  wire gate763_0n;
  wire complete760_0n;
  wire gate759_0n;
  wire complete756_0n;
  wire gate755_0n;
  wire complete752_0n;
  wire complete751_0n;
  wire complete750_0n;
  wire selcomp_0n;
  wire selcomp_1n;
  wire selcomp_2n;
  assign i_2a = complete768_0n;
  OR2 I1 (complete768_0n, ifint_2n, itint_2n);
  INV I2 (gate767_0n, iaint_2n);
  C2RI I3 (itint_2n, i_2r1d, gate767_0n, initialise);
  C2RI I4 (ifint_2n, i_2r0d, gate767_0n, initialise);
  assign i_1a = complete764_0n;
  OR2 I6 (complete764_0n, ifint_1n, itint_1n);
  INV I7 (gate763_0n, iaint_1n);
  C2RI I8 (itint_1n, i_1r1d, gate763_0n, initialise);
  C2RI I9 (ifint_1n, i_1r0d, gate763_0n, initialise);
  assign i_0a = complete760_0n;
  OR2 I11 (complete760_0n, ifint_0n, itint_0n);
  INV I12 (gate759_0n, iaint_0n);
  C2RI I13 (itint_0n, i_0r1d, gate759_0n, initialise);
  C2RI I14 (ifint_0n, i_0r0d, gate759_0n, initialise);
  assign oaint_0n = complete756_0n;
  OR2 I16 (complete756_0n, o_0r0d, o_0r1d);
  INV I17 (gate755_0n, o_0a);
  C2RI I18 (o_0r1d, otint_0n, gate755_0n, initialise);
  C2RI I19 (o_0r0d, ofint_0n, gate755_0n, initialise);
  C2RI I20 (iaint_0n, sel_0n[0], oaint_0n, initialise);
  C2RI I21 (iaint_1n, sel_0n[1], oaint_0n, initialise);
  C2RI I22 (iaint_2n, sel_0n[2], oaint_0n, initialise);
  assign gate_0n[0] = sel_0n[0];
  assign gate_0n[1] = sel_0n[1];
  assign gate_0n[2] = sel_0n[2];
  assign sel_0n[0] = selcomp_0n;
  assign sel_0n[1] = selcomp_1n;
  assign sel_0n[2] = selcomp_2n;
  assign selcomp_2n = complete752_0n;
  OR2 I30 (complete752_0n, ifint_2n, itint_2n);
  assign selcomp_1n = complete751_0n;
  OR2 I32 (complete751_0n, ifint_1n, itint_1n);
  assign selcomp_0n = complete750_0n;
  OR2 I34 (complete750_0n, ifint_0n, itint_0n);
  AND2 I35 (gfint_0n, gate_0n[0], ifint_0n);
  AND2 I36 (gfint_1n, gate_0n[1], ifint_1n);
  AND2 I37 (gfint_2n, gate_0n[2], ifint_2n);
  AND2 I38 (gtint_0n, gate_0n[0], itint_0n);
  AND2 I39 (gtint_1n, gate_0n[1], itint_1n);
  AND2 I40 (gtint_2n, gate_0n[2], itint_2n);
  OR3 I41 (otint_0n, gtint_0n, gtint_1n, gtint_2n);
  OR3 I42 (ofint_0n, gfint_0n, gfint_1n, gfint_2n);
endmodule

module BrzM_2_2 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [1:0] i_0r0d;
  input [1:0] i_0r1d;
  output i_0a;
  input [1:0] i_1r0d;
  input [1:0] i_1r1d;
  output i_1a;
  output [1:0] o_0r0d;
  output [1:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [1:0] sel_0n;
  wire [1:0] ofint_0n;
  wire [1:0] otint_0n;
  wire oaint_0n;
  wire [1:0] ifint_0n;
  wire [1:0] ifint_1n;
  wire [1:0] itint_0n;
  wire [1:0] itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [1:0] gate_0n;
  wire [1:0] gfint_0n;
  wire [1:0] gfint_1n;
  wire [1:0] gtint_0n;
  wire [1:0] gtint_1n;
  wire [1:0] complete782_0n;
  wire gate781_0n;
  wire [1:0] complete778_0n;
  wire gate777_0n;
  wire [1:0] complete774_0n;
  wire gate773_0n;
  wire [1:0] complete770_0n;
  wire [1:0] complete769_0n;
  wire selcomp_0n;
  wire selcomp_1n;
  C2 I0 (i_1a, complete782_0n[0], complete782_0n[1]);
  OR2 I1 (complete782_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I2 (complete782_0n[1], ifint_1n[1], itint_1n[1]);
  INV I3 (gate781_0n, iaint_1n);
  C2RI I4 (itint_1n[0], i_1r1d[0], gate781_0n, initialise);
  C2RI I5 (itint_1n[1], i_1r1d[1], gate781_0n, initialise);
  C2RI I6 (ifint_1n[0], i_1r0d[0], gate781_0n, initialise);
  C2RI I7 (ifint_1n[1], i_1r0d[1], gate781_0n, initialise);
  C2 I8 (i_0a, complete778_0n[0], complete778_0n[1]);
  OR2 I9 (complete778_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I10 (complete778_0n[1], ifint_0n[1], itint_0n[1]);
  INV I11 (gate777_0n, iaint_0n);
  C2RI I12 (itint_0n[0], i_0r1d[0], gate777_0n, initialise);
  C2RI I13 (itint_0n[1], i_0r1d[1], gate777_0n, initialise);
  C2RI I14 (ifint_0n[0], i_0r0d[0], gate777_0n, initialise);
  C2RI I15 (ifint_0n[1], i_0r0d[1], gate777_0n, initialise);
  C2 I16 (oaint_0n, complete774_0n[0], complete774_0n[1]);
  OR2 I17 (complete774_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I18 (complete774_0n[1], o_0r0d[1], o_0r1d[1]);
  INV I19 (gate773_0n, o_0a);
  C2RI I20 (o_0r1d[0], otint_0n[0], gate773_0n, initialise);
  C2RI I21 (o_0r1d[1], otint_0n[1], gate773_0n, initialise);
  C2RI I22 (o_0r0d[0], ofint_0n[0], gate773_0n, initialise);
  C2RI I23 (o_0r0d[1], ofint_0n[1], gate773_0n, initialise);
  C2RI I24 (iaint_0n, sel_0n[0], oaint_0n, initialise);
  C2RI I25 (iaint_1n, sel_0n[1], oaint_0n, initialise);
  assign gate_0n[0] = sel_0n[0];
  assign gate_0n[1] = sel_0n[1];
  assign sel_0n[0] = selcomp_0n;
  assign sel_0n[1] = selcomp_1n;
  C2 I30 (selcomp_1n, complete770_0n[0], complete770_0n[1]);
  OR2 I31 (complete770_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I32 (complete770_0n[1], ifint_1n[1], itint_1n[1]);
  C2 I33 (selcomp_0n, complete769_0n[0], complete769_0n[1]);
  OR2 I34 (complete769_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I35 (complete769_0n[1], ifint_0n[1], itint_0n[1]);
  AND2 I36 (gfint_0n[0], gate_0n[0], ifint_0n[0]);
  AND2 I37 (gfint_0n[1], gate_0n[0], ifint_0n[1]);
  AND2 I38 (gfint_1n[0], gate_0n[1], ifint_1n[0]);
  AND2 I39 (gfint_1n[1], gate_0n[1], ifint_1n[1]);
  AND2 I40 (gtint_0n[0], gate_0n[0], itint_0n[0]);
  AND2 I41 (gtint_0n[1], gate_0n[0], itint_0n[1]);
  AND2 I42 (gtint_1n[0], gate_0n[1], itint_1n[0]);
  AND2 I43 (gtint_1n[1], gate_0n[1], itint_1n[1]);
  OR2 I44 (otint_0n[0], gtint_0n[0], gtint_1n[0]);
  OR2 I45 (otint_0n[1], gtint_0n[1], gtint_1n[1]);
  OR2 I46 (ofint_0n[0], gfint_0n[0], gfint_1n[0]);
  OR2 I47 (ofint_0n[1], gfint_0n[1], gfint_1n[1]);
endmodule

module BrzM_3_3 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  i_2r0d, i_2r1d, i_2a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [2:0] i_0r0d;
  input [2:0] i_0r1d;
  output i_0a;
  input [2:0] i_1r0d;
  input [2:0] i_1r1d;
  output i_1a;
  input [2:0] i_2r0d;
  input [2:0] i_2r1d;
  output i_2a;
  output [2:0] o_0r0d;
  output [2:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [2:0] sel_0n;
  wire [2:0] ofint_0n;
  wire [2:0] otint_0n;
  wire oaint_0n;
  wire [2:0] ifint_0n;
  wire [2:0] ifint_1n;
  wire [2:0] ifint_2n;
  wire [2:0] itint_0n;
  wire [2:0] itint_1n;
  wire [2:0] itint_2n;
  wire iaint_0n;
  wire iaint_1n;
  wire iaint_2n;
  wire [2:0] gate_0n;
  wire [2:0] gfint_0n;
  wire [2:0] gfint_1n;
  wire [2:0] gfint_2n;
  wire [2:0] gtint_0n;
  wire [2:0] gtint_1n;
  wire [2:0] gtint_2n;
  wire [2:0] complete801_0n;
  wire gate800_0n;
  wire [2:0] complete797_0n;
  wire gate796_0n;
  wire [2:0] complete793_0n;
  wire gate792_0n;
  wire [2:0] complete789_0n;
  wire gate788_0n;
  wire [2:0] complete785_0n;
  wire [2:0] complete784_0n;
  wire [2:0] complete783_0n;
  wire selcomp_0n;
  wire selcomp_1n;
  wire selcomp_2n;
  C3 I0 (i_2a, complete801_0n[0], complete801_0n[1], complete801_0n[2]);
  OR2 I1 (complete801_0n[0], ifint_2n[0], itint_2n[0]);
  OR2 I2 (complete801_0n[1], ifint_2n[1], itint_2n[1]);
  OR2 I3 (complete801_0n[2], ifint_2n[2], itint_2n[2]);
  INV I4 (gate800_0n, iaint_2n);
  C2RI I5 (itint_2n[0], i_2r1d[0], gate800_0n, initialise);
  C2RI I6 (itint_2n[1], i_2r1d[1], gate800_0n, initialise);
  C2RI I7 (itint_2n[2], i_2r1d[2], gate800_0n, initialise);
  C2RI I8 (ifint_2n[0], i_2r0d[0], gate800_0n, initialise);
  C2RI I9 (ifint_2n[1], i_2r0d[1], gate800_0n, initialise);
  C2RI I10 (ifint_2n[2], i_2r0d[2], gate800_0n, initialise);
  C3 I11 (i_1a, complete797_0n[0], complete797_0n[1], complete797_0n[2]);
  OR2 I12 (complete797_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I13 (complete797_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I14 (complete797_0n[2], ifint_1n[2], itint_1n[2]);
  INV I15 (gate796_0n, iaint_1n);
  C2RI I16 (itint_1n[0], i_1r1d[0], gate796_0n, initialise);
  C2RI I17 (itint_1n[1], i_1r1d[1], gate796_0n, initialise);
  C2RI I18 (itint_1n[2], i_1r1d[2], gate796_0n, initialise);
  C2RI I19 (ifint_1n[0], i_1r0d[0], gate796_0n, initialise);
  C2RI I20 (ifint_1n[1], i_1r0d[1], gate796_0n, initialise);
  C2RI I21 (ifint_1n[2], i_1r0d[2], gate796_0n, initialise);
  C3 I22 (i_0a, complete793_0n[0], complete793_0n[1], complete793_0n[2]);
  OR2 I23 (complete793_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I24 (complete793_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I25 (complete793_0n[2], ifint_0n[2], itint_0n[2]);
  INV I26 (gate792_0n, iaint_0n);
  C2RI I27 (itint_0n[0], i_0r1d[0], gate792_0n, initialise);
  C2RI I28 (itint_0n[1], i_0r1d[1], gate792_0n, initialise);
  C2RI I29 (itint_0n[2], i_0r1d[2], gate792_0n, initialise);
  C2RI I30 (ifint_0n[0], i_0r0d[0], gate792_0n, initialise);
  C2RI I31 (ifint_0n[1], i_0r0d[1], gate792_0n, initialise);
  C2RI I32 (ifint_0n[2], i_0r0d[2], gate792_0n, initialise);
  C3 I33 (oaint_0n, complete789_0n[0], complete789_0n[1], complete789_0n[2]);
  OR2 I34 (complete789_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I35 (complete789_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I36 (complete789_0n[2], o_0r0d[2], o_0r1d[2]);
  INV I37 (gate788_0n, o_0a);
  C2RI I38 (o_0r1d[0], otint_0n[0], gate788_0n, initialise);
  C2RI I39 (o_0r1d[1], otint_0n[1], gate788_0n, initialise);
  C2RI I40 (o_0r1d[2], otint_0n[2], gate788_0n, initialise);
  C2RI I41 (o_0r0d[0], ofint_0n[0], gate788_0n, initialise);
  C2RI I42 (o_0r0d[1], ofint_0n[1], gate788_0n, initialise);
  C2RI I43 (o_0r0d[2], ofint_0n[2], gate788_0n, initialise);
  C2RI I44 (iaint_0n, sel_0n[0], oaint_0n, initialise);
  C2RI I45 (iaint_1n, sel_0n[1], oaint_0n, initialise);
  C2RI I46 (iaint_2n, sel_0n[2], oaint_0n, initialise);
  assign gate_0n[0] = sel_0n[0];
  assign gate_0n[1] = sel_0n[1];
  assign gate_0n[2] = sel_0n[2];
  assign sel_0n[0] = selcomp_0n;
  assign sel_0n[1] = selcomp_1n;
  assign sel_0n[2] = selcomp_2n;
  C3 I53 (selcomp_2n, complete785_0n[0], complete785_0n[1], complete785_0n[2]);
  OR2 I54 (complete785_0n[0], ifint_2n[0], itint_2n[0]);
  OR2 I55 (complete785_0n[1], ifint_2n[1], itint_2n[1]);
  OR2 I56 (complete785_0n[2], ifint_2n[2], itint_2n[2]);
  C3 I57 (selcomp_1n, complete784_0n[0], complete784_0n[1], complete784_0n[2]);
  OR2 I58 (complete784_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I59 (complete784_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I60 (complete784_0n[2], ifint_1n[2], itint_1n[2]);
  C3 I61 (selcomp_0n, complete783_0n[0], complete783_0n[1], complete783_0n[2]);
  OR2 I62 (complete783_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I63 (complete783_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I64 (complete783_0n[2], ifint_0n[2], itint_0n[2]);
  AND2 I65 (gfint_0n[0], gate_0n[0], ifint_0n[0]);
  AND2 I66 (gfint_0n[1], gate_0n[0], ifint_0n[1]);
  AND2 I67 (gfint_0n[2], gate_0n[0], ifint_0n[2]);
  AND2 I68 (gfint_1n[0], gate_0n[1], ifint_1n[0]);
  AND2 I69 (gfint_1n[1], gate_0n[1], ifint_1n[1]);
  AND2 I70 (gfint_1n[2], gate_0n[1], ifint_1n[2]);
  AND2 I71 (gfint_2n[0], gate_0n[2], ifint_2n[0]);
  AND2 I72 (gfint_2n[1], gate_0n[2], ifint_2n[1]);
  AND2 I73 (gfint_2n[2], gate_0n[2], ifint_2n[2]);
  AND2 I74 (gtint_0n[0], gate_0n[0], itint_0n[0]);
  AND2 I75 (gtint_0n[1], gate_0n[0], itint_0n[1]);
  AND2 I76 (gtint_0n[2], gate_0n[0], itint_0n[2]);
  AND2 I77 (gtint_1n[0], gate_0n[1], itint_1n[0]);
  AND2 I78 (gtint_1n[1], gate_0n[1], itint_1n[1]);
  AND2 I79 (gtint_1n[2], gate_0n[1], itint_1n[2]);
  AND2 I80 (gtint_2n[0], gate_0n[2], itint_2n[0]);
  AND2 I81 (gtint_2n[1], gate_0n[2], itint_2n[1]);
  AND2 I82 (gtint_2n[2], gate_0n[2], itint_2n[2]);
  OR3 I83 (otint_0n[0], gtint_0n[0], gtint_1n[0], gtint_2n[0]);
  OR3 I84 (otint_0n[1], gtint_0n[1], gtint_1n[1], gtint_2n[1]);
  OR3 I85 (otint_0n[2], gtint_0n[2], gtint_1n[2], gtint_2n[2]);
  OR3 I86 (ofint_0n[0], gfint_0n[0], gfint_1n[0], gfint_2n[0]);
  OR3 I87 (ofint_0n[1], gfint_0n[1], gfint_1n[1], gfint_2n[1]);
  OR3 I88 (ofint_0n[2], gfint_0n[2], gfint_1n[2], gfint_2n[2]);
endmodule

module BrzM_9_9 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  i_2r0d, i_2r1d, i_2a,
  i_3r0d, i_3r1d, i_3a,
  i_4r0d, i_4r1d, i_4a,
  i_5r0d, i_5r1d, i_5a,
  i_6r0d, i_6r1d, i_6a,
  i_7r0d, i_7r1d, i_7a,
  i_8r0d, i_8r1d, i_8a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [8:0] i_0r0d;
  input [8:0] i_0r1d;
  output i_0a;
  input [8:0] i_1r0d;
  input [8:0] i_1r1d;
  output i_1a;
  input [8:0] i_2r0d;
  input [8:0] i_2r1d;
  output i_2a;
  input [8:0] i_3r0d;
  input [8:0] i_3r1d;
  output i_3a;
  input [8:0] i_4r0d;
  input [8:0] i_4r1d;
  output i_4a;
  input [8:0] i_5r0d;
  input [8:0] i_5r1d;
  output i_5a;
  input [8:0] i_6r0d;
  input [8:0] i_6r1d;
  output i_6a;
  input [8:0] i_7r0d;
  input [8:0] i_7r1d;
  output i_7a;
  input [8:0] i_8r0d;
  input [8:0] i_8r1d;
  output i_8a;
  output [8:0] o_0r0d;
  output [8:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [110:0] internal_0n;
  wire [8:0] sel_0n;
  wire [8:0] ofint_0n;
  wire [8:0] otint_0n;
  wire oaint_0n;
  wire [8:0] ifint_0n;
  wire [8:0] ifint_1n;
  wire [8:0] ifint_2n;
  wire [8:0] ifint_3n;
  wire [8:0] ifint_4n;
  wire [8:0] ifint_5n;
  wire [8:0] ifint_6n;
  wire [8:0] ifint_7n;
  wire [8:0] ifint_8n;
  wire [8:0] itint_0n;
  wire [8:0] itint_1n;
  wire [8:0] itint_2n;
  wire [8:0] itint_3n;
  wire [8:0] itint_4n;
  wire [8:0] itint_5n;
  wire [8:0] itint_6n;
  wire [8:0] itint_7n;
  wire [8:0] itint_8n;
  wire iaint_0n;
  wire iaint_1n;
  wire iaint_2n;
  wire iaint_3n;
  wire iaint_4n;
  wire iaint_5n;
  wire iaint_6n;
  wire iaint_7n;
  wire iaint_8n;
  wire [8:0] gate_0n;
  wire [8:0] gfint_0n;
  wire [8:0] gfint_1n;
  wire [8:0] gfint_2n;
  wire [8:0] gfint_3n;
  wire [8:0] gfint_4n;
  wire [8:0] gfint_5n;
  wire [8:0] gfint_6n;
  wire [8:0] gfint_7n;
  wire [8:0] gfint_8n;
  wire [8:0] gtint_0n;
  wire [8:0] gtint_1n;
  wire [8:0] gtint_2n;
  wire [8:0] gtint_3n;
  wire [8:0] gtint_4n;
  wire [8:0] gtint_5n;
  wire [8:0] gtint_6n;
  wire [8:0] gtint_7n;
  wire [8:0] gtint_8n;
  wire [8:0] complete850_0n;
  wire gate849_0n;
  wire [8:0] complete846_0n;
  wire gate845_0n;
  wire [8:0] complete842_0n;
  wire gate841_0n;
  wire [8:0] complete838_0n;
  wire gate837_0n;
  wire [8:0] complete834_0n;
  wire gate833_0n;
  wire [8:0] complete830_0n;
  wire gate829_0n;
  wire [8:0] complete826_0n;
  wire gate825_0n;
  wire [8:0] complete822_0n;
  wire gate821_0n;
  wire [8:0] complete818_0n;
  wire gate817_0n;
  wire [8:0] complete814_0n;
  wire gate813_0n;
  wire [8:0] complete810_0n;
  wire [8:0] complete809_0n;
  wire [8:0] complete808_0n;
  wire [8:0] complete807_0n;
  wire [8:0] complete806_0n;
  wire [8:0] complete805_0n;
  wire [8:0] complete804_0n;
  wire [8:0] complete803_0n;
  wire [8:0] complete802_0n;
  wire selcomp_0n;
  wire selcomp_1n;
  wire selcomp_2n;
  wire selcomp_3n;
  wire selcomp_4n;
  wire selcomp_5n;
  wire selcomp_6n;
  wire selcomp_7n;
  wire selcomp_8n;
  C3 I0 (internal_0n[0], complete850_0n[0], complete850_0n[1], complete850_0n[2]);
  C3 I1 (internal_0n[1], complete850_0n[3], complete850_0n[4], complete850_0n[5]);
  C3 I2 (internal_0n[2], complete850_0n[6], complete850_0n[7], complete850_0n[8]);
  C3 I3 (i_8a, internal_0n[0], internal_0n[1], internal_0n[2]);
  OR2 I4 (complete850_0n[0], ifint_8n[0], itint_8n[0]);
  OR2 I5 (complete850_0n[1], ifint_8n[1], itint_8n[1]);
  OR2 I6 (complete850_0n[2], ifint_8n[2], itint_8n[2]);
  OR2 I7 (complete850_0n[3], ifint_8n[3], itint_8n[3]);
  OR2 I8 (complete850_0n[4], ifint_8n[4], itint_8n[4]);
  OR2 I9 (complete850_0n[5], ifint_8n[5], itint_8n[5]);
  OR2 I10 (complete850_0n[6], ifint_8n[6], itint_8n[6]);
  OR2 I11 (complete850_0n[7], ifint_8n[7], itint_8n[7]);
  OR2 I12 (complete850_0n[8], ifint_8n[8], itint_8n[8]);
  INV I13 (gate849_0n, iaint_8n);
  C2RI I14 (itint_8n[0], i_8r1d[0], gate849_0n, initialise);
  C2RI I15 (itint_8n[1], i_8r1d[1], gate849_0n, initialise);
  C2RI I16 (itint_8n[2], i_8r1d[2], gate849_0n, initialise);
  C2RI I17 (itint_8n[3], i_8r1d[3], gate849_0n, initialise);
  C2RI I18 (itint_8n[4], i_8r1d[4], gate849_0n, initialise);
  C2RI I19 (itint_8n[5], i_8r1d[5], gate849_0n, initialise);
  C2RI I20 (itint_8n[6], i_8r1d[6], gate849_0n, initialise);
  C2RI I21 (itint_8n[7], i_8r1d[7], gate849_0n, initialise);
  C2RI I22 (itint_8n[8], i_8r1d[8], gate849_0n, initialise);
  C2RI I23 (ifint_8n[0], i_8r0d[0], gate849_0n, initialise);
  C2RI I24 (ifint_8n[1], i_8r0d[1], gate849_0n, initialise);
  C2RI I25 (ifint_8n[2], i_8r0d[2], gate849_0n, initialise);
  C2RI I26 (ifint_8n[3], i_8r0d[3], gate849_0n, initialise);
  C2RI I27 (ifint_8n[4], i_8r0d[4], gate849_0n, initialise);
  C2RI I28 (ifint_8n[5], i_8r0d[5], gate849_0n, initialise);
  C2RI I29 (ifint_8n[6], i_8r0d[6], gate849_0n, initialise);
  C2RI I30 (ifint_8n[7], i_8r0d[7], gate849_0n, initialise);
  C2RI I31 (ifint_8n[8], i_8r0d[8], gate849_0n, initialise);
  C3 I32 (internal_0n[3], complete846_0n[0], complete846_0n[1], complete846_0n[2]);
  C3 I33 (internal_0n[4], complete846_0n[3], complete846_0n[4], complete846_0n[5]);
  C3 I34 (internal_0n[5], complete846_0n[6], complete846_0n[7], complete846_0n[8]);
  C3 I35 (i_7a, internal_0n[3], internal_0n[4], internal_0n[5]);
  OR2 I36 (complete846_0n[0], ifint_7n[0], itint_7n[0]);
  OR2 I37 (complete846_0n[1], ifint_7n[1], itint_7n[1]);
  OR2 I38 (complete846_0n[2], ifint_7n[2], itint_7n[2]);
  OR2 I39 (complete846_0n[3], ifint_7n[3], itint_7n[3]);
  OR2 I40 (complete846_0n[4], ifint_7n[4], itint_7n[4]);
  OR2 I41 (complete846_0n[5], ifint_7n[5], itint_7n[5]);
  OR2 I42 (complete846_0n[6], ifint_7n[6], itint_7n[6]);
  OR2 I43 (complete846_0n[7], ifint_7n[7], itint_7n[7]);
  OR2 I44 (complete846_0n[8], ifint_7n[8], itint_7n[8]);
  INV I45 (gate845_0n, iaint_7n);
  C2RI I46 (itint_7n[0], i_7r1d[0], gate845_0n, initialise);
  C2RI I47 (itint_7n[1], i_7r1d[1], gate845_0n, initialise);
  C2RI I48 (itint_7n[2], i_7r1d[2], gate845_0n, initialise);
  C2RI I49 (itint_7n[3], i_7r1d[3], gate845_0n, initialise);
  C2RI I50 (itint_7n[4], i_7r1d[4], gate845_0n, initialise);
  C2RI I51 (itint_7n[5], i_7r1d[5], gate845_0n, initialise);
  C2RI I52 (itint_7n[6], i_7r1d[6], gate845_0n, initialise);
  C2RI I53 (itint_7n[7], i_7r1d[7], gate845_0n, initialise);
  C2RI I54 (itint_7n[8], i_7r1d[8], gate845_0n, initialise);
  C2RI I55 (ifint_7n[0], i_7r0d[0], gate845_0n, initialise);
  C2RI I56 (ifint_7n[1], i_7r0d[1], gate845_0n, initialise);
  C2RI I57 (ifint_7n[2], i_7r0d[2], gate845_0n, initialise);
  C2RI I58 (ifint_7n[3], i_7r0d[3], gate845_0n, initialise);
  C2RI I59 (ifint_7n[4], i_7r0d[4], gate845_0n, initialise);
  C2RI I60 (ifint_7n[5], i_7r0d[5], gate845_0n, initialise);
  C2RI I61 (ifint_7n[6], i_7r0d[6], gate845_0n, initialise);
  C2RI I62 (ifint_7n[7], i_7r0d[7], gate845_0n, initialise);
  C2RI I63 (ifint_7n[8], i_7r0d[8], gate845_0n, initialise);
  C3 I64 (internal_0n[6], complete842_0n[0], complete842_0n[1], complete842_0n[2]);
  C3 I65 (internal_0n[7], complete842_0n[3], complete842_0n[4], complete842_0n[5]);
  C3 I66 (internal_0n[8], complete842_0n[6], complete842_0n[7], complete842_0n[8]);
  C3 I67 (i_6a, internal_0n[6], internal_0n[7], internal_0n[8]);
  OR2 I68 (complete842_0n[0], ifint_6n[0], itint_6n[0]);
  OR2 I69 (complete842_0n[1], ifint_6n[1], itint_6n[1]);
  OR2 I70 (complete842_0n[2], ifint_6n[2], itint_6n[2]);
  OR2 I71 (complete842_0n[3], ifint_6n[3], itint_6n[3]);
  OR2 I72 (complete842_0n[4], ifint_6n[4], itint_6n[4]);
  OR2 I73 (complete842_0n[5], ifint_6n[5], itint_6n[5]);
  OR2 I74 (complete842_0n[6], ifint_6n[6], itint_6n[6]);
  OR2 I75 (complete842_0n[7], ifint_6n[7], itint_6n[7]);
  OR2 I76 (complete842_0n[8], ifint_6n[8], itint_6n[8]);
  INV I77 (gate841_0n, iaint_6n);
  C2RI I78 (itint_6n[0], i_6r1d[0], gate841_0n, initialise);
  C2RI I79 (itint_6n[1], i_6r1d[1], gate841_0n, initialise);
  C2RI I80 (itint_6n[2], i_6r1d[2], gate841_0n, initialise);
  C2RI I81 (itint_6n[3], i_6r1d[3], gate841_0n, initialise);
  C2RI I82 (itint_6n[4], i_6r1d[4], gate841_0n, initialise);
  C2RI I83 (itint_6n[5], i_6r1d[5], gate841_0n, initialise);
  C2RI I84 (itint_6n[6], i_6r1d[6], gate841_0n, initialise);
  C2RI I85 (itint_6n[7], i_6r1d[7], gate841_0n, initialise);
  C2RI I86 (itint_6n[8], i_6r1d[8], gate841_0n, initialise);
  C2RI I87 (ifint_6n[0], i_6r0d[0], gate841_0n, initialise);
  C2RI I88 (ifint_6n[1], i_6r0d[1], gate841_0n, initialise);
  C2RI I89 (ifint_6n[2], i_6r0d[2], gate841_0n, initialise);
  C2RI I90 (ifint_6n[3], i_6r0d[3], gate841_0n, initialise);
  C2RI I91 (ifint_6n[4], i_6r0d[4], gate841_0n, initialise);
  C2RI I92 (ifint_6n[5], i_6r0d[5], gate841_0n, initialise);
  C2RI I93 (ifint_6n[6], i_6r0d[6], gate841_0n, initialise);
  C2RI I94 (ifint_6n[7], i_6r0d[7], gate841_0n, initialise);
  C2RI I95 (ifint_6n[8], i_6r0d[8], gate841_0n, initialise);
  C3 I96 (internal_0n[9], complete838_0n[0], complete838_0n[1], complete838_0n[2]);
  C3 I97 (internal_0n[10], complete838_0n[3], complete838_0n[4], complete838_0n[5]);
  C3 I98 (internal_0n[11], complete838_0n[6], complete838_0n[7], complete838_0n[8]);
  C3 I99 (i_5a, internal_0n[9], internal_0n[10], internal_0n[11]);
  OR2 I100 (complete838_0n[0], ifint_5n[0], itint_5n[0]);
  OR2 I101 (complete838_0n[1], ifint_5n[1], itint_5n[1]);
  OR2 I102 (complete838_0n[2], ifint_5n[2], itint_5n[2]);
  OR2 I103 (complete838_0n[3], ifint_5n[3], itint_5n[3]);
  OR2 I104 (complete838_0n[4], ifint_5n[4], itint_5n[4]);
  OR2 I105 (complete838_0n[5], ifint_5n[5], itint_5n[5]);
  OR2 I106 (complete838_0n[6], ifint_5n[6], itint_5n[6]);
  OR2 I107 (complete838_0n[7], ifint_5n[7], itint_5n[7]);
  OR2 I108 (complete838_0n[8], ifint_5n[8], itint_5n[8]);
  INV I109 (gate837_0n, iaint_5n);
  C2RI I110 (itint_5n[0], i_5r1d[0], gate837_0n, initialise);
  C2RI I111 (itint_5n[1], i_5r1d[1], gate837_0n, initialise);
  C2RI I112 (itint_5n[2], i_5r1d[2], gate837_0n, initialise);
  C2RI I113 (itint_5n[3], i_5r1d[3], gate837_0n, initialise);
  C2RI I114 (itint_5n[4], i_5r1d[4], gate837_0n, initialise);
  C2RI I115 (itint_5n[5], i_5r1d[5], gate837_0n, initialise);
  C2RI I116 (itint_5n[6], i_5r1d[6], gate837_0n, initialise);
  C2RI I117 (itint_5n[7], i_5r1d[7], gate837_0n, initialise);
  C2RI I118 (itint_5n[8], i_5r1d[8], gate837_0n, initialise);
  C2RI I119 (ifint_5n[0], i_5r0d[0], gate837_0n, initialise);
  C2RI I120 (ifint_5n[1], i_5r0d[1], gate837_0n, initialise);
  C2RI I121 (ifint_5n[2], i_5r0d[2], gate837_0n, initialise);
  C2RI I122 (ifint_5n[3], i_5r0d[3], gate837_0n, initialise);
  C2RI I123 (ifint_5n[4], i_5r0d[4], gate837_0n, initialise);
  C2RI I124 (ifint_5n[5], i_5r0d[5], gate837_0n, initialise);
  C2RI I125 (ifint_5n[6], i_5r0d[6], gate837_0n, initialise);
  C2RI I126 (ifint_5n[7], i_5r0d[7], gate837_0n, initialise);
  C2RI I127 (ifint_5n[8], i_5r0d[8], gate837_0n, initialise);
  C3 I128 (internal_0n[12], complete834_0n[0], complete834_0n[1], complete834_0n[2]);
  C3 I129 (internal_0n[13], complete834_0n[3], complete834_0n[4], complete834_0n[5]);
  C3 I130 (internal_0n[14], complete834_0n[6], complete834_0n[7], complete834_0n[8]);
  C3 I131 (i_4a, internal_0n[12], internal_0n[13], internal_0n[14]);
  OR2 I132 (complete834_0n[0], ifint_4n[0], itint_4n[0]);
  OR2 I133 (complete834_0n[1], ifint_4n[1], itint_4n[1]);
  OR2 I134 (complete834_0n[2], ifint_4n[2], itint_4n[2]);
  OR2 I135 (complete834_0n[3], ifint_4n[3], itint_4n[3]);
  OR2 I136 (complete834_0n[4], ifint_4n[4], itint_4n[4]);
  OR2 I137 (complete834_0n[5], ifint_4n[5], itint_4n[5]);
  OR2 I138 (complete834_0n[6], ifint_4n[6], itint_4n[6]);
  OR2 I139 (complete834_0n[7], ifint_4n[7], itint_4n[7]);
  OR2 I140 (complete834_0n[8], ifint_4n[8], itint_4n[8]);
  INV I141 (gate833_0n, iaint_4n);
  C2RI I142 (itint_4n[0], i_4r1d[0], gate833_0n, initialise);
  C2RI I143 (itint_4n[1], i_4r1d[1], gate833_0n, initialise);
  C2RI I144 (itint_4n[2], i_4r1d[2], gate833_0n, initialise);
  C2RI I145 (itint_4n[3], i_4r1d[3], gate833_0n, initialise);
  C2RI I146 (itint_4n[4], i_4r1d[4], gate833_0n, initialise);
  C2RI I147 (itint_4n[5], i_4r1d[5], gate833_0n, initialise);
  C2RI I148 (itint_4n[6], i_4r1d[6], gate833_0n, initialise);
  C2RI I149 (itint_4n[7], i_4r1d[7], gate833_0n, initialise);
  C2RI I150 (itint_4n[8], i_4r1d[8], gate833_0n, initialise);
  C2RI I151 (ifint_4n[0], i_4r0d[0], gate833_0n, initialise);
  C2RI I152 (ifint_4n[1], i_4r0d[1], gate833_0n, initialise);
  C2RI I153 (ifint_4n[2], i_4r0d[2], gate833_0n, initialise);
  C2RI I154 (ifint_4n[3], i_4r0d[3], gate833_0n, initialise);
  C2RI I155 (ifint_4n[4], i_4r0d[4], gate833_0n, initialise);
  C2RI I156 (ifint_4n[5], i_4r0d[5], gate833_0n, initialise);
  C2RI I157 (ifint_4n[6], i_4r0d[6], gate833_0n, initialise);
  C2RI I158 (ifint_4n[7], i_4r0d[7], gate833_0n, initialise);
  C2RI I159 (ifint_4n[8], i_4r0d[8], gate833_0n, initialise);
  C3 I160 (internal_0n[15], complete830_0n[0], complete830_0n[1], complete830_0n[2]);
  C3 I161 (internal_0n[16], complete830_0n[3], complete830_0n[4], complete830_0n[5]);
  C3 I162 (internal_0n[17], complete830_0n[6], complete830_0n[7], complete830_0n[8]);
  C3 I163 (i_3a, internal_0n[15], internal_0n[16], internal_0n[17]);
  OR2 I164 (complete830_0n[0], ifint_3n[0], itint_3n[0]);
  OR2 I165 (complete830_0n[1], ifint_3n[1], itint_3n[1]);
  OR2 I166 (complete830_0n[2], ifint_3n[2], itint_3n[2]);
  OR2 I167 (complete830_0n[3], ifint_3n[3], itint_3n[3]);
  OR2 I168 (complete830_0n[4], ifint_3n[4], itint_3n[4]);
  OR2 I169 (complete830_0n[5], ifint_3n[5], itint_3n[5]);
  OR2 I170 (complete830_0n[6], ifint_3n[6], itint_3n[6]);
  OR2 I171 (complete830_0n[7], ifint_3n[7], itint_3n[7]);
  OR2 I172 (complete830_0n[8], ifint_3n[8], itint_3n[8]);
  INV I173 (gate829_0n, iaint_3n);
  C2RI I174 (itint_3n[0], i_3r1d[0], gate829_0n, initialise);
  C2RI I175 (itint_3n[1], i_3r1d[1], gate829_0n, initialise);
  C2RI I176 (itint_3n[2], i_3r1d[2], gate829_0n, initialise);
  C2RI I177 (itint_3n[3], i_3r1d[3], gate829_0n, initialise);
  C2RI I178 (itint_3n[4], i_3r1d[4], gate829_0n, initialise);
  C2RI I179 (itint_3n[5], i_3r1d[5], gate829_0n, initialise);
  C2RI I180 (itint_3n[6], i_3r1d[6], gate829_0n, initialise);
  C2RI I181 (itint_3n[7], i_3r1d[7], gate829_0n, initialise);
  C2RI I182 (itint_3n[8], i_3r1d[8], gate829_0n, initialise);
  C2RI I183 (ifint_3n[0], i_3r0d[0], gate829_0n, initialise);
  C2RI I184 (ifint_3n[1], i_3r0d[1], gate829_0n, initialise);
  C2RI I185 (ifint_3n[2], i_3r0d[2], gate829_0n, initialise);
  C2RI I186 (ifint_3n[3], i_3r0d[3], gate829_0n, initialise);
  C2RI I187 (ifint_3n[4], i_3r0d[4], gate829_0n, initialise);
  C2RI I188 (ifint_3n[5], i_3r0d[5], gate829_0n, initialise);
  C2RI I189 (ifint_3n[6], i_3r0d[6], gate829_0n, initialise);
  C2RI I190 (ifint_3n[7], i_3r0d[7], gate829_0n, initialise);
  C2RI I191 (ifint_3n[8], i_3r0d[8], gate829_0n, initialise);
  C3 I192 (internal_0n[18], complete826_0n[0], complete826_0n[1], complete826_0n[2]);
  C3 I193 (internal_0n[19], complete826_0n[3], complete826_0n[4], complete826_0n[5]);
  C3 I194 (internal_0n[20], complete826_0n[6], complete826_0n[7], complete826_0n[8]);
  C3 I195 (i_2a, internal_0n[18], internal_0n[19], internal_0n[20]);
  OR2 I196 (complete826_0n[0], ifint_2n[0], itint_2n[0]);
  OR2 I197 (complete826_0n[1], ifint_2n[1], itint_2n[1]);
  OR2 I198 (complete826_0n[2], ifint_2n[2], itint_2n[2]);
  OR2 I199 (complete826_0n[3], ifint_2n[3], itint_2n[3]);
  OR2 I200 (complete826_0n[4], ifint_2n[4], itint_2n[4]);
  OR2 I201 (complete826_0n[5], ifint_2n[5], itint_2n[5]);
  OR2 I202 (complete826_0n[6], ifint_2n[6], itint_2n[6]);
  OR2 I203 (complete826_0n[7], ifint_2n[7], itint_2n[7]);
  OR2 I204 (complete826_0n[8], ifint_2n[8], itint_2n[8]);
  INV I205 (gate825_0n, iaint_2n);
  C2RI I206 (itint_2n[0], i_2r1d[0], gate825_0n, initialise);
  C2RI I207 (itint_2n[1], i_2r1d[1], gate825_0n, initialise);
  C2RI I208 (itint_2n[2], i_2r1d[2], gate825_0n, initialise);
  C2RI I209 (itint_2n[3], i_2r1d[3], gate825_0n, initialise);
  C2RI I210 (itint_2n[4], i_2r1d[4], gate825_0n, initialise);
  C2RI I211 (itint_2n[5], i_2r1d[5], gate825_0n, initialise);
  C2RI I212 (itint_2n[6], i_2r1d[6], gate825_0n, initialise);
  C2RI I213 (itint_2n[7], i_2r1d[7], gate825_0n, initialise);
  C2RI I214 (itint_2n[8], i_2r1d[8], gate825_0n, initialise);
  C2RI I215 (ifint_2n[0], i_2r0d[0], gate825_0n, initialise);
  C2RI I216 (ifint_2n[1], i_2r0d[1], gate825_0n, initialise);
  C2RI I217 (ifint_2n[2], i_2r0d[2], gate825_0n, initialise);
  C2RI I218 (ifint_2n[3], i_2r0d[3], gate825_0n, initialise);
  C2RI I219 (ifint_2n[4], i_2r0d[4], gate825_0n, initialise);
  C2RI I220 (ifint_2n[5], i_2r0d[5], gate825_0n, initialise);
  C2RI I221 (ifint_2n[6], i_2r0d[6], gate825_0n, initialise);
  C2RI I222 (ifint_2n[7], i_2r0d[7], gate825_0n, initialise);
  C2RI I223 (ifint_2n[8], i_2r0d[8], gate825_0n, initialise);
  C3 I224 (internal_0n[21], complete822_0n[0], complete822_0n[1], complete822_0n[2]);
  C3 I225 (internal_0n[22], complete822_0n[3], complete822_0n[4], complete822_0n[5]);
  C3 I226 (internal_0n[23], complete822_0n[6], complete822_0n[7], complete822_0n[8]);
  C3 I227 (i_1a, internal_0n[21], internal_0n[22], internal_0n[23]);
  OR2 I228 (complete822_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I229 (complete822_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I230 (complete822_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I231 (complete822_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I232 (complete822_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I233 (complete822_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I234 (complete822_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I235 (complete822_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I236 (complete822_0n[8], ifint_1n[8], itint_1n[8]);
  INV I237 (gate821_0n, iaint_1n);
  C2RI I238 (itint_1n[0], i_1r1d[0], gate821_0n, initialise);
  C2RI I239 (itint_1n[1], i_1r1d[1], gate821_0n, initialise);
  C2RI I240 (itint_1n[2], i_1r1d[2], gate821_0n, initialise);
  C2RI I241 (itint_1n[3], i_1r1d[3], gate821_0n, initialise);
  C2RI I242 (itint_1n[4], i_1r1d[4], gate821_0n, initialise);
  C2RI I243 (itint_1n[5], i_1r1d[5], gate821_0n, initialise);
  C2RI I244 (itint_1n[6], i_1r1d[6], gate821_0n, initialise);
  C2RI I245 (itint_1n[7], i_1r1d[7], gate821_0n, initialise);
  C2RI I246 (itint_1n[8], i_1r1d[8], gate821_0n, initialise);
  C2RI I247 (ifint_1n[0], i_1r0d[0], gate821_0n, initialise);
  C2RI I248 (ifint_1n[1], i_1r0d[1], gate821_0n, initialise);
  C2RI I249 (ifint_1n[2], i_1r0d[2], gate821_0n, initialise);
  C2RI I250 (ifint_1n[3], i_1r0d[3], gate821_0n, initialise);
  C2RI I251 (ifint_1n[4], i_1r0d[4], gate821_0n, initialise);
  C2RI I252 (ifint_1n[5], i_1r0d[5], gate821_0n, initialise);
  C2RI I253 (ifint_1n[6], i_1r0d[6], gate821_0n, initialise);
  C2RI I254 (ifint_1n[7], i_1r0d[7], gate821_0n, initialise);
  C2RI I255 (ifint_1n[8], i_1r0d[8], gate821_0n, initialise);
  C3 I256 (internal_0n[24], complete818_0n[0], complete818_0n[1], complete818_0n[2]);
  C3 I257 (internal_0n[25], complete818_0n[3], complete818_0n[4], complete818_0n[5]);
  C3 I258 (internal_0n[26], complete818_0n[6], complete818_0n[7], complete818_0n[8]);
  C3 I259 (i_0a, internal_0n[24], internal_0n[25], internal_0n[26]);
  OR2 I260 (complete818_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I261 (complete818_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I262 (complete818_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I263 (complete818_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I264 (complete818_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I265 (complete818_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I266 (complete818_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I267 (complete818_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I268 (complete818_0n[8], ifint_0n[8], itint_0n[8]);
  INV I269 (gate817_0n, iaint_0n);
  C2RI I270 (itint_0n[0], i_0r1d[0], gate817_0n, initialise);
  C2RI I271 (itint_0n[1], i_0r1d[1], gate817_0n, initialise);
  C2RI I272 (itint_0n[2], i_0r1d[2], gate817_0n, initialise);
  C2RI I273 (itint_0n[3], i_0r1d[3], gate817_0n, initialise);
  C2RI I274 (itint_0n[4], i_0r1d[4], gate817_0n, initialise);
  C2RI I275 (itint_0n[5], i_0r1d[5], gate817_0n, initialise);
  C2RI I276 (itint_0n[6], i_0r1d[6], gate817_0n, initialise);
  C2RI I277 (itint_0n[7], i_0r1d[7], gate817_0n, initialise);
  C2RI I278 (itint_0n[8], i_0r1d[8], gate817_0n, initialise);
  C2RI I279 (ifint_0n[0], i_0r0d[0], gate817_0n, initialise);
  C2RI I280 (ifint_0n[1], i_0r0d[1], gate817_0n, initialise);
  C2RI I281 (ifint_0n[2], i_0r0d[2], gate817_0n, initialise);
  C2RI I282 (ifint_0n[3], i_0r0d[3], gate817_0n, initialise);
  C2RI I283 (ifint_0n[4], i_0r0d[4], gate817_0n, initialise);
  C2RI I284 (ifint_0n[5], i_0r0d[5], gate817_0n, initialise);
  C2RI I285 (ifint_0n[6], i_0r0d[6], gate817_0n, initialise);
  C2RI I286 (ifint_0n[7], i_0r0d[7], gate817_0n, initialise);
  C2RI I287 (ifint_0n[8], i_0r0d[8], gate817_0n, initialise);
  C3 I288 (internal_0n[27], complete814_0n[0], complete814_0n[1], complete814_0n[2]);
  C3 I289 (internal_0n[28], complete814_0n[3], complete814_0n[4], complete814_0n[5]);
  C3 I290 (internal_0n[29], complete814_0n[6], complete814_0n[7], complete814_0n[8]);
  C3 I291 (oaint_0n, internal_0n[27], internal_0n[28], internal_0n[29]);
  OR2 I292 (complete814_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I293 (complete814_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I294 (complete814_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I295 (complete814_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I296 (complete814_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I297 (complete814_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I298 (complete814_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I299 (complete814_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I300 (complete814_0n[8], o_0r0d[8], o_0r1d[8]);
  INV I301 (gate813_0n, o_0a);
  C2RI I302 (o_0r1d[0], otint_0n[0], gate813_0n, initialise);
  C2RI I303 (o_0r1d[1], otint_0n[1], gate813_0n, initialise);
  C2RI I304 (o_0r1d[2], otint_0n[2], gate813_0n, initialise);
  C2RI I305 (o_0r1d[3], otint_0n[3], gate813_0n, initialise);
  C2RI I306 (o_0r1d[4], otint_0n[4], gate813_0n, initialise);
  C2RI I307 (o_0r1d[5], otint_0n[5], gate813_0n, initialise);
  C2RI I308 (o_0r1d[6], otint_0n[6], gate813_0n, initialise);
  C2RI I309 (o_0r1d[7], otint_0n[7], gate813_0n, initialise);
  C2RI I310 (o_0r1d[8], otint_0n[8], gate813_0n, initialise);
  C2RI I311 (o_0r0d[0], ofint_0n[0], gate813_0n, initialise);
  C2RI I312 (o_0r0d[1], ofint_0n[1], gate813_0n, initialise);
  C2RI I313 (o_0r0d[2], ofint_0n[2], gate813_0n, initialise);
  C2RI I314 (o_0r0d[3], ofint_0n[3], gate813_0n, initialise);
  C2RI I315 (o_0r0d[4], ofint_0n[4], gate813_0n, initialise);
  C2RI I316 (o_0r0d[5], ofint_0n[5], gate813_0n, initialise);
  C2RI I317 (o_0r0d[6], ofint_0n[6], gate813_0n, initialise);
  C2RI I318 (o_0r0d[7], ofint_0n[7], gate813_0n, initialise);
  C2RI I319 (o_0r0d[8], ofint_0n[8], gate813_0n, initialise);
  C2RI I320 (iaint_0n, sel_0n[0], oaint_0n, initialise);
  C2RI I321 (iaint_1n, sel_0n[1], oaint_0n, initialise);
  C2RI I322 (iaint_2n, sel_0n[2], oaint_0n, initialise);
  C2RI I323 (iaint_3n, sel_0n[3], oaint_0n, initialise);
  C2RI I324 (iaint_4n, sel_0n[4], oaint_0n, initialise);
  C2RI I325 (iaint_5n, sel_0n[5], oaint_0n, initialise);
  C2RI I326 (iaint_6n, sel_0n[6], oaint_0n, initialise);
  C2RI I327 (iaint_7n, sel_0n[7], oaint_0n, initialise);
  C2RI I328 (iaint_8n, sel_0n[8], oaint_0n, initialise);
  assign gate_0n[0] = sel_0n[0];
  assign gate_0n[1] = sel_0n[1];
  assign gate_0n[2] = sel_0n[2];
  assign gate_0n[3] = sel_0n[3];
  assign gate_0n[4] = sel_0n[4];
  assign gate_0n[5] = sel_0n[5];
  assign gate_0n[6] = sel_0n[6];
  assign gate_0n[7] = sel_0n[7];
  assign gate_0n[8] = sel_0n[8];
  assign sel_0n[0] = selcomp_0n;
  assign sel_0n[1] = selcomp_1n;
  assign sel_0n[2] = selcomp_2n;
  assign sel_0n[3] = selcomp_3n;
  assign sel_0n[4] = selcomp_4n;
  assign sel_0n[5] = selcomp_5n;
  assign sel_0n[6] = selcomp_6n;
  assign sel_0n[7] = selcomp_7n;
  assign sel_0n[8] = selcomp_8n;
  C3 I347 (internal_0n[30], complete810_0n[0], complete810_0n[1], complete810_0n[2]);
  C3 I348 (internal_0n[31], complete810_0n[3], complete810_0n[4], complete810_0n[5]);
  C3 I349 (internal_0n[32], complete810_0n[6], complete810_0n[7], complete810_0n[8]);
  C3 I350 (selcomp_8n, internal_0n[30], internal_0n[31], internal_0n[32]);
  OR2 I351 (complete810_0n[0], ifint_8n[0], itint_8n[0]);
  OR2 I352 (complete810_0n[1], ifint_8n[1], itint_8n[1]);
  OR2 I353 (complete810_0n[2], ifint_8n[2], itint_8n[2]);
  OR2 I354 (complete810_0n[3], ifint_8n[3], itint_8n[3]);
  OR2 I355 (complete810_0n[4], ifint_8n[4], itint_8n[4]);
  OR2 I356 (complete810_0n[5], ifint_8n[5], itint_8n[5]);
  OR2 I357 (complete810_0n[6], ifint_8n[6], itint_8n[6]);
  OR2 I358 (complete810_0n[7], ifint_8n[7], itint_8n[7]);
  OR2 I359 (complete810_0n[8], ifint_8n[8], itint_8n[8]);
  C3 I360 (internal_0n[33], complete809_0n[0], complete809_0n[1], complete809_0n[2]);
  C3 I361 (internal_0n[34], complete809_0n[3], complete809_0n[4], complete809_0n[5]);
  C3 I362 (internal_0n[35], complete809_0n[6], complete809_0n[7], complete809_0n[8]);
  C3 I363 (selcomp_7n, internal_0n[33], internal_0n[34], internal_0n[35]);
  OR2 I364 (complete809_0n[0], ifint_7n[0], itint_7n[0]);
  OR2 I365 (complete809_0n[1], ifint_7n[1], itint_7n[1]);
  OR2 I366 (complete809_0n[2], ifint_7n[2], itint_7n[2]);
  OR2 I367 (complete809_0n[3], ifint_7n[3], itint_7n[3]);
  OR2 I368 (complete809_0n[4], ifint_7n[4], itint_7n[4]);
  OR2 I369 (complete809_0n[5], ifint_7n[5], itint_7n[5]);
  OR2 I370 (complete809_0n[6], ifint_7n[6], itint_7n[6]);
  OR2 I371 (complete809_0n[7], ifint_7n[7], itint_7n[7]);
  OR2 I372 (complete809_0n[8], ifint_7n[8], itint_7n[8]);
  C3 I373 (internal_0n[36], complete808_0n[0], complete808_0n[1], complete808_0n[2]);
  C3 I374 (internal_0n[37], complete808_0n[3], complete808_0n[4], complete808_0n[5]);
  C3 I375 (internal_0n[38], complete808_0n[6], complete808_0n[7], complete808_0n[8]);
  C3 I376 (selcomp_6n, internal_0n[36], internal_0n[37], internal_0n[38]);
  OR2 I377 (complete808_0n[0], ifint_6n[0], itint_6n[0]);
  OR2 I378 (complete808_0n[1], ifint_6n[1], itint_6n[1]);
  OR2 I379 (complete808_0n[2], ifint_6n[2], itint_6n[2]);
  OR2 I380 (complete808_0n[3], ifint_6n[3], itint_6n[3]);
  OR2 I381 (complete808_0n[4], ifint_6n[4], itint_6n[4]);
  OR2 I382 (complete808_0n[5], ifint_6n[5], itint_6n[5]);
  OR2 I383 (complete808_0n[6], ifint_6n[6], itint_6n[6]);
  OR2 I384 (complete808_0n[7], ifint_6n[7], itint_6n[7]);
  OR2 I385 (complete808_0n[8], ifint_6n[8], itint_6n[8]);
  C3 I386 (internal_0n[39], complete807_0n[0], complete807_0n[1], complete807_0n[2]);
  C3 I387 (internal_0n[40], complete807_0n[3], complete807_0n[4], complete807_0n[5]);
  C3 I388 (internal_0n[41], complete807_0n[6], complete807_0n[7], complete807_0n[8]);
  C3 I389 (selcomp_5n, internal_0n[39], internal_0n[40], internal_0n[41]);
  OR2 I390 (complete807_0n[0], ifint_5n[0], itint_5n[0]);
  OR2 I391 (complete807_0n[1], ifint_5n[1], itint_5n[1]);
  OR2 I392 (complete807_0n[2], ifint_5n[2], itint_5n[2]);
  OR2 I393 (complete807_0n[3], ifint_5n[3], itint_5n[3]);
  OR2 I394 (complete807_0n[4], ifint_5n[4], itint_5n[4]);
  OR2 I395 (complete807_0n[5], ifint_5n[5], itint_5n[5]);
  OR2 I396 (complete807_0n[6], ifint_5n[6], itint_5n[6]);
  OR2 I397 (complete807_0n[7], ifint_5n[7], itint_5n[7]);
  OR2 I398 (complete807_0n[8], ifint_5n[8], itint_5n[8]);
  C3 I399 (internal_0n[42], complete806_0n[0], complete806_0n[1], complete806_0n[2]);
  C3 I400 (internal_0n[43], complete806_0n[3], complete806_0n[4], complete806_0n[5]);
  C3 I401 (internal_0n[44], complete806_0n[6], complete806_0n[7], complete806_0n[8]);
  C3 I402 (selcomp_4n, internal_0n[42], internal_0n[43], internal_0n[44]);
  OR2 I403 (complete806_0n[0], ifint_4n[0], itint_4n[0]);
  OR2 I404 (complete806_0n[1], ifint_4n[1], itint_4n[1]);
  OR2 I405 (complete806_0n[2], ifint_4n[2], itint_4n[2]);
  OR2 I406 (complete806_0n[3], ifint_4n[3], itint_4n[3]);
  OR2 I407 (complete806_0n[4], ifint_4n[4], itint_4n[4]);
  OR2 I408 (complete806_0n[5], ifint_4n[5], itint_4n[5]);
  OR2 I409 (complete806_0n[6], ifint_4n[6], itint_4n[6]);
  OR2 I410 (complete806_0n[7], ifint_4n[7], itint_4n[7]);
  OR2 I411 (complete806_0n[8], ifint_4n[8], itint_4n[8]);
  C3 I412 (internal_0n[45], complete805_0n[0], complete805_0n[1], complete805_0n[2]);
  C3 I413 (internal_0n[46], complete805_0n[3], complete805_0n[4], complete805_0n[5]);
  C3 I414 (internal_0n[47], complete805_0n[6], complete805_0n[7], complete805_0n[8]);
  C3 I415 (selcomp_3n, internal_0n[45], internal_0n[46], internal_0n[47]);
  OR2 I416 (complete805_0n[0], ifint_3n[0], itint_3n[0]);
  OR2 I417 (complete805_0n[1], ifint_3n[1], itint_3n[1]);
  OR2 I418 (complete805_0n[2], ifint_3n[2], itint_3n[2]);
  OR2 I419 (complete805_0n[3], ifint_3n[3], itint_3n[3]);
  OR2 I420 (complete805_0n[4], ifint_3n[4], itint_3n[4]);
  OR2 I421 (complete805_0n[5], ifint_3n[5], itint_3n[5]);
  OR2 I422 (complete805_0n[6], ifint_3n[6], itint_3n[6]);
  OR2 I423 (complete805_0n[7], ifint_3n[7], itint_3n[7]);
  OR2 I424 (complete805_0n[8], ifint_3n[8], itint_3n[8]);
  C3 I425 (internal_0n[48], complete804_0n[0], complete804_0n[1], complete804_0n[2]);
  C3 I426 (internal_0n[49], complete804_0n[3], complete804_0n[4], complete804_0n[5]);
  C3 I427 (internal_0n[50], complete804_0n[6], complete804_0n[7], complete804_0n[8]);
  C3 I428 (selcomp_2n, internal_0n[48], internal_0n[49], internal_0n[50]);
  OR2 I429 (complete804_0n[0], ifint_2n[0], itint_2n[0]);
  OR2 I430 (complete804_0n[1], ifint_2n[1], itint_2n[1]);
  OR2 I431 (complete804_0n[2], ifint_2n[2], itint_2n[2]);
  OR2 I432 (complete804_0n[3], ifint_2n[3], itint_2n[3]);
  OR2 I433 (complete804_0n[4], ifint_2n[4], itint_2n[4]);
  OR2 I434 (complete804_0n[5], ifint_2n[5], itint_2n[5]);
  OR2 I435 (complete804_0n[6], ifint_2n[6], itint_2n[6]);
  OR2 I436 (complete804_0n[7], ifint_2n[7], itint_2n[7]);
  OR2 I437 (complete804_0n[8], ifint_2n[8], itint_2n[8]);
  C3 I438 (internal_0n[51], complete803_0n[0], complete803_0n[1], complete803_0n[2]);
  C3 I439 (internal_0n[52], complete803_0n[3], complete803_0n[4], complete803_0n[5]);
  C3 I440 (internal_0n[53], complete803_0n[6], complete803_0n[7], complete803_0n[8]);
  C3 I441 (selcomp_1n, internal_0n[51], internal_0n[52], internal_0n[53]);
  OR2 I442 (complete803_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I443 (complete803_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I444 (complete803_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I445 (complete803_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I446 (complete803_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I447 (complete803_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I448 (complete803_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I449 (complete803_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I450 (complete803_0n[8], ifint_1n[8], itint_1n[8]);
  C3 I451 (internal_0n[54], complete802_0n[0], complete802_0n[1], complete802_0n[2]);
  C3 I452 (internal_0n[55], complete802_0n[3], complete802_0n[4], complete802_0n[5]);
  C3 I453 (internal_0n[56], complete802_0n[6], complete802_0n[7], complete802_0n[8]);
  C3 I454 (selcomp_0n, internal_0n[54], internal_0n[55], internal_0n[56]);
  OR2 I455 (complete802_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I456 (complete802_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I457 (complete802_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I458 (complete802_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I459 (complete802_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I460 (complete802_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I461 (complete802_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I462 (complete802_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I463 (complete802_0n[8], ifint_0n[8], itint_0n[8]);
  AND2 I464 (gfint_0n[0], gate_0n[0], ifint_0n[0]);
  AND2 I465 (gfint_0n[1], gate_0n[0], ifint_0n[1]);
  AND2 I466 (gfint_0n[2], gate_0n[0], ifint_0n[2]);
  AND2 I467 (gfint_0n[3], gate_0n[0], ifint_0n[3]);
  AND2 I468 (gfint_0n[4], gate_0n[0], ifint_0n[4]);
  AND2 I469 (gfint_0n[5], gate_0n[0], ifint_0n[5]);
  AND2 I470 (gfint_0n[6], gate_0n[0], ifint_0n[6]);
  AND2 I471 (gfint_0n[7], gate_0n[0], ifint_0n[7]);
  AND2 I472 (gfint_0n[8], gate_0n[0], ifint_0n[8]);
  AND2 I473 (gfint_1n[0], gate_0n[1], ifint_1n[0]);
  AND2 I474 (gfint_1n[1], gate_0n[1], ifint_1n[1]);
  AND2 I475 (gfint_1n[2], gate_0n[1], ifint_1n[2]);
  AND2 I476 (gfint_1n[3], gate_0n[1], ifint_1n[3]);
  AND2 I477 (gfint_1n[4], gate_0n[1], ifint_1n[4]);
  AND2 I478 (gfint_1n[5], gate_0n[1], ifint_1n[5]);
  AND2 I479 (gfint_1n[6], gate_0n[1], ifint_1n[6]);
  AND2 I480 (gfint_1n[7], gate_0n[1], ifint_1n[7]);
  AND2 I481 (gfint_1n[8], gate_0n[1], ifint_1n[8]);
  AND2 I482 (gfint_2n[0], gate_0n[2], ifint_2n[0]);
  AND2 I483 (gfint_2n[1], gate_0n[2], ifint_2n[1]);
  AND2 I484 (gfint_2n[2], gate_0n[2], ifint_2n[2]);
  AND2 I485 (gfint_2n[3], gate_0n[2], ifint_2n[3]);
  AND2 I486 (gfint_2n[4], gate_0n[2], ifint_2n[4]);
  AND2 I487 (gfint_2n[5], gate_0n[2], ifint_2n[5]);
  AND2 I488 (gfint_2n[6], gate_0n[2], ifint_2n[6]);
  AND2 I489 (gfint_2n[7], gate_0n[2], ifint_2n[7]);
  AND2 I490 (gfint_2n[8], gate_0n[2], ifint_2n[8]);
  AND2 I491 (gfint_3n[0], gate_0n[3], ifint_3n[0]);
  AND2 I492 (gfint_3n[1], gate_0n[3], ifint_3n[1]);
  AND2 I493 (gfint_3n[2], gate_0n[3], ifint_3n[2]);
  AND2 I494 (gfint_3n[3], gate_0n[3], ifint_3n[3]);
  AND2 I495 (gfint_3n[4], gate_0n[3], ifint_3n[4]);
  AND2 I496 (gfint_3n[5], gate_0n[3], ifint_3n[5]);
  AND2 I497 (gfint_3n[6], gate_0n[3], ifint_3n[6]);
  AND2 I498 (gfint_3n[7], gate_0n[3], ifint_3n[7]);
  AND2 I499 (gfint_3n[8], gate_0n[3], ifint_3n[8]);
  AND2 I500 (gfint_4n[0], gate_0n[4], ifint_4n[0]);
  AND2 I501 (gfint_4n[1], gate_0n[4], ifint_4n[1]);
  AND2 I502 (gfint_4n[2], gate_0n[4], ifint_4n[2]);
  AND2 I503 (gfint_4n[3], gate_0n[4], ifint_4n[3]);
  AND2 I504 (gfint_4n[4], gate_0n[4], ifint_4n[4]);
  AND2 I505 (gfint_4n[5], gate_0n[4], ifint_4n[5]);
  AND2 I506 (gfint_4n[6], gate_0n[4], ifint_4n[6]);
  AND2 I507 (gfint_4n[7], gate_0n[4], ifint_4n[7]);
  AND2 I508 (gfint_4n[8], gate_0n[4], ifint_4n[8]);
  AND2 I509 (gfint_5n[0], gate_0n[5], ifint_5n[0]);
  AND2 I510 (gfint_5n[1], gate_0n[5], ifint_5n[1]);
  AND2 I511 (gfint_5n[2], gate_0n[5], ifint_5n[2]);
  AND2 I512 (gfint_5n[3], gate_0n[5], ifint_5n[3]);
  AND2 I513 (gfint_5n[4], gate_0n[5], ifint_5n[4]);
  AND2 I514 (gfint_5n[5], gate_0n[5], ifint_5n[5]);
  AND2 I515 (gfint_5n[6], gate_0n[5], ifint_5n[6]);
  AND2 I516 (gfint_5n[7], gate_0n[5], ifint_5n[7]);
  AND2 I517 (gfint_5n[8], gate_0n[5], ifint_5n[8]);
  AND2 I518 (gfint_6n[0], gate_0n[6], ifint_6n[0]);
  AND2 I519 (gfint_6n[1], gate_0n[6], ifint_6n[1]);
  AND2 I520 (gfint_6n[2], gate_0n[6], ifint_6n[2]);
  AND2 I521 (gfint_6n[3], gate_0n[6], ifint_6n[3]);
  AND2 I522 (gfint_6n[4], gate_0n[6], ifint_6n[4]);
  AND2 I523 (gfint_6n[5], gate_0n[6], ifint_6n[5]);
  AND2 I524 (gfint_6n[6], gate_0n[6], ifint_6n[6]);
  AND2 I525 (gfint_6n[7], gate_0n[6], ifint_6n[7]);
  AND2 I526 (gfint_6n[8], gate_0n[6], ifint_6n[8]);
  AND2 I527 (gfint_7n[0], gate_0n[7], ifint_7n[0]);
  AND2 I528 (gfint_7n[1], gate_0n[7], ifint_7n[1]);
  AND2 I529 (gfint_7n[2], gate_0n[7], ifint_7n[2]);
  AND2 I530 (gfint_7n[3], gate_0n[7], ifint_7n[3]);
  AND2 I531 (gfint_7n[4], gate_0n[7], ifint_7n[4]);
  AND2 I532 (gfint_7n[5], gate_0n[7], ifint_7n[5]);
  AND2 I533 (gfint_7n[6], gate_0n[7], ifint_7n[6]);
  AND2 I534 (gfint_7n[7], gate_0n[7], ifint_7n[7]);
  AND2 I535 (gfint_7n[8], gate_0n[7], ifint_7n[8]);
  AND2 I536 (gfint_8n[0], gate_0n[8], ifint_8n[0]);
  AND2 I537 (gfint_8n[1], gate_0n[8], ifint_8n[1]);
  AND2 I538 (gfint_8n[2], gate_0n[8], ifint_8n[2]);
  AND2 I539 (gfint_8n[3], gate_0n[8], ifint_8n[3]);
  AND2 I540 (gfint_8n[4], gate_0n[8], ifint_8n[4]);
  AND2 I541 (gfint_8n[5], gate_0n[8], ifint_8n[5]);
  AND2 I542 (gfint_8n[6], gate_0n[8], ifint_8n[6]);
  AND2 I543 (gfint_8n[7], gate_0n[8], ifint_8n[7]);
  AND2 I544 (gfint_8n[8], gate_0n[8], ifint_8n[8]);
  AND2 I545 (gtint_0n[0], gate_0n[0], itint_0n[0]);
  AND2 I546 (gtint_0n[1], gate_0n[0], itint_0n[1]);
  AND2 I547 (gtint_0n[2], gate_0n[0], itint_0n[2]);
  AND2 I548 (gtint_0n[3], gate_0n[0], itint_0n[3]);
  AND2 I549 (gtint_0n[4], gate_0n[0], itint_0n[4]);
  AND2 I550 (gtint_0n[5], gate_0n[0], itint_0n[5]);
  AND2 I551 (gtint_0n[6], gate_0n[0], itint_0n[6]);
  AND2 I552 (gtint_0n[7], gate_0n[0], itint_0n[7]);
  AND2 I553 (gtint_0n[8], gate_0n[0], itint_0n[8]);
  AND2 I554 (gtint_1n[0], gate_0n[1], itint_1n[0]);
  AND2 I555 (gtint_1n[1], gate_0n[1], itint_1n[1]);
  AND2 I556 (gtint_1n[2], gate_0n[1], itint_1n[2]);
  AND2 I557 (gtint_1n[3], gate_0n[1], itint_1n[3]);
  AND2 I558 (gtint_1n[4], gate_0n[1], itint_1n[4]);
  AND2 I559 (gtint_1n[5], gate_0n[1], itint_1n[5]);
  AND2 I560 (gtint_1n[6], gate_0n[1], itint_1n[6]);
  AND2 I561 (gtint_1n[7], gate_0n[1], itint_1n[7]);
  AND2 I562 (gtint_1n[8], gate_0n[1], itint_1n[8]);
  AND2 I563 (gtint_2n[0], gate_0n[2], itint_2n[0]);
  AND2 I564 (gtint_2n[1], gate_0n[2], itint_2n[1]);
  AND2 I565 (gtint_2n[2], gate_0n[2], itint_2n[2]);
  AND2 I566 (gtint_2n[3], gate_0n[2], itint_2n[3]);
  AND2 I567 (gtint_2n[4], gate_0n[2], itint_2n[4]);
  AND2 I568 (gtint_2n[5], gate_0n[2], itint_2n[5]);
  AND2 I569 (gtint_2n[6], gate_0n[2], itint_2n[6]);
  AND2 I570 (gtint_2n[7], gate_0n[2], itint_2n[7]);
  AND2 I571 (gtint_2n[8], gate_0n[2], itint_2n[8]);
  AND2 I572 (gtint_3n[0], gate_0n[3], itint_3n[0]);
  AND2 I573 (gtint_3n[1], gate_0n[3], itint_3n[1]);
  AND2 I574 (gtint_3n[2], gate_0n[3], itint_3n[2]);
  AND2 I575 (gtint_3n[3], gate_0n[3], itint_3n[3]);
  AND2 I576 (gtint_3n[4], gate_0n[3], itint_3n[4]);
  AND2 I577 (gtint_3n[5], gate_0n[3], itint_3n[5]);
  AND2 I578 (gtint_3n[6], gate_0n[3], itint_3n[6]);
  AND2 I579 (gtint_3n[7], gate_0n[3], itint_3n[7]);
  AND2 I580 (gtint_3n[8], gate_0n[3], itint_3n[8]);
  AND2 I581 (gtint_4n[0], gate_0n[4], itint_4n[0]);
  AND2 I582 (gtint_4n[1], gate_0n[4], itint_4n[1]);
  AND2 I583 (gtint_4n[2], gate_0n[4], itint_4n[2]);
  AND2 I584 (gtint_4n[3], gate_0n[4], itint_4n[3]);
  AND2 I585 (gtint_4n[4], gate_0n[4], itint_4n[4]);
  AND2 I586 (gtint_4n[5], gate_0n[4], itint_4n[5]);
  AND2 I587 (gtint_4n[6], gate_0n[4], itint_4n[6]);
  AND2 I588 (gtint_4n[7], gate_0n[4], itint_4n[7]);
  AND2 I589 (gtint_4n[8], gate_0n[4], itint_4n[8]);
  AND2 I590 (gtint_5n[0], gate_0n[5], itint_5n[0]);
  AND2 I591 (gtint_5n[1], gate_0n[5], itint_5n[1]);
  AND2 I592 (gtint_5n[2], gate_0n[5], itint_5n[2]);
  AND2 I593 (gtint_5n[3], gate_0n[5], itint_5n[3]);
  AND2 I594 (gtint_5n[4], gate_0n[5], itint_5n[4]);
  AND2 I595 (gtint_5n[5], gate_0n[5], itint_5n[5]);
  AND2 I596 (gtint_5n[6], gate_0n[5], itint_5n[6]);
  AND2 I597 (gtint_5n[7], gate_0n[5], itint_5n[7]);
  AND2 I598 (gtint_5n[8], gate_0n[5], itint_5n[8]);
  AND2 I599 (gtint_6n[0], gate_0n[6], itint_6n[0]);
  AND2 I600 (gtint_6n[1], gate_0n[6], itint_6n[1]);
  AND2 I601 (gtint_6n[2], gate_0n[6], itint_6n[2]);
  AND2 I602 (gtint_6n[3], gate_0n[6], itint_6n[3]);
  AND2 I603 (gtint_6n[4], gate_0n[6], itint_6n[4]);
  AND2 I604 (gtint_6n[5], gate_0n[6], itint_6n[5]);
  AND2 I605 (gtint_6n[6], gate_0n[6], itint_6n[6]);
  AND2 I606 (gtint_6n[7], gate_0n[6], itint_6n[7]);
  AND2 I607 (gtint_6n[8], gate_0n[6], itint_6n[8]);
  AND2 I608 (gtint_7n[0], gate_0n[7], itint_7n[0]);
  AND2 I609 (gtint_7n[1], gate_0n[7], itint_7n[1]);
  AND2 I610 (gtint_7n[2], gate_0n[7], itint_7n[2]);
  AND2 I611 (gtint_7n[3], gate_0n[7], itint_7n[3]);
  AND2 I612 (gtint_7n[4], gate_0n[7], itint_7n[4]);
  AND2 I613 (gtint_7n[5], gate_0n[7], itint_7n[5]);
  AND2 I614 (gtint_7n[6], gate_0n[7], itint_7n[6]);
  AND2 I615 (gtint_7n[7], gate_0n[7], itint_7n[7]);
  AND2 I616 (gtint_7n[8], gate_0n[7], itint_7n[8]);
  AND2 I617 (gtint_8n[0], gate_0n[8], itint_8n[0]);
  AND2 I618 (gtint_8n[1], gate_0n[8], itint_8n[1]);
  AND2 I619 (gtint_8n[2], gate_0n[8], itint_8n[2]);
  AND2 I620 (gtint_8n[3], gate_0n[8], itint_8n[3]);
  AND2 I621 (gtint_8n[4], gate_0n[8], itint_8n[4]);
  AND2 I622 (gtint_8n[5], gate_0n[8], itint_8n[5]);
  AND2 I623 (gtint_8n[6], gate_0n[8], itint_8n[6]);
  AND2 I624 (gtint_8n[7], gate_0n[8], itint_8n[7]);
  AND2 I625 (gtint_8n[8], gate_0n[8], itint_8n[8]);
  NOR3 I626 (internal_0n[57], gtint_0n[0], gtint_1n[0], gtint_2n[0]);
  NOR3 I627 (internal_0n[58], gtint_3n[0], gtint_4n[0], gtint_5n[0]);
  NOR3 I628 (internal_0n[59], gtint_6n[0], gtint_7n[0], gtint_8n[0]);
  NAND3 I629 (otint_0n[0], internal_0n[57], internal_0n[58], internal_0n[59]);
  NOR3 I630 (internal_0n[60], gtint_0n[1], gtint_1n[1], gtint_2n[1]);
  NOR3 I631 (internal_0n[61], gtint_3n[1], gtint_4n[1], gtint_5n[1]);
  NOR3 I632 (internal_0n[62], gtint_6n[1], gtint_7n[1], gtint_8n[1]);
  NAND3 I633 (otint_0n[1], internal_0n[60], internal_0n[61], internal_0n[62]);
  NOR3 I634 (internal_0n[63], gtint_0n[2], gtint_1n[2], gtint_2n[2]);
  NOR3 I635 (internal_0n[64], gtint_3n[2], gtint_4n[2], gtint_5n[2]);
  NOR3 I636 (internal_0n[65], gtint_6n[2], gtint_7n[2], gtint_8n[2]);
  NAND3 I637 (otint_0n[2], internal_0n[63], internal_0n[64], internal_0n[65]);
  NOR3 I638 (internal_0n[66], gtint_0n[3], gtint_1n[3], gtint_2n[3]);
  NOR3 I639 (internal_0n[67], gtint_3n[3], gtint_4n[3], gtint_5n[3]);
  NOR3 I640 (internal_0n[68], gtint_6n[3], gtint_7n[3], gtint_8n[3]);
  NAND3 I641 (otint_0n[3], internal_0n[66], internal_0n[67], internal_0n[68]);
  NOR3 I642 (internal_0n[69], gtint_0n[4], gtint_1n[4], gtint_2n[4]);
  NOR3 I643 (internal_0n[70], gtint_3n[4], gtint_4n[4], gtint_5n[4]);
  NOR3 I644 (internal_0n[71], gtint_6n[4], gtint_7n[4], gtint_8n[4]);
  NAND3 I645 (otint_0n[4], internal_0n[69], internal_0n[70], internal_0n[71]);
  NOR3 I646 (internal_0n[72], gtint_0n[5], gtint_1n[5], gtint_2n[5]);
  NOR3 I647 (internal_0n[73], gtint_3n[5], gtint_4n[5], gtint_5n[5]);
  NOR3 I648 (internal_0n[74], gtint_6n[5], gtint_7n[5], gtint_8n[5]);
  NAND3 I649 (otint_0n[5], internal_0n[72], internal_0n[73], internal_0n[74]);
  NOR3 I650 (internal_0n[75], gtint_0n[6], gtint_1n[6], gtint_2n[6]);
  NOR3 I651 (internal_0n[76], gtint_3n[6], gtint_4n[6], gtint_5n[6]);
  NOR3 I652 (internal_0n[77], gtint_6n[6], gtint_7n[6], gtint_8n[6]);
  NAND3 I653 (otint_0n[6], internal_0n[75], internal_0n[76], internal_0n[77]);
  NOR3 I654 (internal_0n[78], gtint_0n[7], gtint_1n[7], gtint_2n[7]);
  NOR3 I655 (internal_0n[79], gtint_3n[7], gtint_4n[7], gtint_5n[7]);
  NOR3 I656 (internal_0n[80], gtint_6n[7], gtint_7n[7], gtint_8n[7]);
  NAND3 I657 (otint_0n[7], internal_0n[78], internal_0n[79], internal_0n[80]);
  NOR3 I658 (internal_0n[81], gtint_0n[8], gtint_1n[8], gtint_2n[8]);
  NOR3 I659 (internal_0n[82], gtint_3n[8], gtint_4n[8], gtint_5n[8]);
  NOR3 I660 (internal_0n[83], gtint_6n[8], gtint_7n[8], gtint_8n[8]);
  NAND3 I661 (otint_0n[8], internal_0n[81], internal_0n[82], internal_0n[83]);
  NOR3 I662 (internal_0n[84], gfint_0n[0], gfint_1n[0], gfint_2n[0]);
  NOR3 I663 (internal_0n[85], gfint_3n[0], gfint_4n[0], gfint_5n[0]);
  NOR3 I664 (internal_0n[86], gfint_6n[0], gfint_7n[0], gfint_8n[0]);
  NAND3 I665 (ofint_0n[0], internal_0n[84], internal_0n[85], internal_0n[86]);
  NOR3 I666 (internal_0n[87], gfint_0n[1], gfint_1n[1], gfint_2n[1]);
  NOR3 I667 (internal_0n[88], gfint_3n[1], gfint_4n[1], gfint_5n[1]);
  NOR3 I668 (internal_0n[89], gfint_6n[1], gfint_7n[1], gfint_8n[1]);
  NAND3 I669 (ofint_0n[1], internal_0n[87], internal_0n[88], internal_0n[89]);
  NOR3 I670 (internal_0n[90], gfint_0n[2], gfint_1n[2], gfint_2n[2]);
  NOR3 I671 (internal_0n[91], gfint_3n[2], gfint_4n[2], gfint_5n[2]);
  NOR3 I672 (internal_0n[92], gfint_6n[2], gfint_7n[2], gfint_8n[2]);
  NAND3 I673 (ofint_0n[2], internal_0n[90], internal_0n[91], internal_0n[92]);
  NOR3 I674 (internal_0n[93], gfint_0n[3], gfint_1n[3], gfint_2n[3]);
  NOR3 I675 (internal_0n[94], gfint_3n[3], gfint_4n[3], gfint_5n[3]);
  NOR3 I676 (internal_0n[95], gfint_6n[3], gfint_7n[3], gfint_8n[3]);
  NAND3 I677 (ofint_0n[3], internal_0n[93], internal_0n[94], internal_0n[95]);
  NOR3 I678 (internal_0n[96], gfint_0n[4], gfint_1n[4], gfint_2n[4]);
  NOR3 I679 (internal_0n[97], gfint_3n[4], gfint_4n[4], gfint_5n[4]);
  NOR3 I680 (internal_0n[98], gfint_6n[4], gfint_7n[4], gfint_8n[4]);
  NAND3 I681 (ofint_0n[4], internal_0n[96], internal_0n[97], internal_0n[98]);
  NOR3 I682 (internal_0n[99], gfint_0n[5], gfint_1n[5], gfint_2n[5]);
  NOR3 I683 (internal_0n[100], gfint_3n[5], gfint_4n[5], gfint_5n[5]);
  NOR3 I684 (internal_0n[101], gfint_6n[5], gfint_7n[5], gfint_8n[5]);
  NAND3 I685 (ofint_0n[5], internal_0n[99], internal_0n[100], internal_0n[101]);
  NOR3 I686 (internal_0n[102], gfint_0n[6], gfint_1n[6], gfint_2n[6]);
  NOR3 I687 (internal_0n[103], gfint_3n[6], gfint_4n[6], gfint_5n[6]);
  NOR3 I688 (internal_0n[104], gfint_6n[6], gfint_7n[6], gfint_8n[6]);
  NAND3 I689 (ofint_0n[6], internal_0n[102], internal_0n[103], internal_0n[104]);
  NOR3 I690 (internal_0n[105], gfint_0n[7], gfint_1n[7], gfint_2n[7]);
  NOR3 I691 (internal_0n[106], gfint_3n[7], gfint_4n[7], gfint_5n[7]);
  NOR3 I692 (internal_0n[107], gfint_6n[7], gfint_7n[7], gfint_8n[7]);
  NAND3 I693 (ofint_0n[7], internal_0n[105], internal_0n[106], internal_0n[107]);
  NOR3 I694 (internal_0n[108], gfint_0n[8], gfint_1n[8], gfint_2n[8]);
  NOR3 I695 (internal_0n[109], gfint_3n[8], gfint_4n[8], gfint_5n[8]);
  NOR3 I696 (internal_0n[110], gfint_6n[8], gfint_7n[8], gfint_8n[8]);
  NAND3 I697 (ofint_0n[8], internal_0n[108], internal_0n[109], internal_0n[110]);
endmodule

module BrzM_32_2 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [31:0] i_0r0d;
  input [31:0] i_0r1d;
  output i_0a;
  input [31:0] i_1r0d;
  input [31:0] i_1r1d;
  output i_1a;
  output [31:0] o_0r0d;
  output [31:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [84:0] internal_0n;
  wire [1:0] sel_0n;
  wire [31:0] ofint_0n;
  wire [31:0] otint_0n;
  wire oaint_0n;
  wire [31:0] ifint_0n;
  wire [31:0] ifint_1n;
  wire [31:0] itint_0n;
  wire [31:0] itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [1:0] gate_0n;
  wire [31:0] gfint_0n;
  wire [31:0] gfint_1n;
  wire [31:0] gtint_0n;
  wire [31:0] gtint_1n;
  wire [31:0] complete864_0n;
  wire gate863_0n;
  wire [31:0] complete860_0n;
  wire gate859_0n;
  wire [31:0] complete856_0n;
  wire gate855_0n;
  wire [31:0] complete852_0n;
  wire [31:0] complete851_0n;
  wire selcomp_0n;
  wire selcomp_1n;
  C3 I0 (internal_0n[0], complete864_0n[0], complete864_0n[1], complete864_0n[2]);
  C3 I1 (internal_0n[1], complete864_0n[3], complete864_0n[4], complete864_0n[5]);
  C3 I2 (internal_0n[2], complete864_0n[6], complete864_0n[7], complete864_0n[8]);
  C3 I3 (internal_0n[3], complete864_0n[9], complete864_0n[10], complete864_0n[11]);
  C3 I4 (internal_0n[4], complete864_0n[12], complete864_0n[13], complete864_0n[14]);
  C3 I5 (internal_0n[5], complete864_0n[15], complete864_0n[16], complete864_0n[17]);
  C3 I6 (internal_0n[6], complete864_0n[18], complete864_0n[19], complete864_0n[20]);
  C3 I7 (internal_0n[7], complete864_0n[21], complete864_0n[22], complete864_0n[23]);
  C3 I8 (internal_0n[8], complete864_0n[24], complete864_0n[25], complete864_0n[26]);
  C3 I9 (internal_0n[9], complete864_0n[27], complete864_0n[28], complete864_0n[29]);
  C2 I10 (internal_0n[10], complete864_0n[30], complete864_0n[31]);
  C3 I11 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I12 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I13 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I14 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I15 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I16 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I17 (i_1a, internal_0n[15], internal_0n[16]);
  OR2 I18 (complete864_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I19 (complete864_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I20 (complete864_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I21 (complete864_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I22 (complete864_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I23 (complete864_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I24 (complete864_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I25 (complete864_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I26 (complete864_0n[8], ifint_1n[8], itint_1n[8]);
  OR2 I27 (complete864_0n[9], ifint_1n[9], itint_1n[9]);
  OR2 I28 (complete864_0n[10], ifint_1n[10], itint_1n[10]);
  OR2 I29 (complete864_0n[11], ifint_1n[11], itint_1n[11]);
  OR2 I30 (complete864_0n[12], ifint_1n[12], itint_1n[12]);
  OR2 I31 (complete864_0n[13], ifint_1n[13], itint_1n[13]);
  OR2 I32 (complete864_0n[14], ifint_1n[14], itint_1n[14]);
  OR2 I33 (complete864_0n[15], ifint_1n[15], itint_1n[15]);
  OR2 I34 (complete864_0n[16], ifint_1n[16], itint_1n[16]);
  OR2 I35 (complete864_0n[17], ifint_1n[17], itint_1n[17]);
  OR2 I36 (complete864_0n[18], ifint_1n[18], itint_1n[18]);
  OR2 I37 (complete864_0n[19], ifint_1n[19], itint_1n[19]);
  OR2 I38 (complete864_0n[20], ifint_1n[20], itint_1n[20]);
  OR2 I39 (complete864_0n[21], ifint_1n[21], itint_1n[21]);
  OR2 I40 (complete864_0n[22], ifint_1n[22], itint_1n[22]);
  OR2 I41 (complete864_0n[23], ifint_1n[23], itint_1n[23]);
  OR2 I42 (complete864_0n[24], ifint_1n[24], itint_1n[24]);
  OR2 I43 (complete864_0n[25], ifint_1n[25], itint_1n[25]);
  OR2 I44 (complete864_0n[26], ifint_1n[26], itint_1n[26]);
  OR2 I45 (complete864_0n[27], ifint_1n[27], itint_1n[27]);
  OR2 I46 (complete864_0n[28], ifint_1n[28], itint_1n[28]);
  OR2 I47 (complete864_0n[29], ifint_1n[29], itint_1n[29]);
  OR2 I48 (complete864_0n[30], ifint_1n[30], itint_1n[30]);
  OR2 I49 (complete864_0n[31], ifint_1n[31], itint_1n[31]);
  INV I50 (gate863_0n, iaint_1n);
  C2RI I51 (itint_1n[0], i_1r1d[0], gate863_0n, initialise);
  C2RI I52 (itint_1n[1], i_1r1d[1], gate863_0n, initialise);
  C2RI I53 (itint_1n[2], i_1r1d[2], gate863_0n, initialise);
  C2RI I54 (itint_1n[3], i_1r1d[3], gate863_0n, initialise);
  C2RI I55 (itint_1n[4], i_1r1d[4], gate863_0n, initialise);
  C2RI I56 (itint_1n[5], i_1r1d[5], gate863_0n, initialise);
  C2RI I57 (itint_1n[6], i_1r1d[6], gate863_0n, initialise);
  C2RI I58 (itint_1n[7], i_1r1d[7], gate863_0n, initialise);
  C2RI I59 (itint_1n[8], i_1r1d[8], gate863_0n, initialise);
  C2RI I60 (itint_1n[9], i_1r1d[9], gate863_0n, initialise);
  C2RI I61 (itint_1n[10], i_1r1d[10], gate863_0n, initialise);
  C2RI I62 (itint_1n[11], i_1r1d[11], gate863_0n, initialise);
  C2RI I63 (itint_1n[12], i_1r1d[12], gate863_0n, initialise);
  C2RI I64 (itint_1n[13], i_1r1d[13], gate863_0n, initialise);
  C2RI I65 (itint_1n[14], i_1r1d[14], gate863_0n, initialise);
  C2RI I66 (itint_1n[15], i_1r1d[15], gate863_0n, initialise);
  C2RI I67 (itint_1n[16], i_1r1d[16], gate863_0n, initialise);
  C2RI I68 (itint_1n[17], i_1r1d[17], gate863_0n, initialise);
  C2RI I69 (itint_1n[18], i_1r1d[18], gate863_0n, initialise);
  C2RI I70 (itint_1n[19], i_1r1d[19], gate863_0n, initialise);
  C2RI I71 (itint_1n[20], i_1r1d[20], gate863_0n, initialise);
  C2RI I72 (itint_1n[21], i_1r1d[21], gate863_0n, initialise);
  C2RI I73 (itint_1n[22], i_1r1d[22], gate863_0n, initialise);
  C2RI I74 (itint_1n[23], i_1r1d[23], gate863_0n, initialise);
  C2RI I75 (itint_1n[24], i_1r1d[24], gate863_0n, initialise);
  C2RI I76 (itint_1n[25], i_1r1d[25], gate863_0n, initialise);
  C2RI I77 (itint_1n[26], i_1r1d[26], gate863_0n, initialise);
  C2RI I78 (itint_1n[27], i_1r1d[27], gate863_0n, initialise);
  C2RI I79 (itint_1n[28], i_1r1d[28], gate863_0n, initialise);
  C2RI I80 (itint_1n[29], i_1r1d[29], gate863_0n, initialise);
  C2RI I81 (itint_1n[30], i_1r1d[30], gate863_0n, initialise);
  C2RI I82 (itint_1n[31], i_1r1d[31], gate863_0n, initialise);
  C2RI I83 (ifint_1n[0], i_1r0d[0], gate863_0n, initialise);
  C2RI I84 (ifint_1n[1], i_1r0d[1], gate863_0n, initialise);
  C2RI I85 (ifint_1n[2], i_1r0d[2], gate863_0n, initialise);
  C2RI I86 (ifint_1n[3], i_1r0d[3], gate863_0n, initialise);
  C2RI I87 (ifint_1n[4], i_1r0d[4], gate863_0n, initialise);
  C2RI I88 (ifint_1n[5], i_1r0d[5], gate863_0n, initialise);
  C2RI I89 (ifint_1n[6], i_1r0d[6], gate863_0n, initialise);
  C2RI I90 (ifint_1n[7], i_1r0d[7], gate863_0n, initialise);
  C2RI I91 (ifint_1n[8], i_1r0d[8], gate863_0n, initialise);
  C2RI I92 (ifint_1n[9], i_1r0d[9], gate863_0n, initialise);
  C2RI I93 (ifint_1n[10], i_1r0d[10], gate863_0n, initialise);
  C2RI I94 (ifint_1n[11], i_1r0d[11], gate863_0n, initialise);
  C2RI I95 (ifint_1n[12], i_1r0d[12], gate863_0n, initialise);
  C2RI I96 (ifint_1n[13], i_1r0d[13], gate863_0n, initialise);
  C2RI I97 (ifint_1n[14], i_1r0d[14], gate863_0n, initialise);
  C2RI I98 (ifint_1n[15], i_1r0d[15], gate863_0n, initialise);
  C2RI I99 (ifint_1n[16], i_1r0d[16], gate863_0n, initialise);
  C2RI I100 (ifint_1n[17], i_1r0d[17], gate863_0n, initialise);
  C2RI I101 (ifint_1n[18], i_1r0d[18], gate863_0n, initialise);
  C2RI I102 (ifint_1n[19], i_1r0d[19], gate863_0n, initialise);
  C2RI I103 (ifint_1n[20], i_1r0d[20], gate863_0n, initialise);
  C2RI I104 (ifint_1n[21], i_1r0d[21], gate863_0n, initialise);
  C2RI I105 (ifint_1n[22], i_1r0d[22], gate863_0n, initialise);
  C2RI I106 (ifint_1n[23], i_1r0d[23], gate863_0n, initialise);
  C2RI I107 (ifint_1n[24], i_1r0d[24], gate863_0n, initialise);
  C2RI I108 (ifint_1n[25], i_1r0d[25], gate863_0n, initialise);
  C2RI I109 (ifint_1n[26], i_1r0d[26], gate863_0n, initialise);
  C2RI I110 (ifint_1n[27], i_1r0d[27], gate863_0n, initialise);
  C2RI I111 (ifint_1n[28], i_1r0d[28], gate863_0n, initialise);
  C2RI I112 (ifint_1n[29], i_1r0d[29], gate863_0n, initialise);
  C2RI I113 (ifint_1n[30], i_1r0d[30], gate863_0n, initialise);
  C2RI I114 (ifint_1n[31], i_1r0d[31], gate863_0n, initialise);
  C3 I115 (internal_0n[17], complete860_0n[0], complete860_0n[1], complete860_0n[2]);
  C3 I116 (internal_0n[18], complete860_0n[3], complete860_0n[4], complete860_0n[5]);
  C3 I117 (internal_0n[19], complete860_0n[6], complete860_0n[7], complete860_0n[8]);
  C3 I118 (internal_0n[20], complete860_0n[9], complete860_0n[10], complete860_0n[11]);
  C3 I119 (internal_0n[21], complete860_0n[12], complete860_0n[13], complete860_0n[14]);
  C3 I120 (internal_0n[22], complete860_0n[15], complete860_0n[16], complete860_0n[17]);
  C3 I121 (internal_0n[23], complete860_0n[18], complete860_0n[19], complete860_0n[20]);
  C3 I122 (internal_0n[24], complete860_0n[21], complete860_0n[22], complete860_0n[23]);
  C3 I123 (internal_0n[25], complete860_0n[24], complete860_0n[25], complete860_0n[26]);
  C3 I124 (internal_0n[26], complete860_0n[27], complete860_0n[28], complete860_0n[29]);
  C2 I125 (internal_0n[27], complete860_0n[30], complete860_0n[31]);
  C3 I126 (internal_0n[28], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I127 (internal_0n[29], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I128 (internal_0n[30], internal_0n[23], internal_0n[24], internal_0n[25]);
  C2 I129 (internal_0n[31], internal_0n[26], internal_0n[27]);
  C2 I130 (internal_0n[32], internal_0n[28], internal_0n[29]);
  C2 I131 (internal_0n[33], internal_0n[30], internal_0n[31]);
  C2 I132 (i_0a, internal_0n[32], internal_0n[33]);
  OR2 I133 (complete860_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I134 (complete860_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I135 (complete860_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I136 (complete860_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I137 (complete860_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I138 (complete860_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I139 (complete860_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I140 (complete860_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I141 (complete860_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I142 (complete860_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I143 (complete860_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I144 (complete860_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I145 (complete860_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I146 (complete860_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I147 (complete860_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I148 (complete860_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I149 (complete860_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I150 (complete860_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I151 (complete860_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I152 (complete860_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I153 (complete860_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I154 (complete860_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I155 (complete860_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I156 (complete860_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I157 (complete860_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I158 (complete860_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I159 (complete860_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I160 (complete860_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I161 (complete860_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I162 (complete860_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I163 (complete860_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I164 (complete860_0n[31], ifint_0n[31], itint_0n[31]);
  INV I165 (gate859_0n, iaint_0n);
  C2RI I166 (itint_0n[0], i_0r1d[0], gate859_0n, initialise);
  C2RI I167 (itint_0n[1], i_0r1d[1], gate859_0n, initialise);
  C2RI I168 (itint_0n[2], i_0r1d[2], gate859_0n, initialise);
  C2RI I169 (itint_0n[3], i_0r1d[3], gate859_0n, initialise);
  C2RI I170 (itint_0n[4], i_0r1d[4], gate859_0n, initialise);
  C2RI I171 (itint_0n[5], i_0r1d[5], gate859_0n, initialise);
  C2RI I172 (itint_0n[6], i_0r1d[6], gate859_0n, initialise);
  C2RI I173 (itint_0n[7], i_0r1d[7], gate859_0n, initialise);
  C2RI I174 (itint_0n[8], i_0r1d[8], gate859_0n, initialise);
  C2RI I175 (itint_0n[9], i_0r1d[9], gate859_0n, initialise);
  C2RI I176 (itint_0n[10], i_0r1d[10], gate859_0n, initialise);
  C2RI I177 (itint_0n[11], i_0r1d[11], gate859_0n, initialise);
  C2RI I178 (itint_0n[12], i_0r1d[12], gate859_0n, initialise);
  C2RI I179 (itint_0n[13], i_0r1d[13], gate859_0n, initialise);
  C2RI I180 (itint_0n[14], i_0r1d[14], gate859_0n, initialise);
  C2RI I181 (itint_0n[15], i_0r1d[15], gate859_0n, initialise);
  C2RI I182 (itint_0n[16], i_0r1d[16], gate859_0n, initialise);
  C2RI I183 (itint_0n[17], i_0r1d[17], gate859_0n, initialise);
  C2RI I184 (itint_0n[18], i_0r1d[18], gate859_0n, initialise);
  C2RI I185 (itint_0n[19], i_0r1d[19], gate859_0n, initialise);
  C2RI I186 (itint_0n[20], i_0r1d[20], gate859_0n, initialise);
  C2RI I187 (itint_0n[21], i_0r1d[21], gate859_0n, initialise);
  C2RI I188 (itint_0n[22], i_0r1d[22], gate859_0n, initialise);
  C2RI I189 (itint_0n[23], i_0r1d[23], gate859_0n, initialise);
  C2RI I190 (itint_0n[24], i_0r1d[24], gate859_0n, initialise);
  C2RI I191 (itint_0n[25], i_0r1d[25], gate859_0n, initialise);
  C2RI I192 (itint_0n[26], i_0r1d[26], gate859_0n, initialise);
  C2RI I193 (itint_0n[27], i_0r1d[27], gate859_0n, initialise);
  C2RI I194 (itint_0n[28], i_0r1d[28], gate859_0n, initialise);
  C2RI I195 (itint_0n[29], i_0r1d[29], gate859_0n, initialise);
  C2RI I196 (itint_0n[30], i_0r1d[30], gate859_0n, initialise);
  C2RI I197 (itint_0n[31], i_0r1d[31], gate859_0n, initialise);
  C2RI I198 (ifint_0n[0], i_0r0d[0], gate859_0n, initialise);
  C2RI I199 (ifint_0n[1], i_0r0d[1], gate859_0n, initialise);
  C2RI I200 (ifint_0n[2], i_0r0d[2], gate859_0n, initialise);
  C2RI I201 (ifint_0n[3], i_0r0d[3], gate859_0n, initialise);
  C2RI I202 (ifint_0n[4], i_0r0d[4], gate859_0n, initialise);
  C2RI I203 (ifint_0n[5], i_0r0d[5], gate859_0n, initialise);
  C2RI I204 (ifint_0n[6], i_0r0d[6], gate859_0n, initialise);
  C2RI I205 (ifint_0n[7], i_0r0d[7], gate859_0n, initialise);
  C2RI I206 (ifint_0n[8], i_0r0d[8], gate859_0n, initialise);
  C2RI I207 (ifint_0n[9], i_0r0d[9], gate859_0n, initialise);
  C2RI I208 (ifint_0n[10], i_0r0d[10], gate859_0n, initialise);
  C2RI I209 (ifint_0n[11], i_0r0d[11], gate859_0n, initialise);
  C2RI I210 (ifint_0n[12], i_0r0d[12], gate859_0n, initialise);
  C2RI I211 (ifint_0n[13], i_0r0d[13], gate859_0n, initialise);
  C2RI I212 (ifint_0n[14], i_0r0d[14], gate859_0n, initialise);
  C2RI I213 (ifint_0n[15], i_0r0d[15], gate859_0n, initialise);
  C2RI I214 (ifint_0n[16], i_0r0d[16], gate859_0n, initialise);
  C2RI I215 (ifint_0n[17], i_0r0d[17], gate859_0n, initialise);
  C2RI I216 (ifint_0n[18], i_0r0d[18], gate859_0n, initialise);
  C2RI I217 (ifint_0n[19], i_0r0d[19], gate859_0n, initialise);
  C2RI I218 (ifint_0n[20], i_0r0d[20], gate859_0n, initialise);
  C2RI I219 (ifint_0n[21], i_0r0d[21], gate859_0n, initialise);
  C2RI I220 (ifint_0n[22], i_0r0d[22], gate859_0n, initialise);
  C2RI I221 (ifint_0n[23], i_0r0d[23], gate859_0n, initialise);
  C2RI I222 (ifint_0n[24], i_0r0d[24], gate859_0n, initialise);
  C2RI I223 (ifint_0n[25], i_0r0d[25], gate859_0n, initialise);
  C2RI I224 (ifint_0n[26], i_0r0d[26], gate859_0n, initialise);
  C2RI I225 (ifint_0n[27], i_0r0d[27], gate859_0n, initialise);
  C2RI I226 (ifint_0n[28], i_0r0d[28], gate859_0n, initialise);
  C2RI I227 (ifint_0n[29], i_0r0d[29], gate859_0n, initialise);
  C2RI I228 (ifint_0n[30], i_0r0d[30], gate859_0n, initialise);
  C2RI I229 (ifint_0n[31], i_0r0d[31], gate859_0n, initialise);
  C3 I230 (internal_0n[34], complete856_0n[0], complete856_0n[1], complete856_0n[2]);
  C3 I231 (internal_0n[35], complete856_0n[3], complete856_0n[4], complete856_0n[5]);
  C3 I232 (internal_0n[36], complete856_0n[6], complete856_0n[7], complete856_0n[8]);
  C3 I233 (internal_0n[37], complete856_0n[9], complete856_0n[10], complete856_0n[11]);
  C3 I234 (internal_0n[38], complete856_0n[12], complete856_0n[13], complete856_0n[14]);
  C3 I235 (internal_0n[39], complete856_0n[15], complete856_0n[16], complete856_0n[17]);
  C3 I236 (internal_0n[40], complete856_0n[18], complete856_0n[19], complete856_0n[20]);
  C3 I237 (internal_0n[41], complete856_0n[21], complete856_0n[22], complete856_0n[23]);
  C3 I238 (internal_0n[42], complete856_0n[24], complete856_0n[25], complete856_0n[26]);
  C3 I239 (internal_0n[43], complete856_0n[27], complete856_0n[28], complete856_0n[29]);
  C2 I240 (internal_0n[44], complete856_0n[30], complete856_0n[31]);
  C3 I241 (internal_0n[45], internal_0n[34], internal_0n[35], internal_0n[36]);
  C3 I242 (internal_0n[46], internal_0n[37], internal_0n[38], internal_0n[39]);
  C3 I243 (internal_0n[47], internal_0n[40], internal_0n[41], internal_0n[42]);
  C2 I244 (internal_0n[48], internal_0n[43], internal_0n[44]);
  C2 I245 (internal_0n[49], internal_0n[45], internal_0n[46]);
  C2 I246 (internal_0n[50], internal_0n[47], internal_0n[48]);
  C2 I247 (oaint_0n, internal_0n[49], internal_0n[50]);
  OR2 I248 (complete856_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I249 (complete856_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I250 (complete856_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I251 (complete856_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I252 (complete856_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I253 (complete856_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I254 (complete856_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I255 (complete856_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I256 (complete856_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I257 (complete856_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I258 (complete856_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I259 (complete856_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I260 (complete856_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I261 (complete856_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I262 (complete856_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I263 (complete856_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I264 (complete856_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I265 (complete856_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I266 (complete856_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I267 (complete856_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I268 (complete856_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I269 (complete856_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I270 (complete856_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I271 (complete856_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I272 (complete856_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I273 (complete856_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I274 (complete856_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I275 (complete856_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I276 (complete856_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I277 (complete856_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I278 (complete856_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I279 (complete856_0n[31], o_0r0d[31], o_0r1d[31]);
  INV I280 (gate855_0n, o_0a);
  C2RI I281 (o_0r1d[0], otint_0n[0], gate855_0n, initialise);
  C2RI I282 (o_0r1d[1], otint_0n[1], gate855_0n, initialise);
  C2RI I283 (o_0r1d[2], otint_0n[2], gate855_0n, initialise);
  C2RI I284 (o_0r1d[3], otint_0n[3], gate855_0n, initialise);
  C2RI I285 (o_0r1d[4], otint_0n[4], gate855_0n, initialise);
  C2RI I286 (o_0r1d[5], otint_0n[5], gate855_0n, initialise);
  C2RI I287 (o_0r1d[6], otint_0n[6], gate855_0n, initialise);
  C2RI I288 (o_0r1d[7], otint_0n[7], gate855_0n, initialise);
  C2RI I289 (o_0r1d[8], otint_0n[8], gate855_0n, initialise);
  C2RI I290 (o_0r1d[9], otint_0n[9], gate855_0n, initialise);
  C2RI I291 (o_0r1d[10], otint_0n[10], gate855_0n, initialise);
  C2RI I292 (o_0r1d[11], otint_0n[11], gate855_0n, initialise);
  C2RI I293 (o_0r1d[12], otint_0n[12], gate855_0n, initialise);
  C2RI I294 (o_0r1d[13], otint_0n[13], gate855_0n, initialise);
  C2RI I295 (o_0r1d[14], otint_0n[14], gate855_0n, initialise);
  C2RI I296 (o_0r1d[15], otint_0n[15], gate855_0n, initialise);
  C2RI I297 (o_0r1d[16], otint_0n[16], gate855_0n, initialise);
  C2RI I298 (o_0r1d[17], otint_0n[17], gate855_0n, initialise);
  C2RI I299 (o_0r1d[18], otint_0n[18], gate855_0n, initialise);
  C2RI I300 (o_0r1d[19], otint_0n[19], gate855_0n, initialise);
  C2RI I301 (o_0r1d[20], otint_0n[20], gate855_0n, initialise);
  C2RI I302 (o_0r1d[21], otint_0n[21], gate855_0n, initialise);
  C2RI I303 (o_0r1d[22], otint_0n[22], gate855_0n, initialise);
  C2RI I304 (o_0r1d[23], otint_0n[23], gate855_0n, initialise);
  C2RI I305 (o_0r1d[24], otint_0n[24], gate855_0n, initialise);
  C2RI I306 (o_0r1d[25], otint_0n[25], gate855_0n, initialise);
  C2RI I307 (o_0r1d[26], otint_0n[26], gate855_0n, initialise);
  C2RI I308 (o_0r1d[27], otint_0n[27], gate855_0n, initialise);
  C2RI I309 (o_0r1d[28], otint_0n[28], gate855_0n, initialise);
  C2RI I310 (o_0r1d[29], otint_0n[29], gate855_0n, initialise);
  C2RI I311 (o_0r1d[30], otint_0n[30], gate855_0n, initialise);
  C2RI I312 (o_0r1d[31], otint_0n[31], gate855_0n, initialise);
  C2RI I313 (o_0r0d[0], ofint_0n[0], gate855_0n, initialise);
  C2RI I314 (o_0r0d[1], ofint_0n[1], gate855_0n, initialise);
  C2RI I315 (o_0r0d[2], ofint_0n[2], gate855_0n, initialise);
  C2RI I316 (o_0r0d[3], ofint_0n[3], gate855_0n, initialise);
  C2RI I317 (o_0r0d[4], ofint_0n[4], gate855_0n, initialise);
  C2RI I318 (o_0r0d[5], ofint_0n[5], gate855_0n, initialise);
  C2RI I319 (o_0r0d[6], ofint_0n[6], gate855_0n, initialise);
  C2RI I320 (o_0r0d[7], ofint_0n[7], gate855_0n, initialise);
  C2RI I321 (o_0r0d[8], ofint_0n[8], gate855_0n, initialise);
  C2RI I322 (o_0r0d[9], ofint_0n[9], gate855_0n, initialise);
  C2RI I323 (o_0r0d[10], ofint_0n[10], gate855_0n, initialise);
  C2RI I324 (o_0r0d[11], ofint_0n[11], gate855_0n, initialise);
  C2RI I325 (o_0r0d[12], ofint_0n[12], gate855_0n, initialise);
  C2RI I326 (o_0r0d[13], ofint_0n[13], gate855_0n, initialise);
  C2RI I327 (o_0r0d[14], ofint_0n[14], gate855_0n, initialise);
  C2RI I328 (o_0r0d[15], ofint_0n[15], gate855_0n, initialise);
  C2RI I329 (o_0r0d[16], ofint_0n[16], gate855_0n, initialise);
  C2RI I330 (o_0r0d[17], ofint_0n[17], gate855_0n, initialise);
  C2RI I331 (o_0r0d[18], ofint_0n[18], gate855_0n, initialise);
  C2RI I332 (o_0r0d[19], ofint_0n[19], gate855_0n, initialise);
  C2RI I333 (o_0r0d[20], ofint_0n[20], gate855_0n, initialise);
  C2RI I334 (o_0r0d[21], ofint_0n[21], gate855_0n, initialise);
  C2RI I335 (o_0r0d[22], ofint_0n[22], gate855_0n, initialise);
  C2RI I336 (o_0r0d[23], ofint_0n[23], gate855_0n, initialise);
  C2RI I337 (o_0r0d[24], ofint_0n[24], gate855_0n, initialise);
  C2RI I338 (o_0r0d[25], ofint_0n[25], gate855_0n, initialise);
  C2RI I339 (o_0r0d[26], ofint_0n[26], gate855_0n, initialise);
  C2RI I340 (o_0r0d[27], ofint_0n[27], gate855_0n, initialise);
  C2RI I341 (o_0r0d[28], ofint_0n[28], gate855_0n, initialise);
  C2RI I342 (o_0r0d[29], ofint_0n[29], gate855_0n, initialise);
  C2RI I343 (o_0r0d[30], ofint_0n[30], gate855_0n, initialise);
  C2RI I344 (o_0r0d[31], ofint_0n[31], gate855_0n, initialise);
  C2RI I345 (iaint_0n, sel_0n[0], oaint_0n, initialise);
  C2RI I346 (iaint_1n, sel_0n[1], oaint_0n, initialise);
  assign gate_0n[0] = sel_0n[0];
  assign gate_0n[1] = sel_0n[1];
  assign sel_0n[0] = selcomp_0n;
  assign sel_0n[1] = selcomp_1n;
  C3 I351 (internal_0n[51], complete852_0n[0], complete852_0n[1], complete852_0n[2]);
  C3 I352 (internal_0n[52], complete852_0n[3], complete852_0n[4], complete852_0n[5]);
  C3 I353 (internal_0n[53], complete852_0n[6], complete852_0n[7], complete852_0n[8]);
  C3 I354 (internal_0n[54], complete852_0n[9], complete852_0n[10], complete852_0n[11]);
  C3 I355 (internal_0n[55], complete852_0n[12], complete852_0n[13], complete852_0n[14]);
  C3 I356 (internal_0n[56], complete852_0n[15], complete852_0n[16], complete852_0n[17]);
  C3 I357 (internal_0n[57], complete852_0n[18], complete852_0n[19], complete852_0n[20]);
  C3 I358 (internal_0n[58], complete852_0n[21], complete852_0n[22], complete852_0n[23]);
  C3 I359 (internal_0n[59], complete852_0n[24], complete852_0n[25], complete852_0n[26]);
  C3 I360 (internal_0n[60], complete852_0n[27], complete852_0n[28], complete852_0n[29]);
  C2 I361 (internal_0n[61], complete852_0n[30], complete852_0n[31]);
  C3 I362 (internal_0n[62], internal_0n[51], internal_0n[52], internal_0n[53]);
  C3 I363 (internal_0n[63], internal_0n[54], internal_0n[55], internal_0n[56]);
  C3 I364 (internal_0n[64], internal_0n[57], internal_0n[58], internal_0n[59]);
  C2 I365 (internal_0n[65], internal_0n[60], internal_0n[61]);
  C2 I366 (internal_0n[66], internal_0n[62], internal_0n[63]);
  C2 I367 (internal_0n[67], internal_0n[64], internal_0n[65]);
  C2 I368 (selcomp_1n, internal_0n[66], internal_0n[67]);
  OR2 I369 (complete852_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I370 (complete852_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I371 (complete852_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I372 (complete852_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I373 (complete852_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I374 (complete852_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I375 (complete852_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I376 (complete852_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I377 (complete852_0n[8], ifint_1n[8], itint_1n[8]);
  OR2 I378 (complete852_0n[9], ifint_1n[9], itint_1n[9]);
  OR2 I379 (complete852_0n[10], ifint_1n[10], itint_1n[10]);
  OR2 I380 (complete852_0n[11], ifint_1n[11], itint_1n[11]);
  OR2 I381 (complete852_0n[12], ifint_1n[12], itint_1n[12]);
  OR2 I382 (complete852_0n[13], ifint_1n[13], itint_1n[13]);
  OR2 I383 (complete852_0n[14], ifint_1n[14], itint_1n[14]);
  OR2 I384 (complete852_0n[15], ifint_1n[15], itint_1n[15]);
  OR2 I385 (complete852_0n[16], ifint_1n[16], itint_1n[16]);
  OR2 I386 (complete852_0n[17], ifint_1n[17], itint_1n[17]);
  OR2 I387 (complete852_0n[18], ifint_1n[18], itint_1n[18]);
  OR2 I388 (complete852_0n[19], ifint_1n[19], itint_1n[19]);
  OR2 I389 (complete852_0n[20], ifint_1n[20], itint_1n[20]);
  OR2 I390 (complete852_0n[21], ifint_1n[21], itint_1n[21]);
  OR2 I391 (complete852_0n[22], ifint_1n[22], itint_1n[22]);
  OR2 I392 (complete852_0n[23], ifint_1n[23], itint_1n[23]);
  OR2 I393 (complete852_0n[24], ifint_1n[24], itint_1n[24]);
  OR2 I394 (complete852_0n[25], ifint_1n[25], itint_1n[25]);
  OR2 I395 (complete852_0n[26], ifint_1n[26], itint_1n[26]);
  OR2 I396 (complete852_0n[27], ifint_1n[27], itint_1n[27]);
  OR2 I397 (complete852_0n[28], ifint_1n[28], itint_1n[28]);
  OR2 I398 (complete852_0n[29], ifint_1n[29], itint_1n[29]);
  OR2 I399 (complete852_0n[30], ifint_1n[30], itint_1n[30]);
  OR2 I400 (complete852_0n[31], ifint_1n[31], itint_1n[31]);
  C3 I401 (internal_0n[68], complete851_0n[0], complete851_0n[1], complete851_0n[2]);
  C3 I402 (internal_0n[69], complete851_0n[3], complete851_0n[4], complete851_0n[5]);
  C3 I403 (internal_0n[70], complete851_0n[6], complete851_0n[7], complete851_0n[8]);
  C3 I404 (internal_0n[71], complete851_0n[9], complete851_0n[10], complete851_0n[11]);
  C3 I405 (internal_0n[72], complete851_0n[12], complete851_0n[13], complete851_0n[14]);
  C3 I406 (internal_0n[73], complete851_0n[15], complete851_0n[16], complete851_0n[17]);
  C3 I407 (internal_0n[74], complete851_0n[18], complete851_0n[19], complete851_0n[20]);
  C3 I408 (internal_0n[75], complete851_0n[21], complete851_0n[22], complete851_0n[23]);
  C3 I409 (internal_0n[76], complete851_0n[24], complete851_0n[25], complete851_0n[26]);
  C3 I410 (internal_0n[77], complete851_0n[27], complete851_0n[28], complete851_0n[29]);
  C2 I411 (internal_0n[78], complete851_0n[30], complete851_0n[31]);
  C3 I412 (internal_0n[79], internal_0n[68], internal_0n[69], internal_0n[70]);
  C3 I413 (internal_0n[80], internal_0n[71], internal_0n[72], internal_0n[73]);
  C3 I414 (internal_0n[81], internal_0n[74], internal_0n[75], internal_0n[76]);
  C2 I415 (internal_0n[82], internal_0n[77], internal_0n[78]);
  C2 I416 (internal_0n[83], internal_0n[79], internal_0n[80]);
  C2 I417 (internal_0n[84], internal_0n[81], internal_0n[82]);
  C2 I418 (selcomp_0n, internal_0n[83], internal_0n[84]);
  OR2 I419 (complete851_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I420 (complete851_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I421 (complete851_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I422 (complete851_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I423 (complete851_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I424 (complete851_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I425 (complete851_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I426 (complete851_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I427 (complete851_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I428 (complete851_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I429 (complete851_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I430 (complete851_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I431 (complete851_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I432 (complete851_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I433 (complete851_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I434 (complete851_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I435 (complete851_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I436 (complete851_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I437 (complete851_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I438 (complete851_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I439 (complete851_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I440 (complete851_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I441 (complete851_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I442 (complete851_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I443 (complete851_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I444 (complete851_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I445 (complete851_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I446 (complete851_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I447 (complete851_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I448 (complete851_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I449 (complete851_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I450 (complete851_0n[31], ifint_0n[31], itint_0n[31]);
  AND2 I451 (gfint_0n[0], gate_0n[0], ifint_0n[0]);
  AND2 I452 (gfint_0n[1], gate_0n[0], ifint_0n[1]);
  AND2 I453 (gfint_0n[2], gate_0n[0], ifint_0n[2]);
  AND2 I454 (gfint_0n[3], gate_0n[0], ifint_0n[3]);
  AND2 I455 (gfint_0n[4], gate_0n[0], ifint_0n[4]);
  AND2 I456 (gfint_0n[5], gate_0n[0], ifint_0n[5]);
  AND2 I457 (gfint_0n[6], gate_0n[0], ifint_0n[6]);
  AND2 I458 (gfint_0n[7], gate_0n[0], ifint_0n[7]);
  AND2 I459 (gfint_0n[8], gate_0n[0], ifint_0n[8]);
  AND2 I460 (gfint_0n[9], gate_0n[0], ifint_0n[9]);
  AND2 I461 (gfint_0n[10], gate_0n[0], ifint_0n[10]);
  AND2 I462 (gfint_0n[11], gate_0n[0], ifint_0n[11]);
  AND2 I463 (gfint_0n[12], gate_0n[0], ifint_0n[12]);
  AND2 I464 (gfint_0n[13], gate_0n[0], ifint_0n[13]);
  AND2 I465 (gfint_0n[14], gate_0n[0], ifint_0n[14]);
  AND2 I466 (gfint_0n[15], gate_0n[0], ifint_0n[15]);
  AND2 I467 (gfint_0n[16], gate_0n[0], ifint_0n[16]);
  AND2 I468 (gfint_0n[17], gate_0n[0], ifint_0n[17]);
  AND2 I469 (gfint_0n[18], gate_0n[0], ifint_0n[18]);
  AND2 I470 (gfint_0n[19], gate_0n[0], ifint_0n[19]);
  AND2 I471 (gfint_0n[20], gate_0n[0], ifint_0n[20]);
  AND2 I472 (gfint_0n[21], gate_0n[0], ifint_0n[21]);
  AND2 I473 (gfint_0n[22], gate_0n[0], ifint_0n[22]);
  AND2 I474 (gfint_0n[23], gate_0n[0], ifint_0n[23]);
  AND2 I475 (gfint_0n[24], gate_0n[0], ifint_0n[24]);
  AND2 I476 (gfint_0n[25], gate_0n[0], ifint_0n[25]);
  AND2 I477 (gfint_0n[26], gate_0n[0], ifint_0n[26]);
  AND2 I478 (gfint_0n[27], gate_0n[0], ifint_0n[27]);
  AND2 I479 (gfint_0n[28], gate_0n[0], ifint_0n[28]);
  AND2 I480 (gfint_0n[29], gate_0n[0], ifint_0n[29]);
  AND2 I481 (gfint_0n[30], gate_0n[0], ifint_0n[30]);
  AND2 I482 (gfint_0n[31], gate_0n[0], ifint_0n[31]);
  AND2 I483 (gfint_1n[0], gate_0n[1], ifint_1n[0]);
  AND2 I484 (gfint_1n[1], gate_0n[1], ifint_1n[1]);
  AND2 I485 (gfint_1n[2], gate_0n[1], ifint_1n[2]);
  AND2 I486 (gfint_1n[3], gate_0n[1], ifint_1n[3]);
  AND2 I487 (gfint_1n[4], gate_0n[1], ifint_1n[4]);
  AND2 I488 (gfint_1n[5], gate_0n[1], ifint_1n[5]);
  AND2 I489 (gfint_1n[6], gate_0n[1], ifint_1n[6]);
  AND2 I490 (gfint_1n[7], gate_0n[1], ifint_1n[7]);
  AND2 I491 (gfint_1n[8], gate_0n[1], ifint_1n[8]);
  AND2 I492 (gfint_1n[9], gate_0n[1], ifint_1n[9]);
  AND2 I493 (gfint_1n[10], gate_0n[1], ifint_1n[10]);
  AND2 I494 (gfint_1n[11], gate_0n[1], ifint_1n[11]);
  AND2 I495 (gfint_1n[12], gate_0n[1], ifint_1n[12]);
  AND2 I496 (gfint_1n[13], gate_0n[1], ifint_1n[13]);
  AND2 I497 (gfint_1n[14], gate_0n[1], ifint_1n[14]);
  AND2 I498 (gfint_1n[15], gate_0n[1], ifint_1n[15]);
  AND2 I499 (gfint_1n[16], gate_0n[1], ifint_1n[16]);
  AND2 I500 (gfint_1n[17], gate_0n[1], ifint_1n[17]);
  AND2 I501 (gfint_1n[18], gate_0n[1], ifint_1n[18]);
  AND2 I502 (gfint_1n[19], gate_0n[1], ifint_1n[19]);
  AND2 I503 (gfint_1n[20], gate_0n[1], ifint_1n[20]);
  AND2 I504 (gfint_1n[21], gate_0n[1], ifint_1n[21]);
  AND2 I505 (gfint_1n[22], gate_0n[1], ifint_1n[22]);
  AND2 I506 (gfint_1n[23], gate_0n[1], ifint_1n[23]);
  AND2 I507 (gfint_1n[24], gate_0n[1], ifint_1n[24]);
  AND2 I508 (gfint_1n[25], gate_0n[1], ifint_1n[25]);
  AND2 I509 (gfint_1n[26], gate_0n[1], ifint_1n[26]);
  AND2 I510 (gfint_1n[27], gate_0n[1], ifint_1n[27]);
  AND2 I511 (gfint_1n[28], gate_0n[1], ifint_1n[28]);
  AND2 I512 (gfint_1n[29], gate_0n[1], ifint_1n[29]);
  AND2 I513 (gfint_1n[30], gate_0n[1], ifint_1n[30]);
  AND2 I514 (gfint_1n[31], gate_0n[1], ifint_1n[31]);
  AND2 I515 (gtint_0n[0], gate_0n[0], itint_0n[0]);
  AND2 I516 (gtint_0n[1], gate_0n[0], itint_0n[1]);
  AND2 I517 (gtint_0n[2], gate_0n[0], itint_0n[2]);
  AND2 I518 (gtint_0n[3], gate_0n[0], itint_0n[3]);
  AND2 I519 (gtint_0n[4], gate_0n[0], itint_0n[4]);
  AND2 I520 (gtint_0n[5], gate_0n[0], itint_0n[5]);
  AND2 I521 (gtint_0n[6], gate_0n[0], itint_0n[6]);
  AND2 I522 (gtint_0n[7], gate_0n[0], itint_0n[7]);
  AND2 I523 (gtint_0n[8], gate_0n[0], itint_0n[8]);
  AND2 I524 (gtint_0n[9], gate_0n[0], itint_0n[9]);
  AND2 I525 (gtint_0n[10], gate_0n[0], itint_0n[10]);
  AND2 I526 (gtint_0n[11], gate_0n[0], itint_0n[11]);
  AND2 I527 (gtint_0n[12], gate_0n[0], itint_0n[12]);
  AND2 I528 (gtint_0n[13], gate_0n[0], itint_0n[13]);
  AND2 I529 (gtint_0n[14], gate_0n[0], itint_0n[14]);
  AND2 I530 (gtint_0n[15], gate_0n[0], itint_0n[15]);
  AND2 I531 (gtint_0n[16], gate_0n[0], itint_0n[16]);
  AND2 I532 (gtint_0n[17], gate_0n[0], itint_0n[17]);
  AND2 I533 (gtint_0n[18], gate_0n[0], itint_0n[18]);
  AND2 I534 (gtint_0n[19], gate_0n[0], itint_0n[19]);
  AND2 I535 (gtint_0n[20], gate_0n[0], itint_0n[20]);
  AND2 I536 (gtint_0n[21], gate_0n[0], itint_0n[21]);
  AND2 I537 (gtint_0n[22], gate_0n[0], itint_0n[22]);
  AND2 I538 (gtint_0n[23], gate_0n[0], itint_0n[23]);
  AND2 I539 (gtint_0n[24], gate_0n[0], itint_0n[24]);
  AND2 I540 (gtint_0n[25], gate_0n[0], itint_0n[25]);
  AND2 I541 (gtint_0n[26], gate_0n[0], itint_0n[26]);
  AND2 I542 (gtint_0n[27], gate_0n[0], itint_0n[27]);
  AND2 I543 (gtint_0n[28], gate_0n[0], itint_0n[28]);
  AND2 I544 (gtint_0n[29], gate_0n[0], itint_0n[29]);
  AND2 I545 (gtint_0n[30], gate_0n[0], itint_0n[30]);
  AND2 I546 (gtint_0n[31], gate_0n[0], itint_0n[31]);
  AND2 I547 (gtint_1n[0], gate_0n[1], itint_1n[0]);
  AND2 I548 (gtint_1n[1], gate_0n[1], itint_1n[1]);
  AND2 I549 (gtint_1n[2], gate_0n[1], itint_1n[2]);
  AND2 I550 (gtint_1n[3], gate_0n[1], itint_1n[3]);
  AND2 I551 (gtint_1n[4], gate_0n[1], itint_1n[4]);
  AND2 I552 (gtint_1n[5], gate_0n[1], itint_1n[5]);
  AND2 I553 (gtint_1n[6], gate_0n[1], itint_1n[6]);
  AND2 I554 (gtint_1n[7], gate_0n[1], itint_1n[7]);
  AND2 I555 (gtint_1n[8], gate_0n[1], itint_1n[8]);
  AND2 I556 (gtint_1n[9], gate_0n[1], itint_1n[9]);
  AND2 I557 (gtint_1n[10], gate_0n[1], itint_1n[10]);
  AND2 I558 (gtint_1n[11], gate_0n[1], itint_1n[11]);
  AND2 I559 (gtint_1n[12], gate_0n[1], itint_1n[12]);
  AND2 I560 (gtint_1n[13], gate_0n[1], itint_1n[13]);
  AND2 I561 (gtint_1n[14], gate_0n[1], itint_1n[14]);
  AND2 I562 (gtint_1n[15], gate_0n[1], itint_1n[15]);
  AND2 I563 (gtint_1n[16], gate_0n[1], itint_1n[16]);
  AND2 I564 (gtint_1n[17], gate_0n[1], itint_1n[17]);
  AND2 I565 (gtint_1n[18], gate_0n[1], itint_1n[18]);
  AND2 I566 (gtint_1n[19], gate_0n[1], itint_1n[19]);
  AND2 I567 (gtint_1n[20], gate_0n[1], itint_1n[20]);
  AND2 I568 (gtint_1n[21], gate_0n[1], itint_1n[21]);
  AND2 I569 (gtint_1n[22], gate_0n[1], itint_1n[22]);
  AND2 I570 (gtint_1n[23], gate_0n[1], itint_1n[23]);
  AND2 I571 (gtint_1n[24], gate_0n[1], itint_1n[24]);
  AND2 I572 (gtint_1n[25], gate_0n[1], itint_1n[25]);
  AND2 I573 (gtint_1n[26], gate_0n[1], itint_1n[26]);
  AND2 I574 (gtint_1n[27], gate_0n[1], itint_1n[27]);
  AND2 I575 (gtint_1n[28], gate_0n[1], itint_1n[28]);
  AND2 I576 (gtint_1n[29], gate_0n[1], itint_1n[29]);
  AND2 I577 (gtint_1n[30], gate_0n[1], itint_1n[30]);
  AND2 I578 (gtint_1n[31], gate_0n[1], itint_1n[31]);
  OR2 I579 (otint_0n[0], gtint_0n[0], gtint_1n[0]);
  OR2 I580 (otint_0n[1], gtint_0n[1], gtint_1n[1]);
  OR2 I581 (otint_0n[2], gtint_0n[2], gtint_1n[2]);
  OR2 I582 (otint_0n[3], gtint_0n[3], gtint_1n[3]);
  OR2 I583 (otint_0n[4], gtint_0n[4], gtint_1n[4]);
  OR2 I584 (otint_0n[5], gtint_0n[5], gtint_1n[5]);
  OR2 I585 (otint_0n[6], gtint_0n[6], gtint_1n[6]);
  OR2 I586 (otint_0n[7], gtint_0n[7], gtint_1n[7]);
  OR2 I587 (otint_0n[8], gtint_0n[8], gtint_1n[8]);
  OR2 I588 (otint_0n[9], gtint_0n[9], gtint_1n[9]);
  OR2 I589 (otint_0n[10], gtint_0n[10], gtint_1n[10]);
  OR2 I590 (otint_0n[11], gtint_0n[11], gtint_1n[11]);
  OR2 I591 (otint_0n[12], gtint_0n[12], gtint_1n[12]);
  OR2 I592 (otint_0n[13], gtint_0n[13], gtint_1n[13]);
  OR2 I593 (otint_0n[14], gtint_0n[14], gtint_1n[14]);
  OR2 I594 (otint_0n[15], gtint_0n[15], gtint_1n[15]);
  OR2 I595 (otint_0n[16], gtint_0n[16], gtint_1n[16]);
  OR2 I596 (otint_0n[17], gtint_0n[17], gtint_1n[17]);
  OR2 I597 (otint_0n[18], gtint_0n[18], gtint_1n[18]);
  OR2 I598 (otint_0n[19], gtint_0n[19], gtint_1n[19]);
  OR2 I599 (otint_0n[20], gtint_0n[20], gtint_1n[20]);
  OR2 I600 (otint_0n[21], gtint_0n[21], gtint_1n[21]);
  OR2 I601 (otint_0n[22], gtint_0n[22], gtint_1n[22]);
  OR2 I602 (otint_0n[23], gtint_0n[23], gtint_1n[23]);
  OR2 I603 (otint_0n[24], gtint_0n[24], gtint_1n[24]);
  OR2 I604 (otint_0n[25], gtint_0n[25], gtint_1n[25]);
  OR2 I605 (otint_0n[26], gtint_0n[26], gtint_1n[26]);
  OR2 I606 (otint_0n[27], gtint_0n[27], gtint_1n[27]);
  OR2 I607 (otint_0n[28], gtint_0n[28], gtint_1n[28]);
  OR2 I608 (otint_0n[29], gtint_0n[29], gtint_1n[29]);
  OR2 I609 (otint_0n[30], gtint_0n[30], gtint_1n[30]);
  OR2 I610 (otint_0n[31], gtint_0n[31], gtint_1n[31]);
  OR2 I611 (ofint_0n[0], gfint_0n[0], gfint_1n[0]);
  OR2 I612 (ofint_0n[1], gfint_0n[1], gfint_1n[1]);
  OR2 I613 (ofint_0n[2], gfint_0n[2], gfint_1n[2]);
  OR2 I614 (ofint_0n[3], gfint_0n[3], gfint_1n[3]);
  OR2 I615 (ofint_0n[4], gfint_0n[4], gfint_1n[4]);
  OR2 I616 (ofint_0n[5], gfint_0n[5], gfint_1n[5]);
  OR2 I617 (ofint_0n[6], gfint_0n[6], gfint_1n[6]);
  OR2 I618 (ofint_0n[7], gfint_0n[7], gfint_1n[7]);
  OR2 I619 (ofint_0n[8], gfint_0n[8], gfint_1n[8]);
  OR2 I620 (ofint_0n[9], gfint_0n[9], gfint_1n[9]);
  OR2 I621 (ofint_0n[10], gfint_0n[10], gfint_1n[10]);
  OR2 I622 (ofint_0n[11], gfint_0n[11], gfint_1n[11]);
  OR2 I623 (ofint_0n[12], gfint_0n[12], gfint_1n[12]);
  OR2 I624 (ofint_0n[13], gfint_0n[13], gfint_1n[13]);
  OR2 I625 (ofint_0n[14], gfint_0n[14], gfint_1n[14]);
  OR2 I626 (ofint_0n[15], gfint_0n[15], gfint_1n[15]);
  OR2 I627 (ofint_0n[16], gfint_0n[16], gfint_1n[16]);
  OR2 I628 (ofint_0n[17], gfint_0n[17], gfint_1n[17]);
  OR2 I629 (ofint_0n[18], gfint_0n[18], gfint_1n[18]);
  OR2 I630 (ofint_0n[19], gfint_0n[19], gfint_1n[19]);
  OR2 I631 (ofint_0n[20], gfint_0n[20], gfint_1n[20]);
  OR2 I632 (ofint_0n[21], gfint_0n[21], gfint_1n[21]);
  OR2 I633 (ofint_0n[22], gfint_0n[22], gfint_1n[22]);
  OR2 I634 (ofint_0n[23], gfint_0n[23], gfint_1n[23]);
  OR2 I635 (ofint_0n[24], gfint_0n[24], gfint_1n[24]);
  OR2 I636 (ofint_0n[25], gfint_0n[25], gfint_1n[25]);
  OR2 I637 (ofint_0n[26], gfint_0n[26], gfint_1n[26]);
  OR2 I638 (ofint_0n[27], gfint_0n[27], gfint_1n[27]);
  OR2 I639 (ofint_0n[28], gfint_0n[28], gfint_1n[28]);
  OR2 I640 (ofint_0n[29], gfint_0n[29], gfint_1n[29]);
  OR2 I641 (ofint_0n[30], gfint_0n[30], gfint_1n[30]);
  OR2 I642 (ofint_0n[31], gfint_0n[31], gfint_1n[31]);
endmodule

module BrzM_32_3 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  i_2r0d, i_2r1d, i_2a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [31:0] i_0r0d;
  input [31:0] i_0r1d;
  output i_0a;
  input [31:0] i_1r0d;
  input [31:0] i_1r1d;
  output i_1a;
  input [31:0] i_2r0d;
  input [31:0] i_2r1d;
  output i_2a;
  output [31:0] o_0r0d;
  output [31:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [118:0] internal_0n;
  wire [2:0] sel_0n;
  wire [31:0] ofint_0n;
  wire [31:0] otint_0n;
  wire oaint_0n;
  wire [31:0] ifint_0n;
  wire [31:0] ifint_1n;
  wire [31:0] ifint_2n;
  wire [31:0] itint_0n;
  wire [31:0] itint_1n;
  wire [31:0] itint_2n;
  wire iaint_0n;
  wire iaint_1n;
  wire iaint_2n;
  wire [2:0] gate_0n;
  wire [31:0] gfint_0n;
  wire [31:0] gfint_1n;
  wire [31:0] gfint_2n;
  wire [31:0] gtint_0n;
  wire [31:0] gtint_1n;
  wire [31:0] gtint_2n;
  wire [31:0] complete883_0n;
  wire gate882_0n;
  wire [31:0] complete879_0n;
  wire gate878_0n;
  wire [31:0] complete875_0n;
  wire gate874_0n;
  wire [31:0] complete871_0n;
  wire gate870_0n;
  wire [31:0] complete867_0n;
  wire [31:0] complete866_0n;
  wire [31:0] complete865_0n;
  wire selcomp_0n;
  wire selcomp_1n;
  wire selcomp_2n;
  C3 I0 (internal_0n[0], complete883_0n[0], complete883_0n[1], complete883_0n[2]);
  C3 I1 (internal_0n[1], complete883_0n[3], complete883_0n[4], complete883_0n[5]);
  C3 I2 (internal_0n[2], complete883_0n[6], complete883_0n[7], complete883_0n[8]);
  C3 I3 (internal_0n[3], complete883_0n[9], complete883_0n[10], complete883_0n[11]);
  C3 I4 (internal_0n[4], complete883_0n[12], complete883_0n[13], complete883_0n[14]);
  C3 I5 (internal_0n[5], complete883_0n[15], complete883_0n[16], complete883_0n[17]);
  C3 I6 (internal_0n[6], complete883_0n[18], complete883_0n[19], complete883_0n[20]);
  C3 I7 (internal_0n[7], complete883_0n[21], complete883_0n[22], complete883_0n[23]);
  C3 I8 (internal_0n[8], complete883_0n[24], complete883_0n[25], complete883_0n[26]);
  C3 I9 (internal_0n[9], complete883_0n[27], complete883_0n[28], complete883_0n[29]);
  C2 I10 (internal_0n[10], complete883_0n[30], complete883_0n[31]);
  C3 I11 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I12 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I13 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I14 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I15 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I16 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I17 (i_2a, internal_0n[15], internal_0n[16]);
  OR2 I18 (complete883_0n[0], ifint_2n[0], itint_2n[0]);
  OR2 I19 (complete883_0n[1], ifint_2n[1], itint_2n[1]);
  OR2 I20 (complete883_0n[2], ifint_2n[2], itint_2n[2]);
  OR2 I21 (complete883_0n[3], ifint_2n[3], itint_2n[3]);
  OR2 I22 (complete883_0n[4], ifint_2n[4], itint_2n[4]);
  OR2 I23 (complete883_0n[5], ifint_2n[5], itint_2n[5]);
  OR2 I24 (complete883_0n[6], ifint_2n[6], itint_2n[6]);
  OR2 I25 (complete883_0n[7], ifint_2n[7], itint_2n[7]);
  OR2 I26 (complete883_0n[8], ifint_2n[8], itint_2n[8]);
  OR2 I27 (complete883_0n[9], ifint_2n[9], itint_2n[9]);
  OR2 I28 (complete883_0n[10], ifint_2n[10], itint_2n[10]);
  OR2 I29 (complete883_0n[11], ifint_2n[11], itint_2n[11]);
  OR2 I30 (complete883_0n[12], ifint_2n[12], itint_2n[12]);
  OR2 I31 (complete883_0n[13], ifint_2n[13], itint_2n[13]);
  OR2 I32 (complete883_0n[14], ifint_2n[14], itint_2n[14]);
  OR2 I33 (complete883_0n[15], ifint_2n[15], itint_2n[15]);
  OR2 I34 (complete883_0n[16], ifint_2n[16], itint_2n[16]);
  OR2 I35 (complete883_0n[17], ifint_2n[17], itint_2n[17]);
  OR2 I36 (complete883_0n[18], ifint_2n[18], itint_2n[18]);
  OR2 I37 (complete883_0n[19], ifint_2n[19], itint_2n[19]);
  OR2 I38 (complete883_0n[20], ifint_2n[20], itint_2n[20]);
  OR2 I39 (complete883_0n[21], ifint_2n[21], itint_2n[21]);
  OR2 I40 (complete883_0n[22], ifint_2n[22], itint_2n[22]);
  OR2 I41 (complete883_0n[23], ifint_2n[23], itint_2n[23]);
  OR2 I42 (complete883_0n[24], ifint_2n[24], itint_2n[24]);
  OR2 I43 (complete883_0n[25], ifint_2n[25], itint_2n[25]);
  OR2 I44 (complete883_0n[26], ifint_2n[26], itint_2n[26]);
  OR2 I45 (complete883_0n[27], ifint_2n[27], itint_2n[27]);
  OR2 I46 (complete883_0n[28], ifint_2n[28], itint_2n[28]);
  OR2 I47 (complete883_0n[29], ifint_2n[29], itint_2n[29]);
  OR2 I48 (complete883_0n[30], ifint_2n[30], itint_2n[30]);
  OR2 I49 (complete883_0n[31], ifint_2n[31], itint_2n[31]);
  INV I50 (gate882_0n, iaint_2n);
  C2RI I51 (itint_2n[0], i_2r1d[0], gate882_0n, initialise);
  C2RI I52 (itint_2n[1], i_2r1d[1], gate882_0n, initialise);
  C2RI I53 (itint_2n[2], i_2r1d[2], gate882_0n, initialise);
  C2RI I54 (itint_2n[3], i_2r1d[3], gate882_0n, initialise);
  C2RI I55 (itint_2n[4], i_2r1d[4], gate882_0n, initialise);
  C2RI I56 (itint_2n[5], i_2r1d[5], gate882_0n, initialise);
  C2RI I57 (itint_2n[6], i_2r1d[6], gate882_0n, initialise);
  C2RI I58 (itint_2n[7], i_2r1d[7], gate882_0n, initialise);
  C2RI I59 (itint_2n[8], i_2r1d[8], gate882_0n, initialise);
  C2RI I60 (itint_2n[9], i_2r1d[9], gate882_0n, initialise);
  C2RI I61 (itint_2n[10], i_2r1d[10], gate882_0n, initialise);
  C2RI I62 (itint_2n[11], i_2r1d[11], gate882_0n, initialise);
  C2RI I63 (itint_2n[12], i_2r1d[12], gate882_0n, initialise);
  C2RI I64 (itint_2n[13], i_2r1d[13], gate882_0n, initialise);
  C2RI I65 (itint_2n[14], i_2r1d[14], gate882_0n, initialise);
  C2RI I66 (itint_2n[15], i_2r1d[15], gate882_0n, initialise);
  C2RI I67 (itint_2n[16], i_2r1d[16], gate882_0n, initialise);
  C2RI I68 (itint_2n[17], i_2r1d[17], gate882_0n, initialise);
  C2RI I69 (itint_2n[18], i_2r1d[18], gate882_0n, initialise);
  C2RI I70 (itint_2n[19], i_2r1d[19], gate882_0n, initialise);
  C2RI I71 (itint_2n[20], i_2r1d[20], gate882_0n, initialise);
  C2RI I72 (itint_2n[21], i_2r1d[21], gate882_0n, initialise);
  C2RI I73 (itint_2n[22], i_2r1d[22], gate882_0n, initialise);
  C2RI I74 (itint_2n[23], i_2r1d[23], gate882_0n, initialise);
  C2RI I75 (itint_2n[24], i_2r1d[24], gate882_0n, initialise);
  C2RI I76 (itint_2n[25], i_2r1d[25], gate882_0n, initialise);
  C2RI I77 (itint_2n[26], i_2r1d[26], gate882_0n, initialise);
  C2RI I78 (itint_2n[27], i_2r1d[27], gate882_0n, initialise);
  C2RI I79 (itint_2n[28], i_2r1d[28], gate882_0n, initialise);
  C2RI I80 (itint_2n[29], i_2r1d[29], gate882_0n, initialise);
  C2RI I81 (itint_2n[30], i_2r1d[30], gate882_0n, initialise);
  C2RI I82 (itint_2n[31], i_2r1d[31], gate882_0n, initialise);
  C2RI I83 (ifint_2n[0], i_2r0d[0], gate882_0n, initialise);
  C2RI I84 (ifint_2n[1], i_2r0d[1], gate882_0n, initialise);
  C2RI I85 (ifint_2n[2], i_2r0d[2], gate882_0n, initialise);
  C2RI I86 (ifint_2n[3], i_2r0d[3], gate882_0n, initialise);
  C2RI I87 (ifint_2n[4], i_2r0d[4], gate882_0n, initialise);
  C2RI I88 (ifint_2n[5], i_2r0d[5], gate882_0n, initialise);
  C2RI I89 (ifint_2n[6], i_2r0d[6], gate882_0n, initialise);
  C2RI I90 (ifint_2n[7], i_2r0d[7], gate882_0n, initialise);
  C2RI I91 (ifint_2n[8], i_2r0d[8], gate882_0n, initialise);
  C2RI I92 (ifint_2n[9], i_2r0d[9], gate882_0n, initialise);
  C2RI I93 (ifint_2n[10], i_2r0d[10], gate882_0n, initialise);
  C2RI I94 (ifint_2n[11], i_2r0d[11], gate882_0n, initialise);
  C2RI I95 (ifint_2n[12], i_2r0d[12], gate882_0n, initialise);
  C2RI I96 (ifint_2n[13], i_2r0d[13], gate882_0n, initialise);
  C2RI I97 (ifint_2n[14], i_2r0d[14], gate882_0n, initialise);
  C2RI I98 (ifint_2n[15], i_2r0d[15], gate882_0n, initialise);
  C2RI I99 (ifint_2n[16], i_2r0d[16], gate882_0n, initialise);
  C2RI I100 (ifint_2n[17], i_2r0d[17], gate882_0n, initialise);
  C2RI I101 (ifint_2n[18], i_2r0d[18], gate882_0n, initialise);
  C2RI I102 (ifint_2n[19], i_2r0d[19], gate882_0n, initialise);
  C2RI I103 (ifint_2n[20], i_2r0d[20], gate882_0n, initialise);
  C2RI I104 (ifint_2n[21], i_2r0d[21], gate882_0n, initialise);
  C2RI I105 (ifint_2n[22], i_2r0d[22], gate882_0n, initialise);
  C2RI I106 (ifint_2n[23], i_2r0d[23], gate882_0n, initialise);
  C2RI I107 (ifint_2n[24], i_2r0d[24], gate882_0n, initialise);
  C2RI I108 (ifint_2n[25], i_2r0d[25], gate882_0n, initialise);
  C2RI I109 (ifint_2n[26], i_2r0d[26], gate882_0n, initialise);
  C2RI I110 (ifint_2n[27], i_2r0d[27], gate882_0n, initialise);
  C2RI I111 (ifint_2n[28], i_2r0d[28], gate882_0n, initialise);
  C2RI I112 (ifint_2n[29], i_2r0d[29], gate882_0n, initialise);
  C2RI I113 (ifint_2n[30], i_2r0d[30], gate882_0n, initialise);
  C2RI I114 (ifint_2n[31], i_2r0d[31], gate882_0n, initialise);
  C3 I115 (internal_0n[17], complete879_0n[0], complete879_0n[1], complete879_0n[2]);
  C3 I116 (internal_0n[18], complete879_0n[3], complete879_0n[4], complete879_0n[5]);
  C3 I117 (internal_0n[19], complete879_0n[6], complete879_0n[7], complete879_0n[8]);
  C3 I118 (internal_0n[20], complete879_0n[9], complete879_0n[10], complete879_0n[11]);
  C3 I119 (internal_0n[21], complete879_0n[12], complete879_0n[13], complete879_0n[14]);
  C3 I120 (internal_0n[22], complete879_0n[15], complete879_0n[16], complete879_0n[17]);
  C3 I121 (internal_0n[23], complete879_0n[18], complete879_0n[19], complete879_0n[20]);
  C3 I122 (internal_0n[24], complete879_0n[21], complete879_0n[22], complete879_0n[23]);
  C3 I123 (internal_0n[25], complete879_0n[24], complete879_0n[25], complete879_0n[26]);
  C3 I124 (internal_0n[26], complete879_0n[27], complete879_0n[28], complete879_0n[29]);
  C2 I125 (internal_0n[27], complete879_0n[30], complete879_0n[31]);
  C3 I126 (internal_0n[28], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I127 (internal_0n[29], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I128 (internal_0n[30], internal_0n[23], internal_0n[24], internal_0n[25]);
  C2 I129 (internal_0n[31], internal_0n[26], internal_0n[27]);
  C2 I130 (internal_0n[32], internal_0n[28], internal_0n[29]);
  C2 I131 (internal_0n[33], internal_0n[30], internal_0n[31]);
  C2 I132 (i_1a, internal_0n[32], internal_0n[33]);
  OR2 I133 (complete879_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I134 (complete879_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I135 (complete879_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I136 (complete879_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I137 (complete879_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I138 (complete879_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I139 (complete879_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I140 (complete879_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I141 (complete879_0n[8], ifint_1n[8], itint_1n[8]);
  OR2 I142 (complete879_0n[9], ifint_1n[9], itint_1n[9]);
  OR2 I143 (complete879_0n[10], ifint_1n[10], itint_1n[10]);
  OR2 I144 (complete879_0n[11], ifint_1n[11], itint_1n[11]);
  OR2 I145 (complete879_0n[12], ifint_1n[12], itint_1n[12]);
  OR2 I146 (complete879_0n[13], ifint_1n[13], itint_1n[13]);
  OR2 I147 (complete879_0n[14], ifint_1n[14], itint_1n[14]);
  OR2 I148 (complete879_0n[15], ifint_1n[15], itint_1n[15]);
  OR2 I149 (complete879_0n[16], ifint_1n[16], itint_1n[16]);
  OR2 I150 (complete879_0n[17], ifint_1n[17], itint_1n[17]);
  OR2 I151 (complete879_0n[18], ifint_1n[18], itint_1n[18]);
  OR2 I152 (complete879_0n[19], ifint_1n[19], itint_1n[19]);
  OR2 I153 (complete879_0n[20], ifint_1n[20], itint_1n[20]);
  OR2 I154 (complete879_0n[21], ifint_1n[21], itint_1n[21]);
  OR2 I155 (complete879_0n[22], ifint_1n[22], itint_1n[22]);
  OR2 I156 (complete879_0n[23], ifint_1n[23], itint_1n[23]);
  OR2 I157 (complete879_0n[24], ifint_1n[24], itint_1n[24]);
  OR2 I158 (complete879_0n[25], ifint_1n[25], itint_1n[25]);
  OR2 I159 (complete879_0n[26], ifint_1n[26], itint_1n[26]);
  OR2 I160 (complete879_0n[27], ifint_1n[27], itint_1n[27]);
  OR2 I161 (complete879_0n[28], ifint_1n[28], itint_1n[28]);
  OR2 I162 (complete879_0n[29], ifint_1n[29], itint_1n[29]);
  OR2 I163 (complete879_0n[30], ifint_1n[30], itint_1n[30]);
  OR2 I164 (complete879_0n[31], ifint_1n[31], itint_1n[31]);
  INV I165 (gate878_0n, iaint_1n);
  C2RI I166 (itint_1n[0], i_1r1d[0], gate878_0n, initialise);
  C2RI I167 (itint_1n[1], i_1r1d[1], gate878_0n, initialise);
  C2RI I168 (itint_1n[2], i_1r1d[2], gate878_0n, initialise);
  C2RI I169 (itint_1n[3], i_1r1d[3], gate878_0n, initialise);
  C2RI I170 (itint_1n[4], i_1r1d[4], gate878_0n, initialise);
  C2RI I171 (itint_1n[5], i_1r1d[5], gate878_0n, initialise);
  C2RI I172 (itint_1n[6], i_1r1d[6], gate878_0n, initialise);
  C2RI I173 (itint_1n[7], i_1r1d[7], gate878_0n, initialise);
  C2RI I174 (itint_1n[8], i_1r1d[8], gate878_0n, initialise);
  C2RI I175 (itint_1n[9], i_1r1d[9], gate878_0n, initialise);
  C2RI I176 (itint_1n[10], i_1r1d[10], gate878_0n, initialise);
  C2RI I177 (itint_1n[11], i_1r1d[11], gate878_0n, initialise);
  C2RI I178 (itint_1n[12], i_1r1d[12], gate878_0n, initialise);
  C2RI I179 (itint_1n[13], i_1r1d[13], gate878_0n, initialise);
  C2RI I180 (itint_1n[14], i_1r1d[14], gate878_0n, initialise);
  C2RI I181 (itint_1n[15], i_1r1d[15], gate878_0n, initialise);
  C2RI I182 (itint_1n[16], i_1r1d[16], gate878_0n, initialise);
  C2RI I183 (itint_1n[17], i_1r1d[17], gate878_0n, initialise);
  C2RI I184 (itint_1n[18], i_1r1d[18], gate878_0n, initialise);
  C2RI I185 (itint_1n[19], i_1r1d[19], gate878_0n, initialise);
  C2RI I186 (itint_1n[20], i_1r1d[20], gate878_0n, initialise);
  C2RI I187 (itint_1n[21], i_1r1d[21], gate878_0n, initialise);
  C2RI I188 (itint_1n[22], i_1r1d[22], gate878_0n, initialise);
  C2RI I189 (itint_1n[23], i_1r1d[23], gate878_0n, initialise);
  C2RI I190 (itint_1n[24], i_1r1d[24], gate878_0n, initialise);
  C2RI I191 (itint_1n[25], i_1r1d[25], gate878_0n, initialise);
  C2RI I192 (itint_1n[26], i_1r1d[26], gate878_0n, initialise);
  C2RI I193 (itint_1n[27], i_1r1d[27], gate878_0n, initialise);
  C2RI I194 (itint_1n[28], i_1r1d[28], gate878_0n, initialise);
  C2RI I195 (itint_1n[29], i_1r1d[29], gate878_0n, initialise);
  C2RI I196 (itint_1n[30], i_1r1d[30], gate878_0n, initialise);
  C2RI I197 (itint_1n[31], i_1r1d[31], gate878_0n, initialise);
  C2RI I198 (ifint_1n[0], i_1r0d[0], gate878_0n, initialise);
  C2RI I199 (ifint_1n[1], i_1r0d[1], gate878_0n, initialise);
  C2RI I200 (ifint_1n[2], i_1r0d[2], gate878_0n, initialise);
  C2RI I201 (ifint_1n[3], i_1r0d[3], gate878_0n, initialise);
  C2RI I202 (ifint_1n[4], i_1r0d[4], gate878_0n, initialise);
  C2RI I203 (ifint_1n[5], i_1r0d[5], gate878_0n, initialise);
  C2RI I204 (ifint_1n[6], i_1r0d[6], gate878_0n, initialise);
  C2RI I205 (ifint_1n[7], i_1r0d[7], gate878_0n, initialise);
  C2RI I206 (ifint_1n[8], i_1r0d[8], gate878_0n, initialise);
  C2RI I207 (ifint_1n[9], i_1r0d[9], gate878_0n, initialise);
  C2RI I208 (ifint_1n[10], i_1r0d[10], gate878_0n, initialise);
  C2RI I209 (ifint_1n[11], i_1r0d[11], gate878_0n, initialise);
  C2RI I210 (ifint_1n[12], i_1r0d[12], gate878_0n, initialise);
  C2RI I211 (ifint_1n[13], i_1r0d[13], gate878_0n, initialise);
  C2RI I212 (ifint_1n[14], i_1r0d[14], gate878_0n, initialise);
  C2RI I213 (ifint_1n[15], i_1r0d[15], gate878_0n, initialise);
  C2RI I214 (ifint_1n[16], i_1r0d[16], gate878_0n, initialise);
  C2RI I215 (ifint_1n[17], i_1r0d[17], gate878_0n, initialise);
  C2RI I216 (ifint_1n[18], i_1r0d[18], gate878_0n, initialise);
  C2RI I217 (ifint_1n[19], i_1r0d[19], gate878_0n, initialise);
  C2RI I218 (ifint_1n[20], i_1r0d[20], gate878_0n, initialise);
  C2RI I219 (ifint_1n[21], i_1r0d[21], gate878_0n, initialise);
  C2RI I220 (ifint_1n[22], i_1r0d[22], gate878_0n, initialise);
  C2RI I221 (ifint_1n[23], i_1r0d[23], gate878_0n, initialise);
  C2RI I222 (ifint_1n[24], i_1r0d[24], gate878_0n, initialise);
  C2RI I223 (ifint_1n[25], i_1r0d[25], gate878_0n, initialise);
  C2RI I224 (ifint_1n[26], i_1r0d[26], gate878_0n, initialise);
  C2RI I225 (ifint_1n[27], i_1r0d[27], gate878_0n, initialise);
  C2RI I226 (ifint_1n[28], i_1r0d[28], gate878_0n, initialise);
  C2RI I227 (ifint_1n[29], i_1r0d[29], gate878_0n, initialise);
  C2RI I228 (ifint_1n[30], i_1r0d[30], gate878_0n, initialise);
  C2RI I229 (ifint_1n[31], i_1r0d[31], gate878_0n, initialise);
  C3 I230 (internal_0n[34], complete875_0n[0], complete875_0n[1], complete875_0n[2]);
  C3 I231 (internal_0n[35], complete875_0n[3], complete875_0n[4], complete875_0n[5]);
  C3 I232 (internal_0n[36], complete875_0n[6], complete875_0n[7], complete875_0n[8]);
  C3 I233 (internal_0n[37], complete875_0n[9], complete875_0n[10], complete875_0n[11]);
  C3 I234 (internal_0n[38], complete875_0n[12], complete875_0n[13], complete875_0n[14]);
  C3 I235 (internal_0n[39], complete875_0n[15], complete875_0n[16], complete875_0n[17]);
  C3 I236 (internal_0n[40], complete875_0n[18], complete875_0n[19], complete875_0n[20]);
  C3 I237 (internal_0n[41], complete875_0n[21], complete875_0n[22], complete875_0n[23]);
  C3 I238 (internal_0n[42], complete875_0n[24], complete875_0n[25], complete875_0n[26]);
  C3 I239 (internal_0n[43], complete875_0n[27], complete875_0n[28], complete875_0n[29]);
  C2 I240 (internal_0n[44], complete875_0n[30], complete875_0n[31]);
  C3 I241 (internal_0n[45], internal_0n[34], internal_0n[35], internal_0n[36]);
  C3 I242 (internal_0n[46], internal_0n[37], internal_0n[38], internal_0n[39]);
  C3 I243 (internal_0n[47], internal_0n[40], internal_0n[41], internal_0n[42]);
  C2 I244 (internal_0n[48], internal_0n[43], internal_0n[44]);
  C2 I245 (internal_0n[49], internal_0n[45], internal_0n[46]);
  C2 I246 (internal_0n[50], internal_0n[47], internal_0n[48]);
  C2 I247 (i_0a, internal_0n[49], internal_0n[50]);
  OR2 I248 (complete875_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I249 (complete875_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I250 (complete875_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I251 (complete875_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I252 (complete875_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I253 (complete875_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I254 (complete875_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I255 (complete875_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I256 (complete875_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I257 (complete875_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I258 (complete875_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I259 (complete875_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I260 (complete875_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I261 (complete875_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I262 (complete875_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I263 (complete875_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I264 (complete875_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I265 (complete875_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I266 (complete875_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I267 (complete875_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I268 (complete875_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I269 (complete875_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I270 (complete875_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I271 (complete875_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I272 (complete875_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I273 (complete875_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I274 (complete875_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I275 (complete875_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I276 (complete875_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I277 (complete875_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I278 (complete875_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I279 (complete875_0n[31], ifint_0n[31], itint_0n[31]);
  INV I280 (gate874_0n, iaint_0n);
  C2RI I281 (itint_0n[0], i_0r1d[0], gate874_0n, initialise);
  C2RI I282 (itint_0n[1], i_0r1d[1], gate874_0n, initialise);
  C2RI I283 (itint_0n[2], i_0r1d[2], gate874_0n, initialise);
  C2RI I284 (itint_0n[3], i_0r1d[3], gate874_0n, initialise);
  C2RI I285 (itint_0n[4], i_0r1d[4], gate874_0n, initialise);
  C2RI I286 (itint_0n[5], i_0r1d[5], gate874_0n, initialise);
  C2RI I287 (itint_0n[6], i_0r1d[6], gate874_0n, initialise);
  C2RI I288 (itint_0n[7], i_0r1d[7], gate874_0n, initialise);
  C2RI I289 (itint_0n[8], i_0r1d[8], gate874_0n, initialise);
  C2RI I290 (itint_0n[9], i_0r1d[9], gate874_0n, initialise);
  C2RI I291 (itint_0n[10], i_0r1d[10], gate874_0n, initialise);
  C2RI I292 (itint_0n[11], i_0r1d[11], gate874_0n, initialise);
  C2RI I293 (itint_0n[12], i_0r1d[12], gate874_0n, initialise);
  C2RI I294 (itint_0n[13], i_0r1d[13], gate874_0n, initialise);
  C2RI I295 (itint_0n[14], i_0r1d[14], gate874_0n, initialise);
  C2RI I296 (itint_0n[15], i_0r1d[15], gate874_0n, initialise);
  C2RI I297 (itint_0n[16], i_0r1d[16], gate874_0n, initialise);
  C2RI I298 (itint_0n[17], i_0r1d[17], gate874_0n, initialise);
  C2RI I299 (itint_0n[18], i_0r1d[18], gate874_0n, initialise);
  C2RI I300 (itint_0n[19], i_0r1d[19], gate874_0n, initialise);
  C2RI I301 (itint_0n[20], i_0r1d[20], gate874_0n, initialise);
  C2RI I302 (itint_0n[21], i_0r1d[21], gate874_0n, initialise);
  C2RI I303 (itint_0n[22], i_0r1d[22], gate874_0n, initialise);
  C2RI I304 (itint_0n[23], i_0r1d[23], gate874_0n, initialise);
  C2RI I305 (itint_0n[24], i_0r1d[24], gate874_0n, initialise);
  C2RI I306 (itint_0n[25], i_0r1d[25], gate874_0n, initialise);
  C2RI I307 (itint_0n[26], i_0r1d[26], gate874_0n, initialise);
  C2RI I308 (itint_0n[27], i_0r1d[27], gate874_0n, initialise);
  C2RI I309 (itint_0n[28], i_0r1d[28], gate874_0n, initialise);
  C2RI I310 (itint_0n[29], i_0r1d[29], gate874_0n, initialise);
  C2RI I311 (itint_0n[30], i_0r1d[30], gate874_0n, initialise);
  C2RI I312 (itint_0n[31], i_0r1d[31], gate874_0n, initialise);
  C2RI I313 (ifint_0n[0], i_0r0d[0], gate874_0n, initialise);
  C2RI I314 (ifint_0n[1], i_0r0d[1], gate874_0n, initialise);
  C2RI I315 (ifint_0n[2], i_0r0d[2], gate874_0n, initialise);
  C2RI I316 (ifint_0n[3], i_0r0d[3], gate874_0n, initialise);
  C2RI I317 (ifint_0n[4], i_0r0d[4], gate874_0n, initialise);
  C2RI I318 (ifint_0n[5], i_0r0d[5], gate874_0n, initialise);
  C2RI I319 (ifint_0n[6], i_0r0d[6], gate874_0n, initialise);
  C2RI I320 (ifint_0n[7], i_0r0d[7], gate874_0n, initialise);
  C2RI I321 (ifint_0n[8], i_0r0d[8], gate874_0n, initialise);
  C2RI I322 (ifint_0n[9], i_0r0d[9], gate874_0n, initialise);
  C2RI I323 (ifint_0n[10], i_0r0d[10], gate874_0n, initialise);
  C2RI I324 (ifint_0n[11], i_0r0d[11], gate874_0n, initialise);
  C2RI I325 (ifint_0n[12], i_0r0d[12], gate874_0n, initialise);
  C2RI I326 (ifint_0n[13], i_0r0d[13], gate874_0n, initialise);
  C2RI I327 (ifint_0n[14], i_0r0d[14], gate874_0n, initialise);
  C2RI I328 (ifint_0n[15], i_0r0d[15], gate874_0n, initialise);
  C2RI I329 (ifint_0n[16], i_0r0d[16], gate874_0n, initialise);
  C2RI I330 (ifint_0n[17], i_0r0d[17], gate874_0n, initialise);
  C2RI I331 (ifint_0n[18], i_0r0d[18], gate874_0n, initialise);
  C2RI I332 (ifint_0n[19], i_0r0d[19], gate874_0n, initialise);
  C2RI I333 (ifint_0n[20], i_0r0d[20], gate874_0n, initialise);
  C2RI I334 (ifint_0n[21], i_0r0d[21], gate874_0n, initialise);
  C2RI I335 (ifint_0n[22], i_0r0d[22], gate874_0n, initialise);
  C2RI I336 (ifint_0n[23], i_0r0d[23], gate874_0n, initialise);
  C2RI I337 (ifint_0n[24], i_0r0d[24], gate874_0n, initialise);
  C2RI I338 (ifint_0n[25], i_0r0d[25], gate874_0n, initialise);
  C2RI I339 (ifint_0n[26], i_0r0d[26], gate874_0n, initialise);
  C2RI I340 (ifint_0n[27], i_0r0d[27], gate874_0n, initialise);
  C2RI I341 (ifint_0n[28], i_0r0d[28], gate874_0n, initialise);
  C2RI I342 (ifint_0n[29], i_0r0d[29], gate874_0n, initialise);
  C2RI I343 (ifint_0n[30], i_0r0d[30], gate874_0n, initialise);
  C2RI I344 (ifint_0n[31], i_0r0d[31], gate874_0n, initialise);
  C3 I345 (internal_0n[51], complete871_0n[0], complete871_0n[1], complete871_0n[2]);
  C3 I346 (internal_0n[52], complete871_0n[3], complete871_0n[4], complete871_0n[5]);
  C3 I347 (internal_0n[53], complete871_0n[6], complete871_0n[7], complete871_0n[8]);
  C3 I348 (internal_0n[54], complete871_0n[9], complete871_0n[10], complete871_0n[11]);
  C3 I349 (internal_0n[55], complete871_0n[12], complete871_0n[13], complete871_0n[14]);
  C3 I350 (internal_0n[56], complete871_0n[15], complete871_0n[16], complete871_0n[17]);
  C3 I351 (internal_0n[57], complete871_0n[18], complete871_0n[19], complete871_0n[20]);
  C3 I352 (internal_0n[58], complete871_0n[21], complete871_0n[22], complete871_0n[23]);
  C3 I353 (internal_0n[59], complete871_0n[24], complete871_0n[25], complete871_0n[26]);
  C3 I354 (internal_0n[60], complete871_0n[27], complete871_0n[28], complete871_0n[29]);
  C2 I355 (internal_0n[61], complete871_0n[30], complete871_0n[31]);
  C3 I356 (internal_0n[62], internal_0n[51], internal_0n[52], internal_0n[53]);
  C3 I357 (internal_0n[63], internal_0n[54], internal_0n[55], internal_0n[56]);
  C3 I358 (internal_0n[64], internal_0n[57], internal_0n[58], internal_0n[59]);
  C2 I359 (internal_0n[65], internal_0n[60], internal_0n[61]);
  C2 I360 (internal_0n[66], internal_0n[62], internal_0n[63]);
  C2 I361 (internal_0n[67], internal_0n[64], internal_0n[65]);
  C2 I362 (oaint_0n, internal_0n[66], internal_0n[67]);
  OR2 I363 (complete871_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I364 (complete871_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I365 (complete871_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I366 (complete871_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I367 (complete871_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I368 (complete871_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I369 (complete871_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I370 (complete871_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I371 (complete871_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I372 (complete871_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I373 (complete871_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I374 (complete871_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I375 (complete871_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I376 (complete871_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I377 (complete871_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I378 (complete871_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I379 (complete871_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I380 (complete871_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I381 (complete871_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I382 (complete871_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I383 (complete871_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I384 (complete871_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I385 (complete871_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I386 (complete871_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I387 (complete871_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I388 (complete871_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I389 (complete871_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I390 (complete871_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I391 (complete871_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I392 (complete871_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I393 (complete871_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I394 (complete871_0n[31], o_0r0d[31], o_0r1d[31]);
  INV I395 (gate870_0n, o_0a);
  C2RI I396 (o_0r1d[0], otint_0n[0], gate870_0n, initialise);
  C2RI I397 (o_0r1d[1], otint_0n[1], gate870_0n, initialise);
  C2RI I398 (o_0r1d[2], otint_0n[2], gate870_0n, initialise);
  C2RI I399 (o_0r1d[3], otint_0n[3], gate870_0n, initialise);
  C2RI I400 (o_0r1d[4], otint_0n[4], gate870_0n, initialise);
  C2RI I401 (o_0r1d[5], otint_0n[5], gate870_0n, initialise);
  C2RI I402 (o_0r1d[6], otint_0n[6], gate870_0n, initialise);
  C2RI I403 (o_0r1d[7], otint_0n[7], gate870_0n, initialise);
  C2RI I404 (o_0r1d[8], otint_0n[8], gate870_0n, initialise);
  C2RI I405 (o_0r1d[9], otint_0n[9], gate870_0n, initialise);
  C2RI I406 (o_0r1d[10], otint_0n[10], gate870_0n, initialise);
  C2RI I407 (o_0r1d[11], otint_0n[11], gate870_0n, initialise);
  C2RI I408 (o_0r1d[12], otint_0n[12], gate870_0n, initialise);
  C2RI I409 (o_0r1d[13], otint_0n[13], gate870_0n, initialise);
  C2RI I410 (o_0r1d[14], otint_0n[14], gate870_0n, initialise);
  C2RI I411 (o_0r1d[15], otint_0n[15], gate870_0n, initialise);
  C2RI I412 (o_0r1d[16], otint_0n[16], gate870_0n, initialise);
  C2RI I413 (o_0r1d[17], otint_0n[17], gate870_0n, initialise);
  C2RI I414 (o_0r1d[18], otint_0n[18], gate870_0n, initialise);
  C2RI I415 (o_0r1d[19], otint_0n[19], gate870_0n, initialise);
  C2RI I416 (o_0r1d[20], otint_0n[20], gate870_0n, initialise);
  C2RI I417 (o_0r1d[21], otint_0n[21], gate870_0n, initialise);
  C2RI I418 (o_0r1d[22], otint_0n[22], gate870_0n, initialise);
  C2RI I419 (o_0r1d[23], otint_0n[23], gate870_0n, initialise);
  C2RI I420 (o_0r1d[24], otint_0n[24], gate870_0n, initialise);
  C2RI I421 (o_0r1d[25], otint_0n[25], gate870_0n, initialise);
  C2RI I422 (o_0r1d[26], otint_0n[26], gate870_0n, initialise);
  C2RI I423 (o_0r1d[27], otint_0n[27], gate870_0n, initialise);
  C2RI I424 (o_0r1d[28], otint_0n[28], gate870_0n, initialise);
  C2RI I425 (o_0r1d[29], otint_0n[29], gate870_0n, initialise);
  C2RI I426 (o_0r1d[30], otint_0n[30], gate870_0n, initialise);
  C2RI I427 (o_0r1d[31], otint_0n[31], gate870_0n, initialise);
  C2RI I428 (o_0r0d[0], ofint_0n[0], gate870_0n, initialise);
  C2RI I429 (o_0r0d[1], ofint_0n[1], gate870_0n, initialise);
  C2RI I430 (o_0r0d[2], ofint_0n[2], gate870_0n, initialise);
  C2RI I431 (o_0r0d[3], ofint_0n[3], gate870_0n, initialise);
  C2RI I432 (o_0r0d[4], ofint_0n[4], gate870_0n, initialise);
  C2RI I433 (o_0r0d[5], ofint_0n[5], gate870_0n, initialise);
  C2RI I434 (o_0r0d[6], ofint_0n[6], gate870_0n, initialise);
  C2RI I435 (o_0r0d[7], ofint_0n[7], gate870_0n, initialise);
  C2RI I436 (o_0r0d[8], ofint_0n[8], gate870_0n, initialise);
  C2RI I437 (o_0r0d[9], ofint_0n[9], gate870_0n, initialise);
  C2RI I438 (o_0r0d[10], ofint_0n[10], gate870_0n, initialise);
  C2RI I439 (o_0r0d[11], ofint_0n[11], gate870_0n, initialise);
  C2RI I440 (o_0r0d[12], ofint_0n[12], gate870_0n, initialise);
  C2RI I441 (o_0r0d[13], ofint_0n[13], gate870_0n, initialise);
  C2RI I442 (o_0r0d[14], ofint_0n[14], gate870_0n, initialise);
  C2RI I443 (o_0r0d[15], ofint_0n[15], gate870_0n, initialise);
  C2RI I444 (o_0r0d[16], ofint_0n[16], gate870_0n, initialise);
  C2RI I445 (o_0r0d[17], ofint_0n[17], gate870_0n, initialise);
  C2RI I446 (o_0r0d[18], ofint_0n[18], gate870_0n, initialise);
  C2RI I447 (o_0r0d[19], ofint_0n[19], gate870_0n, initialise);
  C2RI I448 (o_0r0d[20], ofint_0n[20], gate870_0n, initialise);
  C2RI I449 (o_0r0d[21], ofint_0n[21], gate870_0n, initialise);
  C2RI I450 (o_0r0d[22], ofint_0n[22], gate870_0n, initialise);
  C2RI I451 (o_0r0d[23], ofint_0n[23], gate870_0n, initialise);
  C2RI I452 (o_0r0d[24], ofint_0n[24], gate870_0n, initialise);
  C2RI I453 (o_0r0d[25], ofint_0n[25], gate870_0n, initialise);
  C2RI I454 (o_0r0d[26], ofint_0n[26], gate870_0n, initialise);
  C2RI I455 (o_0r0d[27], ofint_0n[27], gate870_0n, initialise);
  C2RI I456 (o_0r0d[28], ofint_0n[28], gate870_0n, initialise);
  C2RI I457 (o_0r0d[29], ofint_0n[29], gate870_0n, initialise);
  C2RI I458 (o_0r0d[30], ofint_0n[30], gate870_0n, initialise);
  C2RI I459 (o_0r0d[31], ofint_0n[31], gate870_0n, initialise);
  C2RI I460 (iaint_0n, sel_0n[0], oaint_0n, initialise);
  C2RI I461 (iaint_1n, sel_0n[1], oaint_0n, initialise);
  C2RI I462 (iaint_2n, sel_0n[2], oaint_0n, initialise);
  assign gate_0n[0] = sel_0n[0];
  assign gate_0n[1] = sel_0n[1];
  assign gate_0n[2] = sel_0n[2];
  assign sel_0n[0] = selcomp_0n;
  assign sel_0n[1] = selcomp_1n;
  assign sel_0n[2] = selcomp_2n;
  C3 I469 (internal_0n[68], complete867_0n[0], complete867_0n[1], complete867_0n[2]);
  C3 I470 (internal_0n[69], complete867_0n[3], complete867_0n[4], complete867_0n[5]);
  C3 I471 (internal_0n[70], complete867_0n[6], complete867_0n[7], complete867_0n[8]);
  C3 I472 (internal_0n[71], complete867_0n[9], complete867_0n[10], complete867_0n[11]);
  C3 I473 (internal_0n[72], complete867_0n[12], complete867_0n[13], complete867_0n[14]);
  C3 I474 (internal_0n[73], complete867_0n[15], complete867_0n[16], complete867_0n[17]);
  C3 I475 (internal_0n[74], complete867_0n[18], complete867_0n[19], complete867_0n[20]);
  C3 I476 (internal_0n[75], complete867_0n[21], complete867_0n[22], complete867_0n[23]);
  C3 I477 (internal_0n[76], complete867_0n[24], complete867_0n[25], complete867_0n[26]);
  C3 I478 (internal_0n[77], complete867_0n[27], complete867_0n[28], complete867_0n[29]);
  C2 I479 (internal_0n[78], complete867_0n[30], complete867_0n[31]);
  C3 I480 (internal_0n[79], internal_0n[68], internal_0n[69], internal_0n[70]);
  C3 I481 (internal_0n[80], internal_0n[71], internal_0n[72], internal_0n[73]);
  C3 I482 (internal_0n[81], internal_0n[74], internal_0n[75], internal_0n[76]);
  C2 I483 (internal_0n[82], internal_0n[77], internal_0n[78]);
  C2 I484 (internal_0n[83], internal_0n[79], internal_0n[80]);
  C2 I485 (internal_0n[84], internal_0n[81], internal_0n[82]);
  C2 I486 (selcomp_2n, internal_0n[83], internal_0n[84]);
  OR2 I487 (complete867_0n[0], ifint_2n[0], itint_2n[0]);
  OR2 I488 (complete867_0n[1], ifint_2n[1], itint_2n[1]);
  OR2 I489 (complete867_0n[2], ifint_2n[2], itint_2n[2]);
  OR2 I490 (complete867_0n[3], ifint_2n[3], itint_2n[3]);
  OR2 I491 (complete867_0n[4], ifint_2n[4], itint_2n[4]);
  OR2 I492 (complete867_0n[5], ifint_2n[5], itint_2n[5]);
  OR2 I493 (complete867_0n[6], ifint_2n[6], itint_2n[6]);
  OR2 I494 (complete867_0n[7], ifint_2n[7], itint_2n[7]);
  OR2 I495 (complete867_0n[8], ifint_2n[8], itint_2n[8]);
  OR2 I496 (complete867_0n[9], ifint_2n[9], itint_2n[9]);
  OR2 I497 (complete867_0n[10], ifint_2n[10], itint_2n[10]);
  OR2 I498 (complete867_0n[11], ifint_2n[11], itint_2n[11]);
  OR2 I499 (complete867_0n[12], ifint_2n[12], itint_2n[12]);
  OR2 I500 (complete867_0n[13], ifint_2n[13], itint_2n[13]);
  OR2 I501 (complete867_0n[14], ifint_2n[14], itint_2n[14]);
  OR2 I502 (complete867_0n[15], ifint_2n[15], itint_2n[15]);
  OR2 I503 (complete867_0n[16], ifint_2n[16], itint_2n[16]);
  OR2 I504 (complete867_0n[17], ifint_2n[17], itint_2n[17]);
  OR2 I505 (complete867_0n[18], ifint_2n[18], itint_2n[18]);
  OR2 I506 (complete867_0n[19], ifint_2n[19], itint_2n[19]);
  OR2 I507 (complete867_0n[20], ifint_2n[20], itint_2n[20]);
  OR2 I508 (complete867_0n[21], ifint_2n[21], itint_2n[21]);
  OR2 I509 (complete867_0n[22], ifint_2n[22], itint_2n[22]);
  OR2 I510 (complete867_0n[23], ifint_2n[23], itint_2n[23]);
  OR2 I511 (complete867_0n[24], ifint_2n[24], itint_2n[24]);
  OR2 I512 (complete867_0n[25], ifint_2n[25], itint_2n[25]);
  OR2 I513 (complete867_0n[26], ifint_2n[26], itint_2n[26]);
  OR2 I514 (complete867_0n[27], ifint_2n[27], itint_2n[27]);
  OR2 I515 (complete867_0n[28], ifint_2n[28], itint_2n[28]);
  OR2 I516 (complete867_0n[29], ifint_2n[29], itint_2n[29]);
  OR2 I517 (complete867_0n[30], ifint_2n[30], itint_2n[30]);
  OR2 I518 (complete867_0n[31], ifint_2n[31], itint_2n[31]);
  C3 I519 (internal_0n[85], complete866_0n[0], complete866_0n[1], complete866_0n[2]);
  C3 I520 (internal_0n[86], complete866_0n[3], complete866_0n[4], complete866_0n[5]);
  C3 I521 (internal_0n[87], complete866_0n[6], complete866_0n[7], complete866_0n[8]);
  C3 I522 (internal_0n[88], complete866_0n[9], complete866_0n[10], complete866_0n[11]);
  C3 I523 (internal_0n[89], complete866_0n[12], complete866_0n[13], complete866_0n[14]);
  C3 I524 (internal_0n[90], complete866_0n[15], complete866_0n[16], complete866_0n[17]);
  C3 I525 (internal_0n[91], complete866_0n[18], complete866_0n[19], complete866_0n[20]);
  C3 I526 (internal_0n[92], complete866_0n[21], complete866_0n[22], complete866_0n[23]);
  C3 I527 (internal_0n[93], complete866_0n[24], complete866_0n[25], complete866_0n[26]);
  C3 I528 (internal_0n[94], complete866_0n[27], complete866_0n[28], complete866_0n[29]);
  C2 I529 (internal_0n[95], complete866_0n[30], complete866_0n[31]);
  C3 I530 (internal_0n[96], internal_0n[85], internal_0n[86], internal_0n[87]);
  C3 I531 (internal_0n[97], internal_0n[88], internal_0n[89], internal_0n[90]);
  C3 I532 (internal_0n[98], internal_0n[91], internal_0n[92], internal_0n[93]);
  C2 I533 (internal_0n[99], internal_0n[94], internal_0n[95]);
  C2 I534 (internal_0n[100], internal_0n[96], internal_0n[97]);
  C2 I535 (internal_0n[101], internal_0n[98], internal_0n[99]);
  C2 I536 (selcomp_1n, internal_0n[100], internal_0n[101]);
  OR2 I537 (complete866_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I538 (complete866_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I539 (complete866_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I540 (complete866_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I541 (complete866_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I542 (complete866_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I543 (complete866_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I544 (complete866_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I545 (complete866_0n[8], ifint_1n[8], itint_1n[8]);
  OR2 I546 (complete866_0n[9], ifint_1n[9], itint_1n[9]);
  OR2 I547 (complete866_0n[10], ifint_1n[10], itint_1n[10]);
  OR2 I548 (complete866_0n[11], ifint_1n[11], itint_1n[11]);
  OR2 I549 (complete866_0n[12], ifint_1n[12], itint_1n[12]);
  OR2 I550 (complete866_0n[13], ifint_1n[13], itint_1n[13]);
  OR2 I551 (complete866_0n[14], ifint_1n[14], itint_1n[14]);
  OR2 I552 (complete866_0n[15], ifint_1n[15], itint_1n[15]);
  OR2 I553 (complete866_0n[16], ifint_1n[16], itint_1n[16]);
  OR2 I554 (complete866_0n[17], ifint_1n[17], itint_1n[17]);
  OR2 I555 (complete866_0n[18], ifint_1n[18], itint_1n[18]);
  OR2 I556 (complete866_0n[19], ifint_1n[19], itint_1n[19]);
  OR2 I557 (complete866_0n[20], ifint_1n[20], itint_1n[20]);
  OR2 I558 (complete866_0n[21], ifint_1n[21], itint_1n[21]);
  OR2 I559 (complete866_0n[22], ifint_1n[22], itint_1n[22]);
  OR2 I560 (complete866_0n[23], ifint_1n[23], itint_1n[23]);
  OR2 I561 (complete866_0n[24], ifint_1n[24], itint_1n[24]);
  OR2 I562 (complete866_0n[25], ifint_1n[25], itint_1n[25]);
  OR2 I563 (complete866_0n[26], ifint_1n[26], itint_1n[26]);
  OR2 I564 (complete866_0n[27], ifint_1n[27], itint_1n[27]);
  OR2 I565 (complete866_0n[28], ifint_1n[28], itint_1n[28]);
  OR2 I566 (complete866_0n[29], ifint_1n[29], itint_1n[29]);
  OR2 I567 (complete866_0n[30], ifint_1n[30], itint_1n[30]);
  OR2 I568 (complete866_0n[31], ifint_1n[31], itint_1n[31]);
  C3 I569 (internal_0n[102], complete865_0n[0], complete865_0n[1], complete865_0n[2]);
  C3 I570 (internal_0n[103], complete865_0n[3], complete865_0n[4], complete865_0n[5]);
  C3 I571 (internal_0n[104], complete865_0n[6], complete865_0n[7], complete865_0n[8]);
  C3 I572 (internal_0n[105], complete865_0n[9], complete865_0n[10], complete865_0n[11]);
  C3 I573 (internal_0n[106], complete865_0n[12], complete865_0n[13], complete865_0n[14]);
  C3 I574 (internal_0n[107], complete865_0n[15], complete865_0n[16], complete865_0n[17]);
  C3 I575 (internal_0n[108], complete865_0n[18], complete865_0n[19], complete865_0n[20]);
  C3 I576 (internal_0n[109], complete865_0n[21], complete865_0n[22], complete865_0n[23]);
  C3 I577 (internal_0n[110], complete865_0n[24], complete865_0n[25], complete865_0n[26]);
  C3 I578 (internal_0n[111], complete865_0n[27], complete865_0n[28], complete865_0n[29]);
  C2 I579 (internal_0n[112], complete865_0n[30], complete865_0n[31]);
  C3 I580 (internal_0n[113], internal_0n[102], internal_0n[103], internal_0n[104]);
  C3 I581 (internal_0n[114], internal_0n[105], internal_0n[106], internal_0n[107]);
  C3 I582 (internal_0n[115], internal_0n[108], internal_0n[109], internal_0n[110]);
  C2 I583 (internal_0n[116], internal_0n[111], internal_0n[112]);
  C2 I584 (internal_0n[117], internal_0n[113], internal_0n[114]);
  C2 I585 (internal_0n[118], internal_0n[115], internal_0n[116]);
  C2 I586 (selcomp_0n, internal_0n[117], internal_0n[118]);
  OR2 I587 (complete865_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I588 (complete865_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I589 (complete865_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I590 (complete865_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I591 (complete865_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I592 (complete865_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I593 (complete865_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I594 (complete865_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I595 (complete865_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I596 (complete865_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I597 (complete865_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I598 (complete865_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I599 (complete865_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I600 (complete865_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I601 (complete865_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I602 (complete865_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I603 (complete865_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I604 (complete865_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I605 (complete865_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I606 (complete865_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I607 (complete865_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I608 (complete865_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I609 (complete865_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I610 (complete865_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I611 (complete865_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I612 (complete865_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I613 (complete865_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I614 (complete865_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I615 (complete865_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I616 (complete865_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I617 (complete865_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I618 (complete865_0n[31], ifint_0n[31], itint_0n[31]);
  AND2 I619 (gfint_0n[0], gate_0n[0], ifint_0n[0]);
  AND2 I620 (gfint_0n[1], gate_0n[0], ifint_0n[1]);
  AND2 I621 (gfint_0n[2], gate_0n[0], ifint_0n[2]);
  AND2 I622 (gfint_0n[3], gate_0n[0], ifint_0n[3]);
  AND2 I623 (gfint_0n[4], gate_0n[0], ifint_0n[4]);
  AND2 I624 (gfint_0n[5], gate_0n[0], ifint_0n[5]);
  AND2 I625 (gfint_0n[6], gate_0n[0], ifint_0n[6]);
  AND2 I626 (gfint_0n[7], gate_0n[0], ifint_0n[7]);
  AND2 I627 (gfint_0n[8], gate_0n[0], ifint_0n[8]);
  AND2 I628 (gfint_0n[9], gate_0n[0], ifint_0n[9]);
  AND2 I629 (gfint_0n[10], gate_0n[0], ifint_0n[10]);
  AND2 I630 (gfint_0n[11], gate_0n[0], ifint_0n[11]);
  AND2 I631 (gfint_0n[12], gate_0n[0], ifint_0n[12]);
  AND2 I632 (gfint_0n[13], gate_0n[0], ifint_0n[13]);
  AND2 I633 (gfint_0n[14], gate_0n[0], ifint_0n[14]);
  AND2 I634 (gfint_0n[15], gate_0n[0], ifint_0n[15]);
  AND2 I635 (gfint_0n[16], gate_0n[0], ifint_0n[16]);
  AND2 I636 (gfint_0n[17], gate_0n[0], ifint_0n[17]);
  AND2 I637 (gfint_0n[18], gate_0n[0], ifint_0n[18]);
  AND2 I638 (gfint_0n[19], gate_0n[0], ifint_0n[19]);
  AND2 I639 (gfint_0n[20], gate_0n[0], ifint_0n[20]);
  AND2 I640 (gfint_0n[21], gate_0n[0], ifint_0n[21]);
  AND2 I641 (gfint_0n[22], gate_0n[0], ifint_0n[22]);
  AND2 I642 (gfint_0n[23], gate_0n[0], ifint_0n[23]);
  AND2 I643 (gfint_0n[24], gate_0n[0], ifint_0n[24]);
  AND2 I644 (gfint_0n[25], gate_0n[0], ifint_0n[25]);
  AND2 I645 (gfint_0n[26], gate_0n[0], ifint_0n[26]);
  AND2 I646 (gfint_0n[27], gate_0n[0], ifint_0n[27]);
  AND2 I647 (gfint_0n[28], gate_0n[0], ifint_0n[28]);
  AND2 I648 (gfint_0n[29], gate_0n[0], ifint_0n[29]);
  AND2 I649 (gfint_0n[30], gate_0n[0], ifint_0n[30]);
  AND2 I650 (gfint_0n[31], gate_0n[0], ifint_0n[31]);
  AND2 I651 (gfint_1n[0], gate_0n[1], ifint_1n[0]);
  AND2 I652 (gfint_1n[1], gate_0n[1], ifint_1n[1]);
  AND2 I653 (gfint_1n[2], gate_0n[1], ifint_1n[2]);
  AND2 I654 (gfint_1n[3], gate_0n[1], ifint_1n[3]);
  AND2 I655 (gfint_1n[4], gate_0n[1], ifint_1n[4]);
  AND2 I656 (gfint_1n[5], gate_0n[1], ifint_1n[5]);
  AND2 I657 (gfint_1n[6], gate_0n[1], ifint_1n[6]);
  AND2 I658 (gfint_1n[7], gate_0n[1], ifint_1n[7]);
  AND2 I659 (gfint_1n[8], gate_0n[1], ifint_1n[8]);
  AND2 I660 (gfint_1n[9], gate_0n[1], ifint_1n[9]);
  AND2 I661 (gfint_1n[10], gate_0n[1], ifint_1n[10]);
  AND2 I662 (gfint_1n[11], gate_0n[1], ifint_1n[11]);
  AND2 I663 (gfint_1n[12], gate_0n[1], ifint_1n[12]);
  AND2 I664 (gfint_1n[13], gate_0n[1], ifint_1n[13]);
  AND2 I665 (gfint_1n[14], gate_0n[1], ifint_1n[14]);
  AND2 I666 (gfint_1n[15], gate_0n[1], ifint_1n[15]);
  AND2 I667 (gfint_1n[16], gate_0n[1], ifint_1n[16]);
  AND2 I668 (gfint_1n[17], gate_0n[1], ifint_1n[17]);
  AND2 I669 (gfint_1n[18], gate_0n[1], ifint_1n[18]);
  AND2 I670 (gfint_1n[19], gate_0n[1], ifint_1n[19]);
  AND2 I671 (gfint_1n[20], gate_0n[1], ifint_1n[20]);
  AND2 I672 (gfint_1n[21], gate_0n[1], ifint_1n[21]);
  AND2 I673 (gfint_1n[22], gate_0n[1], ifint_1n[22]);
  AND2 I674 (gfint_1n[23], gate_0n[1], ifint_1n[23]);
  AND2 I675 (gfint_1n[24], gate_0n[1], ifint_1n[24]);
  AND2 I676 (gfint_1n[25], gate_0n[1], ifint_1n[25]);
  AND2 I677 (gfint_1n[26], gate_0n[1], ifint_1n[26]);
  AND2 I678 (gfint_1n[27], gate_0n[1], ifint_1n[27]);
  AND2 I679 (gfint_1n[28], gate_0n[1], ifint_1n[28]);
  AND2 I680 (gfint_1n[29], gate_0n[1], ifint_1n[29]);
  AND2 I681 (gfint_1n[30], gate_0n[1], ifint_1n[30]);
  AND2 I682 (gfint_1n[31], gate_0n[1], ifint_1n[31]);
  AND2 I683 (gfint_2n[0], gate_0n[2], ifint_2n[0]);
  AND2 I684 (gfint_2n[1], gate_0n[2], ifint_2n[1]);
  AND2 I685 (gfint_2n[2], gate_0n[2], ifint_2n[2]);
  AND2 I686 (gfint_2n[3], gate_0n[2], ifint_2n[3]);
  AND2 I687 (gfint_2n[4], gate_0n[2], ifint_2n[4]);
  AND2 I688 (gfint_2n[5], gate_0n[2], ifint_2n[5]);
  AND2 I689 (gfint_2n[6], gate_0n[2], ifint_2n[6]);
  AND2 I690 (gfint_2n[7], gate_0n[2], ifint_2n[7]);
  AND2 I691 (gfint_2n[8], gate_0n[2], ifint_2n[8]);
  AND2 I692 (gfint_2n[9], gate_0n[2], ifint_2n[9]);
  AND2 I693 (gfint_2n[10], gate_0n[2], ifint_2n[10]);
  AND2 I694 (gfint_2n[11], gate_0n[2], ifint_2n[11]);
  AND2 I695 (gfint_2n[12], gate_0n[2], ifint_2n[12]);
  AND2 I696 (gfint_2n[13], gate_0n[2], ifint_2n[13]);
  AND2 I697 (gfint_2n[14], gate_0n[2], ifint_2n[14]);
  AND2 I698 (gfint_2n[15], gate_0n[2], ifint_2n[15]);
  AND2 I699 (gfint_2n[16], gate_0n[2], ifint_2n[16]);
  AND2 I700 (gfint_2n[17], gate_0n[2], ifint_2n[17]);
  AND2 I701 (gfint_2n[18], gate_0n[2], ifint_2n[18]);
  AND2 I702 (gfint_2n[19], gate_0n[2], ifint_2n[19]);
  AND2 I703 (gfint_2n[20], gate_0n[2], ifint_2n[20]);
  AND2 I704 (gfint_2n[21], gate_0n[2], ifint_2n[21]);
  AND2 I705 (gfint_2n[22], gate_0n[2], ifint_2n[22]);
  AND2 I706 (gfint_2n[23], gate_0n[2], ifint_2n[23]);
  AND2 I707 (gfint_2n[24], gate_0n[2], ifint_2n[24]);
  AND2 I708 (gfint_2n[25], gate_0n[2], ifint_2n[25]);
  AND2 I709 (gfint_2n[26], gate_0n[2], ifint_2n[26]);
  AND2 I710 (gfint_2n[27], gate_0n[2], ifint_2n[27]);
  AND2 I711 (gfint_2n[28], gate_0n[2], ifint_2n[28]);
  AND2 I712 (gfint_2n[29], gate_0n[2], ifint_2n[29]);
  AND2 I713 (gfint_2n[30], gate_0n[2], ifint_2n[30]);
  AND2 I714 (gfint_2n[31], gate_0n[2], ifint_2n[31]);
  AND2 I715 (gtint_0n[0], gate_0n[0], itint_0n[0]);
  AND2 I716 (gtint_0n[1], gate_0n[0], itint_0n[1]);
  AND2 I717 (gtint_0n[2], gate_0n[0], itint_0n[2]);
  AND2 I718 (gtint_0n[3], gate_0n[0], itint_0n[3]);
  AND2 I719 (gtint_0n[4], gate_0n[0], itint_0n[4]);
  AND2 I720 (gtint_0n[5], gate_0n[0], itint_0n[5]);
  AND2 I721 (gtint_0n[6], gate_0n[0], itint_0n[6]);
  AND2 I722 (gtint_0n[7], gate_0n[0], itint_0n[7]);
  AND2 I723 (gtint_0n[8], gate_0n[0], itint_0n[8]);
  AND2 I724 (gtint_0n[9], gate_0n[0], itint_0n[9]);
  AND2 I725 (gtint_0n[10], gate_0n[0], itint_0n[10]);
  AND2 I726 (gtint_0n[11], gate_0n[0], itint_0n[11]);
  AND2 I727 (gtint_0n[12], gate_0n[0], itint_0n[12]);
  AND2 I728 (gtint_0n[13], gate_0n[0], itint_0n[13]);
  AND2 I729 (gtint_0n[14], gate_0n[0], itint_0n[14]);
  AND2 I730 (gtint_0n[15], gate_0n[0], itint_0n[15]);
  AND2 I731 (gtint_0n[16], gate_0n[0], itint_0n[16]);
  AND2 I732 (gtint_0n[17], gate_0n[0], itint_0n[17]);
  AND2 I733 (gtint_0n[18], gate_0n[0], itint_0n[18]);
  AND2 I734 (gtint_0n[19], gate_0n[0], itint_0n[19]);
  AND2 I735 (gtint_0n[20], gate_0n[0], itint_0n[20]);
  AND2 I736 (gtint_0n[21], gate_0n[0], itint_0n[21]);
  AND2 I737 (gtint_0n[22], gate_0n[0], itint_0n[22]);
  AND2 I738 (gtint_0n[23], gate_0n[0], itint_0n[23]);
  AND2 I739 (gtint_0n[24], gate_0n[0], itint_0n[24]);
  AND2 I740 (gtint_0n[25], gate_0n[0], itint_0n[25]);
  AND2 I741 (gtint_0n[26], gate_0n[0], itint_0n[26]);
  AND2 I742 (gtint_0n[27], gate_0n[0], itint_0n[27]);
  AND2 I743 (gtint_0n[28], gate_0n[0], itint_0n[28]);
  AND2 I744 (gtint_0n[29], gate_0n[0], itint_0n[29]);
  AND2 I745 (gtint_0n[30], gate_0n[0], itint_0n[30]);
  AND2 I746 (gtint_0n[31], gate_0n[0], itint_0n[31]);
  AND2 I747 (gtint_1n[0], gate_0n[1], itint_1n[0]);
  AND2 I748 (gtint_1n[1], gate_0n[1], itint_1n[1]);
  AND2 I749 (gtint_1n[2], gate_0n[1], itint_1n[2]);
  AND2 I750 (gtint_1n[3], gate_0n[1], itint_1n[3]);
  AND2 I751 (gtint_1n[4], gate_0n[1], itint_1n[4]);
  AND2 I752 (gtint_1n[5], gate_0n[1], itint_1n[5]);
  AND2 I753 (gtint_1n[6], gate_0n[1], itint_1n[6]);
  AND2 I754 (gtint_1n[7], gate_0n[1], itint_1n[7]);
  AND2 I755 (gtint_1n[8], gate_0n[1], itint_1n[8]);
  AND2 I756 (gtint_1n[9], gate_0n[1], itint_1n[9]);
  AND2 I757 (gtint_1n[10], gate_0n[1], itint_1n[10]);
  AND2 I758 (gtint_1n[11], gate_0n[1], itint_1n[11]);
  AND2 I759 (gtint_1n[12], gate_0n[1], itint_1n[12]);
  AND2 I760 (gtint_1n[13], gate_0n[1], itint_1n[13]);
  AND2 I761 (gtint_1n[14], gate_0n[1], itint_1n[14]);
  AND2 I762 (gtint_1n[15], gate_0n[1], itint_1n[15]);
  AND2 I763 (gtint_1n[16], gate_0n[1], itint_1n[16]);
  AND2 I764 (gtint_1n[17], gate_0n[1], itint_1n[17]);
  AND2 I765 (gtint_1n[18], gate_0n[1], itint_1n[18]);
  AND2 I766 (gtint_1n[19], gate_0n[1], itint_1n[19]);
  AND2 I767 (gtint_1n[20], gate_0n[1], itint_1n[20]);
  AND2 I768 (gtint_1n[21], gate_0n[1], itint_1n[21]);
  AND2 I769 (gtint_1n[22], gate_0n[1], itint_1n[22]);
  AND2 I770 (gtint_1n[23], gate_0n[1], itint_1n[23]);
  AND2 I771 (gtint_1n[24], gate_0n[1], itint_1n[24]);
  AND2 I772 (gtint_1n[25], gate_0n[1], itint_1n[25]);
  AND2 I773 (gtint_1n[26], gate_0n[1], itint_1n[26]);
  AND2 I774 (gtint_1n[27], gate_0n[1], itint_1n[27]);
  AND2 I775 (gtint_1n[28], gate_0n[1], itint_1n[28]);
  AND2 I776 (gtint_1n[29], gate_0n[1], itint_1n[29]);
  AND2 I777 (gtint_1n[30], gate_0n[1], itint_1n[30]);
  AND2 I778 (gtint_1n[31], gate_0n[1], itint_1n[31]);
  AND2 I779 (gtint_2n[0], gate_0n[2], itint_2n[0]);
  AND2 I780 (gtint_2n[1], gate_0n[2], itint_2n[1]);
  AND2 I781 (gtint_2n[2], gate_0n[2], itint_2n[2]);
  AND2 I782 (gtint_2n[3], gate_0n[2], itint_2n[3]);
  AND2 I783 (gtint_2n[4], gate_0n[2], itint_2n[4]);
  AND2 I784 (gtint_2n[5], gate_0n[2], itint_2n[5]);
  AND2 I785 (gtint_2n[6], gate_0n[2], itint_2n[6]);
  AND2 I786 (gtint_2n[7], gate_0n[2], itint_2n[7]);
  AND2 I787 (gtint_2n[8], gate_0n[2], itint_2n[8]);
  AND2 I788 (gtint_2n[9], gate_0n[2], itint_2n[9]);
  AND2 I789 (gtint_2n[10], gate_0n[2], itint_2n[10]);
  AND2 I790 (gtint_2n[11], gate_0n[2], itint_2n[11]);
  AND2 I791 (gtint_2n[12], gate_0n[2], itint_2n[12]);
  AND2 I792 (gtint_2n[13], gate_0n[2], itint_2n[13]);
  AND2 I793 (gtint_2n[14], gate_0n[2], itint_2n[14]);
  AND2 I794 (gtint_2n[15], gate_0n[2], itint_2n[15]);
  AND2 I795 (gtint_2n[16], gate_0n[2], itint_2n[16]);
  AND2 I796 (gtint_2n[17], gate_0n[2], itint_2n[17]);
  AND2 I797 (gtint_2n[18], gate_0n[2], itint_2n[18]);
  AND2 I798 (gtint_2n[19], gate_0n[2], itint_2n[19]);
  AND2 I799 (gtint_2n[20], gate_0n[2], itint_2n[20]);
  AND2 I800 (gtint_2n[21], gate_0n[2], itint_2n[21]);
  AND2 I801 (gtint_2n[22], gate_0n[2], itint_2n[22]);
  AND2 I802 (gtint_2n[23], gate_0n[2], itint_2n[23]);
  AND2 I803 (gtint_2n[24], gate_0n[2], itint_2n[24]);
  AND2 I804 (gtint_2n[25], gate_0n[2], itint_2n[25]);
  AND2 I805 (gtint_2n[26], gate_0n[2], itint_2n[26]);
  AND2 I806 (gtint_2n[27], gate_0n[2], itint_2n[27]);
  AND2 I807 (gtint_2n[28], gate_0n[2], itint_2n[28]);
  AND2 I808 (gtint_2n[29], gate_0n[2], itint_2n[29]);
  AND2 I809 (gtint_2n[30], gate_0n[2], itint_2n[30]);
  AND2 I810 (gtint_2n[31], gate_0n[2], itint_2n[31]);
  OR3 I811 (otint_0n[0], gtint_0n[0], gtint_1n[0], gtint_2n[0]);
  OR3 I812 (otint_0n[1], gtint_0n[1], gtint_1n[1], gtint_2n[1]);
  OR3 I813 (otint_0n[2], gtint_0n[2], gtint_1n[2], gtint_2n[2]);
  OR3 I814 (otint_0n[3], gtint_0n[3], gtint_1n[3], gtint_2n[3]);
  OR3 I815 (otint_0n[4], gtint_0n[4], gtint_1n[4], gtint_2n[4]);
  OR3 I816 (otint_0n[5], gtint_0n[5], gtint_1n[5], gtint_2n[5]);
  OR3 I817 (otint_0n[6], gtint_0n[6], gtint_1n[6], gtint_2n[6]);
  OR3 I818 (otint_0n[7], gtint_0n[7], gtint_1n[7], gtint_2n[7]);
  OR3 I819 (otint_0n[8], gtint_0n[8], gtint_1n[8], gtint_2n[8]);
  OR3 I820 (otint_0n[9], gtint_0n[9], gtint_1n[9], gtint_2n[9]);
  OR3 I821 (otint_0n[10], gtint_0n[10], gtint_1n[10], gtint_2n[10]);
  OR3 I822 (otint_0n[11], gtint_0n[11], gtint_1n[11], gtint_2n[11]);
  OR3 I823 (otint_0n[12], gtint_0n[12], gtint_1n[12], gtint_2n[12]);
  OR3 I824 (otint_0n[13], gtint_0n[13], gtint_1n[13], gtint_2n[13]);
  OR3 I825 (otint_0n[14], gtint_0n[14], gtint_1n[14], gtint_2n[14]);
  OR3 I826 (otint_0n[15], gtint_0n[15], gtint_1n[15], gtint_2n[15]);
  OR3 I827 (otint_0n[16], gtint_0n[16], gtint_1n[16], gtint_2n[16]);
  OR3 I828 (otint_0n[17], gtint_0n[17], gtint_1n[17], gtint_2n[17]);
  OR3 I829 (otint_0n[18], gtint_0n[18], gtint_1n[18], gtint_2n[18]);
  OR3 I830 (otint_0n[19], gtint_0n[19], gtint_1n[19], gtint_2n[19]);
  OR3 I831 (otint_0n[20], gtint_0n[20], gtint_1n[20], gtint_2n[20]);
  OR3 I832 (otint_0n[21], gtint_0n[21], gtint_1n[21], gtint_2n[21]);
  OR3 I833 (otint_0n[22], gtint_0n[22], gtint_1n[22], gtint_2n[22]);
  OR3 I834 (otint_0n[23], gtint_0n[23], gtint_1n[23], gtint_2n[23]);
  OR3 I835 (otint_0n[24], gtint_0n[24], gtint_1n[24], gtint_2n[24]);
  OR3 I836 (otint_0n[25], gtint_0n[25], gtint_1n[25], gtint_2n[25]);
  OR3 I837 (otint_0n[26], gtint_0n[26], gtint_1n[26], gtint_2n[26]);
  OR3 I838 (otint_0n[27], gtint_0n[27], gtint_1n[27], gtint_2n[27]);
  OR3 I839 (otint_0n[28], gtint_0n[28], gtint_1n[28], gtint_2n[28]);
  OR3 I840 (otint_0n[29], gtint_0n[29], gtint_1n[29], gtint_2n[29]);
  OR3 I841 (otint_0n[30], gtint_0n[30], gtint_1n[30], gtint_2n[30]);
  OR3 I842 (otint_0n[31], gtint_0n[31], gtint_1n[31], gtint_2n[31]);
  OR3 I843 (ofint_0n[0], gfint_0n[0], gfint_1n[0], gfint_2n[0]);
  OR3 I844 (ofint_0n[1], gfint_0n[1], gfint_1n[1], gfint_2n[1]);
  OR3 I845 (ofint_0n[2], gfint_0n[2], gfint_1n[2], gfint_2n[2]);
  OR3 I846 (ofint_0n[3], gfint_0n[3], gfint_1n[3], gfint_2n[3]);
  OR3 I847 (ofint_0n[4], gfint_0n[4], gfint_1n[4], gfint_2n[4]);
  OR3 I848 (ofint_0n[5], gfint_0n[5], gfint_1n[5], gfint_2n[5]);
  OR3 I849 (ofint_0n[6], gfint_0n[6], gfint_1n[6], gfint_2n[6]);
  OR3 I850 (ofint_0n[7], gfint_0n[7], gfint_1n[7], gfint_2n[7]);
  OR3 I851 (ofint_0n[8], gfint_0n[8], gfint_1n[8], gfint_2n[8]);
  OR3 I852 (ofint_0n[9], gfint_0n[9], gfint_1n[9], gfint_2n[9]);
  OR3 I853 (ofint_0n[10], gfint_0n[10], gfint_1n[10], gfint_2n[10]);
  OR3 I854 (ofint_0n[11], gfint_0n[11], gfint_1n[11], gfint_2n[11]);
  OR3 I855 (ofint_0n[12], gfint_0n[12], gfint_1n[12], gfint_2n[12]);
  OR3 I856 (ofint_0n[13], gfint_0n[13], gfint_1n[13], gfint_2n[13]);
  OR3 I857 (ofint_0n[14], gfint_0n[14], gfint_1n[14], gfint_2n[14]);
  OR3 I858 (ofint_0n[15], gfint_0n[15], gfint_1n[15], gfint_2n[15]);
  OR3 I859 (ofint_0n[16], gfint_0n[16], gfint_1n[16], gfint_2n[16]);
  OR3 I860 (ofint_0n[17], gfint_0n[17], gfint_1n[17], gfint_2n[17]);
  OR3 I861 (ofint_0n[18], gfint_0n[18], gfint_1n[18], gfint_2n[18]);
  OR3 I862 (ofint_0n[19], gfint_0n[19], gfint_1n[19], gfint_2n[19]);
  OR3 I863 (ofint_0n[20], gfint_0n[20], gfint_1n[20], gfint_2n[20]);
  OR3 I864 (ofint_0n[21], gfint_0n[21], gfint_1n[21], gfint_2n[21]);
  OR3 I865 (ofint_0n[22], gfint_0n[22], gfint_1n[22], gfint_2n[22]);
  OR3 I866 (ofint_0n[23], gfint_0n[23], gfint_1n[23], gfint_2n[23]);
  OR3 I867 (ofint_0n[24], gfint_0n[24], gfint_1n[24], gfint_2n[24]);
  OR3 I868 (ofint_0n[25], gfint_0n[25], gfint_1n[25], gfint_2n[25]);
  OR3 I869 (ofint_0n[26], gfint_0n[26], gfint_1n[26], gfint_2n[26]);
  OR3 I870 (ofint_0n[27], gfint_0n[27], gfint_1n[27], gfint_2n[27]);
  OR3 I871 (ofint_0n[28], gfint_0n[28], gfint_1n[28], gfint_2n[28]);
  OR3 I872 (ofint_0n[29], gfint_0n[29], gfint_1n[29], gfint_2n[29]);
  OR3 I873 (ofint_0n[30], gfint_0n[30], gfint_1n[30], gfint_2n[30]);
  OR3 I874 (ofint_0n[31], gfint_0n[31], gfint_1n[31], gfint_2n[31]);
endmodule

module BrzM_35_2 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [34:0] i_0r0d;
  input [34:0] i_0r1d;
  output i_0a;
  input [34:0] i_1r0d;
  input [34:0] i_1r1d;
  output i_1a;
  output [34:0] o_0r0d;
  output [34:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [89:0] internal_0n;
  wire [1:0] sel_0n;
  wire [34:0] ofint_0n;
  wire [34:0] otint_0n;
  wire oaint_0n;
  wire [34:0] ifint_0n;
  wire [34:0] ifint_1n;
  wire [34:0] itint_0n;
  wire [34:0] itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [1:0] gate_0n;
  wire [34:0] gfint_0n;
  wire [34:0] gfint_1n;
  wire [34:0] gtint_0n;
  wire [34:0] gtint_1n;
  wire [34:0] complete897_0n;
  wire gate896_0n;
  wire [34:0] complete893_0n;
  wire gate892_0n;
  wire [34:0] complete889_0n;
  wire gate888_0n;
  wire [34:0] complete885_0n;
  wire [34:0] complete884_0n;
  wire selcomp_0n;
  wire selcomp_1n;
  C3 I0 (internal_0n[0], complete897_0n[0], complete897_0n[1], complete897_0n[2]);
  C3 I1 (internal_0n[1], complete897_0n[3], complete897_0n[4], complete897_0n[5]);
  C3 I2 (internal_0n[2], complete897_0n[6], complete897_0n[7], complete897_0n[8]);
  C3 I3 (internal_0n[3], complete897_0n[9], complete897_0n[10], complete897_0n[11]);
  C3 I4 (internal_0n[4], complete897_0n[12], complete897_0n[13], complete897_0n[14]);
  C3 I5 (internal_0n[5], complete897_0n[15], complete897_0n[16], complete897_0n[17]);
  C3 I6 (internal_0n[6], complete897_0n[18], complete897_0n[19], complete897_0n[20]);
  C3 I7 (internal_0n[7], complete897_0n[21], complete897_0n[22], complete897_0n[23]);
  C3 I8 (internal_0n[8], complete897_0n[24], complete897_0n[25], complete897_0n[26]);
  C3 I9 (internal_0n[9], complete897_0n[27], complete897_0n[28], complete897_0n[29]);
  C3 I10 (internal_0n[10], complete897_0n[30], complete897_0n[31], complete897_0n[32]);
  C2 I11 (internal_0n[11], complete897_0n[33], complete897_0n[34]);
  C3 I12 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I13 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I14 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I15 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I16 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I17 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I18 (i_1a, internal_0n[16], internal_0n[17]);
  OR2 I19 (complete897_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I20 (complete897_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I21 (complete897_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I22 (complete897_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I23 (complete897_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I24 (complete897_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I25 (complete897_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I26 (complete897_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I27 (complete897_0n[8], ifint_1n[8], itint_1n[8]);
  OR2 I28 (complete897_0n[9], ifint_1n[9], itint_1n[9]);
  OR2 I29 (complete897_0n[10], ifint_1n[10], itint_1n[10]);
  OR2 I30 (complete897_0n[11], ifint_1n[11], itint_1n[11]);
  OR2 I31 (complete897_0n[12], ifint_1n[12], itint_1n[12]);
  OR2 I32 (complete897_0n[13], ifint_1n[13], itint_1n[13]);
  OR2 I33 (complete897_0n[14], ifint_1n[14], itint_1n[14]);
  OR2 I34 (complete897_0n[15], ifint_1n[15], itint_1n[15]);
  OR2 I35 (complete897_0n[16], ifint_1n[16], itint_1n[16]);
  OR2 I36 (complete897_0n[17], ifint_1n[17], itint_1n[17]);
  OR2 I37 (complete897_0n[18], ifint_1n[18], itint_1n[18]);
  OR2 I38 (complete897_0n[19], ifint_1n[19], itint_1n[19]);
  OR2 I39 (complete897_0n[20], ifint_1n[20], itint_1n[20]);
  OR2 I40 (complete897_0n[21], ifint_1n[21], itint_1n[21]);
  OR2 I41 (complete897_0n[22], ifint_1n[22], itint_1n[22]);
  OR2 I42 (complete897_0n[23], ifint_1n[23], itint_1n[23]);
  OR2 I43 (complete897_0n[24], ifint_1n[24], itint_1n[24]);
  OR2 I44 (complete897_0n[25], ifint_1n[25], itint_1n[25]);
  OR2 I45 (complete897_0n[26], ifint_1n[26], itint_1n[26]);
  OR2 I46 (complete897_0n[27], ifint_1n[27], itint_1n[27]);
  OR2 I47 (complete897_0n[28], ifint_1n[28], itint_1n[28]);
  OR2 I48 (complete897_0n[29], ifint_1n[29], itint_1n[29]);
  OR2 I49 (complete897_0n[30], ifint_1n[30], itint_1n[30]);
  OR2 I50 (complete897_0n[31], ifint_1n[31], itint_1n[31]);
  OR2 I51 (complete897_0n[32], ifint_1n[32], itint_1n[32]);
  OR2 I52 (complete897_0n[33], ifint_1n[33], itint_1n[33]);
  OR2 I53 (complete897_0n[34], ifint_1n[34], itint_1n[34]);
  INV I54 (gate896_0n, iaint_1n);
  C2RI I55 (itint_1n[0], i_1r1d[0], gate896_0n, initialise);
  C2RI I56 (itint_1n[1], i_1r1d[1], gate896_0n, initialise);
  C2RI I57 (itint_1n[2], i_1r1d[2], gate896_0n, initialise);
  C2RI I58 (itint_1n[3], i_1r1d[3], gate896_0n, initialise);
  C2RI I59 (itint_1n[4], i_1r1d[4], gate896_0n, initialise);
  C2RI I60 (itint_1n[5], i_1r1d[5], gate896_0n, initialise);
  C2RI I61 (itint_1n[6], i_1r1d[6], gate896_0n, initialise);
  C2RI I62 (itint_1n[7], i_1r1d[7], gate896_0n, initialise);
  C2RI I63 (itint_1n[8], i_1r1d[8], gate896_0n, initialise);
  C2RI I64 (itint_1n[9], i_1r1d[9], gate896_0n, initialise);
  C2RI I65 (itint_1n[10], i_1r1d[10], gate896_0n, initialise);
  C2RI I66 (itint_1n[11], i_1r1d[11], gate896_0n, initialise);
  C2RI I67 (itint_1n[12], i_1r1d[12], gate896_0n, initialise);
  C2RI I68 (itint_1n[13], i_1r1d[13], gate896_0n, initialise);
  C2RI I69 (itint_1n[14], i_1r1d[14], gate896_0n, initialise);
  C2RI I70 (itint_1n[15], i_1r1d[15], gate896_0n, initialise);
  C2RI I71 (itint_1n[16], i_1r1d[16], gate896_0n, initialise);
  C2RI I72 (itint_1n[17], i_1r1d[17], gate896_0n, initialise);
  C2RI I73 (itint_1n[18], i_1r1d[18], gate896_0n, initialise);
  C2RI I74 (itint_1n[19], i_1r1d[19], gate896_0n, initialise);
  C2RI I75 (itint_1n[20], i_1r1d[20], gate896_0n, initialise);
  C2RI I76 (itint_1n[21], i_1r1d[21], gate896_0n, initialise);
  C2RI I77 (itint_1n[22], i_1r1d[22], gate896_0n, initialise);
  C2RI I78 (itint_1n[23], i_1r1d[23], gate896_0n, initialise);
  C2RI I79 (itint_1n[24], i_1r1d[24], gate896_0n, initialise);
  C2RI I80 (itint_1n[25], i_1r1d[25], gate896_0n, initialise);
  C2RI I81 (itint_1n[26], i_1r1d[26], gate896_0n, initialise);
  C2RI I82 (itint_1n[27], i_1r1d[27], gate896_0n, initialise);
  C2RI I83 (itint_1n[28], i_1r1d[28], gate896_0n, initialise);
  C2RI I84 (itint_1n[29], i_1r1d[29], gate896_0n, initialise);
  C2RI I85 (itint_1n[30], i_1r1d[30], gate896_0n, initialise);
  C2RI I86 (itint_1n[31], i_1r1d[31], gate896_0n, initialise);
  C2RI I87 (itint_1n[32], i_1r1d[32], gate896_0n, initialise);
  C2RI I88 (itint_1n[33], i_1r1d[33], gate896_0n, initialise);
  C2RI I89 (itint_1n[34], i_1r1d[34], gate896_0n, initialise);
  C2RI I90 (ifint_1n[0], i_1r0d[0], gate896_0n, initialise);
  C2RI I91 (ifint_1n[1], i_1r0d[1], gate896_0n, initialise);
  C2RI I92 (ifint_1n[2], i_1r0d[2], gate896_0n, initialise);
  C2RI I93 (ifint_1n[3], i_1r0d[3], gate896_0n, initialise);
  C2RI I94 (ifint_1n[4], i_1r0d[4], gate896_0n, initialise);
  C2RI I95 (ifint_1n[5], i_1r0d[5], gate896_0n, initialise);
  C2RI I96 (ifint_1n[6], i_1r0d[6], gate896_0n, initialise);
  C2RI I97 (ifint_1n[7], i_1r0d[7], gate896_0n, initialise);
  C2RI I98 (ifint_1n[8], i_1r0d[8], gate896_0n, initialise);
  C2RI I99 (ifint_1n[9], i_1r0d[9], gate896_0n, initialise);
  C2RI I100 (ifint_1n[10], i_1r0d[10], gate896_0n, initialise);
  C2RI I101 (ifint_1n[11], i_1r0d[11], gate896_0n, initialise);
  C2RI I102 (ifint_1n[12], i_1r0d[12], gate896_0n, initialise);
  C2RI I103 (ifint_1n[13], i_1r0d[13], gate896_0n, initialise);
  C2RI I104 (ifint_1n[14], i_1r0d[14], gate896_0n, initialise);
  C2RI I105 (ifint_1n[15], i_1r0d[15], gate896_0n, initialise);
  C2RI I106 (ifint_1n[16], i_1r0d[16], gate896_0n, initialise);
  C2RI I107 (ifint_1n[17], i_1r0d[17], gate896_0n, initialise);
  C2RI I108 (ifint_1n[18], i_1r0d[18], gate896_0n, initialise);
  C2RI I109 (ifint_1n[19], i_1r0d[19], gate896_0n, initialise);
  C2RI I110 (ifint_1n[20], i_1r0d[20], gate896_0n, initialise);
  C2RI I111 (ifint_1n[21], i_1r0d[21], gate896_0n, initialise);
  C2RI I112 (ifint_1n[22], i_1r0d[22], gate896_0n, initialise);
  C2RI I113 (ifint_1n[23], i_1r0d[23], gate896_0n, initialise);
  C2RI I114 (ifint_1n[24], i_1r0d[24], gate896_0n, initialise);
  C2RI I115 (ifint_1n[25], i_1r0d[25], gate896_0n, initialise);
  C2RI I116 (ifint_1n[26], i_1r0d[26], gate896_0n, initialise);
  C2RI I117 (ifint_1n[27], i_1r0d[27], gate896_0n, initialise);
  C2RI I118 (ifint_1n[28], i_1r0d[28], gate896_0n, initialise);
  C2RI I119 (ifint_1n[29], i_1r0d[29], gate896_0n, initialise);
  C2RI I120 (ifint_1n[30], i_1r0d[30], gate896_0n, initialise);
  C2RI I121 (ifint_1n[31], i_1r0d[31], gate896_0n, initialise);
  C2RI I122 (ifint_1n[32], i_1r0d[32], gate896_0n, initialise);
  C2RI I123 (ifint_1n[33], i_1r0d[33], gate896_0n, initialise);
  C2RI I124 (ifint_1n[34], i_1r0d[34], gate896_0n, initialise);
  C3 I125 (internal_0n[18], complete893_0n[0], complete893_0n[1], complete893_0n[2]);
  C3 I126 (internal_0n[19], complete893_0n[3], complete893_0n[4], complete893_0n[5]);
  C3 I127 (internal_0n[20], complete893_0n[6], complete893_0n[7], complete893_0n[8]);
  C3 I128 (internal_0n[21], complete893_0n[9], complete893_0n[10], complete893_0n[11]);
  C3 I129 (internal_0n[22], complete893_0n[12], complete893_0n[13], complete893_0n[14]);
  C3 I130 (internal_0n[23], complete893_0n[15], complete893_0n[16], complete893_0n[17]);
  C3 I131 (internal_0n[24], complete893_0n[18], complete893_0n[19], complete893_0n[20]);
  C3 I132 (internal_0n[25], complete893_0n[21], complete893_0n[22], complete893_0n[23]);
  C3 I133 (internal_0n[26], complete893_0n[24], complete893_0n[25], complete893_0n[26]);
  C3 I134 (internal_0n[27], complete893_0n[27], complete893_0n[28], complete893_0n[29]);
  C3 I135 (internal_0n[28], complete893_0n[30], complete893_0n[31], complete893_0n[32]);
  C2 I136 (internal_0n[29], complete893_0n[33], complete893_0n[34]);
  C3 I137 (internal_0n[30], internal_0n[18], internal_0n[19], internal_0n[20]);
  C3 I138 (internal_0n[31], internal_0n[21], internal_0n[22], internal_0n[23]);
  C3 I139 (internal_0n[32], internal_0n[24], internal_0n[25], internal_0n[26]);
  C3 I140 (internal_0n[33], internal_0n[27], internal_0n[28], internal_0n[29]);
  C2 I141 (internal_0n[34], internal_0n[30], internal_0n[31]);
  C2 I142 (internal_0n[35], internal_0n[32], internal_0n[33]);
  C2 I143 (i_0a, internal_0n[34], internal_0n[35]);
  OR2 I144 (complete893_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I145 (complete893_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I146 (complete893_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I147 (complete893_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I148 (complete893_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I149 (complete893_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I150 (complete893_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I151 (complete893_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I152 (complete893_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I153 (complete893_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I154 (complete893_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I155 (complete893_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I156 (complete893_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I157 (complete893_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I158 (complete893_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I159 (complete893_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I160 (complete893_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I161 (complete893_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I162 (complete893_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I163 (complete893_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I164 (complete893_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I165 (complete893_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I166 (complete893_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I167 (complete893_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I168 (complete893_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I169 (complete893_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I170 (complete893_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I171 (complete893_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I172 (complete893_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I173 (complete893_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I174 (complete893_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I175 (complete893_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I176 (complete893_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I177 (complete893_0n[33], ifint_0n[33], itint_0n[33]);
  OR2 I178 (complete893_0n[34], ifint_0n[34], itint_0n[34]);
  INV I179 (gate892_0n, iaint_0n);
  C2RI I180 (itint_0n[0], i_0r1d[0], gate892_0n, initialise);
  C2RI I181 (itint_0n[1], i_0r1d[1], gate892_0n, initialise);
  C2RI I182 (itint_0n[2], i_0r1d[2], gate892_0n, initialise);
  C2RI I183 (itint_0n[3], i_0r1d[3], gate892_0n, initialise);
  C2RI I184 (itint_0n[4], i_0r1d[4], gate892_0n, initialise);
  C2RI I185 (itint_0n[5], i_0r1d[5], gate892_0n, initialise);
  C2RI I186 (itint_0n[6], i_0r1d[6], gate892_0n, initialise);
  C2RI I187 (itint_0n[7], i_0r1d[7], gate892_0n, initialise);
  C2RI I188 (itint_0n[8], i_0r1d[8], gate892_0n, initialise);
  C2RI I189 (itint_0n[9], i_0r1d[9], gate892_0n, initialise);
  C2RI I190 (itint_0n[10], i_0r1d[10], gate892_0n, initialise);
  C2RI I191 (itint_0n[11], i_0r1d[11], gate892_0n, initialise);
  C2RI I192 (itint_0n[12], i_0r1d[12], gate892_0n, initialise);
  C2RI I193 (itint_0n[13], i_0r1d[13], gate892_0n, initialise);
  C2RI I194 (itint_0n[14], i_0r1d[14], gate892_0n, initialise);
  C2RI I195 (itint_0n[15], i_0r1d[15], gate892_0n, initialise);
  C2RI I196 (itint_0n[16], i_0r1d[16], gate892_0n, initialise);
  C2RI I197 (itint_0n[17], i_0r1d[17], gate892_0n, initialise);
  C2RI I198 (itint_0n[18], i_0r1d[18], gate892_0n, initialise);
  C2RI I199 (itint_0n[19], i_0r1d[19], gate892_0n, initialise);
  C2RI I200 (itint_0n[20], i_0r1d[20], gate892_0n, initialise);
  C2RI I201 (itint_0n[21], i_0r1d[21], gate892_0n, initialise);
  C2RI I202 (itint_0n[22], i_0r1d[22], gate892_0n, initialise);
  C2RI I203 (itint_0n[23], i_0r1d[23], gate892_0n, initialise);
  C2RI I204 (itint_0n[24], i_0r1d[24], gate892_0n, initialise);
  C2RI I205 (itint_0n[25], i_0r1d[25], gate892_0n, initialise);
  C2RI I206 (itint_0n[26], i_0r1d[26], gate892_0n, initialise);
  C2RI I207 (itint_0n[27], i_0r1d[27], gate892_0n, initialise);
  C2RI I208 (itint_0n[28], i_0r1d[28], gate892_0n, initialise);
  C2RI I209 (itint_0n[29], i_0r1d[29], gate892_0n, initialise);
  C2RI I210 (itint_0n[30], i_0r1d[30], gate892_0n, initialise);
  C2RI I211 (itint_0n[31], i_0r1d[31], gate892_0n, initialise);
  C2RI I212 (itint_0n[32], i_0r1d[32], gate892_0n, initialise);
  C2RI I213 (itint_0n[33], i_0r1d[33], gate892_0n, initialise);
  C2RI I214 (itint_0n[34], i_0r1d[34], gate892_0n, initialise);
  C2RI I215 (ifint_0n[0], i_0r0d[0], gate892_0n, initialise);
  C2RI I216 (ifint_0n[1], i_0r0d[1], gate892_0n, initialise);
  C2RI I217 (ifint_0n[2], i_0r0d[2], gate892_0n, initialise);
  C2RI I218 (ifint_0n[3], i_0r0d[3], gate892_0n, initialise);
  C2RI I219 (ifint_0n[4], i_0r0d[4], gate892_0n, initialise);
  C2RI I220 (ifint_0n[5], i_0r0d[5], gate892_0n, initialise);
  C2RI I221 (ifint_0n[6], i_0r0d[6], gate892_0n, initialise);
  C2RI I222 (ifint_0n[7], i_0r0d[7], gate892_0n, initialise);
  C2RI I223 (ifint_0n[8], i_0r0d[8], gate892_0n, initialise);
  C2RI I224 (ifint_0n[9], i_0r0d[9], gate892_0n, initialise);
  C2RI I225 (ifint_0n[10], i_0r0d[10], gate892_0n, initialise);
  C2RI I226 (ifint_0n[11], i_0r0d[11], gate892_0n, initialise);
  C2RI I227 (ifint_0n[12], i_0r0d[12], gate892_0n, initialise);
  C2RI I228 (ifint_0n[13], i_0r0d[13], gate892_0n, initialise);
  C2RI I229 (ifint_0n[14], i_0r0d[14], gate892_0n, initialise);
  C2RI I230 (ifint_0n[15], i_0r0d[15], gate892_0n, initialise);
  C2RI I231 (ifint_0n[16], i_0r0d[16], gate892_0n, initialise);
  C2RI I232 (ifint_0n[17], i_0r0d[17], gate892_0n, initialise);
  C2RI I233 (ifint_0n[18], i_0r0d[18], gate892_0n, initialise);
  C2RI I234 (ifint_0n[19], i_0r0d[19], gate892_0n, initialise);
  C2RI I235 (ifint_0n[20], i_0r0d[20], gate892_0n, initialise);
  C2RI I236 (ifint_0n[21], i_0r0d[21], gate892_0n, initialise);
  C2RI I237 (ifint_0n[22], i_0r0d[22], gate892_0n, initialise);
  C2RI I238 (ifint_0n[23], i_0r0d[23], gate892_0n, initialise);
  C2RI I239 (ifint_0n[24], i_0r0d[24], gate892_0n, initialise);
  C2RI I240 (ifint_0n[25], i_0r0d[25], gate892_0n, initialise);
  C2RI I241 (ifint_0n[26], i_0r0d[26], gate892_0n, initialise);
  C2RI I242 (ifint_0n[27], i_0r0d[27], gate892_0n, initialise);
  C2RI I243 (ifint_0n[28], i_0r0d[28], gate892_0n, initialise);
  C2RI I244 (ifint_0n[29], i_0r0d[29], gate892_0n, initialise);
  C2RI I245 (ifint_0n[30], i_0r0d[30], gate892_0n, initialise);
  C2RI I246 (ifint_0n[31], i_0r0d[31], gate892_0n, initialise);
  C2RI I247 (ifint_0n[32], i_0r0d[32], gate892_0n, initialise);
  C2RI I248 (ifint_0n[33], i_0r0d[33], gate892_0n, initialise);
  C2RI I249 (ifint_0n[34], i_0r0d[34], gate892_0n, initialise);
  C3 I250 (internal_0n[36], complete889_0n[0], complete889_0n[1], complete889_0n[2]);
  C3 I251 (internal_0n[37], complete889_0n[3], complete889_0n[4], complete889_0n[5]);
  C3 I252 (internal_0n[38], complete889_0n[6], complete889_0n[7], complete889_0n[8]);
  C3 I253 (internal_0n[39], complete889_0n[9], complete889_0n[10], complete889_0n[11]);
  C3 I254 (internal_0n[40], complete889_0n[12], complete889_0n[13], complete889_0n[14]);
  C3 I255 (internal_0n[41], complete889_0n[15], complete889_0n[16], complete889_0n[17]);
  C3 I256 (internal_0n[42], complete889_0n[18], complete889_0n[19], complete889_0n[20]);
  C3 I257 (internal_0n[43], complete889_0n[21], complete889_0n[22], complete889_0n[23]);
  C3 I258 (internal_0n[44], complete889_0n[24], complete889_0n[25], complete889_0n[26]);
  C3 I259 (internal_0n[45], complete889_0n[27], complete889_0n[28], complete889_0n[29]);
  C3 I260 (internal_0n[46], complete889_0n[30], complete889_0n[31], complete889_0n[32]);
  C2 I261 (internal_0n[47], complete889_0n[33], complete889_0n[34]);
  C3 I262 (internal_0n[48], internal_0n[36], internal_0n[37], internal_0n[38]);
  C3 I263 (internal_0n[49], internal_0n[39], internal_0n[40], internal_0n[41]);
  C3 I264 (internal_0n[50], internal_0n[42], internal_0n[43], internal_0n[44]);
  C3 I265 (internal_0n[51], internal_0n[45], internal_0n[46], internal_0n[47]);
  C2 I266 (internal_0n[52], internal_0n[48], internal_0n[49]);
  C2 I267 (internal_0n[53], internal_0n[50], internal_0n[51]);
  C2 I268 (oaint_0n, internal_0n[52], internal_0n[53]);
  OR2 I269 (complete889_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I270 (complete889_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I271 (complete889_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I272 (complete889_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I273 (complete889_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I274 (complete889_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I275 (complete889_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I276 (complete889_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I277 (complete889_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I278 (complete889_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I279 (complete889_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I280 (complete889_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I281 (complete889_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I282 (complete889_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I283 (complete889_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I284 (complete889_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I285 (complete889_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I286 (complete889_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I287 (complete889_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I288 (complete889_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I289 (complete889_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I290 (complete889_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I291 (complete889_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I292 (complete889_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I293 (complete889_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I294 (complete889_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I295 (complete889_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I296 (complete889_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I297 (complete889_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I298 (complete889_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I299 (complete889_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I300 (complete889_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I301 (complete889_0n[32], o_0r0d[32], o_0r1d[32]);
  OR2 I302 (complete889_0n[33], o_0r0d[33], o_0r1d[33]);
  OR2 I303 (complete889_0n[34], o_0r0d[34], o_0r1d[34]);
  INV I304 (gate888_0n, o_0a);
  C2RI I305 (o_0r1d[0], otint_0n[0], gate888_0n, initialise);
  C2RI I306 (o_0r1d[1], otint_0n[1], gate888_0n, initialise);
  C2RI I307 (o_0r1d[2], otint_0n[2], gate888_0n, initialise);
  C2RI I308 (o_0r1d[3], otint_0n[3], gate888_0n, initialise);
  C2RI I309 (o_0r1d[4], otint_0n[4], gate888_0n, initialise);
  C2RI I310 (o_0r1d[5], otint_0n[5], gate888_0n, initialise);
  C2RI I311 (o_0r1d[6], otint_0n[6], gate888_0n, initialise);
  C2RI I312 (o_0r1d[7], otint_0n[7], gate888_0n, initialise);
  C2RI I313 (o_0r1d[8], otint_0n[8], gate888_0n, initialise);
  C2RI I314 (o_0r1d[9], otint_0n[9], gate888_0n, initialise);
  C2RI I315 (o_0r1d[10], otint_0n[10], gate888_0n, initialise);
  C2RI I316 (o_0r1d[11], otint_0n[11], gate888_0n, initialise);
  C2RI I317 (o_0r1d[12], otint_0n[12], gate888_0n, initialise);
  C2RI I318 (o_0r1d[13], otint_0n[13], gate888_0n, initialise);
  C2RI I319 (o_0r1d[14], otint_0n[14], gate888_0n, initialise);
  C2RI I320 (o_0r1d[15], otint_0n[15], gate888_0n, initialise);
  C2RI I321 (o_0r1d[16], otint_0n[16], gate888_0n, initialise);
  C2RI I322 (o_0r1d[17], otint_0n[17], gate888_0n, initialise);
  C2RI I323 (o_0r1d[18], otint_0n[18], gate888_0n, initialise);
  C2RI I324 (o_0r1d[19], otint_0n[19], gate888_0n, initialise);
  C2RI I325 (o_0r1d[20], otint_0n[20], gate888_0n, initialise);
  C2RI I326 (o_0r1d[21], otint_0n[21], gate888_0n, initialise);
  C2RI I327 (o_0r1d[22], otint_0n[22], gate888_0n, initialise);
  C2RI I328 (o_0r1d[23], otint_0n[23], gate888_0n, initialise);
  C2RI I329 (o_0r1d[24], otint_0n[24], gate888_0n, initialise);
  C2RI I330 (o_0r1d[25], otint_0n[25], gate888_0n, initialise);
  C2RI I331 (o_0r1d[26], otint_0n[26], gate888_0n, initialise);
  C2RI I332 (o_0r1d[27], otint_0n[27], gate888_0n, initialise);
  C2RI I333 (o_0r1d[28], otint_0n[28], gate888_0n, initialise);
  C2RI I334 (o_0r1d[29], otint_0n[29], gate888_0n, initialise);
  C2RI I335 (o_0r1d[30], otint_0n[30], gate888_0n, initialise);
  C2RI I336 (o_0r1d[31], otint_0n[31], gate888_0n, initialise);
  C2RI I337 (o_0r1d[32], otint_0n[32], gate888_0n, initialise);
  C2RI I338 (o_0r1d[33], otint_0n[33], gate888_0n, initialise);
  C2RI I339 (o_0r1d[34], otint_0n[34], gate888_0n, initialise);
  C2RI I340 (o_0r0d[0], ofint_0n[0], gate888_0n, initialise);
  C2RI I341 (o_0r0d[1], ofint_0n[1], gate888_0n, initialise);
  C2RI I342 (o_0r0d[2], ofint_0n[2], gate888_0n, initialise);
  C2RI I343 (o_0r0d[3], ofint_0n[3], gate888_0n, initialise);
  C2RI I344 (o_0r0d[4], ofint_0n[4], gate888_0n, initialise);
  C2RI I345 (o_0r0d[5], ofint_0n[5], gate888_0n, initialise);
  C2RI I346 (o_0r0d[6], ofint_0n[6], gate888_0n, initialise);
  C2RI I347 (o_0r0d[7], ofint_0n[7], gate888_0n, initialise);
  C2RI I348 (o_0r0d[8], ofint_0n[8], gate888_0n, initialise);
  C2RI I349 (o_0r0d[9], ofint_0n[9], gate888_0n, initialise);
  C2RI I350 (o_0r0d[10], ofint_0n[10], gate888_0n, initialise);
  C2RI I351 (o_0r0d[11], ofint_0n[11], gate888_0n, initialise);
  C2RI I352 (o_0r0d[12], ofint_0n[12], gate888_0n, initialise);
  C2RI I353 (o_0r0d[13], ofint_0n[13], gate888_0n, initialise);
  C2RI I354 (o_0r0d[14], ofint_0n[14], gate888_0n, initialise);
  C2RI I355 (o_0r0d[15], ofint_0n[15], gate888_0n, initialise);
  C2RI I356 (o_0r0d[16], ofint_0n[16], gate888_0n, initialise);
  C2RI I357 (o_0r0d[17], ofint_0n[17], gate888_0n, initialise);
  C2RI I358 (o_0r0d[18], ofint_0n[18], gate888_0n, initialise);
  C2RI I359 (o_0r0d[19], ofint_0n[19], gate888_0n, initialise);
  C2RI I360 (o_0r0d[20], ofint_0n[20], gate888_0n, initialise);
  C2RI I361 (o_0r0d[21], ofint_0n[21], gate888_0n, initialise);
  C2RI I362 (o_0r0d[22], ofint_0n[22], gate888_0n, initialise);
  C2RI I363 (o_0r0d[23], ofint_0n[23], gate888_0n, initialise);
  C2RI I364 (o_0r0d[24], ofint_0n[24], gate888_0n, initialise);
  C2RI I365 (o_0r0d[25], ofint_0n[25], gate888_0n, initialise);
  C2RI I366 (o_0r0d[26], ofint_0n[26], gate888_0n, initialise);
  C2RI I367 (o_0r0d[27], ofint_0n[27], gate888_0n, initialise);
  C2RI I368 (o_0r0d[28], ofint_0n[28], gate888_0n, initialise);
  C2RI I369 (o_0r0d[29], ofint_0n[29], gate888_0n, initialise);
  C2RI I370 (o_0r0d[30], ofint_0n[30], gate888_0n, initialise);
  C2RI I371 (o_0r0d[31], ofint_0n[31], gate888_0n, initialise);
  C2RI I372 (o_0r0d[32], ofint_0n[32], gate888_0n, initialise);
  C2RI I373 (o_0r0d[33], ofint_0n[33], gate888_0n, initialise);
  C2RI I374 (o_0r0d[34], ofint_0n[34], gate888_0n, initialise);
  C2RI I375 (iaint_0n, sel_0n[0], oaint_0n, initialise);
  C2RI I376 (iaint_1n, sel_0n[1], oaint_0n, initialise);
  assign gate_0n[0] = sel_0n[0];
  assign gate_0n[1] = sel_0n[1];
  assign sel_0n[0] = selcomp_0n;
  assign sel_0n[1] = selcomp_1n;
  C3 I381 (internal_0n[54], complete885_0n[0], complete885_0n[1], complete885_0n[2]);
  C3 I382 (internal_0n[55], complete885_0n[3], complete885_0n[4], complete885_0n[5]);
  C3 I383 (internal_0n[56], complete885_0n[6], complete885_0n[7], complete885_0n[8]);
  C3 I384 (internal_0n[57], complete885_0n[9], complete885_0n[10], complete885_0n[11]);
  C3 I385 (internal_0n[58], complete885_0n[12], complete885_0n[13], complete885_0n[14]);
  C3 I386 (internal_0n[59], complete885_0n[15], complete885_0n[16], complete885_0n[17]);
  C3 I387 (internal_0n[60], complete885_0n[18], complete885_0n[19], complete885_0n[20]);
  C3 I388 (internal_0n[61], complete885_0n[21], complete885_0n[22], complete885_0n[23]);
  C3 I389 (internal_0n[62], complete885_0n[24], complete885_0n[25], complete885_0n[26]);
  C3 I390 (internal_0n[63], complete885_0n[27], complete885_0n[28], complete885_0n[29]);
  C3 I391 (internal_0n[64], complete885_0n[30], complete885_0n[31], complete885_0n[32]);
  C2 I392 (internal_0n[65], complete885_0n[33], complete885_0n[34]);
  C3 I393 (internal_0n[66], internal_0n[54], internal_0n[55], internal_0n[56]);
  C3 I394 (internal_0n[67], internal_0n[57], internal_0n[58], internal_0n[59]);
  C3 I395 (internal_0n[68], internal_0n[60], internal_0n[61], internal_0n[62]);
  C3 I396 (internal_0n[69], internal_0n[63], internal_0n[64], internal_0n[65]);
  C2 I397 (internal_0n[70], internal_0n[66], internal_0n[67]);
  C2 I398 (internal_0n[71], internal_0n[68], internal_0n[69]);
  C2 I399 (selcomp_1n, internal_0n[70], internal_0n[71]);
  OR2 I400 (complete885_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I401 (complete885_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I402 (complete885_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I403 (complete885_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I404 (complete885_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I405 (complete885_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I406 (complete885_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I407 (complete885_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I408 (complete885_0n[8], ifint_1n[8], itint_1n[8]);
  OR2 I409 (complete885_0n[9], ifint_1n[9], itint_1n[9]);
  OR2 I410 (complete885_0n[10], ifint_1n[10], itint_1n[10]);
  OR2 I411 (complete885_0n[11], ifint_1n[11], itint_1n[11]);
  OR2 I412 (complete885_0n[12], ifint_1n[12], itint_1n[12]);
  OR2 I413 (complete885_0n[13], ifint_1n[13], itint_1n[13]);
  OR2 I414 (complete885_0n[14], ifint_1n[14], itint_1n[14]);
  OR2 I415 (complete885_0n[15], ifint_1n[15], itint_1n[15]);
  OR2 I416 (complete885_0n[16], ifint_1n[16], itint_1n[16]);
  OR2 I417 (complete885_0n[17], ifint_1n[17], itint_1n[17]);
  OR2 I418 (complete885_0n[18], ifint_1n[18], itint_1n[18]);
  OR2 I419 (complete885_0n[19], ifint_1n[19], itint_1n[19]);
  OR2 I420 (complete885_0n[20], ifint_1n[20], itint_1n[20]);
  OR2 I421 (complete885_0n[21], ifint_1n[21], itint_1n[21]);
  OR2 I422 (complete885_0n[22], ifint_1n[22], itint_1n[22]);
  OR2 I423 (complete885_0n[23], ifint_1n[23], itint_1n[23]);
  OR2 I424 (complete885_0n[24], ifint_1n[24], itint_1n[24]);
  OR2 I425 (complete885_0n[25], ifint_1n[25], itint_1n[25]);
  OR2 I426 (complete885_0n[26], ifint_1n[26], itint_1n[26]);
  OR2 I427 (complete885_0n[27], ifint_1n[27], itint_1n[27]);
  OR2 I428 (complete885_0n[28], ifint_1n[28], itint_1n[28]);
  OR2 I429 (complete885_0n[29], ifint_1n[29], itint_1n[29]);
  OR2 I430 (complete885_0n[30], ifint_1n[30], itint_1n[30]);
  OR2 I431 (complete885_0n[31], ifint_1n[31], itint_1n[31]);
  OR2 I432 (complete885_0n[32], ifint_1n[32], itint_1n[32]);
  OR2 I433 (complete885_0n[33], ifint_1n[33], itint_1n[33]);
  OR2 I434 (complete885_0n[34], ifint_1n[34], itint_1n[34]);
  C3 I435 (internal_0n[72], complete884_0n[0], complete884_0n[1], complete884_0n[2]);
  C3 I436 (internal_0n[73], complete884_0n[3], complete884_0n[4], complete884_0n[5]);
  C3 I437 (internal_0n[74], complete884_0n[6], complete884_0n[7], complete884_0n[8]);
  C3 I438 (internal_0n[75], complete884_0n[9], complete884_0n[10], complete884_0n[11]);
  C3 I439 (internal_0n[76], complete884_0n[12], complete884_0n[13], complete884_0n[14]);
  C3 I440 (internal_0n[77], complete884_0n[15], complete884_0n[16], complete884_0n[17]);
  C3 I441 (internal_0n[78], complete884_0n[18], complete884_0n[19], complete884_0n[20]);
  C3 I442 (internal_0n[79], complete884_0n[21], complete884_0n[22], complete884_0n[23]);
  C3 I443 (internal_0n[80], complete884_0n[24], complete884_0n[25], complete884_0n[26]);
  C3 I444 (internal_0n[81], complete884_0n[27], complete884_0n[28], complete884_0n[29]);
  C3 I445 (internal_0n[82], complete884_0n[30], complete884_0n[31], complete884_0n[32]);
  C2 I446 (internal_0n[83], complete884_0n[33], complete884_0n[34]);
  C3 I447 (internal_0n[84], internal_0n[72], internal_0n[73], internal_0n[74]);
  C3 I448 (internal_0n[85], internal_0n[75], internal_0n[76], internal_0n[77]);
  C3 I449 (internal_0n[86], internal_0n[78], internal_0n[79], internal_0n[80]);
  C3 I450 (internal_0n[87], internal_0n[81], internal_0n[82], internal_0n[83]);
  C2 I451 (internal_0n[88], internal_0n[84], internal_0n[85]);
  C2 I452 (internal_0n[89], internal_0n[86], internal_0n[87]);
  C2 I453 (selcomp_0n, internal_0n[88], internal_0n[89]);
  OR2 I454 (complete884_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I455 (complete884_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I456 (complete884_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I457 (complete884_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I458 (complete884_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I459 (complete884_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I460 (complete884_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I461 (complete884_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I462 (complete884_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I463 (complete884_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I464 (complete884_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I465 (complete884_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I466 (complete884_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I467 (complete884_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I468 (complete884_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I469 (complete884_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I470 (complete884_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I471 (complete884_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I472 (complete884_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I473 (complete884_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I474 (complete884_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I475 (complete884_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I476 (complete884_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I477 (complete884_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I478 (complete884_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I479 (complete884_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I480 (complete884_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I481 (complete884_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I482 (complete884_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I483 (complete884_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I484 (complete884_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I485 (complete884_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I486 (complete884_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I487 (complete884_0n[33], ifint_0n[33], itint_0n[33]);
  OR2 I488 (complete884_0n[34], ifint_0n[34], itint_0n[34]);
  AND2 I489 (gfint_0n[0], gate_0n[0], ifint_0n[0]);
  AND2 I490 (gfint_0n[1], gate_0n[0], ifint_0n[1]);
  AND2 I491 (gfint_0n[2], gate_0n[0], ifint_0n[2]);
  AND2 I492 (gfint_0n[3], gate_0n[0], ifint_0n[3]);
  AND2 I493 (gfint_0n[4], gate_0n[0], ifint_0n[4]);
  AND2 I494 (gfint_0n[5], gate_0n[0], ifint_0n[5]);
  AND2 I495 (gfint_0n[6], gate_0n[0], ifint_0n[6]);
  AND2 I496 (gfint_0n[7], gate_0n[0], ifint_0n[7]);
  AND2 I497 (gfint_0n[8], gate_0n[0], ifint_0n[8]);
  AND2 I498 (gfint_0n[9], gate_0n[0], ifint_0n[9]);
  AND2 I499 (gfint_0n[10], gate_0n[0], ifint_0n[10]);
  AND2 I500 (gfint_0n[11], gate_0n[0], ifint_0n[11]);
  AND2 I501 (gfint_0n[12], gate_0n[0], ifint_0n[12]);
  AND2 I502 (gfint_0n[13], gate_0n[0], ifint_0n[13]);
  AND2 I503 (gfint_0n[14], gate_0n[0], ifint_0n[14]);
  AND2 I504 (gfint_0n[15], gate_0n[0], ifint_0n[15]);
  AND2 I505 (gfint_0n[16], gate_0n[0], ifint_0n[16]);
  AND2 I506 (gfint_0n[17], gate_0n[0], ifint_0n[17]);
  AND2 I507 (gfint_0n[18], gate_0n[0], ifint_0n[18]);
  AND2 I508 (gfint_0n[19], gate_0n[0], ifint_0n[19]);
  AND2 I509 (gfint_0n[20], gate_0n[0], ifint_0n[20]);
  AND2 I510 (gfint_0n[21], gate_0n[0], ifint_0n[21]);
  AND2 I511 (gfint_0n[22], gate_0n[0], ifint_0n[22]);
  AND2 I512 (gfint_0n[23], gate_0n[0], ifint_0n[23]);
  AND2 I513 (gfint_0n[24], gate_0n[0], ifint_0n[24]);
  AND2 I514 (gfint_0n[25], gate_0n[0], ifint_0n[25]);
  AND2 I515 (gfint_0n[26], gate_0n[0], ifint_0n[26]);
  AND2 I516 (gfint_0n[27], gate_0n[0], ifint_0n[27]);
  AND2 I517 (gfint_0n[28], gate_0n[0], ifint_0n[28]);
  AND2 I518 (gfint_0n[29], gate_0n[0], ifint_0n[29]);
  AND2 I519 (gfint_0n[30], gate_0n[0], ifint_0n[30]);
  AND2 I520 (gfint_0n[31], gate_0n[0], ifint_0n[31]);
  AND2 I521 (gfint_0n[32], gate_0n[0], ifint_0n[32]);
  AND2 I522 (gfint_0n[33], gate_0n[0], ifint_0n[33]);
  AND2 I523 (gfint_0n[34], gate_0n[0], ifint_0n[34]);
  AND2 I524 (gfint_1n[0], gate_0n[1], ifint_1n[0]);
  AND2 I525 (gfint_1n[1], gate_0n[1], ifint_1n[1]);
  AND2 I526 (gfint_1n[2], gate_0n[1], ifint_1n[2]);
  AND2 I527 (gfint_1n[3], gate_0n[1], ifint_1n[3]);
  AND2 I528 (gfint_1n[4], gate_0n[1], ifint_1n[4]);
  AND2 I529 (gfint_1n[5], gate_0n[1], ifint_1n[5]);
  AND2 I530 (gfint_1n[6], gate_0n[1], ifint_1n[6]);
  AND2 I531 (gfint_1n[7], gate_0n[1], ifint_1n[7]);
  AND2 I532 (gfint_1n[8], gate_0n[1], ifint_1n[8]);
  AND2 I533 (gfint_1n[9], gate_0n[1], ifint_1n[9]);
  AND2 I534 (gfint_1n[10], gate_0n[1], ifint_1n[10]);
  AND2 I535 (gfint_1n[11], gate_0n[1], ifint_1n[11]);
  AND2 I536 (gfint_1n[12], gate_0n[1], ifint_1n[12]);
  AND2 I537 (gfint_1n[13], gate_0n[1], ifint_1n[13]);
  AND2 I538 (gfint_1n[14], gate_0n[1], ifint_1n[14]);
  AND2 I539 (gfint_1n[15], gate_0n[1], ifint_1n[15]);
  AND2 I540 (gfint_1n[16], gate_0n[1], ifint_1n[16]);
  AND2 I541 (gfint_1n[17], gate_0n[1], ifint_1n[17]);
  AND2 I542 (gfint_1n[18], gate_0n[1], ifint_1n[18]);
  AND2 I543 (gfint_1n[19], gate_0n[1], ifint_1n[19]);
  AND2 I544 (gfint_1n[20], gate_0n[1], ifint_1n[20]);
  AND2 I545 (gfint_1n[21], gate_0n[1], ifint_1n[21]);
  AND2 I546 (gfint_1n[22], gate_0n[1], ifint_1n[22]);
  AND2 I547 (gfint_1n[23], gate_0n[1], ifint_1n[23]);
  AND2 I548 (gfint_1n[24], gate_0n[1], ifint_1n[24]);
  AND2 I549 (gfint_1n[25], gate_0n[1], ifint_1n[25]);
  AND2 I550 (gfint_1n[26], gate_0n[1], ifint_1n[26]);
  AND2 I551 (gfint_1n[27], gate_0n[1], ifint_1n[27]);
  AND2 I552 (gfint_1n[28], gate_0n[1], ifint_1n[28]);
  AND2 I553 (gfint_1n[29], gate_0n[1], ifint_1n[29]);
  AND2 I554 (gfint_1n[30], gate_0n[1], ifint_1n[30]);
  AND2 I555 (gfint_1n[31], gate_0n[1], ifint_1n[31]);
  AND2 I556 (gfint_1n[32], gate_0n[1], ifint_1n[32]);
  AND2 I557 (gfint_1n[33], gate_0n[1], ifint_1n[33]);
  AND2 I558 (gfint_1n[34], gate_0n[1], ifint_1n[34]);
  AND2 I559 (gtint_0n[0], gate_0n[0], itint_0n[0]);
  AND2 I560 (gtint_0n[1], gate_0n[0], itint_0n[1]);
  AND2 I561 (gtint_0n[2], gate_0n[0], itint_0n[2]);
  AND2 I562 (gtint_0n[3], gate_0n[0], itint_0n[3]);
  AND2 I563 (gtint_0n[4], gate_0n[0], itint_0n[4]);
  AND2 I564 (gtint_0n[5], gate_0n[0], itint_0n[5]);
  AND2 I565 (gtint_0n[6], gate_0n[0], itint_0n[6]);
  AND2 I566 (gtint_0n[7], gate_0n[0], itint_0n[7]);
  AND2 I567 (gtint_0n[8], gate_0n[0], itint_0n[8]);
  AND2 I568 (gtint_0n[9], gate_0n[0], itint_0n[9]);
  AND2 I569 (gtint_0n[10], gate_0n[0], itint_0n[10]);
  AND2 I570 (gtint_0n[11], gate_0n[0], itint_0n[11]);
  AND2 I571 (gtint_0n[12], gate_0n[0], itint_0n[12]);
  AND2 I572 (gtint_0n[13], gate_0n[0], itint_0n[13]);
  AND2 I573 (gtint_0n[14], gate_0n[0], itint_0n[14]);
  AND2 I574 (gtint_0n[15], gate_0n[0], itint_0n[15]);
  AND2 I575 (gtint_0n[16], gate_0n[0], itint_0n[16]);
  AND2 I576 (gtint_0n[17], gate_0n[0], itint_0n[17]);
  AND2 I577 (gtint_0n[18], gate_0n[0], itint_0n[18]);
  AND2 I578 (gtint_0n[19], gate_0n[0], itint_0n[19]);
  AND2 I579 (gtint_0n[20], gate_0n[0], itint_0n[20]);
  AND2 I580 (gtint_0n[21], gate_0n[0], itint_0n[21]);
  AND2 I581 (gtint_0n[22], gate_0n[0], itint_0n[22]);
  AND2 I582 (gtint_0n[23], gate_0n[0], itint_0n[23]);
  AND2 I583 (gtint_0n[24], gate_0n[0], itint_0n[24]);
  AND2 I584 (gtint_0n[25], gate_0n[0], itint_0n[25]);
  AND2 I585 (gtint_0n[26], gate_0n[0], itint_0n[26]);
  AND2 I586 (gtint_0n[27], gate_0n[0], itint_0n[27]);
  AND2 I587 (gtint_0n[28], gate_0n[0], itint_0n[28]);
  AND2 I588 (gtint_0n[29], gate_0n[0], itint_0n[29]);
  AND2 I589 (gtint_0n[30], gate_0n[0], itint_0n[30]);
  AND2 I590 (gtint_0n[31], gate_0n[0], itint_0n[31]);
  AND2 I591 (gtint_0n[32], gate_0n[0], itint_0n[32]);
  AND2 I592 (gtint_0n[33], gate_0n[0], itint_0n[33]);
  AND2 I593 (gtint_0n[34], gate_0n[0], itint_0n[34]);
  AND2 I594 (gtint_1n[0], gate_0n[1], itint_1n[0]);
  AND2 I595 (gtint_1n[1], gate_0n[1], itint_1n[1]);
  AND2 I596 (gtint_1n[2], gate_0n[1], itint_1n[2]);
  AND2 I597 (gtint_1n[3], gate_0n[1], itint_1n[3]);
  AND2 I598 (gtint_1n[4], gate_0n[1], itint_1n[4]);
  AND2 I599 (gtint_1n[5], gate_0n[1], itint_1n[5]);
  AND2 I600 (gtint_1n[6], gate_0n[1], itint_1n[6]);
  AND2 I601 (gtint_1n[7], gate_0n[1], itint_1n[7]);
  AND2 I602 (gtint_1n[8], gate_0n[1], itint_1n[8]);
  AND2 I603 (gtint_1n[9], gate_0n[1], itint_1n[9]);
  AND2 I604 (gtint_1n[10], gate_0n[1], itint_1n[10]);
  AND2 I605 (gtint_1n[11], gate_0n[1], itint_1n[11]);
  AND2 I606 (gtint_1n[12], gate_0n[1], itint_1n[12]);
  AND2 I607 (gtint_1n[13], gate_0n[1], itint_1n[13]);
  AND2 I608 (gtint_1n[14], gate_0n[1], itint_1n[14]);
  AND2 I609 (gtint_1n[15], gate_0n[1], itint_1n[15]);
  AND2 I610 (gtint_1n[16], gate_0n[1], itint_1n[16]);
  AND2 I611 (gtint_1n[17], gate_0n[1], itint_1n[17]);
  AND2 I612 (gtint_1n[18], gate_0n[1], itint_1n[18]);
  AND2 I613 (gtint_1n[19], gate_0n[1], itint_1n[19]);
  AND2 I614 (gtint_1n[20], gate_0n[1], itint_1n[20]);
  AND2 I615 (gtint_1n[21], gate_0n[1], itint_1n[21]);
  AND2 I616 (gtint_1n[22], gate_0n[1], itint_1n[22]);
  AND2 I617 (gtint_1n[23], gate_0n[1], itint_1n[23]);
  AND2 I618 (gtint_1n[24], gate_0n[1], itint_1n[24]);
  AND2 I619 (gtint_1n[25], gate_0n[1], itint_1n[25]);
  AND2 I620 (gtint_1n[26], gate_0n[1], itint_1n[26]);
  AND2 I621 (gtint_1n[27], gate_0n[1], itint_1n[27]);
  AND2 I622 (gtint_1n[28], gate_0n[1], itint_1n[28]);
  AND2 I623 (gtint_1n[29], gate_0n[1], itint_1n[29]);
  AND2 I624 (gtint_1n[30], gate_0n[1], itint_1n[30]);
  AND2 I625 (gtint_1n[31], gate_0n[1], itint_1n[31]);
  AND2 I626 (gtint_1n[32], gate_0n[1], itint_1n[32]);
  AND2 I627 (gtint_1n[33], gate_0n[1], itint_1n[33]);
  AND2 I628 (gtint_1n[34], gate_0n[1], itint_1n[34]);
  OR2 I629 (otint_0n[0], gtint_0n[0], gtint_1n[0]);
  OR2 I630 (otint_0n[1], gtint_0n[1], gtint_1n[1]);
  OR2 I631 (otint_0n[2], gtint_0n[2], gtint_1n[2]);
  OR2 I632 (otint_0n[3], gtint_0n[3], gtint_1n[3]);
  OR2 I633 (otint_0n[4], gtint_0n[4], gtint_1n[4]);
  OR2 I634 (otint_0n[5], gtint_0n[5], gtint_1n[5]);
  OR2 I635 (otint_0n[6], gtint_0n[6], gtint_1n[6]);
  OR2 I636 (otint_0n[7], gtint_0n[7], gtint_1n[7]);
  OR2 I637 (otint_0n[8], gtint_0n[8], gtint_1n[8]);
  OR2 I638 (otint_0n[9], gtint_0n[9], gtint_1n[9]);
  OR2 I639 (otint_0n[10], gtint_0n[10], gtint_1n[10]);
  OR2 I640 (otint_0n[11], gtint_0n[11], gtint_1n[11]);
  OR2 I641 (otint_0n[12], gtint_0n[12], gtint_1n[12]);
  OR2 I642 (otint_0n[13], gtint_0n[13], gtint_1n[13]);
  OR2 I643 (otint_0n[14], gtint_0n[14], gtint_1n[14]);
  OR2 I644 (otint_0n[15], gtint_0n[15], gtint_1n[15]);
  OR2 I645 (otint_0n[16], gtint_0n[16], gtint_1n[16]);
  OR2 I646 (otint_0n[17], gtint_0n[17], gtint_1n[17]);
  OR2 I647 (otint_0n[18], gtint_0n[18], gtint_1n[18]);
  OR2 I648 (otint_0n[19], gtint_0n[19], gtint_1n[19]);
  OR2 I649 (otint_0n[20], gtint_0n[20], gtint_1n[20]);
  OR2 I650 (otint_0n[21], gtint_0n[21], gtint_1n[21]);
  OR2 I651 (otint_0n[22], gtint_0n[22], gtint_1n[22]);
  OR2 I652 (otint_0n[23], gtint_0n[23], gtint_1n[23]);
  OR2 I653 (otint_0n[24], gtint_0n[24], gtint_1n[24]);
  OR2 I654 (otint_0n[25], gtint_0n[25], gtint_1n[25]);
  OR2 I655 (otint_0n[26], gtint_0n[26], gtint_1n[26]);
  OR2 I656 (otint_0n[27], gtint_0n[27], gtint_1n[27]);
  OR2 I657 (otint_0n[28], gtint_0n[28], gtint_1n[28]);
  OR2 I658 (otint_0n[29], gtint_0n[29], gtint_1n[29]);
  OR2 I659 (otint_0n[30], gtint_0n[30], gtint_1n[30]);
  OR2 I660 (otint_0n[31], gtint_0n[31], gtint_1n[31]);
  OR2 I661 (otint_0n[32], gtint_0n[32], gtint_1n[32]);
  OR2 I662 (otint_0n[33], gtint_0n[33], gtint_1n[33]);
  OR2 I663 (otint_0n[34], gtint_0n[34], gtint_1n[34]);
  OR2 I664 (ofint_0n[0], gfint_0n[0], gfint_1n[0]);
  OR2 I665 (ofint_0n[1], gfint_0n[1], gfint_1n[1]);
  OR2 I666 (ofint_0n[2], gfint_0n[2], gfint_1n[2]);
  OR2 I667 (ofint_0n[3], gfint_0n[3], gfint_1n[3]);
  OR2 I668 (ofint_0n[4], gfint_0n[4], gfint_1n[4]);
  OR2 I669 (ofint_0n[5], gfint_0n[5], gfint_1n[5]);
  OR2 I670 (ofint_0n[6], gfint_0n[6], gfint_1n[6]);
  OR2 I671 (ofint_0n[7], gfint_0n[7], gfint_1n[7]);
  OR2 I672 (ofint_0n[8], gfint_0n[8], gfint_1n[8]);
  OR2 I673 (ofint_0n[9], gfint_0n[9], gfint_1n[9]);
  OR2 I674 (ofint_0n[10], gfint_0n[10], gfint_1n[10]);
  OR2 I675 (ofint_0n[11], gfint_0n[11], gfint_1n[11]);
  OR2 I676 (ofint_0n[12], gfint_0n[12], gfint_1n[12]);
  OR2 I677 (ofint_0n[13], gfint_0n[13], gfint_1n[13]);
  OR2 I678 (ofint_0n[14], gfint_0n[14], gfint_1n[14]);
  OR2 I679 (ofint_0n[15], gfint_0n[15], gfint_1n[15]);
  OR2 I680 (ofint_0n[16], gfint_0n[16], gfint_1n[16]);
  OR2 I681 (ofint_0n[17], gfint_0n[17], gfint_1n[17]);
  OR2 I682 (ofint_0n[18], gfint_0n[18], gfint_1n[18]);
  OR2 I683 (ofint_0n[19], gfint_0n[19], gfint_1n[19]);
  OR2 I684 (ofint_0n[20], gfint_0n[20], gfint_1n[20]);
  OR2 I685 (ofint_0n[21], gfint_0n[21], gfint_1n[21]);
  OR2 I686 (ofint_0n[22], gfint_0n[22], gfint_1n[22]);
  OR2 I687 (ofint_0n[23], gfint_0n[23], gfint_1n[23]);
  OR2 I688 (ofint_0n[24], gfint_0n[24], gfint_1n[24]);
  OR2 I689 (ofint_0n[25], gfint_0n[25], gfint_1n[25]);
  OR2 I690 (ofint_0n[26], gfint_0n[26], gfint_1n[26]);
  OR2 I691 (ofint_0n[27], gfint_0n[27], gfint_1n[27]);
  OR2 I692 (ofint_0n[28], gfint_0n[28], gfint_1n[28]);
  OR2 I693 (ofint_0n[29], gfint_0n[29], gfint_1n[29]);
  OR2 I694 (ofint_0n[30], gfint_0n[30], gfint_1n[30]);
  OR2 I695 (ofint_0n[31], gfint_0n[31], gfint_1n[31]);
  OR2 I696 (ofint_0n[32], gfint_0n[32], gfint_1n[32]);
  OR2 I697 (ofint_0n[33], gfint_0n[33], gfint_1n[33]);
  OR2 I698 (ofint_0n[34], gfint_0n[34], gfint_1n[34]);
endmodule

module BrzM_35_9 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  i_2r0d, i_2r1d, i_2a,
  i_3r0d, i_3r1d, i_3a,
  i_4r0d, i_4r1d, i_4a,
  i_5r0d, i_5r1d, i_5a,
  i_6r0d, i_6r1d, i_6a,
  i_7r0d, i_7r1d, i_7a,
  i_8r0d, i_8r1d, i_8a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [34:0] i_0r0d;
  input [34:0] i_0r1d;
  output i_0a;
  input [34:0] i_1r0d;
  input [34:0] i_1r1d;
  output i_1a;
  input [34:0] i_2r0d;
  input [34:0] i_2r1d;
  output i_2a;
  input [34:0] i_3r0d;
  input [34:0] i_3r1d;
  output i_3a;
  input [34:0] i_4r0d;
  input [34:0] i_4r1d;
  output i_4a;
  input [34:0] i_5r0d;
  input [34:0] i_5r1d;
  output i_5a;
  input [34:0] i_6r0d;
  input [34:0] i_6r1d;
  output i_6a;
  input [34:0] i_7r0d;
  input [34:0] i_7r1d;
  output i_7a;
  input [34:0] i_8r0d;
  input [34:0] i_8r1d;
  output i_8a;
  output [34:0] o_0r0d;
  output [34:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [551:0] internal_0n;
  wire [8:0] sel_0n;
  wire [34:0] ofint_0n;
  wire [34:0] otint_0n;
  wire oaint_0n;
  wire [34:0] ifint_0n;
  wire [34:0] ifint_1n;
  wire [34:0] ifint_2n;
  wire [34:0] ifint_3n;
  wire [34:0] ifint_4n;
  wire [34:0] ifint_5n;
  wire [34:0] ifint_6n;
  wire [34:0] ifint_7n;
  wire [34:0] ifint_8n;
  wire [34:0] itint_0n;
  wire [34:0] itint_1n;
  wire [34:0] itint_2n;
  wire [34:0] itint_3n;
  wire [34:0] itint_4n;
  wire [34:0] itint_5n;
  wire [34:0] itint_6n;
  wire [34:0] itint_7n;
  wire [34:0] itint_8n;
  wire iaint_0n;
  wire iaint_1n;
  wire iaint_2n;
  wire iaint_3n;
  wire iaint_4n;
  wire iaint_5n;
  wire iaint_6n;
  wire iaint_7n;
  wire iaint_8n;
  wire [8:0] gate_0n;
  wire [34:0] gfint_0n;
  wire [34:0] gfint_1n;
  wire [34:0] gfint_2n;
  wire [34:0] gfint_3n;
  wire [34:0] gfint_4n;
  wire [34:0] gfint_5n;
  wire [34:0] gfint_6n;
  wire [34:0] gfint_7n;
  wire [34:0] gfint_8n;
  wire [34:0] gtint_0n;
  wire [34:0] gtint_1n;
  wire [34:0] gtint_2n;
  wire [34:0] gtint_3n;
  wire [34:0] gtint_4n;
  wire [34:0] gtint_5n;
  wire [34:0] gtint_6n;
  wire [34:0] gtint_7n;
  wire [34:0] gtint_8n;
  wire [34:0] complete946_0n;
  wire gate945_0n;
  wire [34:0] complete942_0n;
  wire gate941_0n;
  wire [34:0] complete938_0n;
  wire gate937_0n;
  wire [34:0] complete934_0n;
  wire gate933_0n;
  wire [34:0] complete930_0n;
  wire gate929_0n;
  wire [34:0] complete926_0n;
  wire gate925_0n;
  wire [34:0] complete922_0n;
  wire gate921_0n;
  wire [34:0] complete918_0n;
  wire gate917_0n;
  wire [34:0] complete914_0n;
  wire gate913_0n;
  wire [34:0] complete910_0n;
  wire gate909_0n;
  wire [34:0] complete906_0n;
  wire [34:0] complete905_0n;
  wire [34:0] complete904_0n;
  wire [34:0] complete903_0n;
  wire [34:0] complete902_0n;
  wire [34:0] complete901_0n;
  wire [34:0] complete900_0n;
  wire [34:0] complete899_0n;
  wire [34:0] complete898_0n;
  wire selcomp_0n;
  wire selcomp_1n;
  wire selcomp_2n;
  wire selcomp_3n;
  wire selcomp_4n;
  wire selcomp_5n;
  wire selcomp_6n;
  wire selcomp_7n;
  wire selcomp_8n;
  C3 I0 (internal_0n[0], complete946_0n[0], complete946_0n[1], complete946_0n[2]);
  C3 I1 (internal_0n[1], complete946_0n[3], complete946_0n[4], complete946_0n[5]);
  C3 I2 (internal_0n[2], complete946_0n[6], complete946_0n[7], complete946_0n[8]);
  C3 I3 (internal_0n[3], complete946_0n[9], complete946_0n[10], complete946_0n[11]);
  C3 I4 (internal_0n[4], complete946_0n[12], complete946_0n[13], complete946_0n[14]);
  C3 I5 (internal_0n[5], complete946_0n[15], complete946_0n[16], complete946_0n[17]);
  C3 I6 (internal_0n[6], complete946_0n[18], complete946_0n[19], complete946_0n[20]);
  C3 I7 (internal_0n[7], complete946_0n[21], complete946_0n[22], complete946_0n[23]);
  C3 I8 (internal_0n[8], complete946_0n[24], complete946_0n[25], complete946_0n[26]);
  C3 I9 (internal_0n[9], complete946_0n[27], complete946_0n[28], complete946_0n[29]);
  C3 I10 (internal_0n[10], complete946_0n[30], complete946_0n[31], complete946_0n[32]);
  C2 I11 (internal_0n[11], complete946_0n[33], complete946_0n[34]);
  C3 I12 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I13 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I14 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I15 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I16 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I17 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I18 (i_8a, internal_0n[16], internal_0n[17]);
  OR2 I19 (complete946_0n[0], ifint_8n[0], itint_8n[0]);
  OR2 I20 (complete946_0n[1], ifint_8n[1], itint_8n[1]);
  OR2 I21 (complete946_0n[2], ifint_8n[2], itint_8n[2]);
  OR2 I22 (complete946_0n[3], ifint_8n[3], itint_8n[3]);
  OR2 I23 (complete946_0n[4], ifint_8n[4], itint_8n[4]);
  OR2 I24 (complete946_0n[5], ifint_8n[5], itint_8n[5]);
  OR2 I25 (complete946_0n[6], ifint_8n[6], itint_8n[6]);
  OR2 I26 (complete946_0n[7], ifint_8n[7], itint_8n[7]);
  OR2 I27 (complete946_0n[8], ifint_8n[8], itint_8n[8]);
  OR2 I28 (complete946_0n[9], ifint_8n[9], itint_8n[9]);
  OR2 I29 (complete946_0n[10], ifint_8n[10], itint_8n[10]);
  OR2 I30 (complete946_0n[11], ifint_8n[11], itint_8n[11]);
  OR2 I31 (complete946_0n[12], ifint_8n[12], itint_8n[12]);
  OR2 I32 (complete946_0n[13], ifint_8n[13], itint_8n[13]);
  OR2 I33 (complete946_0n[14], ifint_8n[14], itint_8n[14]);
  OR2 I34 (complete946_0n[15], ifint_8n[15], itint_8n[15]);
  OR2 I35 (complete946_0n[16], ifint_8n[16], itint_8n[16]);
  OR2 I36 (complete946_0n[17], ifint_8n[17], itint_8n[17]);
  OR2 I37 (complete946_0n[18], ifint_8n[18], itint_8n[18]);
  OR2 I38 (complete946_0n[19], ifint_8n[19], itint_8n[19]);
  OR2 I39 (complete946_0n[20], ifint_8n[20], itint_8n[20]);
  OR2 I40 (complete946_0n[21], ifint_8n[21], itint_8n[21]);
  OR2 I41 (complete946_0n[22], ifint_8n[22], itint_8n[22]);
  OR2 I42 (complete946_0n[23], ifint_8n[23], itint_8n[23]);
  OR2 I43 (complete946_0n[24], ifint_8n[24], itint_8n[24]);
  OR2 I44 (complete946_0n[25], ifint_8n[25], itint_8n[25]);
  OR2 I45 (complete946_0n[26], ifint_8n[26], itint_8n[26]);
  OR2 I46 (complete946_0n[27], ifint_8n[27], itint_8n[27]);
  OR2 I47 (complete946_0n[28], ifint_8n[28], itint_8n[28]);
  OR2 I48 (complete946_0n[29], ifint_8n[29], itint_8n[29]);
  OR2 I49 (complete946_0n[30], ifint_8n[30], itint_8n[30]);
  OR2 I50 (complete946_0n[31], ifint_8n[31], itint_8n[31]);
  OR2 I51 (complete946_0n[32], ifint_8n[32], itint_8n[32]);
  OR2 I52 (complete946_0n[33], ifint_8n[33], itint_8n[33]);
  OR2 I53 (complete946_0n[34], ifint_8n[34], itint_8n[34]);
  INV I54 (gate945_0n, iaint_8n);
  C2RI I55 (itint_8n[0], i_8r1d[0], gate945_0n, initialise);
  C2RI I56 (itint_8n[1], i_8r1d[1], gate945_0n, initialise);
  C2RI I57 (itint_8n[2], i_8r1d[2], gate945_0n, initialise);
  C2RI I58 (itint_8n[3], i_8r1d[3], gate945_0n, initialise);
  C2RI I59 (itint_8n[4], i_8r1d[4], gate945_0n, initialise);
  C2RI I60 (itint_8n[5], i_8r1d[5], gate945_0n, initialise);
  C2RI I61 (itint_8n[6], i_8r1d[6], gate945_0n, initialise);
  C2RI I62 (itint_8n[7], i_8r1d[7], gate945_0n, initialise);
  C2RI I63 (itint_8n[8], i_8r1d[8], gate945_0n, initialise);
  C2RI I64 (itint_8n[9], i_8r1d[9], gate945_0n, initialise);
  C2RI I65 (itint_8n[10], i_8r1d[10], gate945_0n, initialise);
  C2RI I66 (itint_8n[11], i_8r1d[11], gate945_0n, initialise);
  C2RI I67 (itint_8n[12], i_8r1d[12], gate945_0n, initialise);
  C2RI I68 (itint_8n[13], i_8r1d[13], gate945_0n, initialise);
  C2RI I69 (itint_8n[14], i_8r1d[14], gate945_0n, initialise);
  C2RI I70 (itint_8n[15], i_8r1d[15], gate945_0n, initialise);
  C2RI I71 (itint_8n[16], i_8r1d[16], gate945_0n, initialise);
  C2RI I72 (itint_8n[17], i_8r1d[17], gate945_0n, initialise);
  C2RI I73 (itint_8n[18], i_8r1d[18], gate945_0n, initialise);
  C2RI I74 (itint_8n[19], i_8r1d[19], gate945_0n, initialise);
  C2RI I75 (itint_8n[20], i_8r1d[20], gate945_0n, initialise);
  C2RI I76 (itint_8n[21], i_8r1d[21], gate945_0n, initialise);
  C2RI I77 (itint_8n[22], i_8r1d[22], gate945_0n, initialise);
  C2RI I78 (itint_8n[23], i_8r1d[23], gate945_0n, initialise);
  C2RI I79 (itint_8n[24], i_8r1d[24], gate945_0n, initialise);
  C2RI I80 (itint_8n[25], i_8r1d[25], gate945_0n, initialise);
  C2RI I81 (itint_8n[26], i_8r1d[26], gate945_0n, initialise);
  C2RI I82 (itint_8n[27], i_8r1d[27], gate945_0n, initialise);
  C2RI I83 (itint_8n[28], i_8r1d[28], gate945_0n, initialise);
  C2RI I84 (itint_8n[29], i_8r1d[29], gate945_0n, initialise);
  C2RI I85 (itint_8n[30], i_8r1d[30], gate945_0n, initialise);
  C2RI I86 (itint_8n[31], i_8r1d[31], gate945_0n, initialise);
  C2RI I87 (itint_8n[32], i_8r1d[32], gate945_0n, initialise);
  C2RI I88 (itint_8n[33], i_8r1d[33], gate945_0n, initialise);
  C2RI I89 (itint_8n[34], i_8r1d[34], gate945_0n, initialise);
  C2RI I90 (ifint_8n[0], i_8r0d[0], gate945_0n, initialise);
  C2RI I91 (ifint_8n[1], i_8r0d[1], gate945_0n, initialise);
  C2RI I92 (ifint_8n[2], i_8r0d[2], gate945_0n, initialise);
  C2RI I93 (ifint_8n[3], i_8r0d[3], gate945_0n, initialise);
  C2RI I94 (ifint_8n[4], i_8r0d[4], gate945_0n, initialise);
  C2RI I95 (ifint_8n[5], i_8r0d[5], gate945_0n, initialise);
  C2RI I96 (ifint_8n[6], i_8r0d[6], gate945_0n, initialise);
  C2RI I97 (ifint_8n[7], i_8r0d[7], gate945_0n, initialise);
  C2RI I98 (ifint_8n[8], i_8r0d[8], gate945_0n, initialise);
  C2RI I99 (ifint_8n[9], i_8r0d[9], gate945_0n, initialise);
  C2RI I100 (ifint_8n[10], i_8r0d[10], gate945_0n, initialise);
  C2RI I101 (ifint_8n[11], i_8r0d[11], gate945_0n, initialise);
  C2RI I102 (ifint_8n[12], i_8r0d[12], gate945_0n, initialise);
  C2RI I103 (ifint_8n[13], i_8r0d[13], gate945_0n, initialise);
  C2RI I104 (ifint_8n[14], i_8r0d[14], gate945_0n, initialise);
  C2RI I105 (ifint_8n[15], i_8r0d[15], gate945_0n, initialise);
  C2RI I106 (ifint_8n[16], i_8r0d[16], gate945_0n, initialise);
  C2RI I107 (ifint_8n[17], i_8r0d[17], gate945_0n, initialise);
  C2RI I108 (ifint_8n[18], i_8r0d[18], gate945_0n, initialise);
  C2RI I109 (ifint_8n[19], i_8r0d[19], gate945_0n, initialise);
  C2RI I110 (ifint_8n[20], i_8r0d[20], gate945_0n, initialise);
  C2RI I111 (ifint_8n[21], i_8r0d[21], gate945_0n, initialise);
  C2RI I112 (ifint_8n[22], i_8r0d[22], gate945_0n, initialise);
  C2RI I113 (ifint_8n[23], i_8r0d[23], gate945_0n, initialise);
  C2RI I114 (ifint_8n[24], i_8r0d[24], gate945_0n, initialise);
  C2RI I115 (ifint_8n[25], i_8r0d[25], gate945_0n, initialise);
  C2RI I116 (ifint_8n[26], i_8r0d[26], gate945_0n, initialise);
  C2RI I117 (ifint_8n[27], i_8r0d[27], gate945_0n, initialise);
  C2RI I118 (ifint_8n[28], i_8r0d[28], gate945_0n, initialise);
  C2RI I119 (ifint_8n[29], i_8r0d[29], gate945_0n, initialise);
  C2RI I120 (ifint_8n[30], i_8r0d[30], gate945_0n, initialise);
  C2RI I121 (ifint_8n[31], i_8r0d[31], gate945_0n, initialise);
  C2RI I122 (ifint_8n[32], i_8r0d[32], gate945_0n, initialise);
  C2RI I123 (ifint_8n[33], i_8r0d[33], gate945_0n, initialise);
  C2RI I124 (ifint_8n[34], i_8r0d[34], gate945_0n, initialise);
  C3 I125 (internal_0n[18], complete942_0n[0], complete942_0n[1], complete942_0n[2]);
  C3 I126 (internal_0n[19], complete942_0n[3], complete942_0n[4], complete942_0n[5]);
  C3 I127 (internal_0n[20], complete942_0n[6], complete942_0n[7], complete942_0n[8]);
  C3 I128 (internal_0n[21], complete942_0n[9], complete942_0n[10], complete942_0n[11]);
  C3 I129 (internal_0n[22], complete942_0n[12], complete942_0n[13], complete942_0n[14]);
  C3 I130 (internal_0n[23], complete942_0n[15], complete942_0n[16], complete942_0n[17]);
  C3 I131 (internal_0n[24], complete942_0n[18], complete942_0n[19], complete942_0n[20]);
  C3 I132 (internal_0n[25], complete942_0n[21], complete942_0n[22], complete942_0n[23]);
  C3 I133 (internal_0n[26], complete942_0n[24], complete942_0n[25], complete942_0n[26]);
  C3 I134 (internal_0n[27], complete942_0n[27], complete942_0n[28], complete942_0n[29]);
  C3 I135 (internal_0n[28], complete942_0n[30], complete942_0n[31], complete942_0n[32]);
  C2 I136 (internal_0n[29], complete942_0n[33], complete942_0n[34]);
  C3 I137 (internal_0n[30], internal_0n[18], internal_0n[19], internal_0n[20]);
  C3 I138 (internal_0n[31], internal_0n[21], internal_0n[22], internal_0n[23]);
  C3 I139 (internal_0n[32], internal_0n[24], internal_0n[25], internal_0n[26]);
  C3 I140 (internal_0n[33], internal_0n[27], internal_0n[28], internal_0n[29]);
  C2 I141 (internal_0n[34], internal_0n[30], internal_0n[31]);
  C2 I142 (internal_0n[35], internal_0n[32], internal_0n[33]);
  C2 I143 (i_7a, internal_0n[34], internal_0n[35]);
  OR2 I144 (complete942_0n[0], ifint_7n[0], itint_7n[0]);
  OR2 I145 (complete942_0n[1], ifint_7n[1], itint_7n[1]);
  OR2 I146 (complete942_0n[2], ifint_7n[2], itint_7n[2]);
  OR2 I147 (complete942_0n[3], ifint_7n[3], itint_7n[3]);
  OR2 I148 (complete942_0n[4], ifint_7n[4], itint_7n[4]);
  OR2 I149 (complete942_0n[5], ifint_7n[5], itint_7n[5]);
  OR2 I150 (complete942_0n[6], ifint_7n[6], itint_7n[6]);
  OR2 I151 (complete942_0n[7], ifint_7n[7], itint_7n[7]);
  OR2 I152 (complete942_0n[8], ifint_7n[8], itint_7n[8]);
  OR2 I153 (complete942_0n[9], ifint_7n[9], itint_7n[9]);
  OR2 I154 (complete942_0n[10], ifint_7n[10], itint_7n[10]);
  OR2 I155 (complete942_0n[11], ifint_7n[11], itint_7n[11]);
  OR2 I156 (complete942_0n[12], ifint_7n[12], itint_7n[12]);
  OR2 I157 (complete942_0n[13], ifint_7n[13], itint_7n[13]);
  OR2 I158 (complete942_0n[14], ifint_7n[14], itint_7n[14]);
  OR2 I159 (complete942_0n[15], ifint_7n[15], itint_7n[15]);
  OR2 I160 (complete942_0n[16], ifint_7n[16], itint_7n[16]);
  OR2 I161 (complete942_0n[17], ifint_7n[17], itint_7n[17]);
  OR2 I162 (complete942_0n[18], ifint_7n[18], itint_7n[18]);
  OR2 I163 (complete942_0n[19], ifint_7n[19], itint_7n[19]);
  OR2 I164 (complete942_0n[20], ifint_7n[20], itint_7n[20]);
  OR2 I165 (complete942_0n[21], ifint_7n[21], itint_7n[21]);
  OR2 I166 (complete942_0n[22], ifint_7n[22], itint_7n[22]);
  OR2 I167 (complete942_0n[23], ifint_7n[23], itint_7n[23]);
  OR2 I168 (complete942_0n[24], ifint_7n[24], itint_7n[24]);
  OR2 I169 (complete942_0n[25], ifint_7n[25], itint_7n[25]);
  OR2 I170 (complete942_0n[26], ifint_7n[26], itint_7n[26]);
  OR2 I171 (complete942_0n[27], ifint_7n[27], itint_7n[27]);
  OR2 I172 (complete942_0n[28], ifint_7n[28], itint_7n[28]);
  OR2 I173 (complete942_0n[29], ifint_7n[29], itint_7n[29]);
  OR2 I174 (complete942_0n[30], ifint_7n[30], itint_7n[30]);
  OR2 I175 (complete942_0n[31], ifint_7n[31], itint_7n[31]);
  OR2 I176 (complete942_0n[32], ifint_7n[32], itint_7n[32]);
  OR2 I177 (complete942_0n[33], ifint_7n[33], itint_7n[33]);
  OR2 I178 (complete942_0n[34], ifint_7n[34], itint_7n[34]);
  INV I179 (gate941_0n, iaint_7n);
  C2RI I180 (itint_7n[0], i_7r1d[0], gate941_0n, initialise);
  C2RI I181 (itint_7n[1], i_7r1d[1], gate941_0n, initialise);
  C2RI I182 (itint_7n[2], i_7r1d[2], gate941_0n, initialise);
  C2RI I183 (itint_7n[3], i_7r1d[3], gate941_0n, initialise);
  C2RI I184 (itint_7n[4], i_7r1d[4], gate941_0n, initialise);
  C2RI I185 (itint_7n[5], i_7r1d[5], gate941_0n, initialise);
  C2RI I186 (itint_7n[6], i_7r1d[6], gate941_0n, initialise);
  C2RI I187 (itint_7n[7], i_7r1d[7], gate941_0n, initialise);
  C2RI I188 (itint_7n[8], i_7r1d[8], gate941_0n, initialise);
  C2RI I189 (itint_7n[9], i_7r1d[9], gate941_0n, initialise);
  C2RI I190 (itint_7n[10], i_7r1d[10], gate941_0n, initialise);
  C2RI I191 (itint_7n[11], i_7r1d[11], gate941_0n, initialise);
  C2RI I192 (itint_7n[12], i_7r1d[12], gate941_0n, initialise);
  C2RI I193 (itint_7n[13], i_7r1d[13], gate941_0n, initialise);
  C2RI I194 (itint_7n[14], i_7r1d[14], gate941_0n, initialise);
  C2RI I195 (itint_7n[15], i_7r1d[15], gate941_0n, initialise);
  C2RI I196 (itint_7n[16], i_7r1d[16], gate941_0n, initialise);
  C2RI I197 (itint_7n[17], i_7r1d[17], gate941_0n, initialise);
  C2RI I198 (itint_7n[18], i_7r1d[18], gate941_0n, initialise);
  C2RI I199 (itint_7n[19], i_7r1d[19], gate941_0n, initialise);
  C2RI I200 (itint_7n[20], i_7r1d[20], gate941_0n, initialise);
  C2RI I201 (itint_7n[21], i_7r1d[21], gate941_0n, initialise);
  C2RI I202 (itint_7n[22], i_7r1d[22], gate941_0n, initialise);
  C2RI I203 (itint_7n[23], i_7r1d[23], gate941_0n, initialise);
  C2RI I204 (itint_7n[24], i_7r1d[24], gate941_0n, initialise);
  C2RI I205 (itint_7n[25], i_7r1d[25], gate941_0n, initialise);
  C2RI I206 (itint_7n[26], i_7r1d[26], gate941_0n, initialise);
  C2RI I207 (itint_7n[27], i_7r1d[27], gate941_0n, initialise);
  C2RI I208 (itint_7n[28], i_7r1d[28], gate941_0n, initialise);
  C2RI I209 (itint_7n[29], i_7r1d[29], gate941_0n, initialise);
  C2RI I210 (itint_7n[30], i_7r1d[30], gate941_0n, initialise);
  C2RI I211 (itint_7n[31], i_7r1d[31], gate941_0n, initialise);
  C2RI I212 (itint_7n[32], i_7r1d[32], gate941_0n, initialise);
  C2RI I213 (itint_7n[33], i_7r1d[33], gate941_0n, initialise);
  C2RI I214 (itint_7n[34], i_7r1d[34], gate941_0n, initialise);
  C2RI I215 (ifint_7n[0], i_7r0d[0], gate941_0n, initialise);
  C2RI I216 (ifint_7n[1], i_7r0d[1], gate941_0n, initialise);
  C2RI I217 (ifint_7n[2], i_7r0d[2], gate941_0n, initialise);
  C2RI I218 (ifint_7n[3], i_7r0d[3], gate941_0n, initialise);
  C2RI I219 (ifint_7n[4], i_7r0d[4], gate941_0n, initialise);
  C2RI I220 (ifint_7n[5], i_7r0d[5], gate941_0n, initialise);
  C2RI I221 (ifint_7n[6], i_7r0d[6], gate941_0n, initialise);
  C2RI I222 (ifint_7n[7], i_7r0d[7], gate941_0n, initialise);
  C2RI I223 (ifint_7n[8], i_7r0d[8], gate941_0n, initialise);
  C2RI I224 (ifint_7n[9], i_7r0d[9], gate941_0n, initialise);
  C2RI I225 (ifint_7n[10], i_7r0d[10], gate941_0n, initialise);
  C2RI I226 (ifint_7n[11], i_7r0d[11], gate941_0n, initialise);
  C2RI I227 (ifint_7n[12], i_7r0d[12], gate941_0n, initialise);
  C2RI I228 (ifint_7n[13], i_7r0d[13], gate941_0n, initialise);
  C2RI I229 (ifint_7n[14], i_7r0d[14], gate941_0n, initialise);
  C2RI I230 (ifint_7n[15], i_7r0d[15], gate941_0n, initialise);
  C2RI I231 (ifint_7n[16], i_7r0d[16], gate941_0n, initialise);
  C2RI I232 (ifint_7n[17], i_7r0d[17], gate941_0n, initialise);
  C2RI I233 (ifint_7n[18], i_7r0d[18], gate941_0n, initialise);
  C2RI I234 (ifint_7n[19], i_7r0d[19], gate941_0n, initialise);
  C2RI I235 (ifint_7n[20], i_7r0d[20], gate941_0n, initialise);
  C2RI I236 (ifint_7n[21], i_7r0d[21], gate941_0n, initialise);
  C2RI I237 (ifint_7n[22], i_7r0d[22], gate941_0n, initialise);
  C2RI I238 (ifint_7n[23], i_7r0d[23], gate941_0n, initialise);
  C2RI I239 (ifint_7n[24], i_7r0d[24], gate941_0n, initialise);
  C2RI I240 (ifint_7n[25], i_7r0d[25], gate941_0n, initialise);
  C2RI I241 (ifint_7n[26], i_7r0d[26], gate941_0n, initialise);
  C2RI I242 (ifint_7n[27], i_7r0d[27], gate941_0n, initialise);
  C2RI I243 (ifint_7n[28], i_7r0d[28], gate941_0n, initialise);
  C2RI I244 (ifint_7n[29], i_7r0d[29], gate941_0n, initialise);
  C2RI I245 (ifint_7n[30], i_7r0d[30], gate941_0n, initialise);
  C2RI I246 (ifint_7n[31], i_7r0d[31], gate941_0n, initialise);
  C2RI I247 (ifint_7n[32], i_7r0d[32], gate941_0n, initialise);
  C2RI I248 (ifint_7n[33], i_7r0d[33], gate941_0n, initialise);
  C2RI I249 (ifint_7n[34], i_7r0d[34], gate941_0n, initialise);
  C3 I250 (internal_0n[36], complete938_0n[0], complete938_0n[1], complete938_0n[2]);
  C3 I251 (internal_0n[37], complete938_0n[3], complete938_0n[4], complete938_0n[5]);
  C3 I252 (internal_0n[38], complete938_0n[6], complete938_0n[7], complete938_0n[8]);
  C3 I253 (internal_0n[39], complete938_0n[9], complete938_0n[10], complete938_0n[11]);
  C3 I254 (internal_0n[40], complete938_0n[12], complete938_0n[13], complete938_0n[14]);
  C3 I255 (internal_0n[41], complete938_0n[15], complete938_0n[16], complete938_0n[17]);
  C3 I256 (internal_0n[42], complete938_0n[18], complete938_0n[19], complete938_0n[20]);
  C3 I257 (internal_0n[43], complete938_0n[21], complete938_0n[22], complete938_0n[23]);
  C3 I258 (internal_0n[44], complete938_0n[24], complete938_0n[25], complete938_0n[26]);
  C3 I259 (internal_0n[45], complete938_0n[27], complete938_0n[28], complete938_0n[29]);
  C3 I260 (internal_0n[46], complete938_0n[30], complete938_0n[31], complete938_0n[32]);
  C2 I261 (internal_0n[47], complete938_0n[33], complete938_0n[34]);
  C3 I262 (internal_0n[48], internal_0n[36], internal_0n[37], internal_0n[38]);
  C3 I263 (internal_0n[49], internal_0n[39], internal_0n[40], internal_0n[41]);
  C3 I264 (internal_0n[50], internal_0n[42], internal_0n[43], internal_0n[44]);
  C3 I265 (internal_0n[51], internal_0n[45], internal_0n[46], internal_0n[47]);
  C2 I266 (internal_0n[52], internal_0n[48], internal_0n[49]);
  C2 I267 (internal_0n[53], internal_0n[50], internal_0n[51]);
  C2 I268 (i_6a, internal_0n[52], internal_0n[53]);
  OR2 I269 (complete938_0n[0], ifint_6n[0], itint_6n[0]);
  OR2 I270 (complete938_0n[1], ifint_6n[1], itint_6n[1]);
  OR2 I271 (complete938_0n[2], ifint_6n[2], itint_6n[2]);
  OR2 I272 (complete938_0n[3], ifint_6n[3], itint_6n[3]);
  OR2 I273 (complete938_0n[4], ifint_6n[4], itint_6n[4]);
  OR2 I274 (complete938_0n[5], ifint_6n[5], itint_6n[5]);
  OR2 I275 (complete938_0n[6], ifint_6n[6], itint_6n[6]);
  OR2 I276 (complete938_0n[7], ifint_6n[7], itint_6n[7]);
  OR2 I277 (complete938_0n[8], ifint_6n[8], itint_6n[8]);
  OR2 I278 (complete938_0n[9], ifint_6n[9], itint_6n[9]);
  OR2 I279 (complete938_0n[10], ifint_6n[10], itint_6n[10]);
  OR2 I280 (complete938_0n[11], ifint_6n[11], itint_6n[11]);
  OR2 I281 (complete938_0n[12], ifint_6n[12], itint_6n[12]);
  OR2 I282 (complete938_0n[13], ifint_6n[13], itint_6n[13]);
  OR2 I283 (complete938_0n[14], ifint_6n[14], itint_6n[14]);
  OR2 I284 (complete938_0n[15], ifint_6n[15], itint_6n[15]);
  OR2 I285 (complete938_0n[16], ifint_6n[16], itint_6n[16]);
  OR2 I286 (complete938_0n[17], ifint_6n[17], itint_6n[17]);
  OR2 I287 (complete938_0n[18], ifint_6n[18], itint_6n[18]);
  OR2 I288 (complete938_0n[19], ifint_6n[19], itint_6n[19]);
  OR2 I289 (complete938_0n[20], ifint_6n[20], itint_6n[20]);
  OR2 I290 (complete938_0n[21], ifint_6n[21], itint_6n[21]);
  OR2 I291 (complete938_0n[22], ifint_6n[22], itint_6n[22]);
  OR2 I292 (complete938_0n[23], ifint_6n[23], itint_6n[23]);
  OR2 I293 (complete938_0n[24], ifint_6n[24], itint_6n[24]);
  OR2 I294 (complete938_0n[25], ifint_6n[25], itint_6n[25]);
  OR2 I295 (complete938_0n[26], ifint_6n[26], itint_6n[26]);
  OR2 I296 (complete938_0n[27], ifint_6n[27], itint_6n[27]);
  OR2 I297 (complete938_0n[28], ifint_6n[28], itint_6n[28]);
  OR2 I298 (complete938_0n[29], ifint_6n[29], itint_6n[29]);
  OR2 I299 (complete938_0n[30], ifint_6n[30], itint_6n[30]);
  OR2 I300 (complete938_0n[31], ifint_6n[31], itint_6n[31]);
  OR2 I301 (complete938_0n[32], ifint_6n[32], itint_6n[32]);
  OR2 I302 (complete938_0n[33], ifint_6n[33], itint_6n[33]);
  OR2 I303 (complete938_0n[34], ifint_6n[34], itint_6n[34]);
  INV I304 (gate937_0n, iaint_6n);
  C2RI I305 (itint_6n[0], i_6r1d[0], gate937_0n, initialise);
  C2RI I306 (itint_6n[1], i_6r1d[1], gate937_0n, initialise);
  C2RI I307 (itint_6n[2], i_6r1d[2], gate937_0n, initialise);
  C2RI I308 (itint_6n[3], i_6r1d[3], gate937_0n, initialise);
  C2RI I309 (itint_6n[4], i_6r1d[4], gate937_0n, initialise);
  C2RI I310 (itint_6n[5], i_6r1d[5], gate937_0n, initialise);
  C2RI I311 (itint_6n[6], i_6r1d[6], gate937_0n, initialise);
  C2RI I312 (itint_6n[7], i_6r1d[7], gate937_0n, initialise);
  C2RI I313 (itint_6n[8], i_6r1d[8], gate937_0n, initialise);
  C2RI I314 (itint_6n[9], i_6r1d[9], gate937_0n, initialise);
  C2RI I315 (itint_6n[10], i_6r1d[10], gate937_0n, initialise);
  C2RI I316 (itint_6n[11], i_6r1d[11], gate937_0n, initialise);
  C2RI I317 (itint_6n[12], i_6r1d[12], gate937_0n, initialise);
  C2RI I318 (itint_6n[13], i_6r1d[13], gate937_0n, initialise);
  C2RI I319 (itint_6n[14], i_6r1d[14], gate937_0n, initialise);
  C2RI I320 (itint_6n[15], i_6r1d[15], gate937_0n, initialise);
  C2RI I321 (itint_6n[16], i_6r1d[16], gate937_0n, initialise);
  C2RI I322 (itint_6n[17], i_6r1d[17], gate937_0n, initialise);
  C2RI I323 (itint_6n[18], i_6r1d[18], gate937_0n, initialise);
  C2RI I324 (itint_6n[19], i_6r1d[19], gate937_0n, initialise);
  C2RI I325 (itint_6n[20], i_6r1d[20], gate937_0n, initialise);
  C2RI I326 (itint_6n[21], i_6r1d[21], gate937_0n, initialise);
  C2RI I327 (itint_6n[22], i_6r1d[22], gate937_0n, initialise);
  C2RI I328 (itint_6n[23], i_6r1d[23], gate937_0n, initialise);
  C2RI I329 (itint_6n[24], i_6r1d[24], gate937_0n, initialise);
  C2RI I330 (itint_6n[25], i_6r1d[25], gate937_0n, initialise);
  C2RI I331 (itint_6n[26], i_6r1d[26], gate937_0n, initialise);
  C2RI I332 (itint_6n[27], i_6r1d[27], gate937_0n, initialise);
  C2RI I333 (itint_6n[28], i_6r1d[28], gate937_0n, initialise);
  C2RI I334 (itint_6n[29], i_6r1d[29], gate937_0n, initialise);
  C2RI I335 (itint_6n[30], i_6r1d[30], gate937_0n, initialise);
  C2RI I336 (itint_6n[31], i_6r1d[31], gate937_0n, initialise);
  C2RI I337 (itint_6n[32], i_6r1d[32], gate937_0n, initialise);
  C2RI I338 (itint_6n[33], i_6r1d[33], gate937_0n, initialise);
  C2RI I339 (itint_6n[34], i_6r1d[34], gate937_0n, initialise);
  C2RI I340 (ifint_6n[0], i_6r0d[0], gate937_0n, initialise);
  C2RI I341 (ifint_6n[1], i_6r0d[1], gate937_0n, initialise);
  C2RI I342 (ifint_6n[2], i_6r0d[2], gate937_0n, initialise);
  C2RI I343 (ifint_6n[3], i_6r0d[3], gate937_0n, initialise);
  C2RI I344 (ifint_6n[4], i_6r0d[4], gate937_0n, initialise);
  C2RI I345 (ifint_6n[5], i_6r0d[5], gate937_0n, initialise);
  C2RI I346 (ifint_6n[6], i_6r0d[6], gate937_0n, initialise);
  C2RI I347 (ifint_6n[7], i_6r0d[7], gate937_0n, initialise);
  C2RI I348 (ifint_6n[8], i_6r0d[8], gate937_0n, initialise);
  C2RI I349 (ifint_6n[9], i_6r0d[9], gate937_0n, initialise);
  C2RI I350 (ifint_6n[10], i_6r0d[10], gate937_0n, initialise);
  C2RI I351 (ifint_6n[11], i_6r0d[11], gate937_0n, initialise);
  C2RI I352 (ifint_6n[12], i_6r0d[12], gate937_0n, initialise);
  C2RI I353 (ifint_6n[13], i_6r0d[13], gate937_0n, initialise);
  C2RI I354 (ifint_6n[14], i_6r0d[14], gate937_0n, initialise);
  C2RI I355 (ifint_6n[15], i_6r0d[15], gate937_0n, initialise);
  C2RI I356 (ifint_6n[16], i_6r0d[16], gate937_0n, initialise);
  C2RI I357 (ifint_6n[17], i_6r0d[17], gate937_0n, initialise);
  C2RI I358 (ifint_6n[18], i_6r0d[18], gate937_0n, initialise);
  C2RI I359 (ifint_6n[19], i_6r0d[19], gate937_0n, initialise);
  C2RI I360 (ifint_6n[20], i_6r0d[20], gate937_0n, initialise);
  C2RI I361 (ifint_6n[21], i_6r0d[21], gate937_0n, initialise);
  C2RI I362 (ifint_6n[22], i_6r0d[22], gate937_0n, initialise);
  C2RI I363 (ifint_6n[23], i_6r0d[23], gate937_0n, initialise);
  C2RI I364 (ifint_6n[24], i_6r0d[24], gate937_0n, initialise);
  C2RI I365 (ifint_6n[25], i_6r0d[25], gate937_0n, initialise);
  C2RI I366 (ifint_6n[26], i_6r0d[26], gate937_0n, initialise);
  C2RI I367 (ifint_6n[27], i_6r0d[27], gate937_0n, initialise);
  C2RI I368 (ifint_6n[28], i_6r0d[28], gate937_0n, initialise);
  C2RI I369 (ifint_6n[29], i_6r0d[29], gate937_0n, initialise);
  C2RI I370 (ifint_6n[30], i_6r0d[30], gate937_0n, initialise);
  C2RI I371 (ifint_6n[31], i_6r0d[31], gate937_0n, initialise);
  C2RI I372 (ifint_6n[32], i_6r0d[32], gate937_0n, initialise);
  C2RI I373 (ifint_6n[33], i_6r0d[33], gate937_0n, initialise);
  C2RI I374 (ifint_6n[34], i_6r0d[34], gate937_0n, initialise);
  C3 I375 (internal_0n[54], complete934_0n[0], complete934_0n[1], complete934_0n[2]);
  C3 I376 (internal_0n[55], complete934_0n[3], complete934_0n[4], complete934_0n[5]);
  C3 I377 (internal_0n[56], complete934_0n[6], complete934_0n[7], complete934_0n[8]);
  C3 I378 (internal_0n[57], complete934_0n[9], complete934_0n[10], complete934_0n[11]);
  C3 I379 (internal_0n[58], complete934_0n[12], complete934_0n[13], complete934_0n[14]);
  C3 I380 (internal_0n[59], complete934_0n[15], complete934_0n[16], complete934_0n[17]);
  C3 I381 (internal_0n[60], complete934_0n[18], complete934_0n[19], complete934_0n[20]);
  C3 I382 (internal_0n[61], complete934_0n[21], complete934_0n[22], complete934_0n[23]);
  C3 I383 (internal_0n[62], complete934_0n[24], complete934_0n[25], complete934_0n[26]);
  C3 I384 (internal_0n[63], complete934_0n[27], complete934_0n[28], complete934_0n[29]);
  C3 I385 (internal_0n[64], complete934_0n[30], complete934_0n[31], complete934_0n[32]);
  C2 I386 (internal_0n[65], complete934_0n[33], complete934_0n[34]);
  C3 I387 (internal_0n[66], internal_0n[54], internal_0n[55], internal_0n[56]);
  C3 I388 (internal_0n[67], internal_0n[57], internal_0n[58], internal_0n[59]);
  C3 I389 (internal_0n[68], internal_0n[60], internal_0n[61], internal_0n[62]);
  C3 I390 (internal_0n[69], internal_0n[63], internal_0n[64], internal_0n[65]);
  C2 I391 (internal_0n[70], internal_0n[66], internal_0n[67]);
  C2 I392 (internal_0n[71], internal_0n[68], internal_0n[69]);
  C2 I393 (i_5a, internal_0n[70], internal_0n[71]);
  OR2 I394 (complete934_0n[0], ifint_5n[0], itint_5n[0]);
  OR2 I395 (complete934_0n[1], ifint_5n[1], itint_5n[1]);
  OR2 I396 (complete934_0n[2], ifint_5n[2], itint_5n[2]);
  OR2 I397 (complete934_0n[3], ifint_5n[3], itint_5n[3]);
  OR2 I398 (complete934_0n[4], ifint_5n[4], itint_5n[4]);
  OR2 I399 (complete934_0n[5], ifint_5n[5], itint_5n[5]);
  OR2 I400 (complete934_0n[6], ifint_5n[6], itint_5n[6]);
  OR2 I401 (complete934_0n[7], ifint_5n[7], itint_5n[7]);
  OR2 I402 (complete934_0n[8], ifint_5n[8], itint_5n[8]);
  OR2 I403 (complete934_0n[9], ifint_5n[9], itint_5n[9]);
  OR2 I404 (complete934_0n[10], ifint_5n[10], itint_5n[10]);
  OR2 I405 (complete934_0n[11], ifint_5n[11], itint_5n[11]);
  OR2 I406 (complete934_0n[12], ifint_5n[12], itint_5n[12]);
  OR2 I407 (complete934_0n[13], ifint_5n[13], itint_5n[13]);
  OR2 I408 (complete934_0n[14], ifint_5n[14], itint_5n[14]);
  OR2 I409 (complete934_0n[15], ifint_5n[15], itint_5n[15]);
  OR2 I410 (complete934_0n[16], ifint_5n[16], itint_5n[16]);
  OR2 I411 (complete934_0n[17], ifint_5n[17], itint_5n[17]);
  OR2 I412 (complete934_0n[18], ifint_5n[18], itint_5n[18]);
  OR2 I413 (complete934_0n[19], ifint_5n[19], itint_5n[19]);
  OR2 I414 (complete934_0n[20], ifint_5n[20], itint_5n[20]);
  OR2 I415 (complete934_0n[21], ifint_5n[21], itint_5n[21]);
  OR2 I416 (complete934_0n[22], ifint_5n[22], itint_5n[22]);
  OR2 I417 (complete934_0n[23], ifint_5n[23], itint_5n[23]);
  OR2 I418 (complete934_0n[24], ifint_5n[24], itint_5n[24]);
  OR2 I419 (complete934_0n[25], ifint_5n[25], itint_5n[25]);
  OR2 I420 (complete934_0n[26], ifint_5n[26], itint_5n[26]);
  OR2 I421 (complete934_0n[27], ifint_5n[27], itint_5n[27]);
  OR2 I422 (complete934_0n[28], ifint_5n[28], itint_5n[28]);
  OR2 I423 (complete934_0n[29], ifint_5n[29], itint_5n[29]);
  OR2 I424 (complete934_0n[30], ifint_5n[30], itint_5n[30]);
  OR2 I425 (complete934_0n[31], ifint_5n[31], itint_5n[31]);
  OR2 I426 (complete934_0n[32], ifint_5n[32], itint_5n[32]);
  OR2 I427 (complete934_0n[33], ifint_5n[33], itint_5n[33]);
  OR2 I428 (complete934_0n[34], ifint_5n[34], itint_5n[34]);
  INV I429 (gate933_0n, iaint_5n);
  C2RI I430 (itint_5n[0], i_5r1d[0], gate933_0n, initialise);
  C2RI I431 (itint_5n[1], i_5r1d[1], gate933_0n, initialise);
  C2RI I432 (itint_5n[2], i_5r1d[2], gate933_0n, initialise);
  C2RI I433 (itint_5n[3], i_5r1d[3], gate933_0n, initialise);
  C2RI I434 (itint_5n[4], i_5r1d[4], gate933_0n, initialise);
  C2RI I435 (itint_5n[5], i_5r1d[5], gate933_0n, initialise);
  C2RI I436 (itint_5n[6], i_5r1d[6], gate933_0n, initialise);
  C2RI I437 (itint_5n[7], i_5r1d[7], gate933_0n, initialise);
  C2RI I438 (itint_5n[8], i_5r1d[8], gate933_0n, initialise);
  C2RI I439 (itint_5n[9], i_5r1d[9], gate933_0n, initialise);
  C2RI I440 (itint_5n[10], i_5r1d[10], gate933_0n, initialise);
  C2RI I441 (itint_5n[11], i_5r1d[11], gate933_0n, initialise);
  C2RI I442 (itint_5n[12], i_5r1d[12], gate933_0n, initialise);
  C2RI I443 (itint_5n[13], i_5r1d[13], gate933_0n, initialise);
  C2RI I444 (itint_5n[14], i_5r1d[14], gate933_0n, initialise);
  C2RI I445 (itint_5n[15], i_5r1d[15], gate933_0n, initialise);
  C2RI I446 (itint_5n[16], i_5r1d[16], gate933_0n, initialise);
  C2RI I447 (itint_5n[17], i_5r1d[17], gate933_0n, initialise);
  C2RI I448 (itint_5n[18], i_5r1d[18], gate933_0n, initialise);
  C2RI I449 (itint_5n[19], i_5r1d[19], gate933_0n, initialise);
  C2RI I450 (itint_5n[20], i_5r1d[20], gate933_0n, initialise);
  C2RI I451 (itint_5n[21], i_5r1d[21], gate933_0n, initialise);
  C2RI I452 (itint_5n[22], i_5r1d[22], gate933_0n, initialise);
  C2RI I453 (itint_5n[23], i_5r1d[23], gate933_0n, initialise);
  C2RI I454 (itint_5n[24], i_5r1d[24], gate933_0n, initialise);
  C2RI I455 (itint_5n[25], i_5r1d[25], gate933_0n, initialise);
  C2RI I456 (itint_5n[26], i_5r1d[26], gate933_0n, initialise);
  C2RI I457 (itint_5n[27], i_5r1d[27], gate933_0n, initialise);
  C2RI I458 (itint_5n[28], i_5r1d[28], gate933_0n, initialise);
  C2RI I459 (itint_5n[29], i_5r1d[29], gate933_0n, initialise);
  C2RI I460 (itint_5n[30], i_5r1d[30], gate933_0n, initialise);
  C2RI I461 (itint_5n[31], i_5r1d[31], gate933_0n, initialise);
  C2RI I462 (itint_5n[32], i_5r1d[32], gate933_0n, initialise);
  C2RI I463 (itint_5n[33], i_5r1d[33], gate933_0n, initialise);
  C2RI I464 (itint_5n[34], i_5r1d[34], gate933_0n, initialise);
  C2RI I465 (ifint_5n[0], i_5r0d[0], gate933_0n, initialise);
  C2RI I466 (ifint_5n[1], i_5r0d[1], gate933_0n, initialise);
  C2RI I467 (ifint_5n[2], i_5r0d[2], gate933_0n, initialise);
  C2RI I468 (ifint_5n[3], i_5r0d[3], gate933_0n, initialise);
  C2RI I469 (ifint_5n[4], i_5r0d[4], gate933_0n, initialise);
  C2RI I470 (ifint_5n[5], i_5r0d[5], gate933_0n, initialise);
  C2RI I471 (ifint_5n[6], i_5r0d[6], gate933_0n, initialise);
  C2RI I472 (ifint_5n[7], i_5r0d[7], gate933_0n, initialise);
  C2RI I473 (ifint_5n[8], i_5r0d[8], gate933_0n, initialise);
  C2RI I474 (ifint_5n[9], i_5r0d[9], gate933_0n, initialise);
  C2RI I475 (ifint_5n[10], i_5r0d[10], gate933_0n, initialise);
  C2RI I476 (ifint_5n[11], i_5r0d[11], gate933_0n, initialise);
  C2RI I477 (ifint_5n[12], i_5r0d[12], gate933_0n, initialise);
  C2RI I478 (ifint_5n[13], i_5r0d[13], gate933_0n, initialise);
  C2RI I479 (ifint_5n[14], i_5r0d[14], gate933_0n, initialise);
  C2RI I480 (ifint_5n[15], i_5r0d[15], gate933_0n, initialise);
  C2RI I481 (ifint_5n[16], i_5r0d[16], gate933_0n, initialise);
  C2RI I482 (ifint_5n[17], i_5r0d[17], gate933_0n, initialise);
  C2RI I483 (ifint_5n[18], i_5r0d[18], gate933_0n, initialise);
  C2RI I484 (ifint_5n[19], i_5r0d[19], gate933_0n, initialise);
  C2RI I485 (ifint_5n[20], i_5r0d[20], gate933_0n, initialise);
  C2RI I486 (ifint_5n[21], i_5r0d[21], gate933_0n, initialise);
  C2RI I487 (ifint_5n[22], i_5r0d[22], gate933_0n, initialise);
  C2RI I488 (ifint_5n[23], i_5r0d[23], gate933_0n, initialise);
  C2RI I489 (ifint_5n[24], i_5r0d[24], gate933_0n, initialise);
  C2RI I490 (ifint_5n[25], i_5r0d[25], gate933_0n, initialise);
  C2RI I491 (ifint_5n[26], i_5r0d[26], gate933_0n, initialise);
  C2RI I492 (ifint_5n[27], i_5r0d[27], gate933_0n, initialise);
  C2RI I493 (ifint_5n[28], i_5r0d[28], gate933_0n, initialise);
  C2RI I494 (ifint_5n[29], i_5r0d[29], gate933_0n, initialise);
  C2RI I495 (ifint_5n[30], i_5r0d[30], gate933_0n, initialise);
  C2RI I496 (ifint_5n[31], i_5r0d[31], gate933_0n, initialise);
  C2RI I497 (ifint_5n[32], i_5r0d[32], gate933_0n, initialise);
  C2RI I498 (ifint_5n[33], i_5r0d[33], gate933_0n, initialise);
  C2RI I499 (ifint_5n[34], i_5r0d[34], gate933_0n, initialise);
  C3 I500 (internal_0n[72], complete930_0n[0], complete930_0n[1], complete930_0n[2]);
  C3 I501 (internal_0n[73], complete930_0n[3], complete930_0n[4], complete930_0n[5]);
  C3 I502 (internal_0n[74], complete930_0n[6], complete930_0n[7], complete930_0n[8]);
  C3 I503 (internal_0n[75], complete930_0n[9], complete930_0n[10], complete930_0n[11]);
  C3 I504 (internal_0n[76], complete930_0n[12], complete930_0n[13], complete930_0n[14]);
  C3 I505 (internal_0n[77], complete930_0n[15], complete930_0n[16], complete930_0n[17]);
  C3 I506 (internal_0n[78], complete930_0n[18], complete930_0n[19], complete930_0n[20]);
  C3 I507 (internal_0n[79], complete930_0n[21], complete930_0n[22], complete930_0n[23]);
  C3 I508 (internal_0n[80], complete930_0n[24], complete930_0n[25], complete930_0n[26]);
  C3 I509 (internal_0n[81], complete930_0n[27], complete930_0n[28], complete930_0n[29]);
  C3 I510 (internal_0n[82], complete930_0n[30], complete930_0n[31], complete930_0n[32]);
  C2 I511 (internal_0n[83], complete930_0n[33], complete930_0n[34]);
  C3 I512 (internal_0n[84], internal_0n[72], internal_0n[73], internal_0n[74]);
  C3 I513 (internal_0n[85], internal_0n[75], internal_0n[76], internal_0n[77]);
  C3 I514 (internal_0n[86], internal_0n[78], internal_0n[79], internal_0n[80]);
  C3 I515 (internal_0n[87], internal_0n[81], internal_0n[82], internal_0n[83]);
  C2 I516 (internal_0n[88], internal_0n[84], internal_0n[85]);
  C2 I517 (internal_0n[89], internal_0n[86], internal_0n[87]);
  C2 I518 (i_4a, internal_0n[88], internal_0n[89]);
  OR2 I519 (complete930_0n[0], ifint_4n[0], itint_4n[0]);
  OR2 I520 (complete930_0n[1], ifint_4n[1], itint_4n[1]);
  OR2 I521 (complete930_0n[2], ifint_4n[2], itint_4n[2]);
  OR2 I522 (complete930_0n[3], ifint_4n[3], itint_4n[3]);
  OR2 I523 (complete930_0n[4], ifint_4n[4], itint_4n[4]);
  OR2 I524 (complete930_0n[5], ifint_4n[5], itint_4n[5]);
  OR2 I525 (complete930_0n[6], ifint_4n[6], itint_4n[6]);
  OR2 I526 (complete930_0n[7], ifint_4n[7], itint_4n[7]);
  OR2 I527 (complete930_0n[8], ifint_4n[8], itint_4n[8]);
  OR2 I528 (complete930_0n[9], ifint_4n[9], itint_4n[9]);
  OR2 I529 (complete930_0n[10], ifint_4n[10], itint_4n[10]);
  OR2 I530 (complete930_0n[11], ifint_4n[11], itint_4n[11]);
  OR2 I531 (complete930_0n[12], ifint_4n[12], itint_4n[12]);
  OR2 I532 (complete930_0n[13], ifint_4n[13], itint_4n[13]);
  OR2 I533 (complete930_0n[14], ifint_4n[14], itint_4n[14]);
  OR2 I534 (complete930_0n[15], ifint_4n[15], itint_4n[15]);
  OR2 I535 (complete930_0n[16], ifint_4n[16], itint_4n[16]);
  OR2 I536 (complete930_0n[17], ifint_4n[17], itint_4n[17]);
  OR2 I537 (complete930_0n[18], ifint_4n[18], itint_4n[18]);
  OR2 I538 (complete930_0n[19], ifint_4n[19], itint_4n[19]);
  OR2 I539 (complete930_0n[20], ifint_4n[20], itint_4n[20]);
  OR2 I540 (complete930_0n[21], ifint_4n[21], itint_4n[21]);
  OR2 I541 (complete930_0n[22], ifint_4n[22], itint_4n[22]);
  OR2 I542 (complete930_0n[23], ifint_4n[23], itint_4n[23]);
  OR2 I543 (complete930_0n[24], ifint_4n[24], itint_4n[24]);
  OR2 I544 (complete930_0n[25], ifint_4n[25], itint_4n[25]);
  OR2 I545 (complete930_0n[26], ifint_4n[26], itint_4n[26]);
  OR2 I546 (complete930_0n[27], ifint_4n[27], itint_4n[27]);
  OR2 I547 (complete930_0n[28], ifint_4n[28], itint_4n[28]);
  OR2 I548 (complete930_0n[29], ifint_4n[29], itint_4n[29]);
  OR2 I549 (complete930_0n[30], ifint_4n[30], itint_4n[30]);
  OR2 I550 (complete930_0n[31], ifint_4n[31], itint_4n[31]);
  OR2 I551 (complete930_0n[32], ifint_4n[32], itint_4n[32]);
  OR2 I552 (complete930_0n[33], ifint_4n[33], itint_4n[33]);
  OR2 I553 (complete930_0n[34], ifint_4n[34], itint_4n[34]);
  INV I554 (gate929_0n, iaint_4n);
  C2RI I555 (itint_4n[0], i_4r1d[0], gate929_0n, initialise);
  C2RI I556 (itint_4n[1], i_4r1d[1], gate929_0n, initialise);
  C2RI I557 (itint_4n[2], i_4r1d[2], gate929_0n, initialise);
  C2RI I558 (itint_4n[3], i_4r1d[3], gate929_0n, initialise);
  C2RI I559 (itint_4n[4], i_4r1d[4], gate929_0n, initialise);
  C2RI I560 (itint_4n[5], i_4r1d[5], gate929_0n, initialise);
  C2RI I561 (itint_4n[6], i_4r1d[6], gate929_0n, initialise);
  C2RI I562 (itint_4n[7], i_4r1d[7], gate929_0n, initialise);
  C2RI I563 (itint_4n[8], i_4r1d[8], gate929_0n, initialise);
  C2RI I564 (itint_4n[9], i_4r1d[9], gate929_0n, initialise);
  C2RI I565 (itint_4n[10], i_4r1d[10], gate929_0n, initialise);
  C2RI I566 (itint_4n[11], i_4r1d[11], gate929_0n, initialise);
  C2RI I567 (itint_4n[12], i_4r1d[12], gate929_0n, initialise);
  C2RI I568 (itint_4n[13], i_4r1d[13], gate929_0n, initialise);
  C2RI I569 (itint_4n[14], i_4r1d[14], gate929_0n, initialise);
  C2RI I570 (itint_4n[15], i_4r1d[15], gate929_0n, initialise);
  C2RI I571 (itint_4n[16], i_4r1d[16], gate929_0n, initialise);
  C2RI I572 (itint_4n[17], i_4r1d[17], gate929_0n, initialise);
  C2RI I573 (itint_4n[18], i_4r1d[18], gate929_0n, initialise);
  C2RI I574 (itint_4n[19], i_4r1d[19], gate929_0n, initialise);
  C2RI I575 (itint_4n[20], i_4r1d[20], gate929_0n, initialise);
  C2RI I576 (itint_4n[21], i_4r1d[21], gate929_0n, initialise);
  C2RI I577 (itint_4n[22], i_4r1d[22], gate929_0n, initialise);
  C2RI I578 (itint_4n[23], i_4r1d[23], gate929_0n, initialise);
  C2RI I579 (itint_4n[24], i_4r1d[24], gate929_0n, initialise);
  C2RI I580 (itint_4n[25], i_4r1d[25], gate929_0n, initialise);
  C2RI I581 (itint_4n[26], i_4r1d[26], gate929_0n, initialise);
  C2RI I582 (itint_4n[27], i_4r1d[27], gate929_0n, initialise);
  C2RI I583 (itint_4n[28], i_4r1d[28], gate929_0n, initialise);
  C2RI I584 (itint_4n[29], i_4r1d[29], gate929_0n, initialise);
  C2RI I585 (itint_4n[30], i_4r1d[30], gate929_0n, initialise);
  C2RI I586 (itint_4n[31], i_4r1d[31], gate929_0n, initialise);
  C2RI I587 (itint_4n[32], i_4r1d[32], gate929_0n, initialise);
  C2RI I588 (itint_4n[33], i_4r1d[33], gate929_0n, initialise);
  C2RI I589 (itint_4n[34], i_4r1d[34], gate929_0n, initialise);
  C2RI I590 (ifint_4n[0], i_4r0d[0], gate929_0n, initialise);
  C2RI I591 (ifint_4n[1], i_4r0d[1], gate929_0n, initialise);
  C2RI I592 (ifint_4n[2], i_4r0d[2], gate929_0n, initialise);
  C2RI I593 (ifint_4n[3], i_4r0d[3], gate929_0n, initialise);
  C2RI I594 (ifint_4n[4], i_4r0d[4], gate929_0n, initialise);
  C2RI I595 (ifint_4n[5], i_4r0d[5], gate929_0n, initialise);
  C2RI I596 (ifint_4n[6], i_4r0d[6], gate929_0n, initialise);
  C2RI I597 (ifint_4n[7], i_4r0d[7], gate929_0n, initialise);
  C2RI I598 (ifint_4n[8], i_4r0d[8], gate929_0n, initialise);
  C2RI I599 (ifint_4n[9], i_4r0d[9], gate929_0n, initialise);
  C2RI I600 (ifint_4n[10], i_4r0d[10], gate929_0n, initialise);
  C2RI I601 (ifint_4n[11], i_4r0d[11], gate929_0n, initialise);
  C2RI I602 (ifint_4n[12], i_4r0d[12], gate929_0n, initialise);
  C2RI I603 (ifint_4n[13], i_4r0d[13], gate929_0n, initialise);
  C2RI I604 (ifint_4n[14], i_4r0d[14], gate929_0n, initialise);
  C2RI I605 (ifint_4n[15], i_4r0d[15], gate929_0n, initialise);
  C2RI I606 (ifint_4n[16], i_4r0d[16], gate929_0n, initialise);
  C2RI I607 (ifint_4n[17], i_4r0d[17], gate929_0n, initialise);
  C2RI I608 (ifint_4n[18], i_4r0d[18], gate929_0n, initialise);
  C2RI I609 (ifint_4n[19], i_4r0d[19], gate929_0n, initialise);
  C2RI I610 (ifint_4n[20], i_4r0d[20], gate929_0n, initialise);
  C2RI I611 (ifint_4n[21], i_4r0d[21], gate929_0n, initialise);
  C2RI I612 (ifint_4n[22], i_4r0d[22], gate929_0n, initialise);
  C2RI I613 (ifint_4n[23], i_4r0d[23], gate929_0n, initialise);
  C2RI I614 (ifint_4n[24], i_4r0d[24], gate929_0n, initialise);
  C2RI I615 (ifint_4n[25], i_4r0d[25], gate929_0n, initialise);
  C2RI I616 (ifint_4n[26], i_4r0d[26], gate929_0n, initialise);
  C2RI I617 (ifint_4n[27], i_4r0d[27], gate929_0n, initialise);
  C2RI I618 (ifint_4n[28], i_4r0d[28], gate929_0n, initialise);
  C2RI I619 (ifint_4n[29], i_4r0d[29], gate929_0n, initialise);
  C2RI I620 (ifint_4n[30], i_4r0d[30], gate929_0n, initialise);
  C2RI I621 (ifint_4n[31], i_4r0d[31], gate929_0n, initialise);
  C2RI I622 (ifint_4n[32], i_4r0d[32], gate929_0n, initialise);
  C2RI I623 (ifint_4n[33], i_4r0d[33], gate929_0n, initialise);
  C2RI I624 (ifint_4n[34], i_4r0d[34], gate929_0n, initialise);
  C3 I625 (internal_0n[90], complete926_0n[0], complete926_0n[1], complete926_0n[2]);
  C3 I626 (internal_0n[91], complete926_0n[3], complete926_0n[4], complete926_0n[5]);
  C3 I627 (internal_0n[92], complete926_0n[6], complete926_0n[7], complete926_0n[8]);
  C3 I628 (internal_0n[93], complete926_0n[9], complete926_0n[10], complete926_0n[11]);
  C3 I629 (internal_0n[94], complete926_0n[12], complete926_0n[13], complete926_0n[14]);
  C3 I630 (internal_0n[95], complete926_0n[15], complete926_0n[16], complete926_0n[17]);
  C3 I631 (internal_0n[96], complete926_0n[18], complete926_0n[19], complete926_0n[20]);
  C3 I632 (internal_0n[97], complete926_0n[21], complete926_0n[22], complete926_0n[23]);
  C3 I633 (internal_0n[98], complete926_0n[24], complete926_0n[25], complete926_0n[26]);
  C3 I634 (internal_0n[99], complete926_0n[27], complete926_0n[28], complete926_0n[29]);
  C3 I635 (internal_0n[100], complete926_0n[30], complete926_0n[31], complete926_0n[32]);
  C2 I636 (internal_0n[101], complete926_0n[33], complete926_0n[34]);
  C3 I637 (internal_0n[102], internal_0n[90], internal_0n[91], internal_0n[92]);
  C3 I638 (internal_0n[103], internal_0n[93], internal_0n[94], internal_0n[95]);
  C3 I639 (internal_0n[104], internal_0n[96], internal_0n[97], internal_0n[98]);
  C3 I640 (internal_0n[105], internal_0n[99], internal_0n[100], internal_0n[101]);
  C2 I641 (internal_0n[106], internal_0n[102], internal_0n[103]);
  C2 I642 (internal_0n[107], internal_0n[104], internal_0n[105]);
  C2 I643 (i_3a, internal_0n[106], internal_0n[107]);
  OR2 I644 (complete926_0n[0], ifint_3n[0], itint_3n[0]);
  OR2 I645 (complete926_0n[1], ifint_3n[1], itint_3n[1]);
  OR2 I646 (complete926_0n[2], ifint_3n[2], itint_3n[2]);
  OR2 I647 (complete926_0n[3], ifint_3n[3], itint_3n[3]);
  OR2 I648 (complete926_0n[4], ifint_3n[4], itint_3n[4]);
  OR2 I649 (complete926_0n[5], ifint_3n[5], itint_3n[5]);
  OR2 I650 (complete926_0n[6], ifint_3n[6], itint_3n[6]);
  OR2 I651 (complete926_0n[7], ifint_3n[7], itint_3n[7]);
  OR2 I652 (complete926_0n[8], ifint_3n[8], itint_3n[8]);
  OR2 I653 (complete926_0n[9], ifint_3n[9], itint_3n[9]);
  OR2 I654 (complete926_0n[10], ifint_3n[10], itint_3n[10]);
  OR2 I655 (complete926_0n[11], ifint_3n[11], itint_3n[11]);
  OR2 I656 (complete926_0n[12], ifint_3n[12], itint_3n[12]);
  OR2 I657 (complete926_0n[13], ifint_3n[13], itint_3n[13]);
  OR2 I658 (complete926_0n[14], ifint_3n[14], itint_3n[14]);
  OR2 I659 (complete926_0n[15], ifint_3n[15], itint_3n[15]);
  OR2 I660 (complete926_0n[16], ifint_3n[16], itint_3n[16]);
  OR2 I661 (complete926_0n[17], ifint_3n[17], itint_3n[17]);
  OR2 I662 (complete926_0n[18], ifint_3n[18], itint_3n[18]);
  OR2 I663 (complete926_0n[19], ifint_3n[19], itint_3n[19]);
  OR2 I664 (complete926_0n[20], ifint_3n[20], itint_3n[20]);
  OR2 I665 (complete926_0n[21], ifint_3n[21], itint_3n[21]);
  OR2 I666 (complete926_0n[22], ifint_3n[22], itint_3n[22]);
  OR2 I667 (complete926_0n[23], ifint_3n[23], itint_3n[23]);
  OR2 I668 (complete926_0n[24], ifint_3n[24], itint_3n[24]);
  OR2 I669 (complete926_0n[25], ifint_3n[25], itint_3n[25]);
  OR2 I670 (complete926_0n[26], ifint_3n[26], itint_3n[26]);
  OR2 I671 (complete926_0n[27], ifint_3n[27], itint_3n[27]);
  OR2 I672 (complete926_0n[28], ifint_3n[28], itint_3n[28]);
  OR2 I673 (complete926_0n[29], ifint_3n[29], itint_3n[29]);
  OR2 I674 (complete926_0n[30], ifint_3n[30], itint_3n[30]);
  OR2 I675 (complete926_0n[31], ifint_3n[31], itint_3n[31]);
  OR2 I676 (complete926_0n[32], ifint_3n[32], itint_3n[32]);
  OR2 I677 (complete926_0n[33], ifint_3n[33], itint_3n[33]);
  OR2 I678 (complete926_0n[34], ifint_3n[34], itint_3n[34]);
  INV I679 (gate925_0n, iaint_3n);
  C2RI I680 (itint_3n[0], i_3r1d[0], gate925_0n, initialise);
  C2RI I681 (itint_3n[1], i_3r1d[1], gate925_0n, initialise);
  C2RI I682 (itint_3n[2], i_3r1d[2], gate925_0n, initialise);
  C2RI I683 (itint_3n[3], i_3r1d[3], gate925_0n, initialise);
  C2RI I684 (itint_3n[4], i_3r1d[4], gate925_0n, initialise);
  C2RI I685 (itint_3n[5], i_3r1d[5], gate925_0n, initialise);
  C2RI I686 (itint_3n[6], i_3r1d[6], gate925_0n, initialise);
  C2RI I687 (itint_3n[7], i_3r1d[7], gate925_0n, initialise);
  C2RI I688 (itint_3n[8], i_3r1d[8], gate925_0n, initialise);
  C2RI I689 (itint_3n[9], i_3r1d[9], gate925_0n, initialise);
  C2RI I690 (itint_3n[10], i_3r1d[10], gate925_0n, initialise);
  C2RI I691 (itint_3n[11], i_3r1d[11], gate925_0n, initialise);
  C2RI I692 (itint_3n[12], i_3r1d[12], gate925_0n, initialise);
  C2RI I693 (itint_3n[13], i_3r1d[13], gate925_0n, initialise);
  C2RI I694 (itint_3n[14], i_3r1d[14], gate925_0n, initialise);
  C2RI I695 (itint_3n[15], i_3r1d[15], gate925_0n, initialise);
  C2RI I696 (itint_3n[16], i_3r1d[16], gate925_0n, initialise);
  C2RI I697 (itint_3n[17], i_3r1d[17], gate925_0n, initialise);
  C2RI I698 (itint_3n[18], i_3r1d[18], gate925_0n, initialise);
  C2RI I699 (itint_3n[19], i_3r1d[19], gate925_0n, initialise);
  C2RI I700 (itint_3n[20], i_3r1d[20], gate925_0n, initialise);
  C2RI I701 (itint_3n[21], i_3r1d[21], gate925_0n, initialise);
  C2RI I702 (itint_3n[22], i_3r1d[22], gate925_0n, initialise);
  C2RI I703 (itint_3n[23], i_3r1d[23], gate925_0n, initialise);
  C2RI I704 (itint_3n[24], i_3r1d[24], gate925_0n, initialise);
  C2RI I705 (itint_3n[25], i_3r1d[25], gate925_0n, initialise);
  C2RI I706 (itint_3n[26], i_3r1d[26], gate925_0n, initialise);
  C2RI I707 (itint_3n[27], i_3r1d[27], gate925_0n, initialise);
  C2RI I708 (itint_3n[28], i_3r1d[28], gate925_0n, initialise);
  C2RI I709 (itint_3n[29], i_3r1d[29], gate925_0n, initialise);
  C2RI I710 (itint_3n[30], i_3r1d[30], gate925_0n, initialise);
  C2RI I711 (itint_3n[31], i_3r1d[31], gate925_0n, initialise);
  C2RI I712 (itint_3n[32], i_3r1d[32], gate925_0n, initialise);
  C2RI I713 (itint_3n[33], i_3r1d[33], gate925_0n, initialise);
  C2RI I714 (itint_3n[34], i_3r1d[34], gate925_0n, initialise);
  C2RI I715 (ifint_3n[0], i_3r0d[0], gate925_0n, initialise);
  C2RI I716 (ifint_3n[1], i_3r0d[1], gate925_0n, initialise);
  C2RI I717 (ifint_3n[2], i_3r0d[2], gate925_0n, initialise);
  C2RI I718 (ifint_3n[3], i_3r0d[3], gate925_0n, initialise);
  C2RI I719 (ifint_3n[4], i_3r0d[4], gate925_0n, initialise);
  C2RI I720 (ifint_3n[5], i_3r0d[5], gate925_0n, initialise);
  C2RI I721 (ifint_3n[6], i_3r0d[6], gate925_0n, initialise);
  C2RI I722 (ifint_3n[7], i_3r0d[7], gate925_0n, initialise);
  C2RI I723 (ifint_3n[8], i_3r0d[8], gate925_0n, initialise);
  C2RI I724 (ifint_3n[9], i_3r0d[9], gate925_0n, initialise);
  C2RI I725 (ifint_3n[10], i_3r0d[10], gate925_0n, initialise);
  C2RI I726 (ifint_3n[11], i_3r0d[11], gate925_0n, initialise);
  C2RI I727 (ifint_3n[12], i_3r0d[12], gate925_0n, initialise);
  C2RI I728 (ifint_3n[13], i_3r0d[13], gate925_0n, initialise);
  C2RI I729 (ifint_3n[14], i_3r0d[14], gate925_0n, initialise);
  C2RI I730 (ifint_3n[15], i_3r0d[15], gate925_0n, initialise);
  C2RI I731 (ifint_3n[16], i_3r0d[16], gate925_0n, initialise);
  C2RI I732 (ifint_3n[17], i_3r0d[17], gate925_0n, initialise);
  C2RI I733 (ifint_3n[18], i_3r0d[18], gate925_0n, initialise);
  C2RI I734 (ifint_3n[19], i_3r0d[19], gate925_0n, initialise);
  C2RI I735 (ifint_3n[20], i_3r0d[20], gate925_0n, initialise);
  C2RI I736 (ifint_3n[21], i_3r0d[21], gate925_0n, initialise);
  C2RI I737 (ifint_3n[22], i_3r0d[22], gate925_0n, initialise);
  C2RI I738 (ifint_3n[23], i_3r0d[23], gate925_0n, initialise);
  C2RI I739 (ifint_3n[24], i_3r0d[24], gate925_0n, initialise);
  C2RI I740 (ifint_3n[25], i_3r0d[25], gate925_0n, initialise);
  C2RI I741 (ifint_3n[26], i_3r0d[26], gate925_0n, initialise);
  C2RI I742 (ifint_3n[27], i_3r0d[27], gate925_0n, initialise);
  C2RI I743 (ifint_3n[28], i_3r0d[28], gate925_0n, initialise);
  C2RI I744 (ifint_3n[29], i_3r0d[29], gate925_0n, initialise);
  C2RI I745 (ifint_3n[30], i_3r0d[30], gate925_0n, initialise);
  C2RI I746 (ifint_3n[31], i_3r0d[31], gate925_0n, initialise);
  C2RI I747 (ifint_3n[32], i_3r0d[32], gate925_0n, initialise);
  C2RI I748 (ifint_3n[33], i_3r0d[33], gate925_0n, initialise);
  C2RI I749 (ifint_3n[34], i_3r0d[34], gate925_0n, initialise);
  C3 I750 (internal_0n[108], complete922_0n[0], complete922_0n[1], complete922_0n[2]);
  C3 I751 (internal_0n[109], complete922_0n[3], complete922_0n[4], complete922_0n[5]);
  C3 I752 (internal_0n[110], complete922_0n[6], complete922_0n[7], complete922_0n[8]);
  C3 I753 (internal_0n[111], complete922_0n[9], complete922_0n[10], complete922_0n[11]);
  C3 I754 (internal_0n[112], complete922_0n[12], complete922_0n[13], complete922_0n[14]);
  C3 I755 (internal_0n[113], complete922_0n[15], complete922_0n[16], complete922_0n[17]);
  C3 I756 (internal_0n[114], complete922_0n[18], complete922_0n[19], complete922_0n[20]);
  C3 I757 (internal_0n[115], complete922_0n[21], complete922_0n[22], complete922_0n[23]);
  C3 I758 (internal_0n[116], complete922_0n[24], complete922_0n[25], complete922_0n[26]);
  C3 I759 (internal_0n[117], complete922_0n[27], complete922_0n[28], complete922_0n[29]);
  C3 I760 (internal_0n[118], complete922_0n[30], complete922_0n[31], complete922_0n[32]);
  C2 I761 (internal_0n[119], complete922_0n[33], complete922_0n[34]);
  C3 I762 (internal_0n[120], internal_0n[108], internal_0n[109], internal_0n[110]);
  C3 I763 (internal_0n[121], internal_0n[111], internal_0n[112], internal_0n[113]);
  C3 I764 (internal_0n[122], internal_0n[114], internal_0n[115], internal_0n[116]);
  C3 I765 (internal_0n[123], internal_0n[117], internal_0n[118], internal_0n[119]);
  C2 I766 (internal_0n[124], internal_0n[120], internal_0n[121]);
  C2 I767 (internal_0n[125], internal_0n[122], internal_0n[123]);
  C2 I768 (i_2a, internal_0n[124], internal_0n[125]);
  OR2 I769 (complete922_0n[0], ifint_2n[0], itint_2n[0]);
  OR2 I770 (complete922_0n[1], ifint_2n[1], itint_2n[1]);
  OR2 I771 (complete922_0n[2], ifint_2n[2], itint_2n[2]);
  OR2 I772 (complete922_0n[3], ifint_2n[3], itint_2n[3]);
  OR2 I773 (complete922_0n[4], ifint_2n[4], itint_2n[4]);
  OR2 I774 (complete922_0n[5], ifint_2n[5], itint_2n[5]);
  OR2 I775 (complete922_0n[6], ifint_2n[6], itint_2n[6]);
  OR2 I776 (complete922_0n[7], ifint_2n[7], itint_2n[7]);
  OR2 I777 (complete922_0n[8], ifint_2n[8], itint_2n[8]);
  OR2 I778 (complete922_0n[9], ifint_2n[9], itint_2n[9]);
  OR2 I779 (complete922_0n[10], ifint_2n[10], itint_2n[10]);
  OR2 I780 (complete922_0n[11], ifint_2n[11], itint_2n[11]);
  OR2 I781 (complete922_0n[12], ifint_2n[12], itint_2n[12]);
  OR2 I782 (complete922_0n[13], ifint_2n[13], itint_2n[13]);
  OR2 I783 (complete922_0n[14], ifint_2n[14], itint_2n[14]);
  OR2 I784 (complete922_0n[15], ifint_2n[15], itint_2n[15]);
  OR2 I785 (complete922_0n[16], ifint_2n[16], itint_2n[16]);
  OR2 I786 (complete922_0n[17], ifint_2n[17], itint_2n[17]);
  OR2 I787 (complete922_0n[18], ifint_2n[18], itint_2n[18]);
  OR2 I788 (complete922_0n[19], ifint_2n[19], itint_2n[19]);
  OR2 I789 (complete922_0n[20], ifint_2n[20], itint_2n[20]);
  OR2 I790 (complete922_0n[21], ifint_2n[21], itint_2n[21]);
  OR2 I791 (complete922_0n[22], ifint_2n[22], itint_2n[22]);
  OR2 I792 (complete922_0n[23], ifint_2n[23], itint_2n[23]);
  OR2 I793 (complete922_0n[24], ifint_2n[24], itint_2n[24]);
  OR2 I794 (complete922_0n[25], ifint_2n[25], itint_2n[25]);
  OR2 I795 (complete922_0n[26], ifint_2n[26], itint_2n[26]);
  OR2 I796 (complete922_0n[27], ifint_2n[27], itint_2n[27]);
  OR2 I797 (complete922_0n[28], ifint_2n[28], itint_2n[28]);
  OR2 I798 (complete922_0n[29], ifint_2n[29], itint_2n[29]);
  OR2 I799 (complete922_0n[30], ifint_2n[30], itint_2n[30]);
  OR2 I800 (complete922_0n[31], ifint_2n[31], itint_2n[31]);
  OR2 I801 (complete922_0n[32], ifint_2n[32], itint_2n[32]);
  OR2 I802 (complete922_0n[33], ifint_2n[33], itint_2n[33]);
  OR2 I803 (complete922_0n[34], ifint_2n[34], itint_2n[34]);
  INV I804 (gate921_0n, iaint_2n);
  C2RI I805 (itint_2n[0], i_2r1d[0], gate921_0n, initialise);
  C2RI I806 (itint_2n[1], i_2r1d[1], gate921_0n, initialise);
  C2RI I807 (itint_2n[2], i_2r1d[2], gate921_0n, initialise);
  C2RI I808 (itint_2n[3], i_2r1d[3], gate921_0n, initialise);
  C2RI I809 (itint_2n[4], i_2r1d[4], gate921_0n, initialise);
  C2RI I810 (itint_2n[5], i_2r1d[5], gate921_0n, initialise);
  C2RI I811 (itint_2n[6], i_2r1d[6], gate921_0n, initialise);
  C2RI I812 (itint_2n[7], i_2r1d[7], gate921_0n, initialise);
  C2RI I813 (itint_2n[8], i_2r1d[8], gate921_0n, initialise);
  C2RI I814 (itint_2n[9], i_2r1d[9], gate921_0n, initialise);
  C2RI I815 (itint_2n[10], i_2r1d[10], gate921_0n, initialise);
  C2RI I816 (itint_2n[11], i_2r1d[11], gate921_0n, initialise);
  C2RI I817 (itint_2n[12], i_2r1d[12], gate921_0n, initialise);
  C2RI I818 (itint_2n[13], i_2r1d[13], gate921_0n, initialise);
  C2RI I819 (itint_2n[14], i_2r1d[14], gate921_0n, initialise);
  C2RI I820 (itint_2n[15], i_2r1d[15], gate921_0n, initialise);
  C2RI I821 (itint_2n[16], i_2r1d[16], gate921_0n, initialise);
  C2RI I822 (itint_2n[17], i_2r1d[17], gate921_0n, initialise);
  C2RI I823 (itint_2n[18], i_2r1d[18], gate921_0n, initialise);
  C2RI I824 (itint_2n[19], i_2r1d[19], gate921_0n, initialise);
  C2RI I825 (itint_2n[20], i_2r1d[20], gate921_0n, initialise);
  C2RI I826 (itint_2n[21], i_2r1d[21], gate921_0n, initialise);
  C2RI I827 (itint_2n[22], i_2r1d[22], gate921_0n, initialise);
  C2RI I828 (itint_2n[23], i_2r1d[23], gate921_0n, initialise);
  C2RI I829 (itint_2n[24], i_2r1d[24], gate921_0n, initialise);
  C2RI I830 (itint_2n[25], i_2r1d[25], gate921_0n, initialise);
  C2RI I831 (itint_2n[26], i_2r1d[26], gate921_0n, initialise);
  C2RI I832 (itint_2n[27], i_2r1d[27], gate921_0n, initialise);
  C2RI I833 (itint_2n[28], i_2r1d[28], gate921_0n, initialise);
  C2RI I834 (itint_2n[29], i_2r1d[29], gate921_0n, initialise);
  C2RI I835 (itint_2n[30], i_2r1d[30], gate921_0n, initialise);
  C2RI I836 (itint_2n[31], i_2r1d[31], gate921_0n, initialise);
  C2RI I837 (itint_2n[32], i_2r1d[32], gate921_0n, initialise);
  C2RI I838 (itint_2n[33], i_2r1d[33], gate921_0n, initialise);
  C2RI I839 (itint_2n[34], i_2r1d[34], gate921_0n, initialise);
  C2RI I840 (ifint_2n[0], i_2r0d[0], gate921_0n, initialise);
  C2RI I841 (ifint_2n[1], i_2r0d[1], gate921_0n, initialise);
  C2RI I842 (ifint_2n[2], i_2r0d[2], gate921_0n, initialise);
  C2RI I843 (ifint_2n[3], i_2r0d[3], gate921_0n, initialise);
  C2RI I844 (ifint_2n[4], i_2r0d[4], gate921_0n, initialise);
  C2RI I845 (ifint_2n[5], i_2r0d[5], gate921_0n, initialise);
  C2RI I846 (ifint_2n[6], i_2r0d[6], gate921_0n, initialise);
  C2RI I847 (ifint_2n[7], i_2r0d[7], gate921_0n, initialise);
  C2RI I848 (ifint_2n[8], i_2r0d[8], gate921_0n, initialise);
  C2RI I849 (ifint_2n[9], i_2r0d[9], gate921_0n, initialise);
  C2RI I850 (ifint_2n[10], i_2r0d[10], gate921_0n, initialise);
  C2RI I851 (ifint_2n[11], i_2r0d[11], gate921_0n, initialise);
  C2RI I852 (ifint_2n[12], i_2r0d[12], gate921_0n, initialise);
  C2RI I853 (ifint_2n[13], i_2r0d[13], gate921_0n, initialise);
  C2RI I854 (ifint_2n[14], i_2r0d[14], gate921_0n, initialise);
  C2RI I855 (ifint_2n[15], i_2r0d[15], gate921_0n, initialise);
  C2RI I856 (ifint_2n[16], i_2r0d[16], gate921_0n, initialise);
  C2RI I857 (ifint_2n[17], i_2r0d[17], gate921_0n, initialise);
  C2RI I858 (ifint_2n[18], i_2r0d[18], gate921_0n, initialise);
  C2RI I859 (ifint_2n[19], i_2r0d[19], gate921_0n, initialise);
  C2RI I860 (ifint_2n[20], i_2r0d[20], gate921_0n, initialise);
  C2RI I861 (ifint_2n[21], i_2r0d[21], gate921_0n, initialise);
  C2RI I862 (ifint_2n[22], i_2r0d[22], gate921_0n, initialise);
  C2RI I863 (ifint_2n[23], i_2r0d[23], gate921_0n, initialise);
  C2RI I864 (ifint_2n[24], i_2r0d[24], gate921_0n, initialise);
  C2RI I865 (ifint_2n[25], i_2r0d[25], gate921_0n, initialise);
  C2RI I866 (ifint_2n[26], i_2r0d[26], gate921_0n, initialise);
  C2RI I867 (ifint_2n[27], i_2r0d[27], gate921_0n, initialise);
  C2RI I868 (ifint_2n[28], i_2r0d[28], gate921_0n, initialise);
  C2RI I869 (ifint_2n[29], i_2r0d[29], gate921_0n, initialise);
  C2RI I870 (ifint_2n[30], i_2r0d[30], gate921_0n, initialise);
  C2RI I871 (ifint_2n[31], i_2r0d[31], gate921_0n, initialise);
  C2RI I872 (ifint_2n[32], i_2r0d[32], gate921_0n, initialise);
  C2RI I873 (ifint_2n[33], i_2r0d[33], gate921_0n, initialise);
  C2RI I874 (ifint_2n[34], i_2r0d[34], gate921_0n, initialise);
  C3 I875 (internal_0n[126], complete918_0n[0], complete918_0n[1], complete918_0n[2]);
  C3 I876 (internal_0n[127], complete918_0n[3], complete918_0n[4], complete918_0n[5]);
  C3 I877 (internal_0n[128], complete918_0n[6], complete918_0n[7], complete918_0n[8]);
  C3 I878 (internal_0n[129], complete918_0n[9], complete918_0n[10], complete918_0n[11]);
  C3 I879 (internal_0n[130], complete918_0n[12], complete918_0n[13], complete918_0n[14]);
  C3 I880 (internal_0n[131], complete918_0n[15], complete918_0n[16], complete918_0n[17]);
  C3 I881 (internal_0n[132], complete918_0n[18], complete918_0n[19], complete918_0n[20]);
  C3 I882 (internal_0n[133], complete918_0n[21], complete918_0n[22], complete918_0n[23]);
  C3 I883 (internal_0n[134], complete918_0n[24], complete918_0n[25], complete918_0n[26]);
  C3 I884 (internal_0n[135], complete918_0n[27], complete918_0n[28], complete918_0n[29]);
  C3 I885 (internal_0n[136], complete918_0n[30], complete918_0n[31], complete918_0n[32]);
  C2 I886 (internal_0n[137], complete918_0n[33], complete918_0n[34]);
  C3 I887 (internal_0n[138], internal_0n[126], internal_0n[127], internal_0n[128]);
  C3 I888 (internal_0n[139], internal_0n[129], internal_0n[130], internal_0n[131]);
  C3 I889 (internal_0n[140], internal_0n[132], internal_0n[133], internal_0n[134]);
  C3 I890 (internal_0n[141], internal_0n[135], internal_0n[136], internal_0n[137]);
  C2 I891 (internal_0n[142], internal_0n[138], internal_0n[139]);
  C2 I892 (internal_0n[143], internal_0n[140], internal_0n[141]);
  C2 I893 (i_1a, internal_0n[142], internal_0n[143]);
  OR2 I894 (complete918_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I895 (complete918_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I896 (complete918_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I897 (complete918_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I898 (complete918_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I899 (complete918_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I900 (complete918_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I901 (complete918_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I902 (complete918_0n[8], ifint_1n[8], itint_1n[8]);
  OR2 I903 (complete918_0n[9], ifint_1n[9], itint_1n[9]);
  OR2 I904 (complete918_0n[10], ifint_1n[10], itint_1n[10]);
  OR2 I905 (complete918_0n[11], ifint_1n[11], itint_1n[11]);
  OR2 I906 (complete918_0n[12], ifint_1n[12], itint_1n[12]);
  OR2 I907 (complete918_0n[13], ifint_1n[13], itint_1n[13]);
  OR2 I908 (complete918_0n[14], ifint_1n[14], itint_1n[14]);
  OR2 I909 (complete918_0n[15], ifint_1n[15], itint_1n[15]);
  OR2 I910 (complete918_0n[16], ifint_1n[16], itint_1n[16]);
  OR2 I911 (complete918_0n[17], ifint_1n[17], itint_1n[17]);
  OR2 I912 (complete918_0n[18], ifint_1n[18], itint_1n[18]);
  OR2 I913 (complete918_0n[19], ifint_1n[19], itint_1n[19]);
  OR2 I914 (complete918_0n[20], ifint_1n[20], itint_1n[20]);
  OR2 I915 (complete918_0n[21], ifint_1n[21], itint_1n[21]);
  OR2 I916 (complete918_0n[22], ifint_1n[22], itint_1n[22]);
  OR2 I917 (complete918_0n[23], ifint_1n[23], itint_1n[23]);
  OR2 I918 (complete918_0n[24], ifint_1n[24], itint_1n[24]);
  OR2 I919 (complete918_0n[25], ifint_1n[25], itint_1n[25]);
  OR2 I920 (complete918_0n[26], ifint_1n[26], itint_1n[26]);
  OR2 I921 (complete918_0n[27], ifint_1n[27], itint_1n[27]);
  OR2 I922 (complete918_0n[28], ifint_1n[28], itint_1n[28]);
  OR2 I923 (complete918_0n[29], ifint_1n[29], itint_1n[29]);
  OR2 I924 (complete918_0n[30], ifint_1n[30], itint_1n[30]);
  OR2 I925 (complete918_0n[31], ifint_1n[31], itint_1n[31]);
  OR2 I926 (complete918_0n[32], ifint_1n[32], itint_1n[32]);
  OR2 I927 (complete918_0n[33], ifint_1n[33], itint_1n[33]);
  OR2 I928 (complete918_0n[34], ifint_1n[34], itint_1n[34]);
  INV I929 (gate917_0n, iaint_1n);
  C2RI I930 (itint_1n[0], i_1r1d[0], gate917_0n, initialise);
  C2RI I931 (itint_1n[1], i_1r1d[1], gate917_0n, initialise);
  C2RI I932 (itint_1n[2], i_1r1d[2], gate917_0n, initialise);
  C2RI I933 (itint_1n[3], i_1r1d[3], gate917_0n, initialise);
  C2RI I934 (itint_1n[4], i_1r1d[4], gate917_0n, initialise);
  C2RI I935 (itint_1n[5], i_1r1d[5], gate917_0n, initialise);
  C2RI I936 (itint_1n[6], i_1r1d[6], gate917_0n, initialise);
  C2RI I937 (itint_1n[7], i_1r1d[7], gate917_0n, initialise);
  C2RI I938 (itint_1n[8], i_1r1d[8], gate917_0n, initialise);
  C2RI I939 (itint_1n[9], i_1r1d[9], gate917_0n, initialise);
  C2RI I940 (itint_1n[10], i_1r1d[10], gate917_0n, initialise);
  C2RI I941 (itint_1n[11], i_1r1d[11], gate917_0n, initialise);
  C2RI I942 (itint_1n[12], i_1r1d[12], gate917_0n, initialise);
  C2RI I943 (itint_1n[13], i_1r1d[13], gate917_0n, initialise);
  C2RI I944 (itint_1n[14], i_1r1d[14], gate917_0n, initialise);
  C2RI I945 (itint_1n[15], i_1r1d[15], gate917_0n, initialise);
  C2RI I946 (itint_1n[16], i_1r1d[16], gate917_0n, initialise);
  C2RI I947 (itint_1n[17], i_1r1d[17], gate917_0n, initialise);
  C2RI I948 (itint_1n[18], i_1r1d[18], gate917_0n, initialise);
  C2RI I949 (itint_1n[19], i_1r1d[19], gate917_0n, initialise);
  C2RI I950 (itint_1n[20], i_1r1d[20], gate917_0n, initialise);
  C2RI I951 (itint_1n[21], i_1r1d[21], gate917_0n, initialise);
  C2RI I952 (itint_1n[22], i_1r1d[22], gate917_0n, initialise);
  C2RI I953 (itint_1n[23], i_1r1d[23], gate917_0n, initialise);
  C2RI I954 (itint_1n[24], i_1r1d[24], gate917_0n, initialise);
  C2RI I955 (itint_1n[25], i_1r1d[25], gate917_0n, initialise);
  C2RI I956 (itint_1n[26], i_1r1d[26], gate917_0n, initialise);
  C2RI I957 (itint_1n[27], i_1r1d[27], gate917_0n, initialise);
  C2RI I958 (itint_1n[28], i_1r1d[28], gate917_0n, initialise);
  C2RI I959 (itint_1n[29], i_1r1d[29], gate917_0n, initialise);
  C2RI I960 (itint_1n[30], i_1r1d[30], gate917_0n, initialise);
  C2RI I961 (itint_1n[31], i_1r1d[31], gate917_0n, initialise);
  C2RI I962 (itint_1n[32], i_1r1d[32], gate917_0n, initialise);
  C2RI I963 (itint_1n[33], i_1r1d[33], gate917_0n, initialise);
  C2RI I964 (itint_1n[34], i_1r1d[34], gate917_0n, initialise);
  C2RI I965 (ifint_1n[0], i_1r0d[0], gate917_0n, initialise);
  C2RI I966 (ifint_1n[1], i_1r0d[1], gate917_0n, initialise);
  C2RI I967 (ifint_1n[2], i_1r0d[2], gate917_0n, initialise);
  C2RI I968 (ifint_1n[3], i_1r0d[3], gate917_0n, initialise);
  C2RI I969 (ifint_1n[4], i_1r0d[4], gate917_0n, initialise);
  C2RI I970 (ifint_1n[5], i_1r0d[5], gate917_0n, initialise);
  C2RI I971 (ifint_1n[6], i_1r0d[6], gate917_0n, initialise);
  C2RI I972 (ifint_1n[7], i_1r0d[7], gate917_0n, initialise);
  C2RI I973 (ifint_1n[8], i_1r0d[8], gate917_0n, initialise);
  C2RI I974 (ifint_1n[9], i_1r0d[9], gate917_0n, initialise);
  C2RI I975 (ifint_1n[10], i_1r0d[10], gate917_0n, initialise);
  C2RI I976 (ifint_1n[11], i_1r0d[11], gate917_0n, initialise);
  C2RI I977 (ifint_1n[12], i_1r0d[12], gate917_0n, initialise);
  C2RI I978 (ifint_1n[13], i_1r0d[13], gate917_0n, initialise);
  C2RI I979 (ifint_1n[14], i_1r0d[14], gate917_0n, initialise);
  C2RI I980 (ifint_1n[15], i_1r0d[15], gate917_0n, initialise);
  C2RI I981 (ifint_1n[16], i_1r0d[16], gate917_0n, initialise);
  C2RI I982 (ifint_1n[17], i_1r0d[17], gate917_0n, initialise);
  C2RI I983 (ifint_1n[18], i_1r0d[18], gate917_0n, initialise);
  C2RI I984 (ifint_1n[19], i_1r0d[19], gate917_0n, initialise);
  C2RI I985 (ifint_1n[20], i_1r0d[20], gate917_0n, initialise);
  C2RI I986 (ifint_1n[21], i_1r0d[21], gate917_0n, initialise);
  C2RI I987 (ifint_1n[22], i_1r0d[22], gate917_0n, initialise);
  C2RI I988 (ifint_1n[23], i_1r0d[23], gate917_0n, initialise);
  C2RI I989 (ifint_1n[24], i_1r0d[24], gate917_0n, initialise);
  C2RI I990 (ifint_1n[25], i_1r0d[25], gate917_0n, initialise);
  C2RI I991 (ifint_1n[26], i_1r0d[26], gate917_0n, initialise);
  C2RI I992 (ifint_1n[27], i_1r0d[27], gate917_0n, initialise);
  C2RI I993 (ifint_1n[28], i_1r0d[28], gate917_0n, initialise);
  C2RI I994 (ifint_1n[29], i_1r0d[29], gate917_0n, initialise);
  C2RI I995 (ifint_1n[30], i_1r0d[30], gate917_0n, initialise);
  C2RI I996 (ifint_1n[31], i_1r0d[31], gate917_0n, initialise);
  C2RI I997 (ifint_1n[32], i_1r0d[32], gate917_0n, initialise);
  C2RI I998 (ifint_1n[33], i_1r0d[33], gate917_0n, initialise);
  C2RI I999 (ifint_1n[34], i_1r0d[34], gate917_0n, initialise);
  C3 I1000 (internal_0n[144], complete914_0n[0], complete914_0n[1], complete914_0n[2]);
  C3 I1001 (internal_0n[145], complete914_0n[3], complete914_0n[4], complete914_0n[5]);
  C3 I1002 (internal_0n[146], complete914_0n[6], complete914_0n[7], complete914_0n[8]);
  C3 I1003 (internal_0n[147], complete914_0n[9], complete914_0n[10], complete914_0n[11]);
  C3 I1004 (internal_0n[148], complete914_0n[12], complete914_0n[13], complete914_0n[14]);
  C3 I1005 (internal_0n[149], complete914_0n[15], complete914_0n[16], complete914_0n[17]);
  C3 I1006 (internal_0n[150], complete914_0n[18], complete914_0n[19], complete914_0n[20]);
  C3 I1007 (internal_0n[151], complete914_0n[21], complete914_0n[22], complete914_0n[23]);
  C3 I1008 (internal_0n[152], complete914_0n[24], complete914_0n[25], complete914_0n[26]);
  C3 I1009 (internal_0n[153], complete914_0n[27], complete914_0n[28], complete914_0n[29]);
  C3 I1010 (internal_0n[154], complete914_0n[30], complete914_0n[31], complete914_0n[32]);
  C2 I1011 (internal_0n[155], complete914_0n[33], complete914_0n[34]);
  C3 I1012 (internal_0n[156], internal_0n[144], internal_0n[145], internal_0n[146]);
  C3 I1013 (internal_0n[157], internal_0n[147], internal_0n[148], internal_0n[149]);
  C3 I1014 (internal_0n[158], internal_0n[150], internal_0n[151], internal_0n[152]);
  C3 I1015 (internal_0n[159], internal_0n[153], internal_0n[154], internal_0n[155]);
  C2 I1016 (internal_0n[160], internal_0n[156], internal_0n[157]);
  C2 I1017 (internal_0n[161], internal_0n[158], internal_0n[159]);
  C2 I1018 (i_0a, internal_0n[160], internal_0n[161]);
  OR2 I1019 (complete914_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I1020 (complete914_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I1021 (complete914_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I1022 (complete914_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I1023 (complete914_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I1024 (complete914_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I1025 (complete914_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I1026 (complete914_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I1027 (complete914_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I1028 (complete914_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I1029 (complete914_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I1030 (complete914_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I1031 (complete914_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I1032 (complete914_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I1033 (complete914_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I1034 (complete914_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I1035 (complete914_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I1036 (complete914_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I1037 (complete914_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I1038 (complete914_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I1039 (complete914_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I1040 (complete914_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I1041 (complete914_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I1042 (complete914_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I1043 (complete914_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I1044 (complete914_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I1045 (complete914_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I1046 (complete914_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I1047 (complete914_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I1048 (complete914_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I1049 (complete914_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I1050 (complete914_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I1051 (complete914_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I1052 (complete914_0n[33], ifint_0n[33], itint_0n[33]);
  OR2 I1053 (complete914_0n[34], ifint_0n[34], itint_0n[34]);
  INV I1054 (gate913_0n, iaint_0n);
  C2RI I1055 (itint_0n[0], i_0r1d[0], gate913_0n, initialise);
  C2RI I1056 (itint_0n[1], i_0r1d[1], gate913_0n, initialise);
  C2RI I1057 (itint_0n[2], i_0r1d[2], gate913_0n, initialise);
  C2RI I1058 (itint_0n[3], i_0r1d[3], gate913_0n, initialise);
  C2RI I1059 (itint_0n[4], i_0r1d[4], gate913_0n, initialise);
  C2RI I1060 (itint_0n[5], i_0r1d[5], gate913_0n, initialise);
  C2RI I1061 (itint_0n[6], i_0r1d[6], gate913_0n, initialise);
  C2RI I1062 (itint_0n[7], i_0r1d[7], gate913_0n, initialise);
  C2RI I1063 (itint_0n[8], i_0r1d[8], gate913_0n, initialise);
  C2RI I1064 (itint_0n[9], i_0r1d[9], gate913_0n, initialise);
  C2RI I1065 (itint_0n[10], i_0r1d[10], gate913_0n, initialise);
  C2RI I1066 (itint_0n[11], i_0r1d[11], gate913_0n, initialise);
  C2RI I1067 (itint_0n[12], i_0r1d[12], gate913_0n, initialise);
  C2RI I1068 (itint_0n[13], i_0r1d[13], gate913_0n, initialise);
  C2RI I1069 (itint_0n[14], i_0r1d[14], gate913_0n, initialise);
  C2RI I1070 (itint_0n[15], i_0r1d[15], gate913_0n, initialise);
  C2RI I1071 (itint_0n[16], i_0r1d[16], gate913_0n, initialise);
  C2RI I1072 (itint_0n[17], i_0r1d[17], gate913_0n, initialise);
  C2RI I1073 (itint_0n[18], i_0r1d[18], gate913_0n, initialise);
  C2RI I1074 (itint_0n[19], i_0r1d[19], gate913_0n, initialise);
  C2RI I1075 (itint_0n[20], i_0r1d[20], gate913_0n, initialise);
  C2RI I1076 (itint_0n[21], i_0r1d[21], gate913_0n, initialise);
  C2RI I1077 (itint_0n[22], i_0r1d[22], gate913_0n, initialise);
  C2RI I1078 (itint_0n[23], i_0r1d[23], gate913_0n, initialise);
  C2RI I1079 (itint_0n[24], i_0r1d[24], gate913_0n, initialise);
  C2RI I1080 (itint_0n[25], i_0r1d[25], gate913_0n, initialise);
  C2RI I1081 (itint_0n[26], i_0r1d[26], gate913_0n, initialise);
  C2RI I1082 (itint_0n[27], i_0r1d[27], gate913_0n, initialise);
  C2RI I1083 (itint_0n[28], i_0r1d[28], gate913_0n, initialise);
  C2RI I1084 (itint_0n[29], i_0r1d[29], gate913_0n, initialise);
  C2RI I1085 (itint_0n[30], i_0r1d[30], gate913_0n, initialise);
  C2RI I1086 (itint_0n[31], i_0r1d[31], gate913_0n, initialise);
  C2RI I1087 (itint_0n[32], i_0r1d[32], gate913_0n, initialise);
  C2RI I1088 (itint_0n[33], i_0r1d[33], gate913_0n, initialise);
  C2RI I1089 (itint_0n[34], i_0r1d[34], gate913_0n, initialise);
  C2RI I1090 (ifint_0n[0], i_0r0d[0], gate913_0n, initialise);
  C2RI I1091 (ifint_0n[1], i_0r0d[1], gate913_0n, initialise);
  C2RI I1092 (ifint_0n[2], i_0r0d[2], gate913_0n, initialise);
  C2RI I1093 (ifint_0n[3], i_0r0d[3], gate913_0n, initialise);
  C2RI I1094 (ifint_0n[4], i_0r0d[4], gate913_0n, initialise);
  C2RI I1095 (ifint_0n[5], i_0r0d[5], gate913_0n, initialise);
  C2RI I1096 (ifint_0n[6], i_0r0d[6], gate913_0n, initialise);
  C2RI I1097 (ifint_0n[7], i_0r0d[7], gate913_0n, initialise);
  C2RI I1098 (ifint_0n[8], i_0r0d[8], gate913_0n, initialise);
  C2RI I1099 (ifint_0n[9], i_0r0d[9], gate913_0n, initialise);
  C2RI I1100 (ifint_0n[10], i_0r0d[10], gate913_0n, initialise);
  C2RI I1101 (ifint_0n[11], i_0r0d[11], gate913_0n, initialise);
  C2RI I1102 (ifint_0n[12], i_0r0d[12], gate913_0n, initialise);
  C2RI I1103 (ifint_0n[13], i_0r0d[13], gate913_0n, initialise);
  C2RI I1104 (ifint_0n[14], i_0r0d[14], gate913_0n, initialise);
  C2RI I1105 (ifint_0n[15], i_0r0d[15], gate913_0n, initialise);
  C2RI I1106 (ifint_0n[16], i_0r0d[16], gate913_0n, initialise);
  C2RI I1107 (ifint_0n[17], i_0r0d[17], gate913_0n, initialise);
  C2RI I1108 (ifint_0n[18], i_0r0d[18], gate913_0n, initialise);
  C2RI I1109 (ifint_0n[19], i_0r0d[19], gate913_0n, initialise);
  C2RI I1110 (ifint_0n[20], i_0r0d[20], gate913_0n, initialise);
  C2RI I1111 (ifint_0n[21], i_0r0d[21], gate913_0n, initialise);
  C2RI I1112 (ifint_0n[22], i_0r0d[22], gate913_0n, initialise);
  C2RI I1113 (ifint_0n[23], i_0r0d[23], gate913_0n, initialise);
  C2RI I1114 (ifint_0n[24], i_0r0d[24], gate913_0n, initialise);
  C2RI I1115 (ifint_0n[25], i_0r0d[25], gate913_0n, initialise);
  C2RI I1116 (ifint_0n[26], i_0r0d[26], gate913_0n, initialise);
  C2RI I1117 (ifint_0n[27], i_0r0d[27], gate913_0n, initialise);
  C2RI I1118 (ifint_0n[28], i_0r0d[28], gate913_0n, initialise);
  C2RI I1119 (ifint_0n[29], i_0r0d[29], gate913_0n, initialise);
  C2RI I1120 (ifint_0n[30], i_0r0d[30], gate913_0n, initialise);
  C2RI I1121 (ifint_0n[31], i_0r0d[31], gate913_0n, initialise);
  C2RI I1122 (ifint_0n[32], i_0r0d[32], gate913_0n, initialise);
  C2RI I1123 (ifint_0n[33], i_0r0d[33], gate913_0n, initialise);
  C2RI I1124 (ifint_0n[34], i_0r0d[34], gate913_0n, initialise);
  C3 I1125 (internal_0n[162], complete910_0n[0], complete910_0n[1], complete910_0n[2]);
  C3 I1126 (internal_0n[163], complete910_0n[3], complete910_0n[4], complete910_0n[5]);
  C3 I1127 (internal_0n[164], complete910_0n[6], complete910_0n[7], complete910_0n[8]);
  C3 I1128 (internal_0n[165], complete910_0n[9], complete910_0n[10], complete910_0n[11]);
  C3 I1129 (internal_0n[166], complete910_0n[12], complete910_0n[13], complete910_0n[14]);
  C3 I1130 (internal_0n[167], complete910_0n[15], complete910_0n[16], complete910_0n[17]);
  C3 I1131 (internal_0n[168], complete910_0n[18], complete910_0n[19], complete910_0n[20]);
  C3 I1132 (internal_0n[169], complete910_0n[21], complete910_0n[22], complete910_0n[23]);
  C3 I1133 (internal_0n[170], complete910_0n[24], complete910_0n[25], complete910_0n[26]);
  C3 I1134 (internal_0n[171], complete910_0n[27], complete910_0n[28], complete910_0n[29]);
  C3 I1135 (internal_0n[172], complete910_0n[30], complete910_0n[31], complete910_0n[32]);
  C2 I1136 (internal_0n[173], complete910_0n[33], complete910_0n[34]);
  C3 I1137 (internal_0n[174], internal_0n[162], internal_0n[163], internal_0n[164]);
  C3 I1138 (internal_0n[175], internal_0n[165], internal_0n[166], internal_0n[167]);
  C3 I1139 (internal_0n[176], internal_0n[168], internal_0n[169], internal_0n[170]);
  C3 I1140 (internal_0n[177], internal_0n[171], internal_0n[172], internal_0n[173]);
  C2 I1141 (internal_0n[178], internal_0n[174], internal_0n[175]);
  C2 I1142 (internal_0n[179], internal_0n[176], internal_0n[177]);
  C2 I1143 (oaint_0n, internal_0n[178], internal_0n[179]);
  OR2 I1144 (complete910_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I1145 (complete910_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I1146 (complete910_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I1147 (complete910_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I1148 (complete910_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I1149 (complete910_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I1150 (complete910_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I1151 (complete910_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I1152 (complete910_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I1153 (complete910_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I1154 (complete910_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I1155 (complete910_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I1156 (complete910_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I1157 (complete910_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I1158 (complete910_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I1159 (complete910_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I1160 (complete910_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I1161 (complete910_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I1162 (complete910_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I1163 (complete910_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I1164 (complete910_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I1165 (complete910_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I1166 (complete910_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I1167 (complete910_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I1168 (complete910_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I1169 (complete910_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I1170 (complete910_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I1171 (complete910_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I1172 (complete910_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I1173 (complete910_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I1174 (complete910_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I1175 (complete910_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I1176 (complete910_0n[32], o_0r0d[32], o_0r1d[32]);
  OR2 I1177 (complete910_0n[33], o_0r0d[33], o_0r1d[33]);
  OR2 I1178 (complete910_0n[34], o_0r0d[34], o_0r1d[34]);
  INV I1179 (gate909_0n, o_0a);
  C2RI I1180 (o_0r1d[0], otint_0n[0], gate909_0n, initialise);
  C2RI I1181 (o_0r1d[1], otint_0n[1], gate909_0n, initialise);
  C2RI I1182 (o_0r1d[2], otint_0n[2], gate909_0n, initialise);
  C2RI I1183 (o_0r1d[3], otint_0n[3], gate909_0n, initialise);
  C2RI I1184 (o_0r1d[4], otint_0n[4], gate909_0n, initialise);
  C2RI I1185 (o_0r1d[5], otint_0n[5], gate909_0n, initialise);
  C2RI I1186 (o_0r1d[6], otint_0n[6], gate909_0n, initialise);
  C2RI I1187 (o_0r1d[7], otint_0n[7], gate909_0n, initialise);
  C2RI I1188 (o_0r1d[8], otint_0n[8], gate909_0n, initialise);
  C2RI I1189 (o_0r1d[9], otint_0n[9], gate909_0n, initialise);
  C2RI I1190 (o_0r1d[10], otint_0n[10], gate909_0n, initialise);
  C2RI I1191 (o_0r1d[11], otint_0n[11], gate909_0n, initialise);
  C2RI I1192 (o_0r1d[12], otint_0n[12], gate909_0n, initialise);
  C2RI I1193 (o_0r1d[13], otint_0n[13], gate909_0n, initialise);
  C2RI I1194 (o_0r1d[14], otint_0n[14], gate909_0n, initialise);
  C2RI I1195 (o_0r1d[15], otint_0n[15], gate909_0n, initialise);
  C2RI I1196 (o_0r1d[16], otint_0n[16], gate909_0n, initialise);
  C2RI I1197 (o_0r1d[17], otint_0n[17], gate909_0n, initialise);
  C2RI I1198 (o_0r1d[18], otint_0n[18], gate909_0n, initialise);
  C2RI I1199 (o_0r1d[19], otint_0n[19], gate909_0n, initialise);
  C2RI I1200 (o_0r1d[20], otint_0n[20], gate909_0n, initialise);
  C2RI I1201 (o_0r1d[21], otint_0n[21], gate909_0n, initialise);
  C2RI I1202 (o_0r1d[22], otint_0n[22], gate909_0n, initialise);
  C2RI I1203 (o_0r1d[23], otint_0n[23], gate909_0n, initialise);
  C2RI I1204 (o_0r1d[24], otint_0n[24], gate909_0n, initialise);
  C2RI I1205 (o_0r1d[25], otint_0n[25], gate909_0n, initialise);
  C2RI I1206 (o_0r1d[26], otint_0n[26], gate909_0n, initialise);
  C2RI I1207 (o_0r1d[27], otint_0n[27], gate909_0n, initialise);
  C2RI I1208 (o_0r1d[28], otint_0n[28], gate909_0n, initialise);
  C2RI I1209 (o_0r1d[29], otint_0n[29], gate909_0n, initialise);
  C2RI I1210 (o_0r1d[30], otint_0n[30], gate909_0n, initialise);
  C2RI I1211 (o_0r1d[31], otint_0n[31], gate909_0n, initialise);
  C2RI I1212 (o_0r1d[32], otint_0n[32], gate909_0n, initialise);
  C2RI I1213 (o_0r1d[33], otint_0n[33], gate909_0n, initialise);
  C2RI I1214 (o_0r1d[34], otint_0n[34], gate909_0n, initialise);
  C2RI I1215 (o_0r0d[0], ofint_0n[0], gate909_0n, initialise);
  C2RI I1216 (o_0r0d[1], ofint_0n[1], gate909_0n, initialise);
  C2RI I1217 (o_0r0d[2], ofint_0n[2], gate909_0n, initialise);
  C2RI I1218 (o_0r0d[3], ofint_0n[3], gate909_0n, initialise);
  C2RI I1219 (o_0r0d[4], ofint_0n[4], gate909_0n, initialise);
  C2RI I1220 (o_0r0d[5], ofint_0n[5], gate909_0n, initialise);
  C2RI I1221 (o_0r0d[6], ofint_0n[6], gate909_0n, initialise);
  C2RI I1222 (o_0r0d[7], ofint_0n[7], gate909_0n, initialise);
  C2RI I1223 (o_0r0d[8], ofint_0n[8], gate909_0n, initialise);
  C2RI I1224 (o_0r0d[9], ofint_0n[9], gate909_0n, initialise);
  C2RI I1225 (o_0r0d[10], ofint_0n[10], gate909_0n, initialise);
  C2RI I1226 (o_0r0d[11], ofint_0n[11], gate909_0n, initialise);
  C2RI I1227 (o_0r0d[12], ofint_0n[12], gate909_0n, initialise);
  C2RI I1228 (o_0r0d[13], ofint_0n[13], gate909_0n, initialise);
  C2RI I1229 (o_0r0d[14], ofint_0n[14], gate909_0n, initialise);
  C2RI I1230 (o_0r0d[15], ofint_0n[15], gate909_0n, initialise);
  C2RI I1231 (o_0r0d[16], ofint_0n[16], gate909_0n, initialise);
  C2RI I1232 (o_0r0d[17], ofint_0n[17], gate909_0n, initialise);
  C2RI I1233 (o_0r0d[18], ofint_0n[18], gate909_0n, initialise);
  C2RI I1234 (o_0r0d[19], ofint_0n[19], gate909_0n, initialise);
  C2RI I1235 (o_0r0d[20], ofint_0n[20], gate909_0n, initialise);
  C2RI I1236 (o_0r0d[21], ofint_0n[21], gate909_0n, initialise);
  C2RI I1237 (o_0r0d[22], ofint_0n[22], gate909_0n, initialise);
  C2RI I1238 (o_0r0d[23], ofint_0n[23], gate909_0n, initialise);
  C2RI I1239 (o_0r0d[24], ofint_0n[24], gate909_0n, initialise);
  C2RI I1240 (o_0r0d[25], ofint_0n[25], gate909_0n, initialise);
  C2RI I1241 (o_0r0d[26], ofint_0n[26], gate909_0n, initialise);
  C2RI I1242 (o_0r0d[27], ofint_0n[27], gate909_0n, initialise);
  C2RI I1243 (o_0r0d[28], ofint_0n[28], gate909_0n, initialise);
  C2RI I1244 (o_0r0d[29], ofint_0n[29], gate909_0n, initialise);
  C2RI I1245 (o_0r0d[30], ofint_0n[30], gate909_0n, initialise);
  C2RI I1246 (o_0r0d[31], ofint_0n[31], gate909_0n, initialise);
  C2RI I1247 (o_0r0d[32], ofint_0n[32], gate909_0n, initialise);
  C2RI I1248 (o_0r0d[33], ofint_0n[33], gate909_0n, initialise);
  C2RI I1249 (o_0r0d[34], ofint_0n[34], gate909_0n, initialise);
  C2RI I1250 (iaint_0n, sel_0n[0], oaint_0n, initialise);
  C2RI I1251 (iaint_1n, sel_0n[1], oaint_0n, initialise);
  C2RI I1252 (iaint_2n, sel_0n[2], oaint_0n, initialise);
  C2RI I1253 (iaint_3n, sel_0n[3], oaint_0n, initialise);
  C2RI I1254 (iaint_4n, sel_0n[4], oaint_0n, initialise);
  C2RI I1255 (iaint_5n, sel_0n[5], oaint_0n, initialise);
  C2RI I1256 (iaint_6n, sel_0n[6], oaint_0n, initialise);
  C2RI I1257 (iaint_7n, sel_0n[7], oaint_0n, initialise);
  C2RI I1258 (iaint_8n, sel_0n[8], oaint_0n, initialise);
  assign gate_0n[0] = sel_0n[0];
  assign gate_0n[1] = sel_0n[1];
  assign gate_0n[2] = sel_0n[2];
  assign gate_0n[3] = sel_0n[3];
  assign gate_0n[4] = sel_0n[4];
  assign gate_0n[5] = sel_0n[5];
  assign gate_0n[6] = sel_0n[6];
  assign gate_0n[7] = sel_0n[7];
  assign gate_0n[8] = sel_0n[8];
  assign sel_0n[0] = selcomp_0n;
  assign sel_0n[1] = selcomp_1n;
  assign sel_0n[2] = selcomp_2n;
  assign sel_0n[3] = selcomp_3n;
  assign sel_0n[4] = selcomp_4n;
  assign sel_0n[5] = selcomp_5n;
  assign sel_0n[6] = selcomp_6n;
  assign sel_0n[7] = selcomp_7n;
  assign sel_0n[8] = selcomp_8n;
  C3 I1277 (internal_0n[180], complete906_0n[0], complete906_0n[1], complete906_0n[2]);
  C3 I1278 (internal_0n[181], complete906_0n[3], complete906_0n[4], complete906_0n[5]);
  C3 I1279 (internal_0n[182], complete906_0n[6], complete906_0n[7], complete906_0n[8]);
  C3 I1280 (internal_0n[183], complete906_0n[9], complete906_0n[10], complete906_0n[11]);
  C3 I1281 (internal_0n[184], complete906_0n[12], complete906_0n[13], complete906_0n[14]);
  C3 I1282 (internal_0n[185], complete906_0n[15], complete906_0n[16], complete906_0n[17]);
  C3 I1283 (internal_0n[186], complete906_0n[18], complete906_0n[19], complete906_0n[20]);
  C3 I1284 (internal_0n[187], complete906_0n[21], complete906_0n[22], complete906_0n[23]);
  C3 I1285 (internal_0n[188], complete906_0n[24], complete906_0n[25], complete906_0n[26]);
  C3 I1286 (internal_0n[189], complete906_0n[27], complete906_0n[28], complete906_0n[29]);
  C3 I1287 (internal_0n[190], complete906_0n[30], complete906_0n[31], complete906_0n[32]);
  C2 I1288 (internal_0n[191], complete906_0n[33], complete906_0n[34]);
  C3 I1289 (internal_0n[192], internal_0n[180], internal_0n[181], internal_0n[182]);
  C3 I1290 (internal_0n[193], internal_0n[183], internal_0n[184], internal_0n[185]);
  C3 I1291 (internal_0n[194], internal_0n[186], internal_0n[187], internal_0n[188]);
  C3 I1292 (internal_0n[195], internal_0n[189], internal_0n[190], internal_0n[191]);
  C2 I1293 (internal_0n[196], internal_0n[192], internal_0n[193]);
  C2 I1294 (internal_0n[197], internal_0n[194], internal_0n[195]);
  C2 I1295 (selcomp_8n, internal_0n[196], internal_0n[197]);
  OR2 I1296 (complete906_0n[0], ifint_8n[0], itint_8n[0]);
  OR2 I1297 (complete906_0n[1], ifint_8n[1], itint_8n[1]);
  OR2 I1298 (complete906_0n[2], ifint_8n[2], itint_8n[2]);
  OR2 I1299 (complete906_0n[3], ifint_8n[3], itint_8n[3]);
  OR2 I1300 (complete906_0n[4], ifint_8n[4], itint_8n[4]);
  OR2 I1301 (complete906_0n[5], ifint_8n[5], itint_8n[5]);
  OR2 I1302 (complete906_0n[6], ifint_8n[6], itint_8n[6]);
  OR2 I1303 (complete906_0n[7], ifint_8n[7], itint_8n[7]);
  OR2 I1304 (complete906_0n[8], ifint_8n[8], itint_8n[8]);
  OR2 I1305 (complete906_0n[9], ifint_8n[9], itint_8n[9]);
  OR2 I1306 (complete906_0n[10], ifint_8n[10], itint_8n[10]);
  OR2 I1307 (complete906_0n[11], ifint_8n[11], itint_8n[11]);
  OR2 I1308 (complete906_0n[12], ifint_8n[12], itint_8n[12]);
  OR2 I1309 (complete906_0n[13], ifint_8n[13], itint_8n[13]);
  OR2 I1310 (complete906_0n[14], ifint_8n[14], itint_8n[14]);
  OR2 I1311 (complete906_0n[15], ifint_8n[15], itint_8n[15]);
  OR2 I1312 (complete906_0n[16], ifint_8n[16], itint_8n[16]);
  OR2 I1313 (complete906_0n[17], ifint_8n[17], itint_8n[17]);
  OR2 I1314 (complete906_0n[18], ifint_8n[18], itint_8n[18]);
  OR2 I1315 (complete906_0n[19], ifint_8n[19], itint_8n[19]);
  OR2 I1316 (complete906_0n[20], ifint_8n[20], itint_8n[20]);
  OR2 I1317 (complete906_0n[21], ifint_8n[21], itint_8n[21]);
  OR2 I1318 (complete906_0n[22], ifint_8n[22], itint_8n[22]);
  OR2 I1319 (complete906_0n[23], ifint_8n[23], itint_8n[23]);
  OR2 I1320 (complete906_0n[24], ifint_8n[24], itint_8n[24]);
  OR2 I1321 (complete906_0n[25], ifint_8n[25], itint_8n[25]);
  OR2 I1322 (complete906_0n[26], ifint_8n[26], itint_8n[26]);
  OR2 I1323 (complete906_0n[27], ifint_8n[27], itint_8n[27]);
  OR2 I1324 (complete906_0n[28], ifint_8n[28], itint_8n[28]);
  OR2 I1325 (complete906_0n[29], ifint_8n[29], itint_8n[29]);
  OR2 I1326 (complete906_0n[30], ifint_8n[30], itint_8n[30]);
  OR2 I1327 (complete906_0n[31], ifint_8n[31], itint_8n[31]);
  OR2 I1328 (complete906_0n[32], ifint_8n[32], itint_8n[32]);
  OR2 I1329 (complete906_0n[33], ifint_8n[33], itint_8n[33]);
  OR2 I1330 (complete906_0n[34], ifint_8n[34], itint_8n[34]);
  C3 I1331 (internal_0n[198], complete905_0n[0], complete905_0n[1], complete905_0n[2]);
  C3 I1332 (internal_0n[199], complete905_0n[3], complete905_0n[4], complete905_0n[5]);
  C3 I1333 (internal_0n[200], complete905_0n[6], complete905_0n[7], complete905_0n[8]);
  C3 I1334 (internal_0n[201], complete905_0n[9], complete905_0n[10], complete905_0n[11]);
  C3 I1335 (internal_0n[202], complete905_0n[12], complete905_0n[13], complete905_0n[14]);
  C3 I1336 (internal_0n[203], complete905_0n[15], complete905_0n[16], complete905_0n[17]);
  C3 I1337 (internal_0n[204], complete905_0n[18], complete905_0n[19], complete905_0n[20]);
  C3 I1338 (internal_0n[205], complete905_0n[21], complete905_0n[22], complete905_0n[23]);
  C3 I1339 (internal_0n[206], complete905_0n[24], complete905_0n[25], complete905_0n[26]);
  C3 I1340 (internal_0n[207], complete905_0n[27], complete905_0n[28], complete905_0n[29]);
  C3 I1341 (internal_0n[208], complete905_0n[30], complete905_0n[31], complete905_0n[32]);
  C2 I1342 (internal_0n[209], complete905_0n[33], complete905_0n[34]);
  C3 I1343 (internal_0n[210], internal_0n[198], internal_0n[199], internal_0n[200]);
  C3 I1344 (internal_0n[211], internal_0n[201], internal_0n[202], internal_0n[203]);
  C3 I1345 (internal_0n[212], internal_0n[204], internal_0n[205], internal_0n[206]);
  C3 I1346 (internal_0n[213], internal_0n[207], internal_0n[208], internal_0n[209]);
  C2 I1347 (internal_0n[214], internal_0n[210], internal_0n[211]);
  C2 I1348 (internal_0n[215], internal_0n[212], internal_0n[213]);
  C2 I1349 (selcomp_7n, internal_0n[214], internal_0n[215]);
  OR2 I1350 (complete905_0n[0], ifint_7n[0], itint_7n[0]);
  OR2 I1351 (complete905_0n[1], ifint_7n[1], itint_7n[1]);
  OR2 I1352 (complete905_0n[2], ifint_7n[2], itint_7n[2]);
  OR2 I1353 (complete905_0n[3], ifint_7n[3], itint_7n[3]);
  OR2 I1354 (complete905_0n[4], ifint_7n[4], itint_7n[4]);
  OR2 I1355 (complete905_0n[5], ifint_7n[5], itint_7n[5]);
  OR2 I1356 (complete905_0n[6], ifint_7n[6], itint_7n[6]);
  OR2 I1357 (complete905_0n[7], ifint_7n[7], itint_7n[7]);
  OR2 I1358 (complete905_0n[8], ifint_7n[8], itint_7n[8]);
  OR2 I1359 (complete905_0n[9], ifint_7n[9], itint_7n[9]);
  OR2 I1360 (complete905_0n[10], ifint_7n[10], itint_7n[10]);
  OR2 I1361 (complete905_0n[11], ifint_7n[11], itint_7n[11]);
  OR2 I1362 (complete905_0n[12], ifint_7n[12], itint_7n[12]);
  OR2 I1363 (complete905_0n[13], ifint_7n[13], itint_7n[13]);
  OR2 I1364 (complete905_0n[14], ifint_7n[14], itint_7n[14]);
  OR2 I1365 (complete905_0n[15], ifint_7n[15], itint_7n[15]);
  OR2 I1366 (complete905_0n[16], ifint_7n[16], itint_7n[16]);
  OR2 I1367 (complete905_0n[17], ifint_7n[17], itint_7n[17]);
  OR2 I1368 (complete905_0n[18], ifint_7n[18], itint_7n[18]);
  OR2 I1369 (complete905_0n[19], ifint_7n[19], itint_7n[19]);
  OR2 I1370 (complete905_0n[20], ifint_7n[20], itint_7n[20]);
  OR2 I1371 (complete905_0n[21], ifint_7n[21], itint_7n[21]);
  OR2 I1372 (complete905_0n[22], ifint_7n[22], itint_7n[22]);
  OR2 I1373 (complete905_0n[23], ifint_7n[23], itint_7n[23]);
  OR2 I1374 (complete905_0n[24], ifint_7n[24], itint_7n[24]);
  OR2 I1375 (complete905_0n[25], ifint_7n[25], itint_7n[25]);
  OR2 I1376 (complete905_0n[26], ifint_7n[26], itint_7n[26]);
  OR2 I1377 (complete905_0n[27], ifint_7n[27], itint_7n[27]);
  OR2 I1378 (complete905_0n[28], ifint_7n[28], itint_7n[28]);
  OR2 I1379 (complete905_0n[29], ifint_7n[29], itint_7n[29]);
  OR2 I1380 (complete905_0n[30], ifint_7n[30], itint_7n[30]);
  OR2 I1381 (complete905_0n[31], ifint_7n[31], itint_7n[31]);
  OR2 I1382 (complete905_0n[32], ifint_7n[32], itint_7n[32]);
  OR2 I1383 (complete905_0n[33], ifint_7n[33], itint_7n[33]);
  OR2 I1384 (complete905_0n[34], ifint_7n[34], itint_7n[34]);
  C3 I1385 (internal_0n[216], complete904_0n[0], complete904_0n[1], complete904_0n[2]);
  C3 I1386 (internal_0n[217], complete904_0n[3], complete904_0n[4], complete904_0n[5]);
  C3 I1387 (internal_0n[218], complete904_0n[6], complete904_0n[7], complete904_0n[8]);
  C3 I1388 (internal_0n[219], complete904_0n[9], complete904_0n[10], complete904_0n[11]);
  C3 I1389 (internal_0n[220], complete904_0n[12], complete904_0n[13], complete904_0n[14]);
  C3 I1390 (internal_0n[221], complete904_0n[15], complete904_0n[16], complete904_0n[17]);
  C3 I1391 (internal_0n[222], complete904_0n[18], complete904_0n[19], complete904_0n[20]);
  C3 I1392 (internal_0n[223], complete904_0n[21], complete904_0n[22], complete904_0n[23]);
  C3 I1393 (internal_0n[224], complete904_0n[24], complete904_0n[25], complete904_0n[26]);
  C3 I1394 (internal_0n[225], complete904_0n[27], complete904_0n[28], complete904_0n[29]);
  C3 I1395 (internal_0n[226], complete904_0n[30], complete904_0n[31], complete904_0n[32]);
  C2 I1396 (internal_0n[227], complete904_0n[33], complete904_0n[34]);
  C3 I1397 (internal_0n[228], internal_0n[216], internal_0n[217], internal_0n[218]);
  C3 I1398 (internal_0n[229], internal_0n[219], internal_0n[220], internal_0n[221]);
  C3 I1399 (internal_0n[230], internal_0n[222], internal_0n[223], internal_0n[224]);
  C3 I1400 (internal_0n[231], internal_0n[225], internal_0n[226], internal_0n[227]);
  C2 I1401 (internal_0n[232], internal_0n[228], internal_0n[229]);
  C2 I1402 (internal_0n[233], internal_0n[230], internal_0n[231]);
  C2 I1403 (selcomp_6n, internal_0n[232], internal_0n[233]);
  OR2 I1404 (complete904_0n[0], ifint_6n[0], itint_6n[0]);
  OR2 I1405 (complete904_0n[1], ifint_6n[1], itint_6n[1]);
  OR2 I1406 (complete904_0n[2], ifint_6n[2], itint_6n[2]);
  OR2 I1407 (complete904_0n[3], ifint_6n[3], itint_6n[3]);
  OR2 I1408 (complete904_0n[4], ifint_6n[4], itint_6n[4]);
  OR2 I1409 (complete904_0n[5], ifint_6n[5], itint_6n[5]);
  OR2 I1410 (complete904_0n[6], ifint_6n[6], itint_6n[6]);
  OR2 I1411 (complete904_0n[7], ifint_6n[7], itint_6n[7]);
  OR2 I1412 (complete904_0n[8], ifint_6n[8], itint_6n[8]);
  OR2 I1413 (complete904_0n[9], ifint_6n[9], itint_6n[9]);
  OR2 I1414 (complete904_0n[10], ifint_6n[10], itint_6n[10]);
  OR2 I1415 (complete904_0n[11], ifint_6n[11], itint_6n[11]);
  OR2 I1416 (complete904_0n[12], ifint_6n[12], itint_6n[12]);
  OR2 I1417 (complete904_0n[13], ifint_6n[13], itint_6n[13]);
  OR2 I1418 (complete904_0n[14], ifint_6n[14], itint_6n[14]);
  OR2 I1419 (complete904_0n[15], ifint_6n[15], itint_6n[15]);
  OR2 I1420 (complete904_0n[16], ifint_6n[16], itint_6n[16]);
  OR2 I1421 (complete904_0n[17], ifint_6n[17], itint_6n[17]);
  OR2 I1422 (complete904_0n[18], ifint_6n[18], itint_6n[18]);
  OR2 I1423 (complete904_0n[19], ifint_6n[19], itint_6n[19]);
  OR2 I1424 (complete904_0n[20], ifint_6n[20], itint_6n[20]);
  OR2 I1425 (complete904_0n[21], ifint_6n[21], itint_6n[21]);
  OR2 I1426 (complete904_0n[22], ifint_6n[22], itint_6n[22]);
  OR2 I1427 (complete904_0n[23], ifint_6n[23], itint_6n[23]);
  OR2 I1428 (complete904_0n[24], ifint_6n[24], itint_6n[24]);
  OR2 I1429 (complete904_0n[25], ifint_6n[25], itint_6n[25]);
  OR2 I1430 (complete904_0n[26], ifint_6n[26], itint_6n[26]);
  OR2 I1431 (complete904_0n[27], ifint_6n[27], itint_6n[27]);
  OR2 I1432 (complete904_0n[28], ifint_6n[28], itint_6n[28]);
  OR2 I1433 (complete904_0n[29], ifint_6n[29], itint_6n[29]);
  OR2 I1434 (complete904_0n[30], ifint_6n[30], itint_6n[30]);
  OR2 I1435 (complete904_0n[31], ifint_6n[31], itint_6n[31]);
  OR2 I1436 (complete904_0n[32], ifint_6n[32], itint_6n[32]);
  OR2 I1437 (complete904_0n[33], ifint_6n[33], itint_6n[33]);
  OR2 I1438 (complete904_0n[34], ifint_6n[34], itint_6n[34]);
  C3 I1439 (internal_0n[234], complete903_0n[0], complete903_0n[1], complete903_0n[2]);
  C3 I1440 (internal_0n[235], complete903_0n[3], complete903_0n[4], complete903_0n[5]);
  C3 I1441 (internal_0n[236], complete903_0n[6], complete903_0n[7], complete903_0n[8]);
  C3 I1442 (internal_0n[237], complete903_0n[9], complete903_0n[10], complete903_0n[11]);
  C3 I1443 (internal_0n[238], complete903_0n[12], complete903_0n[13], complete903_0n[14]);
  C3 I1444 (internal_0n[239], complete903_0n[15], complete903_0n[16], complete903_0n[17]);
  C3 I1445 (internal_0n[240], complete903_0n[18], complete903_0n[19], complete903_0n[20]);
  C3 I1446 (internal_0n[241], complete903_0n[21], complete903_0n[22], complete903_0n[23]);
  C3 I1447 (internal_0n[242], complete903_0n[24], complete903_0n[25], complete903_0n[26]);
  C3 I1448 (internal_0n[243], complete903_0n[27], complete903_0n[28], complete903_0n[29]);
  C3 I1449 (internal_0n[244], complete903_0n[30], complete903_0n[31], complete903_0n[32]);
  C2 I1450 (internal_0n[245], complete903_0n[33], complete903_0n[34]);
  C3 I1451 (internal_0n[246], internal_0n[234], internal_0n[235], internal_0n[236]);
  C3 I1452 (internal_0n[247], internal_0n[237], internal_0n[238], internal_0n[239]);
  C3 I1453 (internal_0n[248], internal_0n[240], internal_0n[241], internal_0n[242]);
  C3 I1454 (internal_0n[249], internal_0n[243], internal_0n[244], internal_0n[245]);
  C2 I1455 (internal_0n[250], internal_0n[246], internal_0n[247]);
  C2 I1456 (internal_0n[251], internal_0n[248], internal_0n[249]);
  C2 I1457 (selcomp_5n, internal_0n[250], internal_0n[251]);
  OR2 I1458 (complete903_0n[0], ifint_5n[0], itint_5n[0]);
  OR2 I1459 (complete903_0n[1], ifint_5n[1], itint_5n[1]);
  OR2 I1460 (complete903_0n[2], ifint_5n[2], itint_5n[2]);
  OR2 I1461 (complete903_0n[3], ifint_5n[3], itint_5n[3]);
  OR2 I1462 (complete903_0n[4], ifint_5n[4], itint_5n[4]);
  OR2 I1463 (complete903_0n[5], ifint_5n[5], itint_5n[5]);
  OR2 I1464 (complete903_0n[6], ifint_5n[6], itint_5n[6]);
  OR2 I1465 (complete903_0n[7], ifint_5n[7], itint_5n[7]);
  OR2 I1466 (complete903_0n[8], ifint_5n[8], itint_5n[8]);
  OR2 I1467 (complete903_0n[9], ifint_5n[9], itint_5n[9]);
  OR2 I1468 (complete903_0n[10], ifint_5n[10], itint_5n[10]);
  OR2 I1469 (complete903_0n[11], ifint_5n[11], itint_5n[11]);
  OR2 I1470 (complete903_0n[12], ifint_5n[12], itint_5n[12]);
  OR2 I1471 (complete903_0n[13], ifint_5n[13], itint_5n[13]);
  OR2 I1472 (complete903_0n[14], ifint_5n[14], itint_5n[14]);
  OR2 I1473 (complete903_0n[15], ifint_5n[15], itint_5n[15]);
  OR2 I1474 (complete903_0n[16], ifint_5n[16], itint_5n[16]);
  OR2 I1475 (complete903_0n[17], ifint_5n[17], itint_5n[17]);
  OR2 I1476 (complete903_0n[18], ifint_5n[18], itint_5n[18]);
  OR2 I1477 (complete903_0n[19], ifint_5n[19], itint_5n[19]);
  OR2 I1478 (complete903_0n[20], ifint_5n[20], itint_5n[20]);
  OR2 I1479 (complete903_0n[21], ifint_5n[21], itint_5n[21]);
  OR2 I1480 (complete903_0n[22], ifint_5n[22], itint_5n[22]);
  OR2 I1481 (complete903_0n[23], ifint_5n[23], itint_5n[23]);
  OR2 I1482 (complete903_0n[24], ifint_5n[24], itint_5n[24]);
  OR2 I1483 (complete903_0n[25], ifint_5n[25], itint_5n[25]);
  OR2 I1484 (complete903_0n[26], ifint_5n[26], itint_5n[26]);
  OR2 I1485 (complete903_0n[27], ifint_5n[27], itint_5n[27]);
  OR2 I1486 (complete903_0n[28], ifint_5n[28], itint_5n[28]);
  OR2 I1487 (complete903_0n[29], ifint_5n[29], itint_5n[29]);
  OR2 I1488 (complete903_0n[30], ifint_5n[30], itint_5n[30]);
  OR2 I1489 (complete903_0n[31], ifint_5n[31], itint_5n[31]);
  OR2 I1490 (complete903_0n[32], ifint_5n[32], itint_5n[32]);
  OR2 I1491 (complete903_0n[33], ifint_5n[33], itint_5n[33]);
  OR2 I1492 (complete903_0n[34], ifint_5n[34], itint_5n[34]);
  C3 I1493 (internal_0n[252], complete902_0n[0], complete902_0n[1], complete902_0n[2]);
  C3 I1494 (internal_0n[253], complete902_0n[3], complete902_0n[4], complete902_0n[5]);
  C3 I1495 (internal_0n[254], complete902_0n[6], complete902_0n[7], complete902_0n[8]);
  C3 I1496 (internal_0n[255], complete902_0n[9], complete902_0n[10], complete902_0n[11]);
  C3 I1497 (internal_0n[256], complete902_0n[12], complete902_0n[13], complete902_0n[14]);
  C3 I1498 (internal_0n[257], complete902_0n[15], complete902_0n[16], complete902_0n[17]);
  C3 I1499 (internal_0n[258], complete902_0n[18], complete902_0n[19], complete902_0n[20]);
  C3 I1500 (internal_0n[259], complete902_0n[21], complete902_0n[22], complete902_0n[23]);
  C3 I1501 (internal_0n[260], complete902_0n[24], complete902_0n[25], complete902_0n[26]);
  C3 I1502 (internal_0n[261], complete902_0n[27], complete902_0n[28], complete902_0n[29]);
  C3 I1503 (internal_0n[262], complete902_0n[30], complete902_0n[31], complete902_0n[32]);
  C2 I1504 (internal_0n[263], complete902_0n[33], complete902_0n[34]);
  C3 I1505 (internal_0n[264], internal_0n[252], internal_0n[253], internal_0n[254]);
  C3 I1506 (internal_0n[265], internal_0n[255], internal_0n[256], internal_0n[257]);
  C3 I1507 (internal_0n[266], internal_0n[258], internal_0n[259], internal_0n[260]);
  C3 I1508 (internal_0n[267], internal_0n[261], internal_0n[262], internal_0n[263]);
  C2 I1509 (internal_0n[268], internal_0n[264], internal_0n[265]);
  C2 I1510 (internal_0n[269], internal_0n[266], internal_0n[267]);
  C2 I1511 (selcomp_4n, internal_0n[268], internal_0n[269]);
  OR2 I1512 (complete902_0n[0], ifint_4n[0], itint_4n[0]);
  OR2 I1513 (complete902_0n[1], ifint_4n[1], itint_4n[1]);
  OR2 I1514 (complete902_0n[2], ifint_4n[2], itint_4n[2]);
  OR2 I1515 (complete902_0n[3], ifint_4n[3], itint_4n[3]);
  OR2 I1516 (complete902_0n[4], ifint_4n[4], itint_4n[4]);
  OR2 I1517 (complete902_0n[5], ifint_4n[5], itint_4n[5]);
  OR2 I1518 (complete902_0n[6], ifint_4n[6], itint_4n[6]);
  OR2 I1519 (complete902_0n[7], ifint_4n[7], itint_4n[7]);
  OR2 I1520 (complete902_0n[8], ifint_4n[8], itint_4n[8]);
  OR2 I1521 (complete902_0n[9], ifint_4n[9], itint_4n[9]);
  OR2 I1522 (complete902_0n[10], ifint_4n[10], itint_4n[10]);
  OR2 I1523 (complete902_0n[11], ifint_4n[11], itint_4n[11]);
  OR2 I1524 (complete902_0n[12], ifint_4n[12], itint_4n[12]);
  OR2 I1525 (complete902_0n[13], ifint_4n[13], itint_4n[13]);
  OR2 I1526 (complete902_0n[14], ifint_4n[14], itint_4n[14]);
  OR2 I1527 (complete902_0n[15], ifint_4n[15], itint_4n[15]);
  OR2 I1528 (complete902_0n[16], ifint_4n[16], itint_4n[16]);
  OR2 I1529 (complete902_0n[17], ifint_4n[17], itint_4n[17]);
  OR2 I1530 (complete902_0n[18], ifint_4n[18], itint_4n[18]);
  OR2 I1531 (complete902_0n[19], ifint_4n[19], itint_4n[19]);
  OR2 I1532 (complete902_0n[20], ifint_4n[20], itint_4n[20]);
  OR2 I1533 (complete902_0n[21], ifint_4n[21], itint_4n[21]);
  OR2 I1534 (complete902_0n[22], ifint_4n[22], itint_4n[22]);
  OR2 I1535 (complete902_0n[23], ifint_4n[23], itint_4n[23]);
  OR2 I1536 (complete902_0n[24], ifint_4n[24], itint_4n[24]);
  OR2 I1537 (complete902_0n[25], ifint_4n[25], itint_4n[25]);
  OR2 I1538 (complete902_0n[26], ifint_4n[26], itint_4n[26]);
  OR2 I1539 (complete902_0n[27], ifint_4n[27], itint_4n[27]);
  OR2 I1540 (complete902_0n[28], ifint_4n[28], itint_4n[28]);
  OR2 I1541 (complete902_0n[29], ifint_4n[29], itint_4n[29]);
  OR2 I1542 (complete902_0n[30], ifint_4n[30], itint_4n[30]);
  OR2 I1543 (complete902_0n[31], ifint_4n[31], itint_4n[31]);
  OR2 I1544 (complete902_0n[32], ifint_4n[32], itint_4n[32]);
  OR2 I1545 (complete902_0n[33], ifint_4n[33], itint_4n[33]);
  OR2 I1546 (complete902_0n[34], ifint_4n[34], itint_4n[34]);
  C3 I1547 (internal_0n[270], complete901_0n[0], complete901_0n[1], complete901_0n[2]);
  C3 I1548 (internal_0n[271], complete901_0n[3], complete901_0n[4], complete901_0n[5]);
  C3 I1549 (internal_0n[272], complete901_0n[6], complete901_0n[7], complete901_0n[8]);
  C3 I1550 (internal_0n[273], complete901_0n[9], complete901_0n[10], complete901_0n[11]);
  C3 I1551 (internal_0n[274], complete901_0n[12], complete901_0n[13], complete901_0n[14]);
  C3 I1552 (internal_0n[275], complete901_0n[15], complete901_0n[16], complete901_0n[17]);
  C3 I1553 (internal_0n[276], complete901_0n[18], complete901_0n[19], complete901_0n[20]);
  C3 I1554 (internal_0n[277], complete901_0n[21], complete901_0n[22], complete901_0n[23]);
  C3 I1555 (internal_0n[278], complete901_0n[24], complete901_0n[25], complete901_0n[26]);
  C3 I1556 (internal_0n[279], complete901_0n[27], complete901_0n[28], complete901_0n[29]);
  C3 I1557 (internal_0n[280], complete901_0n[30], complete901_0n[31], complete901_0n[32]);
  C2 I1558 (internal_0n[281], complete901_0n[33], complete901_0n[34]);
  C3 I1559 (internal_0n[282], internal_0n[270], internal_0n[271], internal_0n[272]);
  C3 I1560 (internal_0n[283], internal_0n[273], internal_0n[274], internal_0n[275]);
  C3 I1561 (internal_0n[284], internal_0n[276], internal_0n[277], internal_0n[278]);
  C3 I1562 (internal_0n[285], internal_0n[279], internal_0n[280], internal_0n[281]);
  C2 I1563 (internal_0n[286], internal_0n[282], internal_0n[283]);
  C2 I1564 (internal_0n[287], internal_0n[284], internal_0n[285]);
  C2 I1565 (selcomp_3n, internal_0n[286], internal_0n[287]);
  OR2 I1566 (complete901_0n[0], ifint_3n[0], itint_3n[0]);
  OR2 I1567 (complete901_0n[1], ifint_3n[1], itint_3n[1]);
  OR2 I1568 (complete901_0n[2], ifint_3n[2], itint_3n[2]);
  OR2 I1569 (complete901_0n[3], ifint_3n[3], itint_3n[3]);
  OR2 I1570 (complete901_0n[4], ifint_3n[4], itint_3n[4]);
  OR2 I1571 (complete901_0n[5], ifint_3n[5], itint_3n[5]);
  OR2 I1572 (complete901_0n[6], ifint_3n[6], itint_3n[6]);
  OR2 I1573 (complete901_0n[7], ifint_3n[7], itint_3n[7]);
  OR2 I1574 (complete901_0n[8], ifint_3n[8], itint_3n[8]);
  OR2 I1575 (complete901_0n[9], ifint_3n[9], itint_3n[9]);
  OR2 I1576 (complete901_0n[10], ifint_3n[10], itint_3n[10]);
  OR2 I1577 (complete901_0n[11], ifint_3n[11], itint_3n[11]);
  OR2 I1578 (complete901_0n[12], ifint_3n[12], itint_3n[12]);
  OR2 I1579 (complete901_0n[13], ifint_3n[13], itint_3n[13]);
  OR2 I1580 (complete901_0n[14], ifint_3n[14], itint_3n[14]);
  OR2 I1581 (complete901_0n[15], ifint_3n[15], itint_3n[15]);
  OR2 I1582 (complete901_0n[16], ifint_3n[16], itint_3n[16]);
  OR2 I1583 (complete901_0n[17], ifint_3n[17], itint_3n[17]);
  OR2 I1584 (complete901_0n[18], ifint_3n[18], itint_3n[18]);
  OR2 I1585 (complete901_0n[19], ifint_3n[19], itint_3n[19]);
  OR2 I1586 (complete901_0n[20], ifint_3n[20], itint_3n[20]);
  OR2 I1587 (complete901_0n[21], ifint_3n[21], itint_3n[21]);
  OR2 I1588 (complete901_0n[22], ifint_3n[22], itint_3n[22]);
  OR2 I1589 (complete901_0n[23], ifint_3n[23], itint_3n[23]);
  OR2 I1590 (complete901_0n[24], ifint_3n[24], itint_3n[24]);
  OR2 I1591 (complete901_0n[25], ifint_3n[25], itint_3n[25]);
  OR2 I1592 (complete901_0n[26], ifint_3n[26], itint_3n[26]);
  OR2 I1593 (complete901_0n[27], ifint_3n[27], itint_3n[27]);
  OR2 I1594 (complete901_0n[28], ifint_3n[28], itint_3n[28]);
  OR2 I1595 (complete901_0n[29], ifint_3n[29], itint_3n[29]);
  OR2 I1596 (complete901_0n[30], ifint_3n[30], itint_3n[30]);
  OR2 I1597 (complete901_0n[31], ifint_3n[31], itint_3n[31]);
  OR2 I1598 (complete901_0n[32], ifint_3n[32], itint_3n[32]);
  OR2 I1599 (complete901_0n[33], ifint_3n[33], itint_3n[33]);
  OR2 I1600 (complete901_0n[34], ifint_3n[34], itint_3n[34]);
  C3 I1601 (internal_0n[288], complete900_0n[0], complete900_0n[1], complete900_0n[2]);
  C3 I1602 (internal_0n[289], complete900_0n[3], complete900_0n[4], complete900_0n[5]);
  C3 I1603 (internal_0n[290], complete900_0n[6], complete900_0n[7], complete900_0n[8]);
  C3 I1604 (internal_0n[291], complete900_0n[9], complete900_0n[10], complete900_0n[11]);
  C3 I1605 (internal_0n[292], complete900_0n[12], complete900_0n[13], complete900_0n[14]);
  C3 I1606 (internal_0n[293], complete900_0n[15], complete900_0n[16], complete900_0n[17]);
  C3 I1607 (internal_0n[294], complete900_0n[18], complete900_0n[19], complete900_0n[20]);
  C3 I1608 (internal_0n[295], complete900_0n[21], complete900_0n[22], complete900_0n[23]);
  C3 I1609 (internal_0n[296], complete900_0n[24], complete900_0n[25], complete900_0n[26]);
  C3 I1610 (internal_0n[297], complete900_0n[27], complete900_0n[28], complete900_0n[29]);
  C3 I1611 (internal_0n[298], complete900_0n[30], complete900_0n[31], complete900_0n[32]);
  C2 I1612 (internal_0n[299], complete900_0n[33], complete900_0n[34]);
  C3 I1613 (internal_0n[300], internal_0n[288], internal_0n[289], internal_0n[290]);
  C3 I1614 (internal_0n[301], internal_0n[291], internal_0n[292], internal_0n[293]);
  C3 I1615 (internal_0n[302], internal_0n[294], internal_0n[295], internal_0n[296]);
  C3 I1616 (internal_0n[303], internal_0n[297], internal_0n[298], internal_0n[299]);
  C2 I1617 (internal_0n[304], internal_0n[300], internal_0n[301]);
  C2 I1618 (internal_0n[305], internal_0n[302], internal_0n[303]);
  C2 I1619 (selcomp_2n, internal_0n[304], internal_0n[305]);
  OR2 I1620 (complete900_0n[0], ifint_2n[0], itint_2n[0]);
  OR2 I1621 (complete900_0n[1], ifint_2n[1], itint_2n[1]);
  OR2 I1622 (complete900_0n[2], ifint_2n[2], itint_2n[2]);
  OR2 I1623 (complete900_0n[3], ifint_2n[3], itint_2n[3]);
  OR2 I1624 (complete900_0n[4], ifint_2n[4], itint_2n[4]);
  OR2 I1625 (complete900_0n[5], ifint_2n[5], itint_2n[5]);
  OR2 I1626 (complete900_0n[6], ifint_2n[6], itint_2n[6]);
  OR2 I1627 (complete900_0n[7], ifint_2n[7], itint_2n[7]);
  OR2 I1628 (complete900_0n[8], ifint_2n[8], itint_2n[8]);
  OR2 I1629 (complete900_0n[9], ifint_2n[9], itint_2n[9]);
  OR2 I1630 (complete900_0n[10], ifint_2n[10], itint_2n[10]);
  OR2 I1631 (complete900_0n[11], ifint_2n[11], itint_2n[11]);
  OR2 I1632 (complete900_0n[12], ifint_2n[12], itint_2n[12]);
  OR2 I1633 (complete900_0n[13], ifint_2n[13], itint_2n[13]);
  OR2 I1634 (complete900_0n[14], ifint_2n[14], itint_2n[14]);
  OR2 I1635 (complete900_0n[15], ifint_2n[15], itint_2n[15]);
  OR2 I1636 (complete900_0n[16], ifint_2n[16], itint_2n[16]);
  OR2 I1637 (complete900_0n[17], ifint_2n[17], itint_2n[17]);
  OR2 I1638 (complete900_0n[18], ifint_2n[18], itint_2n[18]);
  OR2 I1639 (complete900_0n[19], ifint_2n[19], itint_2n[19]);
  OR2 I1640 (complete900_0n[20], ifint_2n[20], itint_2n[20]);
  OR2 I1641 (complete900_0n[21], ifint_2n[21], itint_2n[21]);
  OR2 I1642 (complete900_0n[22], ifint_2n[22], itint_2n[22]);
  OR2 I1643 (complete900_0n[23], ifint_2n[23], itint_2n[23]);
  OR2 I1644 (complete900_0n[24], ifint_2n[24], itint_2n[24]);
  OR2 I1645 (complete900_0n[25], ifint_2n[25], itint_2n[25]);
  OR2 I1646 (complete900_0n[26], ifint_2n[26], itint_2n[26]);
  OR2 I1647 (complete900_0n[27], ifint_2n[27], itint_2n[27]);
  OR2 I1648 (complete900_0n[28], ifint_2n[28], itint_2n[28]);
  OR2 I1649 (complete900_0n[29], ifint_2n[29], itint_2n[29]);
  OR2 I1650 (complete900_0n[30], ifint_2n[30], itint_2n[30]);
  OR2 I1651 (complete900_0n[31], ifint_2n[31], itint_2n[31]);
  OR2 I1652 (complete900_0n[32], ifint_2n[32], itint_2n[32]);
  OR2 I1653 (complete900_0n[33], ifint_2n[33], itint_2n[33]);
  OR2 I1654 (complete900_0n[34], ifint_2n[34], itint_2n[34]);
  C3 I1655 (internal_0n[306], complete899_0n[0], complete899_0n[1], complete899_0n[2]);
  C3 I1656 (internal_0n[307], complete899_0n[3], complete899_0n[4], complete899_0n[5]);
  C3 I1657 (internal_0n[308], complete899_0n[6], complete899_0n[7], complete899_0n[8]);
  C3 I1658 (internal_0n[309], complete899_0n[9], complete899_0n[10], complete899_0n[11]);
  C3 I1659 (internal_0n[310], complete899_0n[12], complete899_0n[13], complete899_0n[14]);
  C3 I1660 (internal_0n[311], complete899_0n[15], complete899_0n[16], complete899_0n[17]);
  C3 I1661 (internal_0n[312], complete899_0n[18], complete899_0n[19], complete899_0n[20]);
  C3 I1662 (internal_0n[313], complete899_0n[21], complete899_0n[22], complete899_0n[23]);
  C3 I1663 (internal_0n[314], complete899_0n[24], complete899_0n[25], complete899_0n[26]);
  C3 I1664 (internal_0n[315], complete899_0n[27], complete899_0n[28], complete899_0n[29]);
  C3 I1665 (internal_0n[316], complete899_0n[30], complete899_0n[31], complete899_0n[32]);
  C2 I1666 (internal_0n[317], complete899_0n[33], complete899_0n[34]);
  C3 I1667 (internal_0n[318], internal_0n[306], internal_0n[307], internal_0n[308]);
  C3 I1668 (internal_0n[319], internal_0n[309], internal_0n[310], internal_0n[311]);
  C3 I1669 (internal_0n[320], internal_0n[312], internal_0n[313], internal_0n[314]);
  C3 I1670 (internal_0n[321], internal_0n[315], internal_0n[316], internal_0n[317]);
  C2 I1671 (internal_0n[322], internal_0n[318], internal_0n[319]);
  C2 I1672 (internal_0n[323], internal_0n[320], internal_0n[321]);
  C2 I1673 (selcomp_1n, internal_0n[322], internal_0n[323]);
  OR2 I1674 (complete899_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I1675 (complete899_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I1676 (complete899_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I1677 (complete899_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I1678 (complete899_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I1679 (complete899_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I1680 (complete899_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I1681 (complete899_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I1682 (complete899_0n[8], ifint_1n[8], itint_1n[8]);
  OR2 I1683 (complete899_0n[9], ifint_1n[9], itint_1n[9]);
  OR2 I1684 (complete899_0n[10], ifint_1n[10], itint_1n[10]);
  OR2 I1685 (complete899_0n[11], ifint_1n[11], itint_1n[11]);
  OR2 I1686 (complete899_0n[12], ifint_1n[12], itint_1n[12]);
  OR2 I1687 (complete899_0n[13], ifint_1n[13], itint_1n[13]);
  OR2 I1688 (complete899_0n[14], ifint_1n[14], itint_1n[14]);
  OR2 I1689 (complete899_0n[15], ifint_1n[15], itint_1n[15]);
  OR2 I1690 (complete899_0n[16], ifint_1n[16], itint_1n[16]);
  OR2 I1691 (complete899_0n[17], ifint_1n[17], itint_1n[17]);
  OR2 I1692 (complete899_0n[18], ifint_1n[18], itint_1n[18]);
  OR2 I1693 (complete899_0n[19], ifint_1n[19], itint_1n[19]);
  OR2 I1694 (complete899_0n[20], ifint_1n[20], itint_1n[20]);
  OR2 I1695 (complete899_0n[21], ifint_1n[21], itint_1n[21]);
  OR2 I1696 (complete899_0n[22], ifint_1n[22], itint_1n[22]);
  OR2 I1697 (complete899_0n[23], ifint_1n[23], itint_1n[23]);
  OR2 I1698 (complete899_0n[24], ifint_1n[24], itint_1n[24]);
  OR2 I1699 (complete899_0n[25], ifint_1n[25], itint_1n[25]);
  OR2 I1700 (complete899_0n[26], ifint_1n[26], itint_1n[26]);
  OR2 I1701 (complete899_0n[27], ifint_1n[27], itint_1n[27]);
  OR2 I1702 (complete899_0n[28], ifint_1n[28], itint_1n[28]);
  OR2 I1703 (complete899_0n[29], ifint_1n[29], itint_1n[29]);
  OR2 I1704 (complete899_0n[30], ifint_1n[30], itint_1n[30]);
  OR2 I1705 (complete899_0n[31], ifint_1n[31], itint_1n[31]);
  OR2 I1706 (complete899_0n[32], ifint_1n[32], itint_1n[32]);
  OR2 I1707 (complete899_0n[33], ifint_1n[33], itint_1n[33]);
  OR2 I1708 (complete899_0n[34], ifint_1n[34], itint_1n[34]);
  C3 I1709 (internal_0n[324], complete898_0n[0], complete898_0n[1], complete898_0n[2]);
  C3 I1710 (internal_0n[325], complete898_0n[3], complete898_0n[4], complete898_0n[5]);
  C3 I1711 (internal_0n[326], complete898_0n[6], complete898_0n[7], complete898_0n[8]);
  C3 I1712 (internal_0n[327], complete898_0n[9], complete898_0n[10], complete898_0n[11]);
  C3 I1713 (internal_0n[328], complete898_0n[12], complete898_0n[13], complete898_0n[14]);
  C3 I1714 (internal_0n[329], complete898_0n[15], complete898_0n[16], complete898_0n[17]);
  C3 I1715 (internal_0n[330], complete898_0n[18], complete898_0n[19], complete898_0n[20]);
  C3 I1716 (internal_0n[331], complete898_0n[21], complete898_0n[22], complete898_0n[23]);
  C3 I1717 (internal_0n[332], complete898_0n[24], complete898_0n[25], complete898_0n[26]);
  C3 I1718 (internal_0n[333], complete898_0n[27], complete898_0n[28], complete898_0n[29]);
  C3 I1719 (internal_0n[334], complete898_0n[30], complete898_0n[31], complete898_0n[32]);
  C2 I1720 (internal_0n[335], complete898_0n[33], complete898_0n[34]);
  C3 I1721 (internal_0n[336], internal_0n[324], internal_0n[325], internal_0n[326]);
  C3 I1722 (internal_0n[337], internal_0n[327], internal_0n[328], internal_0n[329]);
  C3 I1723 (internal_0n[338], internal_0n[330], internal_0n[331], internal_0n[332]);
  C3 I1724 (internal_0n[339], internal_0n[333], internal_0n[334], internal_0n[335]);
  C2 I1725 (internal_0n[340], internal_0n[336], internal_0n[337]);
  C2 I1726 (internal_0n[341], internal_0n[338], internal_0n[339]);
  C2 I1727 (selcomp_0n, internal_0n[340], internal_0n[341]);
  OR2 I1728 (complete898_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I1729 (complete898_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I1730 (complete898_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I1731 (complete898_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I1732 (complete898_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I1733 (complete898_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I1734 (complete898_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I1735 (complete898_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I1736 (complete898_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I1737 (complete898_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I1738 (complete898_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I1739 (complete898_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I1740 (complete898_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I1741 (complete898_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I1742 (complete898_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I1743 (complete898_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I1744 (complete898_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I1745 (complete898_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I1746 (complete898_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I1747 (complete898_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I1748 (complete898_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I1749 (complete898_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I1750 (complete898_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I1751 (complete898_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I1752 (complete898_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I1753 (complete898_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I1754 (complete898_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I1755 (complete898_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I1756 (complete898_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I1757 (complete898_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I1758 (complete898_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I1759 (complete898_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I1760 (complete898_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I1761 (complete898_0n[33], ifint_0n[33], itint_0n[33]);
  OR2 I1762 (complete898_0n[34], ifint_0n[34], itint_0n[34]);
  AND2 I1763 (gfint_0n[0], gate_0n[0], ifint_0n[0]);
  AND2 I1764 (gfint_0n[1], gate_0n[0], ifint_0n[1]);
  AND2 I1765 (gfint_0n[2], gate_0n[0], ifint_0n[2]);
  AND2 I1766 (gfint_0n[3], gate_0n[0], ifint_0n[3]);
  AND2 I1767 (gfint_0n[4], gate_0n[0], ifint_0n[4]);
  AND2 I1768 (gfint_0n[5], gate_0n[0], ifint_0n[5]);
  AND2 I1769 (gfint_0n[6], gate_0n[0], ifint_0n[6]);
  AND2 I1770 (gfint_0n[7], gate_0n[0], ifint_0n[7]);
  AND2 I1771 (gfint_0n[8], gate_0n[0], ifint_0n[8]);
  AND2 I1772 (gfint_0n[9], gate_0n[0], ifint_0n[9]);
  AND2 I1773 (gfint_0n[10], gate_0n[0], ifint_0n[10]);
  AND2 I1774 (gfint_0n[11], gate_0n[0], ifint_0n[11]);
  AND2 I1775 (gfint_0n[12], gate_0n[0], ifint_0n[12]);
  AND2 I1776 (gfint_0n[13], gate_0n[0], ifint_0n[13]);
  AND2 I1777 (gfint_0n[14], gate_0n[0], ifint_0n[14]);
  AND2 I1778 (gfint_0n[15], gate_0n[0], ifint_0n[15]);
  AND2 I1779 (gfint_0n[16], gate_0n[0], ifint_0n[16]);
  AND2 I1780 (gfint_0n[17], gate_0n[0], ifint_0n[17]);
  AND2 I1781 (gfint_0n[18], gate_0n[0], ifint_0n[18]);
  AND2 I1782 (gfint_0n[19], gate_0n[0], ifint_0n[19]);
  AND2 I1783 (gfint_0n[20], gate_0n[0], ifint_0n[20]);
  AND2 I1784 (gfint_0n[21], gate_0n[0], ifint_0n[21]);
  AND2 I1785 (gfint_0n[22], gate_0n[0], ifint_0n[22]);
  AND2 I1786 (gfint_0n[23], gate_0n[0], ifint_0n[23]);
  AND2 I1787 (gfint_0n[24], gate_0n[0], ifint_0n[24]);
  AND2 I1788 (gfint_0n[25], gate_0n[0], ifint_0n[25]);
  AND2 I1789 (gfint_0n[26], gate_0n[0], ifint_0n[26]);
  AND2 I1790 (gfint_0n[27], gate_0n[0], ifint_0n[27]);
  AND2 I1791 (gfint_0n[28], gate_0n[0], ifint_0n[28]);
  AND2 I1792 (gfint_0n[29], gate_0n[0], ifint_0n[29]);
  AND2 I1793 (gfint_0n[30], gate_0n[0], ifint_0n[30]);
  AND2 I1794 (gfint_0n[31], gate_0n[0], ifint_0n[31]);
  AND2 I1795 (gfint_0n[32], gate_0n[0], ifint_0n[32]);
  AND2 I1796 (gfint_0n[33], gate_0n[0], ifint_0n[33]);
  AND2 I1797 (gfint_0n[34], gate_0n[0], ifint_0n[34]);
  AND2 I1798 (gfint_1n[0], gate_0n[1], ifint_1n[0]);
  AND2 I1799 (gfint_1n[1], gate_0n[1], ifint_1n[1]);
  AND2 I1800 (gfint_1n[2], gate_0n[1], ifint_1n[2]);
  AND2 I1801 (gfint_1n[3], gate_0n[1], ifint_1n[3]);
  AND2 I1802 (gfint_1n[4], gate_0n[1], ifint_1n[4]);
  AND2 I1803 (gfint_1n[5], gate_0n[1], ifint_1n[5]);
  AND2 I1804 (gfint_1n[6], gate_0n[1], ifint_1n[6]);
  AND2 I1805 (gfint_1n[7], gate_0n[1], ifint_1n[7]);
  AND2 I1806 (gfint_1n[8], gate_0n[1], ifint_1n[8]);
  AND2 I1807 (gfint_1n[9], gate_0n[1], ifint_1n[9]);
  AND2 I1808 (gfint_1n[10], gate_0n[1], ifint_1n[10]);
  AND2 I1809 (gfint_1n[11], gate_0n[1], ifint_1n[11]);
  AND2 I1810 (gfint_1n[12], gate_0n[1], ifint_1n[12]);
  AND2 I1811 (gfint_1n[13], gate_0n[1], ifint_1n[13]);
  AND2 I1812 (gfint_1n[14], gate_0n[1], ifint_1n[14]);
  AND2 I1813 (gfint_1n[15], gate_0n[1], ifint_1n[15]);
  AND2 I1814 (gfint_1n[16], gate_0n[1], ifint_1n[16]);
  AND2 I1815 (gfint_1n[17], gate_0n[1], ifint_1n[17]);
  AND2 I1816 (gfint_1n[18], gate_0n[1], ifint_1n[18]);
  AND2 I1817 (gfint_1n[19], gate_0n[1], ifint_1n[19]);
  AND2 I1818 (gfint_1n[20], gate_0n[1], ifint_1n[20]);
  AND2 I1819 (gfint_1n[21], gate_0n[1], ifint_1n[21]);
  AND2 I1820 (gfint_1n[22], gate_0n[1], ifint_1n[22]);
  AND2 I1821 (gfint_1n[23], gate_0n[1], ifint_1n[23]);
  AND2 I1822 (gfint_1n[24], gate_0n[1], ifint_1n[24]);
  AND2 I1823 (gfint_1n[25], gate_0n[1], ifint_1n[25]);
  AND2 I1824 (gfint_1n[26], gate_0n[1], ifint_1n[26]);
  AND2 I1825 (gfint_1n[27], gate_0n[1], ifint_1n[27]);
  AND2 I1826 (gfint_1n[28], gate_0n[1], ifint_1n[28]);
  AND2 I1827 (gfint_1n[29], gate_0n[1], ifint_1n[29]);
  AND2 I1828 (gfint_1n[30], gate_0n[1], ifint_1n[30]);
  AND2 I1829 (gfint_1n[31], gate_0n[1], ifint_1n[31]);
  AND2 I1830 (gfint_1n[32], gate_0n[1], ifint_1n[32]);
  AND2 I1831 (gfint_1n[33], gate_0n[1], ifint_1n[33]);
  AND2 I1832 (gfint_1n[34], gate_0n[1], ifint_1n[34]);
  AND2 I1833 (gfint_2n[0], gate_0n[2], ifint_2n[0]);
  AND2 I1834 (gfint_2n[1], gate_0n[2], ifint_2n[1]);
  AND2 I1835 (gfint_2n[2], gate_0n[2], ifint_2n[2]);
  AND2 I1836 (gfint_2n[3], gate_0n[2], ifint_2n[3]);
  AND2 I1837 (gfint_2n[4], gate_0n[2], ifint_2n[4]);
  AND2 I1838 (gfint_2n[5], gate_0n[2], ifint_2n[5]);
  AND2 I1839 (gfint_2n[6], gate_0n[2], ifint_2n[6]);
  AND2 I1840 (gfint_2n[7], gate_0n[2], ifint_2n[7]);
  AND2 I1841 (gfint_2n[8], gate_0n[2], ifint_2n[8]);
  AND2 I1842 (gfint_2n[9], gate_0n[2], ifint_2n[9]);
  AND2 I1843 (gfint_2n[10], gate_0n[2], ifint_2n[10]);
  AND2 I1844 (gfint_2n[11], gate_0n[2], ifint_2n[11]);
  AND2 I1845 (gfint_2n[12], gate_0n[2], ifint_2n[12]);
  AND2 I1846 (gfint_2n[13], gate_0n[2], ifint_2n[13]);
  AND2 I1847 (gfint_2n[14], gate_0n[2], ifint_2n[14]);
  AND2 I1848 (gfint_2n[15], gate_0n[2], ifint_2n[15]);
  AND2 I1849 (gfint_2n[16], gate_0n[2], ifint_2n[16]);
  AND2 I1850 (gfint_2n[17], gate_0n[2], ifint_2n[17]);
  AND2 I1851 (gfint_2n[18], gate_0n[2], ifint_2n[18]);
  AND2 I1852 (gfint_2n[19], gate_0n[2], ifint_2n[19]);
  AND2 I1853 (gfint_2n[20], gate_0n[2], ifint_2n[20]);
  AND2 I1854 (gfint_2n[21], gate_0n[2], ifint_2n[21]);
  AND2 I1855 (gfint_2n[22], gate_0n[2], ifint_2n[22]);
  AND2 I1856 (gfint_2n[23], gate_0n[2], ifint_2n[23]);
  AND2 I1857 (gfint_2n[24], gate_0n[2], ifint_2n[24]);
  AND2 I1858 (gfint_2n[25], gate_0n[2], ifint_2n[25]);
  AND2 I1859 (gfint_2n[26], gate_0n[2], ifint_2n[26]);
  AND2 I1860 (gfint_2n[27], gate_0n[2], ifint_2n[27]);
  AND2 I1861 (gfint_2n[28], gate_0n[2], ifint_2n[28]);
  AND2 I1862 (gfint_2n[29], gate_0n[2], ifint_2n[29]);
  AND2 I1863 (gfint_2n[30], gate_0n[2], ifint_2n[30]);
  AND2 I1864 (gfint_2n[31], gate_0n[2], ifint_2n[31]);
  AND2 I1865 (gfint_2n[32], gate_0n[2], ifint_2n[32]);
  AND2 I1866 (gfint_2n[33], gate_0n[2], ifint_2n[33]);
  AND2 I1867 (gfint_2n[34], gate_0n[2], ifint_2n[34]);
  AND2 I1868 (gfint_3n[0], gate_0n[3], ifint_3n[0]);
  AND2 I1869 (gfint_3n[1], gate_0n[3], ifint_3n[1]);
  AND2 I1870 (gfint_3n[2], gate_0n[3], ifint_3n[2]);
  AND2 I1871 (gfint_3n[3], gate_0n[3], ifint_3n[3]);
  AND2 I1872 (gfint_3n[4], gate_0n[3], ifint_3n[4]);
  AND2 I1873 (gfint_3n[5], gate_0n[3], ifint_3n[5]);
  AND2 I1874 (gfint_3n[6], gate_0n[3], ifint_3n[6]);
  AND2 I1875 (gfint_3n[7], gate_0n[3], ifint_3n[7]);
  AND2 I1876 (gfint_3n[8], gate_0n[3], ifint_3n[8]);
  AND2 I1877 (gfint_3n[9], gate_0n[3], ifint_3n[9]);
  AND2 I1878 (gfint_3n[10], gate_0n[3], ifint_3n[10]);
  AND2 I1879 (gfint_3n[11], gate_0n[3], ifint_3n[11]);
  AND2 I1880 (gfint_3n[12], gate_0n[3], ifint_3n[12]);
  AND2 I1881 (gfint_3n[13], gate_0n[3], ifint_3n[13]);
  AND2 I1882 (gfint_3n[14], gate_0n[3], ifint_3n[14]);
  AND2 I1883 (gfint_3n[15], gate_0n[3], ifint_3n[15]);
  AND2 I1884 (gfint_3n[16], gate_0n[3], ifint_3n[16]);
  AND2 I1885 (gfint_3n[17], gate_0n[3], ifint_3n[17]);
  AND2 I1886 (gfint_3n[18], gate_0n[3], ifint_3n[18]);
  AND2 I1887 (gfint_3n[19], gate_0n[3], ifint_3n[19]);
  AND2 I1888 (gfint_3n[20], gate_0n[3], ifint_3n[20]);
  AND2 I1889 (gfint_3n[21], gate_0n[3], ifint_3n[21]);
  AND2 I1890 (gfint_3n[22], gate_0n[3], ifint_3n[22]);
  AND2 I1891 (gfint_3n[23], gate_0n[3], ifint_3n[23]);
  AND2 I1892 (gfint_3n[24], gate_0n[3], ifint_3n[24]);
  AND2 I1893 (gfint_3n[25], gate_0n[3], ifint_3n[25]);
  AND2 I1894 (gfint_3n[26], gate_0n[3], ifint_3n[26]);
  AND2 I1895 (gfint_3n[27], gate_0n[3], ifint_3n[27]);
  AND2 I1896 (gfint_3n[28], gate_0n[3], ifint_3n[28]);
  AND2 I1897 (gfint_3n[29], gate_0n[3], ifint_3n[29]);
  AND2 I1898 (gfint_3n[30], gate_0n[3], ifint_3n[30]);
  AND2 I1899 (gfint_3n[31], gate_0n[3], ifint_3n[31]);
  AND2 I1900 (gfint_3n[32], gate_0n[3], ifint_3n[32]);
  AND2 I1901 (gfint_3n[33], gate_0n[3], ifint_3n[33]);
  AND2 I1902 (gfint_3n[34], gate_0n[3], ifint_3n[34]);
  AND2 I1903 (gfint_4n[0], gate_0n[4], ifint_4n[0]);
  AND2 I1904 (gfint_4n[1], gate_0n[4], ifint_4n[1]);
  AND2 I1905 (gfint_4n[2], gate_0n[4], ifint_4n[2]);
  AND2 I1906 (gfint_4n[3], gate_0n[4], ifint_4n[3]);
  AND2 I1907 (gfint_4n[4], gate_0n[4], ifint_4n[4]);
  AND2 I1908 (gfint_4n[5], gate_0n[4], ifint_4n[5]);
  AND2 I1909 (gfint_4n[6], gate_0n[4], ifint_4n[6]);
  AND2 I1910 (gfint_4n[7], gate_0n[4], ifint_4n[7]);
  AND2 I1911 (gfint_4n[8], gate_0n[4], ifint_4n[8]);
  AND2 I1912 (gfint_4n[9], gate_0n[4], ifint_4n[9]);
  AND2 I1913 (gfint_4n[10], gate_0n[4], ifint_4n[10]);
  AND2 I1914 (gfint_4n[11], gate_0n[4], ifint_4n[11]);
  AND2 I1915 (gfint_4n[12], gate_0n[4], ifint_4n[12]);
  AND2 I1916 (gfint_4n[13], gate_0n[4], ifint_4n[13]);
  AND2 I1917 (gfint_4n[14], gate_0n[4], ifint_4n[14]);
  AND2 I1918 (gfint_4n[15], gate_0n[4], ifint_4n[15]);
  AND2 I1919 (gfint_4n[16], gate_0n[4], ifint_4n[16]);
  AND2 I1920 (gfint_4n[17], gate_0n[4], ifint_4n[17]);
  AND2 I1921 (gfint_4n[18], gate_0n[4], ifint_4n[18]);
  AND2 I1922 (gfint_4n[19], gate_0n[4], ifint_4n[19]);
  AND2 I1923 (gfint_4n[20], gate_0n[4], ifint_4n[20]);
  AND2 I1924 (gfint_4n[21], gate_0n[4], ifint_4n[21]);
  AND2 I1925 (gfint_4n[22], gate_0n[4], ifint_4n[22]);
  AND2 I1926 (gfint_4n[23], gate_0n[4], ifint_4n[23]);
  AND2 I1927 (gfint_4n[24], gate_0n[4], ifint_4n[24]);
  AND2 I1928 (gfint_4n[25], gate_0n[4], ifint_4n[25]);
  AND2 I1929 (gfint_4n[26], gate_0n[4], ifint_4n[26]);
  AND2 I1930 (gfint_4n[27], gate_0n[4], ifint_4n[27]);
  AND2 I1931 (gfint_4n[28], gate_0n[4], ifint_4n[28]);
  AND2 I1932 (gfint_4n[29], gate_0n[4], ifint_4n[29]);
  AND2 I1933 (gfint_4n[30], gate_0n[4], ifint_4n[30]);
  AND2 I1934 (gfint_4n[31], gate_0n[4], ifint_4n[31]);
  AND2 I1935 (gfint_4n[32], gate_0n[4], ifint_4n[32]);
  AND2 I1936 (gfint_4n[33], gate_0n[4], ifint_4n[33]);
  AND2 I1937 (gfint_4n[34], gate_0n[4], ifint_4n[34]);
  AND2 I1938 (gfint_5n[0], gate_0n[5], ifint_5n[0]);
  AND2 I1939 (gfint_5n[1], gate_0n[5], ifint_5n[1]);
  AND2 I1940 (gfint_5n[2], gate_0n[5], ifint_5n[2]);
  AND2 I1941 (gfint_5n[3], gate_0n[5], ifint_5n[3]);
  AND2 I1942 (gfint_5n[4], gate_0n[5], ifint_5n[4]);
  AND2 I1943 (gfint_5n[5], gate_0n[5], ifint_5n[5]);
  AND2 I1944 (gfint_5n[6], gate_0n[5], ifint_5n[6]);
  AND2 I1945 (gfint_5n[7], gate_0n[5], ifint_5n[7]);
  AND2 I1946 (gfint_5n[8], gate_0n[5], ifint_5n[8]);
  AND2 I1947 (gfint_5n[9], gate_0n[5], ifint_5n[9]);
  AND2 I1948 (gfint_5n[10], gate_0n[5], ifint_5n[10]);
  AND2 I1949 (gfint_5n[11], gate_0n[5], ifint_5n[11]);
  AND2 I1950 (gfint_5n[12], gate_0n[5], ifint_5n[12]);
  AND2 I1951 (gfint_5n[13], gate_0n[5], ifint_5n[13]);
  AND2 I1952 (gfint_5n[14], gate_0n[5], ifint_5n[14]);
  AND2 I1953 (gfint_5n[15], gate_0n[5], ifint_5n[15]);
  AND2 I1954 (gfint_5n[16], gate_0n[5], ifint_5n[16]);
  AND2 I1955 (gfint_5n[17], gate_0n[5], ifint_5n[17]);
  AND2 I1956 (gfint_5n[18], gate_0n[5], ifint_5n[18]);
  AND2 I1957 (gfint_5n[19], gate_0n[5], ifint_5n[19]);
  AND2 I1958 (gfint_5n[20], gate_0n[5], ifint_5n[20]);
  AND2 I1959 (gfint_5n[21], gate_0n[5], ifint_5n[21]);
  AND2 I1960 (gfint_5n[22], gate_0n[5], ifint_5n[22]);
  AND2 I1961 (gfint_5n[23], gate_0n[5], ifint_5n[23]);
  AND2 I1962 (gfint_5n[24], gate_0n[5], ifint_5n[24]);
  AND2 I1963 (gfint_5n[25], gate_0n[5], ifint_5n[25]);
  AND2 I1964 (gfint_5n[26], gate_0n[5], ifint_5n[26]);
  AND2 I1965 (gfint_5n[27], gate_0n[5], ifint_5n[27]);
  AND2 I1966 (gfint_5n[28], gate_0n[5], ifint_5n[28]);
  AND2 I1967 (gfint_5n[29], gate_0n[5], ifint_5n[29]);
  AND2 I1968 (gfint_5n[30], gate_0n[5], ifint_5n[30]);
  AND2 I1969 (gfint_5n[31], gate_0n[5], ifint_5n[31]);
  AND2 I1970 (gfint_5n[32], gate_0n[5], ifint_5n[32]);
  AND2 I1971 (gfint_5n[33], gate_0n[5], ifint_5n[33]);
  AND2 I1972 (gfint_5n[34], gate_0n[5], ifint_5n[34]);
  AND2 I1973 (gfint_6n[0], gate_0n[6], ifint_6n[0]);
  AND2 I1974 (gfint_6n[1], gate_0n[6], ifint_6n[1]);
  AND2 I1975 (gfint_6n[2], gate_0n[6], ifint_6n[2]);
  AND2 I1976 (gfint_6n[3], gate_0n[6], ifint_6n[3]);
  AND2 I1977 (gfint_6n[4], gate_0n[6], ifint_6n[4]);
  AND2 I1978 (gfint_6n[5], gate_0n[6], ifint_6n[5]);
  AND2 I1979 (gfint_6n[6], gate_0n[6], ifint_6n[6]);
  AND2 I1980 (gfint_6n[7], gate_0n[6], ifint_6n[7]);
  AND2 I1981 (gfint_6n[8], gate_0n[6], ifint_6n[8]);
  AND2 I1982 (gfint_6n[9], gate_0n[6], ifint_6n[9]);
  AND2 I1983 (gfint_6n[10], gate_0n[6], ifint_6n[10]);
  AND2 I1984 (gfint_6n[11], gate_0n[6], ifint_6n[11]);
  AND2 I1985 (gfint_6n[12], gate_0n[6], ifint_6n[12]);
  AND2 I1986 (gfint_6n[13], gate_0n[6], ifint_6n[13]);
  AND2 I1987 (gfint_6n[14], gate_0n[6], ifint_6n[14]);
  AND2 I1988 (gfint_6n[15], gate_0n[6], ifint_6n[15]);
  AND2 I1989 (gfint_6n[16], gate_0n[6], ifint_6n[16]);
  AND2 I1990 (gfint_6n[17], gate_0n[6], ifint_6n[17]);
  AND2 I1991 (gfint_6n[18], gate_0n[6], ifint_6n[18]);
  AND2 I1992 (gfint_6n[19], gate_0n[6], ifint_6n[19]);
  AND2 I1993 (gfint_6n[20], gate_0n[6], ifint_6n[20]);
  AND2 I1994 (gfint_6n[21], gate_0n[6], ifint_6n[21]);
  AND2 I1995 (gfint_6n[22], gate_0n[6], ifint_6n[22]);
  AND2 I1996 (gfint_6n[23], gate_0n[6], ifint_6n[23]);
  AND2 I1997 (gfint_6n[24], gate_0n[6], ifint_6n[24]);
  AND2 I1998 (gfint_6n[25], gate_0n[6], ifint_6n[25]);
  AND2 I1999 (gfint_6n[26], gate_0n[6], ifint_6n[26]);
  AND2 I2000 (gfint_6n[27], gate_0n[6], ifint_6n[27]);
  AND2 I2001 (gfint_6n[28], gate_0n[6], ifint_6n[28]);
  AND2 I2002 (gfint_6n[29], gate_0n[6], ifint_6n[29]);
  AND2 I2003 (gfint_6n[30], gate_0n[6], ifint_6n[30]);
  AND2 I2004 (gfint_6n[31], gate_0n[6], ifint_6n[31]);
  AND2 I2005 (gfint_6n[32], gate_0n[6], ifint_6n[32]);
  AND2 I2006 (gfint_6n[33], gate_0n[6], ifint_6n[33]);
  AND2 I2007 (gfint_6n[34], gate_0n[6], ifint_6n[34]);
  AND2 I2008 (gfint_7n[0], gate_0n[7], ifint_7n[0]);
  AND2 I2009 (gfint_7n[1], gate_0n[7], ifint_7n[1]);
  AND2 I2010 (gfint_7n[2], gate_0n[7], ifint_7n[2]);
  AND2 I2011 (gfint_7n[3], gate_0n[7], ifint_7n[3]);
  AND2 I2012 (gfint_7n[4], gate_0n[7], ifint_7n[4]);
  AND2 I2013 (gfint_7n[5], gate_0n[7], ifint_7n[5]);
  AND2 I2014 (gfint_7n[6], gate_0n[7], ifint_7n[6]);
  AND2 I2015 (gfint_7n[7], gate_0n[7], ifint_7n[7]);
  AND2 I2016 (gfint_7n[8], gate_0n[7], ifint_7n[8]);
  AND2 I2017 (gfint_7n[9], gate_0n[7], ifint_7n[9]);
  AND2 I2018 (gfint_7n[10], gate_0n[7], ifint_7n[10]);
  AND2 I2019 (gfint_7n[11], gate_0n[7], ifint_7n[11]);
  AND2 I2020 (gfint_7n[12], gate_0n[7], ifint_7n[12]);
  AND2 I2021 (gfint_7n[13], gate_0n[7], ifint_7n[13]);
  AND2 I2022 (gfint_7n[14], gate_0n[7], ifint_7n[14]);
  AND2 I2023 (gfint_7n[15], gate_0n[7], ifint_7n[15]);
  AND2 I2024 (gfint_7n[16], gate_0n[7], ifint_7n[16]);
  AND2 I2025 (gfint_7n[17], gate_0n[7], ifint_7n[17]);
  AND2 I2026 (gfint_7n[18], gate_0n[7], ifint_7n[18]);
  AND2 I2027 (gfint_7n[19], gate_0n[7], ifint_7n[19]);
  AND2 I2028 (gfint_7n[20], gate_0n[7], ifint_7n[20]);
  AND2 I2029 (gfint_7n[21], gate_0n[7], ifint_7n[21]);
  AND2 I2030 (gfint_7n[22], gate_0n[7], ifint_7n[22]);
  AND2 I2031 (gfint_7n[23], gate_0n[7], ifint_7n[23]);
  AND2 I2032 (gfint_7n[24], gate_0n[7], ifint_7n[24]);
  AND2 I2033 (gfint_7n[25], gate_0n[7], ifint_7n[25]);
  AND2 I2034 (gfint_7n[26], gate_0n[7], ifint_7n[26]);
  AND2 I2035 (gfint_7n[27], gate_0n[7], ifint_7n[27]);
  AND2 I2036 (gfint_7n[28], gate_0n[7], ifint_7n[28]);
  AND2 I2037 (gfint_7n[29], gate_0n[7], ifint_7n[29]);
  AND2 I2038 (gfint_7n[30], gate_0n[7], ifint_7n[30]);
  AND2 I2039 (gfint_7n[31], gate_0n[7], ifint_7n[31]);
  AND2 I2040 (gfint_7n[32], gate_0n[7], ifint_7n[32]);
  AND2 I2041 (gfint_7n[33], gate_0n[7], ifint_7n[33]);
  AND2 I2042 (gfint_7n[34], gate_0n[7], ifint_7n[34]);
  AND2 I2043 (gfint_8n[0], gate_0n[8], ifint_8n[0]);
  AND2 I2044 (gfint_8n[1], gate_0n[8], ifint_8n[1]);
  AND2 I2045 (gfint_8n[2], gate_0n[8], ifint_8n[2]);
  AND2 I2046 (gfint_8n[3], gate_0n[8], ifint_8n[3]);
  AND2 I2047 (gfint_8n[4], gate_0n[8], ifint_8n[4]);
  AND2 I2048 (gfint_8n[5], gate_0n[8], ifint_8n[5]);
  AND2 I2049 (gfint_8n[6], gate_0n[8], ifint_8n[6]);
  AND2 I2050 (gfint_8n[7], gate_0n[8], ifint_8n[7]);
  AND2 I2051 (gfint_8n[8], gate_0n[8], ifint_8n[8]);
  AND2 I2052 (gfint_8n[9], gate_0n[8], ifint_8n[9]);
  AND2 I2053 (gfint_8n[10], gate_0n[8], ifint_8n[10]);
  AND2 I2054 (gfint_8n[11], gate_0n[8], ifint_8n[11]);
  AND2 I2055 (gfint_8n[12], gate_0n[8], ifint_8n[12]);
  AND2 I2056 (gfint_8n[13], gate_0n[8], ifint_8n[13]);
  AND2 I2057 (gfint_8n[14], gate_0n[8], ifint_8n[14]);
  AND2 I2058 (gfint_8n[15], gate_0n[8], ifint_8n[15]);
  AND2 I2059 (gfint_8n[16], gate_0n[8], ifint_8n[16]);
  AND2 I2060 (gfint_8n[17], gate_0n[8], ifint_8n[17]);
  AND2 I2061 (gfint_8n[18], gate_0n[8], ifint_8n[18]);
  AND2 I2062 (gfint_8n[19], gate_0n[8], ifint_8n[19]);
  AND2 I2063 (gfint_8n[20], gate_0n[8], ifint_8n[20]);
  AND2 I2064 (gfint_8n[21], gate_0n[8], ifint_8n[21]);
  AND2 I2065 (gfint_8n[22], gate_0n[8], ifint_8n[22]);
  AND2 I2066 (gfint_8n[23], gate_0n[8], ifint_8n[23]);
  AND2 I2067 (gfint_8n[24], gate_0n[8], ifint_8n[24]);
  AND2 I2068 (gfint_8n[25], gate_0n[8], ifint_8n[25]);
  AND2 I2069 (gfint_8n[26], gate_0n[8], ifint_8n[26]);
  AND2 I2070 (gfint_8n[27], gate_0n[8], ifint_8n[27]);
  AND2 I2071 (gfint_8n[28], gate_0n[8], ifint_8n[28]);
  AND2 I2072 (gfint_8n[29], gate_0n[8], ifint_8n[29]);
  AND2 I2073 (gfint_8n[30], gate_0n[8], ifint_8n[30]);
  AND2 I2074 (gfint_8n[31], gate_0n[8], ifint_8n[31]);
  AND2 I2075 (gfint_8n[32], gate_0n[8], ifint_8n[32]);
  AND2 I2076 (gfint_8n[33], gate_0n[8], ifint_8n[33]);
  AND2 I2077 (gfint_8n[34], gate_0n[8], ifint_8n[34]);
  AND2 I2078 (gtint_0n[0], gate_0n[0], itint_0n[0]);
  AND2 I2079 (gtint_0n[1], gate_0n[0], itint_0n[1]);
  AND2 I2080 (gtint_0n[2], gate_0n[0], itint_0n[2]);
  AND2 I2081 (gtint_0n[3], gate_0n[0], itint_0n[3]);
  AND2 I2082 (gtint_0n[4], gate_0n[0], itint_0n[4]);
  AND2 I2083 (gtint_0n[5], gate_0n[0], itint_0n[5]);
  AND2 I2084 (gtint_0n[6], gate_0n[0], itint_0n[6]);
  AND2 I2085 (gtint_0n[7], gate_0n[0], itint_0n[7]);
  AND2 I2086 (gtint_0n[8], gate_0n[0], itint_0n[8]);
  AND2 I2087 (gtint_0n[9], gate_0n[0], itint_0n[9]);
  AND2 I2088 (gtint_0n[10], gate_0n[0], itint_0n[10]);
  AND2 I2089 (gtint_0n[11], gate_0n[0], itint_0n[11]);
  AND2 I2090 (gtint_0n[12], gate_0n[0], itint_0n[12]);
  AND2 I2091 (gtint_0n[13], gate_0n[0], itint_0n[13]);
  AND2 I2092 (gtint_0n[14], gate_0n[0], itint_0n[14]);
  AND2 I2093 (gtint_0n[15], gate_0n[0], itint_0n[15]);
  AND2 I2094 (gtint_0n[16], gate_0n[0], itint_0n[16]);
  AND2 I2095 (gtint_0n[17], gate_0n[0], itint_0n[17]);
  AND2 I2096 (gtint_0n[18], gate_0n[0], itint_0n[18]);
  AND2 I2097 (gtint_0n[19], gate_0n[0], itint_0n[19]);
  AND2 I2098 (gtint_0n[20], gate_0n[0], itint_0n[20]);
  AND2 I2099 (gtint_0n[21], gate_0n[0], itint_0n[21]);
  AND2 I2100 (gtint_0n[22], gate_0n[0], itint_0n[22]);
  AND2 I2101 (gtint_0n[23], gate_0n[0], itint_0n[23]);
  AND2 I2102 (gtint_0n[24], gate_0n[0], itint_0n[24]);
  AND2 I2103 (gtint_0n[25], gate_0n[0], itint_0n[25]);
  AND2 I2104 (gtint_0n[26], gate_0n[0], itint_0n[26]);
  AND2 I2105 (gtint_0n[27], gate_0n[0], itint_0n[27]);
  AND2 I2106 (gtint_0n[28], gate_0n[0], itint_0n[28]);
  AND2 I2107 (gtint_0n[29], gate_0n[0], itint_0n[29]);
  AND2 I2108 (gtint_0n[30], gate_0n[0], itint_0n[30]);
  AND2 I2109 (gtint_0n[31], gate_0n[0], itint_0n[31]);
  AND2 I2110 (gtint_0n[32], gate_0n[0], itint_0n[32]);
  AND2 I2111 (gtint_0n[33], gate_0n[0], itint_0n[33]);
  AND2 I2112 (gtint_0n[34], gate_0n[0], itint_0n[34]);
  AND2 I2113 (gtint_1n[0], gate_0n[1], itint_1n[0]);
  AND2 I2114 (gtint_1n[1], gate_0n[1], itint_1n[1]);
  AND2 I2115 (gtint_1n[2], gate_0n[1], itint_1n[2]);
  AND2 I2116 (gtint_1n[3], gate_0n[1], itint_1n[3]);
  AND2 I2117 (gtint_1n[4], gate_0n[1], itint_1n[4]);
  AND2 I2118 (gtint_1n[5], gate_0n[1], itint_1n[5]);
  AND2 I2119 (gtint_1n[6], gate_0n[1], itint_1n[6]);
  AND2 I2120 (gtint_1n[7], gate_0n[1], itint_1n[7]);
  AND2 I2121 (gtint_1n[8], gate_0n[1], itint_1n[8]);
  AND2 I2122 (gtint_1n[9], gate_0n[1], itint_1n[9]);
  AND2 I2123 (gtint_1n[10], gate_0n[1], itint_1n[10]);
  AND2 I2124 (gtint_1n[11], gate_0n[1], itint_1n[11]);
  AND2 I2125 (gtint_1n[12], gate_0n[1], itint_1n[12]);
  AND2 I2126 (gtint_1n[13], gate_0n[1], itint_1n[13]);
  AND2 I2127 (gtint_1n[14], gate_0n[1], itint_1n[14]);
  AND2 I2128 (gtint_1n[15], gate_0n[1], itint_1n[15]);
  AND2 I2129 (gtint_1n[16], gate_0n[1], itint_1n[16]);
  AND2 I2130 (gtint_1n[17], gate_0n[1], itint_1n[17]);
  AND2 I2131 (gtint_1n[18], gate_0n[1], itint_1n[18]);
  AND2 I2132 (gtint_1n[19], gate_0n[1], itint_1n[19]);
  AND2 I2133 (gtint_1n[20], gate_0n[1], itint_1n[20]);
  AND2 I2134 (gtint_1n[21], gate_0n[1], itint_1n[21]);
  AND2 I2135 (gtint_1n[22], gate_0n[1], itint_1n[22]);
  AND2 I2136 (gtint_1n[23], gate_0n[1], itint_1n[23]);
  AND2 I2137 (gtint_1n[24], gate_0n[1], itint_1n[24]);
  AND2 I2138 (gtint_1n[25], gate_0n[1], itint_1n[25]);
  AND2 I2139 (gtint_1n[26], gate_0n[1], itint_1n[26]);
  AND2 I2140 (gtint_1n[27], gate_0n[1], itint_1n[27]);
  AND2 I2141 (gtint_1n[28], gate_0n[1], itint_1n[28]);
  AND2 I2142 (gtint_1n[29], gate_0n[1], itint_1n[29]);
  AND2 I2143 (gtint_1n[30], gate_0n[1], itint_1n[30]);
  AND2 I2144 (gtint_1n[31], gate_0n[1], itint_1n[31]);
  AND2 I2145 (gtint_1n[32], gate_0n[1], itint_1n[32]);
  AND2 I2146 (gtint_1n[33], gate_0n[1], itint_1n[33]);
  AND2 I2147 (gtint_1n[34], gate_0n[1], itint_1n[34]);
  AND2 I2148 (gtint_2n[0], gate_0n[2], itint_2n[0]);
  AND2 I2149 (gtint_2n[1], gate_0n[2], itint_2n[1]);
  AND2 I2150 (gtint_2n[2], gate_0n[2], itint_2n[2]);
  AND2 I2151 (gtint_2n[3], gate_0n[2], itint_2n[3]);
  AND2 I2152 (gtint_2n[4], gate_0n[2], itint_2n[4]);
  AND2 I2153 (gtint_2n[5], gate_0n[2], itint_2n[5]);
  AND2 I2154 (gtint_2n[6], gate_0n[2], itint_2n[6]);
  AND2 I2155 (gtint_2n[7], gate_0n[2], itint_2n[7]);
  AND2 I2156 (gtint_2n[8], gate_0n[2], itint_2n[8]);
  AND2 I2157 (gtint_2n[9], gate_0n[2], itint_2n[9]);
  AND2 I2158 (gtint_2n[10], gate_0n[2], itint_2n[10]);
  AND2 I2159 (gtint_2n[11], gate_0n[2], itint_2n[11]);
  AND2 I2160 (gtint_2n[12], gate_0n[2], itint_2n[12]);
  AND2 I2161 (gtint_2n[13], gate_0n[2], itint_2n[13]);
  AND2 I2162 (gtint_2n[14], gate_0n[2], itint_2n[14]);
  AND2 I2163 (gtint_2n[15], gate_0n[2], itint_2n[15]);
  AND2 I2164 (gtint_2n[16], gate_0n[2], itint_2n[16]);
  AND2 I2165 (gtint_2n[17], gate_0n[2], itint_2n[17]);
  AND2 I2166 (gtint_2n[18], gate_0n[2], itint_2n[18]);
  AND2 I2167 (gtint_2n[19], gate_0n[2], itint_2n[19]);
  AND2 I2168 (gtint_2n[20], gate_0n[2], itint_2n[20]);
  AND2 I2169 (gtint_2n[21], gate_0n[2], itint_2n[21]);
  AND2 I2170 (gtint_2n[22], gate_0n[2], itint_2n[22]);
  AND2 I2171 (gtint_2n[23], gate_0n[2], itint_2n[23]);
  AND2 I2172 (gtint_2n[24], gate_0n[2], itint_2n[24]);
  AND2 I2173 (gtint_2n[25], gate_0n[2], itint_2n[25]);
  AND2 I2174 (gtint_2n[26], gate_0n[2], itint_2n[26]);
  AND2 I2175 (gtint_2n[27], gate_0n[2], itint_2n[27]);
  AND2 I2176 (gtint_2n[28], gate_0n[2], itint_2n[28]);
  AND2 I2177 (gtint_2n[29], gate_0n[2], itint_2n[29]);
  AND2 I2178 (gtint_2n[30], gate_0n[2], itint_2n[30]);
  AND2 I2179 (gtint_2n[31], gate_0n[2], itint_2n[31]);
  AND2 I2180 (gtint_2n[32], gate_0n[2], itint_2n[32]);
  AND2 I2181 (gtint_2n[33], gate_0n[2], itint_2n[33]);
  AND2 I2182 (gtint_2n[34], gate_0n[2], itint_2n[34]);
  AND2 I2183 (gtint_3n[0], gate_0n[3], itint_3n[0]);
  AND2 I2184 (gtint_3n[1], gate_0n[3], itint_3n[1]);
  AND2 I2185 (gtint_3n[2], gate_0n[3], itint_3n[2]);
  AND2 I2186 (gtint_3n[3], gate_0n[3], itint_3n[3]);
  AND2 I2187 (gtint_3n[4], gate_0n[3], itint_3n[4]);
  AND2 I2188 (gtint_3n[5], gate_0n[3], itint_3n[5]);
  AND2 I2189 (gtint_3n[6], gate_0n[3], itint_3n[6]);
  AND2 I2190 (gtint_3n[7], gate_0n[3], itint_3n[7]);
  AND2 I2191 (gtint_3n[8], gate_0n[3], itint_3n[8]);
  AND2 I2192 (gtint_3n[9], gate_0n[3], itint_3n[9]);
  AND2 I2193 (gtint_3n[10], gate_0n[3], itint_3n[10]);
  AND2 I2194 (gtint_3n[11], gate_0n[3], itint_3n[11]);
  AND2 I2195 (gtint_3n[12], gate_0n[3], itint_3n[12]);
  AND2 I2196 (gtint_3n[13], gate_0n[3], itint_3n[13]);
  AND2 I2197 (gtint_3n[14], gate_0n[3], itint_3n[14]);
  AND2 I2198 (gtint_3n[15], gate_0n[3], itint_3n[15]);
  AND2 I2199 (gtint_3n[16], gate_0n[3], itint_3n[16]);
  AND2 I2200 (gtint_3n[17], gate_0n[3], itint_3n[17]);
  AND2 I2201 (gtint_3n[18], gate_0n[3], itint_3n[18]);
  AND2 I2202 (gtint_3n[19], gate_0n[3], itint_3n[19]);
  AND2 I2203 (gtint_3n[20], gate_0n[3], itint_3n[20]);
  AND2 I2204 (gtint_3n[21], gate_0n[3], itint_3n[21]);
  AND2 I2205 (gtint_3n[22], gate_0n[3], itint_3n[22]);
  AND2 I2206 (gtint_3n[23], gate_0n[3], itint_3n[23]);
  AND2 I2207 (gtint_3n[24], gate_0n[3], itint_3n[24]);
  AND2 I2208 (gtint_3n[25], gate_0n[3], itint_3n[25]);
  AND2 I2209 (gtint_3n[26], gate_0n[3], itint_3n[26]);
  AND2 I2210 (gtint_3n[27], gate_0n[3], itint_3n[27]);
  AND2 I2211 (gtint_3n[28], gate_0n[3], itint_3n[28]);
  AND2 I2212 (gtint_3n[29], gate_0n[3], itint_3n[29]);
  AND2 I2213 (gtint_3n[30], gate_0n[3], itint_3n[30]);
  AND2 I2214 (gtint_3n[31], gate_0n[3], itint_3n[31]);
  AND2 I2215 (gtint_3n[32], gate_0n[3], itint_3n[32]);
  AND2 I2216 (gtint_3n[33], gate_0n[3], itint_3n[33]);
  AND2 I2217 (gtint_3n[34], gate_0n[3], itint_3n[34]);
  AND2 I2218 (gtint_4n[0], gate_0n[4], itint_4n[0]);
  AND2 I2219 (gtint_4n[1], gate_0n[4], itint_4n[1]);
  AND2 I2220 (gtint_4n[2], gate_0n[4], itint_4n[2]);
  AND2 I2221 (gtint_4n[3], gate_0n[4], itint_4n[3]);
  AND2 I2222 (gtint_4n[4], gate_0n[4], itint_4n[4]);
  AND2 I2223 (gtint_4n[5], gate_0n[4], itint_4n[5]);
  AND2 I2224 (gtint_4n[6], gate_0n[4], itint_4n[6]);
  AND2 I2225 (gtint_4n[7], gate_0n[4], itint_4n[7]);
  AND2 I2226 (gtint_4n[8], gate_0n[4], itint_4n[8]);
  AND2 I2227 (gtint_4n[9], gate_0n[4], itint_4n[9]);
  AND2 I2228 (gtint_4n[10], gate_0n[4], itint_4n[10]);
  AND2 I2229 (gtint_4n[11], gate_0n[4], itint_4n[11]);
  AND2 I2230 (gtint_4n[12], gate_0n[4], itint_4n[12]);
  AND2 I2231 (gtint_4n[13], gate_0n[4], itint_4n[13]);
  AND2 I2232 (gtint_4n[14], gate_0n[4], itint_4n[14]);
  AND2 I2233 (gtint_4n[15], gate_0n[4], itint_4n[15]);
  AND2 I2234 (gtint_4n[16], gate_0n[4], itint_4n[16]);
  AND2 I2235 (gtint_4n[17], gate_0n[4], itint_4n[17]);
  AND2 I2236 (gtint_4n[18], gate_0n[4], itint_4n[18]);
  AND2 I2237 (gtint_4n[19], gate_0n[4], itint_4n[19]);
  AND2 I2238 (gtint_4n[20], gate_0n[4], itint_4n[20]);
  AND2 I2239 (gtint_4n[21], gate_0n[4], itint_4n[21]);
  AND2 I2240 (gtint_4n[22], gate_0n[4], itint_4n[22]);
  AND2 I2241 (gtint_4n[23], gate_0n[4], itint_4n[23]);
  AND2 I2242 (gtint_4n[24], gate_0n[4], itint_4n[24]);
  AND2 I2243 (gtint_4n[25], gate_0n[4], itint_4n[25]);
  AND2 I2244 (gtint_4n[26], gate_0n[4], itint_4n[26]);
  AND2 I2245 (gtint_4n[27], gate_0n[4], itint_4n[27]);
  AND2 I2246 (gtint_4n[28], gate_0n[4], itint_4n[28]);
  AND2 I2247 (gtint_4n[29], gate_0n[4], itint_4n[29]);
  AND2 I2248 (gtint_4n[30], gate_0n[4], itint_4n[30]);
  AND2 I2249 (gtint_4n[31], gate_0n[4], itint_4n[31]);
  AND2 I2250 (gtint_4n[32], gate_0n[4], itint_4n[32]);
  AND2 I2251 (gtint_4n[33], gate_0n[4], itint_4n[33]);
  AND2 I2252 (gtint_4n[34], gate_0n[4], itint_4n[34]);
  AND2 I2253 (gtint_5n[0], gate_0n[5], itint_5n[0]);
  AND2 I2254 (gtint_5n[1], gate_0n[5], itint_5n[1]);
  AND2 I2255 (gtint_5n[2], gate_0n[5], itint_5n[2]);
  AND2 I2256 (gtint_5n[3], gate_0n[5], itint_5n[3]);
  AND2 I2257 (gtint_5n[4], gate_0n[5], itint_5n[4]);
  AND2 I2258 (gtint_5n[5], gate_0n[5], itint_5n[5]);
  AND2 I2259 (gtint_5n[6], gate_0n[5], itint_5n[6]);
  AND2 I2260 (gtint_5n[7], gate_0n[5], itint_5n[7]);
  AND2 I2261 (gtint_5n[8], gate_0n[5], itint_5n[8]);
  AND2 I2262 (gtint_5n[9], gate_0n[5], itint_5n[9]);
  AND2 I2263 (gtint_5n[10], gate_0n[5], itint_5n[10]);
  AND2 I2264 (gtint_5n[11], gate_0n[5], itint_5n[11]);
  AND2 I2265 (gtint_5n[12], gate_0n[5], itint_5n[12]);
  AND2 I2266 (gtint_5n[13], gate_0n[5], itint_5n[13]);
  AND2 I2267 (gtint_5n[14], gate_0n[5], itint_5n[14]);
  AND2 I2268 (gtint_5n[15], gate_0n[5], itint_5n[15]);
  AND2 I2269 (gtint_5n[16], gate_0n[5], itint_5n[16]);
  AND2 I2270 (gtint_5n[17], gate_0n[5], itint_5n[17]);
  AND2 I2271 (gtint_5n[18], gate_0n[5], itint_5n[18]);
  AND2 I2272 (gtint_5n[19], gate_0n[5], itint_5n[19]);
  AND2 I2273 (gtint_5n[20], gate_0n[5], itint_5n[20]);
  AND2 I2274 (gtint_5n[21], gate_0n[5], itint_5n[21]);
  AND2 I2275 (gtint_5n[22], gate_0n[5], itint_5n[22]);
  AND2 I2276 (gtint_5n[23], gate_0n[5], itint_5n[23]);
  AND2 I2277 (gtint_5n[24], gate_0n[5], itint_5n[24]);
  AND2 I2278 (gtint_5n[25], gate_0n[5], itint_5n[25]);
  AND2 I2279 (gtint_5n[26], gate_0n[5], itint_5n[26]);
  AND2 I2280 (gtint_5n[27], gate_0n[5], itint_5n[27]);
  AND2 I2281 (gtint_5n[28], gate_0n[5], itint_5n[28]);
  AND2 I2282 (gtint_5n[29], gate_0n[5], itint_5n[29]);
  AND2 I2283 (gtint_5n[30], gate_0n[5], itint_5n[30]);
  AND2 I2284 (gtint_5n[31], gate_0n[5], itint_5n[31]);
  AND2 I2285 (gtint_5n[32], gate_0n[5], itint_5n[32]);
  AND2 I2286 (gtint_5n[33], gate_0n[5], itint_5n[33]);
  AND2 I2287 (gtint_5n[34], gate_0n[5], itint_5n[34]);
  AND2 I2288 (gtint_6n[0], gate_0n[6], itint_6n[0]);
  AND2 I2289 (gtint_6n[1], gate_0n[6], itint_6n[1]);
  AND2 I2290 (gtint_6n[2], gate_0n[6], itint_6n[2]);
  AND2 I2291 (gtint_6n[3], gate_0n[6], itint_6n[3]);
  AND2 I2292 (gtint_6n[4], gate_0n[6], itint_6n[4]);
  AND2 I2293 (gtint_6n[5], gate_0n[6], itint_6n[5]);
  AND2 I2294 (gtint_6n[6], gate_0n[6], itint_6n[6]);
  AND2 I2295 (gtint_6n[7], gate_0n[6], itint_6n[7]);
  AND2 I2296 (gtint_6n[8], gate_0n[6], itint_6n[8]);
  AND2 I2297 (gtint_6n[9], gate_0n[6], itint_6n[9]);
  AND2 I2298 (gtint_6n[10], gate_0n[6], itint_6n[10]);
  AND2 I2299 (gtint_6n[11], gate_0n[6], itint_6n[11]);
  AND2 I2300 (gtint_6n[12], gate_0n[6], itint_6n[12]);
  AND2 I2301 (gtint_6n[13], gate_0n[6], itint_6n[13]);
  AND2 I2302 (gtint_6n[14], gate_0n[6], itint_6n[14]);
  AND2 I2303 (gtint_6n[15], gate_0n[6], itint_6n[15]);
  AND2 I2304 (gtint_6n[16], gate_0n[6], itint_6n[16]);
  AND2 I2305 (gtint_6n[17], gate_0n[6], itint_6n[17]);
  AND2 I2306 (gtint_6n[18], gate_0n[6], itint_6n[18]);
  AND2 I2307 (gtint_6n[19], gate_0n[6], itint_6n[19]);
  AND2 I2308 (gtint_6n[20], gate_0n[6], itint_6n[20]);
  AND2 I2309 (gtint_6n[21], gate_0n[6], itint_6n[21]);
  AND2 I2310 (gtint_6n[22], gate_0n[6], itint_6n[22]);
  AND2 I2311 (gtint_6n[23], gate_0n[6], itint_6n[23]);
  AND2 I2312 (gtint_6n[24], gate_0n[6], itint_6n[24]);
  AND2 I2313 (gtint_6n[25], gate_0n[6], itint_6n[25]);
  AND2 I2314 (gtint_6n[26], gate_0n[6], itint_6n[26]);
  AND2 I2315 (gtint_6n[27], gate_0n[6], itint_6n[27]);
  AND2 I2316 (gtint_6n[28], gate_0n[6], itint_6n[28]);
  AND2 I2317 (gtint_6n[29], gate_0n[6], itint_6n[29]);
  AND2 I2318 (gtint_6n[30], gate_0n[6], itint_6n[30]);
  AND2 I2319 (gtint_6n[31], gate_0n[6], itint_6n[31]);
  AND2 I2320 (gtint_6n[32], gate_0n[6], itint_6n[32]);
  AND2 I2321 (gtint_6n[33], gate_0n[6], itint_6n[33]);
  AND2 I2322 (gtint_6n[34], gate_0n[6], itint_6n[34]);
  AND2 I2323 (gtint_7n[0], gate_0n[7], itint_7n[0]);
  AND2 I2324 (gtint_7n[1], gate_0n[7], itint_7n[1]);
  AND2 I2325 (gtint_7n[2], gate_0n[7], itint_7n[2]);
  AND2 I2326 (gtint_7n[3], gate_0n[7], itint_7n[3]);
  AND2 I2327 (gtint_7n[4], gate_0n[7], itint_7n[4]);
  AND2 I2328 (gtint_7n[5], gate_0n[7], itint_7n[5]);
  AND2 I2329 (gtint_7n[6], gate_0n[7], itint_7n[6]);
  AND2 I2330 (gtint_7n[7], gate_0n[7], itint_7n[7]);
  AND2 I2331 (gtint_7n[8], gate_0n[7], itint_7n[8]);
  AND2 I2332 (gtint_7n[9], gate_0n[7], itint_7n[9]);
  AND2 I2333 (gtint_7n[10], gate_0n[7], itint_7n[10]);
  AND2 I2334 (gtint_7n[11], gate_0n[7], itint_7n[11]);
  AND2 I2335 (gtint_7n[12], gate_0n[7], itint_7n[12]);
  AND2 I2336 (gtint_7n[13], gate_0n[7], itint_7n[13]);
  AND2 I2337 (gtint_7n[14], gate_0n[7], itint_7n[14]);
  AND2 I2338 (gtint_7n[15], gate_0n[7], itint_7n[15]);
  AND2 I2339 (gtint_7n[16], gate_0n[7], itint_7n[16]);
  AND2 I2340 (gtint_7n[17], gate_0n[7], itint_7n[17]);
  AND2 I2341 (gtint_7n[18], gate_0n[7], itint_7n[18]);
  AND2 I2342 (gtint_7n[19], gate_0n[7], itint_7n[19]);
  AND2 I2343 (gtint_7n[20], gate_0n[7], itint_7n[20]);
  AND2 I2344 (gtint_7n[21], gate_0n[7], itint_7n[21]);
  AND2 I2345 (gtint_7n[22], gate_0n[7], itint_7n[22]);
  AND2 I2346 (gtint_7n[23], gate_0n[7], itint_7n[23]);
  AND2 I2347 (gtint_7n[24], gate_0n[7], itint_7n[24]);
  AND2 I2348 (gtint_7n[25], gate_0n[7], itint_7n[25]);
  AND2 I2349 (gtint_7n[26], gate_0n[7], itint_7n[26]);
  AND2 I2350 (gtint_7n[27], gate_0n[7], itint_7n[27]);
  AND2 I2351 (gtint_7n[28], gate_0n[7], itint_7n[28]);
  AND2 I2352 (gtint_7n[29], gate_0n[7], itint_7n[29]);
  AND2 I2353 (gtint_7n[30], gate_0n[7], itint_7n[30]);
  AND2 I2354 (gtint_7n[31], gate_0n[7], itint_7n[31]);
  AND2 I2355 (gtint_7n[32], gate_0n[7], itint_7n[32]);
  AND2 I2356 (gtint_7n[33], gate_0n[7], itint_7n[33]);
  AND2 I2357 (gtint_7n[34], gate_0n[7], itint_7n[34]);
  AND2 I2358 (gtint_8n[0], gate_0n[8], itint_8n[0]);
  AND2 I2359 (gtint_8n[1], gate_0n[8], itint_8n[1]);
  AND2 I2360 (gtint_8n[2], gate_0n[8], itint_8n[2]);
  AND2 I2361 (gtint_8n[3], gate_0n[8], itint_8n[3]);
  AND2 I2362 (gtint_8n[4], gate_0n[8], itint_8n[4]);
  AND2 I2363 (gtint_8n[5], gate_0n[8], itint_8n[5]);
  AND2 I2364 (gtint_8n[6], gate_0n[8], itint_8n[6]);
  AND2 I2365 (gtint_8n[7], gate_0n[8], itint_8n[7]);
  AND2 I2366 (gtint_8n[8], gate_0n[8], itint_8n[8]);
  AND2 I2367 (gtint_8n[9], gate_0n[8], itint_8n[9]);
  AND2 I2368 (gtint_8n[10], gate_0n[8], itint_8n[10]);
  AND2 I2369 (gtint_8n[11], gate_0n[8], itint_8n[11]);
  AND2 I2370 (gtint_8n[12], gate_0n[8], itint_8n[12]);
  AND2 I2371 (gtint_8n[13], gate_0n[8], itint_8n[13]);
  AND2 I2372 (gtint_8n[14], gate_0n[8], itint_8n[14]);
  AND2 I2373 (gtint_8n[15], gate_0n[8], itint_8n[15]);
  AND2 I2374 (gtint_8n[16], gate_0n[8], itint_8n[16]);
  AND2 I2375 (gtint_8n[17], gate_0n[8], itint_8n[17]);
  AND2 I2376 (gtint_8n[18], gate_0n[8], itint_8n[18]);
  AND2 I2377 (gtint_8n[19], gate_0n[8], itint_8n[19]);
  AND2 I2378 (gtint_8n[20], gate_0n[8], itint_8n[20]);
  AND2 I2379 (gtint_8n[21], gate_0n[8], itint_8n[21]);
  AND2 I2380 (gtint_8n[22], gate_0n[8], itint_8n[22]);
  AND2 I2381 (gtint_8n[23], gate_0n[8], itint_8n[23]);
  AND2 I2382 (gtint_8n[24], gate_0n[8], itint_8n[24]);
  AND2 I2383 (gtint_8n[25], gate_0n[8], itint_8n[25]);
  AND2 I2384 (gtint_8n[26], gate_0n[8], itint_8n[26]);
  AND2 I2385 (gtint_8n[27], gate_0n[8], itint_8n[27]);
  AND2 I2386 (gtint_8n[28], gate_0n[8], itint_8n[28]);
  AND2 I2387 (gtint_8n[29], gate_0n[8], itint_8n[29]);
  AND2 I2388 (gtint_8n[30], gate_0n[8], itint_8n[30]);
  AND2 I2389 (gtint_8n[31], gate_0n[8], itint_8n[31]);
  AND2 I2390 (gtint_8n[32], gate_0n[8], itint_8n[32]);
  AND2 I2391 (gtint_8n[33], gate_0n[8], itint_8n[33]);
  AND2 I2392 (gtint_8n[34], gate_0n[8], itint_8n[34]);
  NOR3 I2393 (internal_0n[342], gtint_0n[0], gtint_1n[0], gtint_2n[0]);
  NOR3 I2394 (internal_0n[343], gtint_3n[0], gtint_4n[0], gtint_5n[0]);
  NOR3 I2395 (internal_0n[344], gtint_6n[0], gtint_7n[0], gtint_8n[0]);
  NAND3 I2396 (otint_0n[0], internal_0n[342], internal_0n[343], internal_0n[344]);
  NOR3 I2397 (internal_0n[345], gtint_0n[1], gtint_1n[1], gtint_2n[1]);
  NOR3 I2398 (internal_0n[346], gtint_3n[1], gtint_4n[1], gtint_5n[1]);
  NOR3 I2399 (internal_0n[347], gtint_6n[1], gtint_7n[1], gtint_8n[1]);
  NAND3 I2400 (otint_0n[1], internal_0n[345], internal_0n[346], internal_0n[347]);
  NOR3 I2401 (internal_0n[348], gtint_0n[2], gtint_1n[2], gtint_2n[2]);
  NOR3 I2402 (internal_0n[349], gtint_3n[2], gtint_4n[2], gtint_5n[2]);
  NOR3 I2403 (internal_0n[350], gtint_6n[2], gtint_7n[2], gtint_8n[2]);
  NAND3 I2404 (otint_0n[2], internal_0n[348], internal_0n[349], internal_0n[350]);
  NOR3 I2405 (internal_0n[351], gtint_0n[3], gtint_1n[3], gtint_2n[3]);
  NOR3 I2406 (internal_0n[352], gtint_3n[3], gtint_4n[3], gtint_5n[3]);
  NOR3 I2407 (internal_0n[353], gtint_6n[3], gtint_7n[3], gtint_8n[3]);
  NAND3 I2408 (otint_0n[3], internal_0n[351], internal_0n[352], internal_0n[353]);
  NOR3 I2409 (internal_0n[354], gtint_0n[4], gtint_1n[4], gtint_2n[4]);
  NOR3 I2410 (internal_0n[355], gtint_3n[4], gtint_4n[4], gtint_5n[4]);
  NOR3 I2411 (internal_0n[356], gtint_6n[4], gtint_7n[4], gtint_8n[4]);
  NAND3 I2412 (otint_0n[4], internal_0n[354], internal_0n[355], internal_0n[356]);
  NOR3 I2413 (internal_0n[357], gtint_0n[5], gtint_1n[5], gtint_2n[5]);
  NOR3 I2414 (internal_0n[358], gtint_3n[5], gtint_4n[5], gtint_5n[5]);
  NOR3 I2415 (internal_0n[359], gtint_6n[5], gtint_7n[5], gtint_8n[5]);
  NAND3 I2416 (otint_0n[5], internal_0n[357], internal_0n[358], internal_0n[359]);
  NOR3 I2417 (internal_0n[360], gtint_0n[6], gtint_1n[6], gtint_2n[6]);
  NOR3 I2418 (internal_0n[361], gtint_3n[6], gtint_4n[6], gtint_5n[6]);
  NOR3 I2419 (internal_0n[362], gtint_6n[6], gtint_7n[6], gtint_8n[6]);
  NAND3 I2420 (otint_0n[6], internal_0n[360], internal_0n[361], internal_0n[362]);
  NOR3 I2421 (internal_0n[363], gtint_0n[7], gtint_1n[7], gtint_2n[7]);
  NOR3 I2422 (internal_0n[364], gtint_3n[7], gtint_4n[7], gtint_5n[7]);
  NOR3 I2423 (internal_0n[365], gtint_6n[7], gtint_7n[7], gtint_8n[7]);
  NAND3 I2424 (otint_0n[7], internal_0n[363], internal_0n[364], internal_0n[365]);
  NOR3 I2425 (internal_0n[366], gtint_0n[8], gtint_1n[8], gtint_2n[8]);
  NOR3 I2426 (internal_0n[367], gtint_3n[8], gtint_4n[8], gtint_5n[8]);
  NOR3 I2427 (internal_0n[368], gtint_6n[8], gtint_7n[8], gtint_8n[8]);
  NAND3 I2428 (otint_0n[8], internal_0n[366], internal_0n[367], internal_0n[368]);
  NOR3 I2429 (internal_0n[369], gtint_0n[9], gtint_1n[9], gtint_2n[9]);
  NOR3 I2430 (internal_0n[370], gtint_3n[9], gtint_4n[9], gtint_5n[9]);
  NOR3 I2431 (internal_0n[371], gtint_6n[9], gtint_7n[9], gtint_8n[9]);
  NAND3 I2432 (otint_0n[9], internal_0n[369], internal_0n[370], internal_0n[371]);
  NOR3 I2433 (internal_0n[372], gtint_0n[10], gtint_1n[10], gtint_2n[10]);
  NOR3 I2434 (internal_0n[373], gtint_3n[10], gtint_4n[10], gtint_5n[10]);
  NOR3 I2435 (internal_0n[374], gtint_6n[10], gtint_7n[10], gtint_8n[10]);
  NAND3 I2436 (otint_0n[10], internal_0n[372], internal_0n[373], internal_0n[374]);
  NOR3 I2437 (internal_0n[375], gtint_0n[11], gtint_1n[11], gtint_2n[11]);
  NOR3 I2438 (internal_0n[376], gtint_3n[11], gtint_4n[11], gtint_5n[11]);
  NOR3 I2439 (internal_0n[377], gtint_6n[11], gtint_7n[11], gtint_8n[11]);
  NAND3 I2440 (otint_0n[11], internal_0n[375], internal_0n[376], internal_0n[377]);
  NOR3 I2441 (internal_0n[378], gtint_0n[12], gtint_1n[12], gtint_2n[12]);
  NOR3 I2442 (internal_0n[379], gtint_3n[12], gtint_4n[12], gtint_5n[12]);
  NOR3 I2443 (internal_0n[380], gtint_6n[12], gtint_7n[12], gtint_8n[12]);
  NAND3 I2444 (otint_0n[12], internal_0n[378], internal_0n[379], internal_0n[380]);
  NOR3 I2445 (internal_0n[381], gtint_0n[13], gtint_1n[13], gtint_2n[13]);
  NOR3 I2446 (internal_0n[382], gtint_3n[13], gtint_4n[13], gtint_5n[13]);
  NOR3 I2447 (internal_0n[383], gtint_6n[13], gtint_7n[13], gtint_8n[13]);
  NAND3 I2448 (otint_0n[13], internal_0n[381], internal_0n[382], internal_0n[383]);
  NOR3 I2449 (internal_0n[384], gtint_0n[14], gtint_1n[14], gtint_2n[14]);
  NOR3 I2450 (internal_0n[385], gtint_3n[14], gtint_4n[14], gtint_5n[14]);
  NOR3 I2451 (internal_0n[386], gtint_6n[14], gtint_7n[14], gtint_8n[14]);
  NAND3 I2452 (otint_0n[14], internal_0n[384], internal_0n[385], internal_0n[386]);
  NOR3 I2453 (internal_0n[387], gtint_0n[15], gtint_1n[15], gtint_2n[15]);
  NOR3 I2454 (internal_0n[388], gtint_3n[15], gtint_4n[15], gtint_5n[15]);
  NOR3 I2455 (internal_0n[389], gtint_6n[15], gtint_7n[15], gtint_8n[15]);
  NAND3 I2456 (otint_0n[15], internal_0n[387], internal_0n[388], internal_0n[389]);
  NOR3 I2457 (internal_0n[390], gtint_0n[16], gtint_1n[16], gtint_2n[16]);
  NOR3 I2458 (internal_0n[391], gtint_3n[16], gtint_4n[16], gtint_5n[16]);
  NOR3 I2459 (internal_0n[392], gtint_6n[16], gtint_7n[16], gtint_8n[16]);
  NAND3 I2460 (otint_0n[16], internal_0n[390], internal_0n[391], internal_0n[392]);
  NOR3 I2461 (internal_0n[393], gtint_0n[17], gtint_1n[17], gtint_2n[17]);
  NOR3 I2462 (internal_0n[394], gtint_3n[17], gtint_4n[17], gtint_5n[17]);
  NOR3 I2463 (internal_0n[395], gtint_6n[17], gtint_7n[17], gtint_8n[17]);
  NAND3 I2464 (otint_0n[17], internal_0n[393], internal_0n[394], internal_0n[395]);
  NOR3 I2465 (internal_0n[396], gtint_0n[18], gtint_1n[18], gtint_2n[18]);
  NOR3 I2466 (internal_0n[397], gtint_3n[18], gtint_4n[18], gtint_5n[18]);
  NOR3 I2467 (internal_0n[398], gtint_6n[18], gtint_7n[18], gtint_8n[18]);
  NAND3 I2468 (otint_0n[18], internal_0n[396], internal_0n[397], internal_0n[398]);
  NOR3 I2469 (internal_0n[399], gtint_0n[19], gtint_1n[19], gtint_2n[19]);
  NOR3 I2470 (internal_0n[400], gtint_3n[19], gtint_4n[19], gtint_5n[19]);
  NOR3 I2471 (internal_0n[401], gtint_6n[19], gtint_7n[19], gtint_8n[19]);
  NAND3 I2472 (otint_0n[19], internal_0n[399], internal_0n[400], internal_0n[401]);
  NOR3 I2473 (internal_0n[402], gtint_0n[20], gtint_1n[20], gtint_2n[20]);
  NOR3 I2474 (internal_0n[403], gtint_3n[20], gtint_4n[20], gtint_5n[20]);
  NOR3 I2475 (internal_0n[404], gtint_6n[20], gtint_7n[20], gtint_8n[20]);
  NAND3 I2476 (otint_0n[20], internal_0n[402], internal_0n[403], internal_0n[404]);
  NOR3 I2477 (internal_0n[405], gtint_0n[21], gtint_1n[21], gtint_2n[21]);
  NOR3 I2478 (internal_0n[406], gtint_3n[21], gtint_4n[21], gtint_5n[21]);
  NOR3 I2479 (internal_0n[407], gtint_6n[21], gtint_7n[21], gtint_8n[21]);
  NAND3 I2480 (otint_0n[21], internal_0n[405], internal_0n[406], internal_0n[407]);
  NOR3 I2481 (internal_0n[408], gtint_0n[22], gtint_1n[22], gtint_2n[22]);
  NOR3 I2482 (internal_0n[409], gtint_3n[22], gtint_4n[22], gtint_5n[22]);
  NOR3 I2483 (internal_0n[410], gtint_6n[22], gtint_7n[22], gtint_8n[22]);
  NAND3 I2484 (otint_0n[22], internal_0n[408], internal_0n[409], internal_0n[410]);
  NOR3 I2485 (internal_0n[411], gtint_0n[23], gtint_1n[23], gtint_2n[23]);
  NOR3 I2486 (internal_0n[412], gtint_3n[23], gtint_4n[23], gtint_5n[23]);
  NOR3 I2487 (internal_0n[413], gtint_6n[23], gtint_7n[23], gtint_8n[23]);
  NAND3 I2488 (otint_0n[23], internal_0n[411], internal_0n[412], internal_0n[413]);
  NOR3 I2489 (internal_0n[414], gtint_0n[24], gtint_1n[24], gtint_2n[24]);
  NOR3 I2490 (internal_0n[415], gtint_3n[24], gtint_4n[24], gtint_5n[24]);
  NOR3 I2491 (internal_0n[416], gtint_6n[24], gtint_7n[24], gtint_8n[24]);
  NAND3 I2492 (otint_0n[24], internal_0n[414], internal_0n[415], internal_0n[416]);
  NOR3 I2493 (internal_0n[417], gtint_0n[25], gtint_1n[25], gtint_2n[25]);
  NOR3 I2494 (internal_0n[418], gtint_3n[25], gtint_4n[25], gtint_5n[25]);
  NOR3 I2495 (internal_0n[419], gtint_6n[25], gtint_7n[25], gtint_8n[25]);
  NAND3 I2496 (otint_0n[25], internal_0n[417], internal_0n[418], internal_0n[419]);
  NOR3 I2497 (internal_0n[420], gtint_0n[26], gtint_1n[26], gtint_2n[26]);
  NOR3 I2498 (internal_0n[421], gtint_3n[26], gtint_4n[26], gtint_5n[26]);
  NOR3 I2499 (internal_0n[422], gtint_6n[26], gtint_7n[26], gtint_8n[26]);
  NAND3 I2500 (otint_0n[26], internal_0n[420], internal_0n[421], internal_0n[422]);
  NOR3 I2501 (internal_0n[423], gtint_0n[27], gtint_1n[27], gtint_2n[27]);
  NOR3 I2502 (internal_0n[424], gtint_3n[27], gtint_4n[27], gtint_5n[27]);
  NOR3 I2503 (internal_0n[425], gtint_6n[27], gtint_7n[27], gtint_8n[27]);
  NAND3 I2504 (otint_0n[27], internal_0n[423], internal_0n[424], internal_0n[425]);
  NOR3 I2505 (internal_0n[426], gtint_0n[28], gtint_1n[28], gtint_2n[28]);
  NOR3 I2506 (internal_0n[427], gtint_3n[28], gtint_4n[28], gtint_5n[28]);
  NOR3 I2507 (internal_0n[428], gtint_6n[28], gtint_7n[28], gtint_8n[28]);
  NAND3 I2508 (otint_0n[28], internal_0n[426], internal_0n[427], internal_0n[428]);
  NOR3 I2509 (internal_0n[429], gtint_0n[29], gtint_1n[29], gtint_2n[29]);
  NOR3 I2510 (internal_0n[430], gtint_3n[29], gtint_4n[29], gtint_5n[29]);
  NOR3 I2511 (internal_0n[431], gtint_6n[29], gtint_7n[29], gtint_8n[29]);
  NAND3 I2512 (otint_0n[29], internal_0n[429], internal_0n[430], internal_0n[431]);
  NOR3 I2513 (internal_0n[432], gtint_0n[30], gtint_1n[30], gtint_2n[30]);
  NOR3 I2514 (internal_0n[433], gtint_3n[30], gtint_4n[30], gtint_5n[30]);
  NOR3 I2515 (internal_0n[434], gtint_6n[30], gtint_7n[30], gtint_8n[30]);
  NAND3 I2516 (otint_0n[30], internal_0n[432], internal_0n[433], internal_0n[434]);
  NOR3 I2517 (internal_0n[435], gtint_0n[31], gtint_1n[31], gtint_2n[31]);
  NOR3 I2518 (internal_0n[436], gtint_3n[31], gtint_4n[31], gtint_5n[31]);
  NOR3 I2519 (internal_0n[437], gtint_6n[31], gtint_7n[31], gtint_8n[31]);
  NAND3 I2520 (otint_0n[31], internal_0n[435], internal_0n[436], internal_0n[437]);
  NOR3 I2521 (internal_0n[438], gtint_0n[32], gtint_1n[32], gtint_2n[32]);
  NOR3 I2522 (internal_0n[439], gtint_3n[32], gtint_4n[32], gtint_5n[32]);
  NOR3 I2523 (internal_0n[440], gtint_6n[32], gtint_7n[32], gtint_8n[32]);
  NAND3 I2524 (otint_0n[32], internal_0n[438], internal_0n[439], internal_0n[440]);
  NOR3 I2525 (internal_0n[441], gtint_0n[33], gtint_1n[33], gtint_2n[33]);
  NOR3 I2526 (internal_0n[442], gtint_3n[33], gtint_4n[33], gtint_5n[33]);
  NOR3 I2527 (internal_0n[443], gtint_6n[33], gtint_7n[33], gtint_8n[33]);
  NAND3 I2528 (otint_0n[33], internal_0n[441], internal_0n[442], internal_0n[443]);
  NOR3 I2529 (internal_0n[444], gtint_0n[34], gtint_1n[34], gtint_2n[34]);
  NOR3 I2530 (internal_0n[445], gtint_3n[34], gtint_4n[34], gtint_5n[34]);
  NOR3 I2531 (internal_0n[446], gtint_6n[34], gtint_7n[34], gtint_8n[34]);
  NAND3 I2532 (otint_0n[34], internal_0n[444], internal_0n[445], internal_0n[446]);
  NOR3 I2533 (internal_0n[447], gfint_0n[0], gfint_1n[0], gfint_2n[0]);
  NOR3 I2534 (internal_0n[448], gfint_3n[0], gfint_4n[0], gfint_5n[0]);
  NOR3 I2535 (internal_0n[449], gfint_6n[0], gfint_7n[0], gfint_8n[0]);
  NAND3 I2536 (ofint_0n[0], internal_0n[447], internal_0n[448], internal_0n[449]);
  NOR3 I2537 (internal_0n[450], gfint_0n[1], gfint_1n[1], gfint_2n[1]);
  NOR3 I2538 (internal_0n[451], gfint_3n[1], gfint_4n[1], gfint_5n[1]);
  NOR3 I2539 (internal_0n[452], gfint_6n[1], gfint_7n[1], gfint_8n[1]);
  NAND3 I2540 (ofint_0n[1], internal_0n[450], internal_0n[451], internal_0n[452]);
  NOR3 I2541 (internal_0n[453], gfint_0n[2], gfint_1n[2], gfint_2n[2]);
  NOR3 I2542 (internal_0n[454], gfint_3n[2], gfint_4n[2], gfint_5n[2]);
  NOR3 I2543 (internal_0n[455], gfint_6n[2], gfint_7n[2], gfint_8n[2]);
  NAND3 I2544 (ofint_0n[2], internal_0n[453], internal_0n[454], internal_0n[455]);
  NOR3 I2545 (internal_0n[456], gfint_0n[3], gfint_1n[3], gfint_2n[3]);
  NOR3 I2546 (internal_0n[457], gfint_3n[3], gfint_4n[3], gfint_5n[3]);
  NOR3 I2547 (internal_0n[458], gfint_6n[3], gfint_7n[3], gfint_8n[3]);
  NAND3 I2548 (ofint_0n[3], internal_0n[456], internal_0n[457], internal_0n[458]);
  NOR3 I2549 (internal_0n[459], gfint_0n[4], gfint_1n[4], gfint_2n[4]);
  NOR3 I2550 (internal_0n[460], gfint_3n[4], gfint_4n[4], gfint_5n[4]);
  NOR3 I2551 (internal_0n[461], gfint_6n[4], gfint_7n[4], gfint_8n[4]);
  NAND3 I2552 (ofint_0n[4], internal_0n[459], internal_0n[460], internal_0n[461]);
  NOR3 I2553 (internal_0n[462], gfint_0n[5], gfint_1n[5], gfint_2n[5]);
  NOR3 I2554 (internal_0n[463], gfint_3n[5], gfint_4n[5], gfint_5n[5]);
  NOR3 I2555 (internal_0n[464], gfint_6n[5], gfint_7n[5], gfint_8n[5]);
  NAND3 I2556 (ofint_0n[5], internal_0n[462], internal_0n[463], internal_0n[464]);
  NOR3 I2557 (internal_0n[465], gfint_0n[6], gfint_1n[6], gfint_2n[6]);
  NOR3 I2558 (internal_0n[466], gfint_3n[6], gfint_4n[6], gfint_5n[6]);
  NOR3 I2559 (internal_0n[467], gfint_6n[6], gfint_7n[6], gfint_8n[6]);
  NAND3 I2560 (ofint_0n[6], internal_0n[465], internal_0n[466], internal_0n[467]);
  NOR3 I2561 (internal_0n[468], gfint_0n[7], gfint_1n[7], gfint_2n[7]);
  NOR3 I2562 (internal_0n[469], gfint_3n[7], gfint_4n[7], gfint_5n[7]);
  NOR3 I2563 (internal_0n[470], gfint_6n[7], gfint_7n[7], gfint_8n[7]);
  NAND3 I2564 (ofint_0n[7], internal_0n[468], internal_0n[469], internal_0n[470]);
  NOR3 I2565 (internal_0n[471], gfint_0n[8], gfint_1n[8], gfint_2n[8]);
  NOR3 I2566 (internal_0n[472], gfint_3n[8], gfint_4n[8], gfint_5n[8]);
  NOR3 I2567 (internal_0n[473], gfint_6n[8], gfint_7n[8], gfint_8n[8]);
  NAND3 I2568 (ofint_0n[8], internal_0n[471], internal_0n[472], internal_0n[473]);
  NOR3 I2569 (internal_0n[474], gfint_0n[9], gfint_1n[9], gfint_2n[9]);
  NOR3 I2570 (internal_0n[475], gfint_3n[9], gfint_4n[9], gfint_5n[9]);
  NOR3 I2571 (internal_0n[476], gfint_6n[9], gfint_7n[9], gfint_8n[9]);
  NAND3 I2572 (ofint_0n[9], internal_0n[474], internal_0n[475], internal_0n[476]);
  NOR3 I2573 (internal_0n[477], gfint_0n[10], gfint_1n[10], gfint_2n[10]);
  NOR3 I2574 (internal_0n[478], gfint_3n[10], gfint_4n[10], gfint_5n[10]);
  NOR3 I2575 (internal_0n[479], gfint_6n[10], gfint_7n[10], gfint_8n[10]);
  NAND3 I2576 (ofint_0n[10], internal_0n[477], internal_0n[478], internal_0n[479]);
  NOR3 I2577 (internal_0n[480], gfint_0n[11], gfint_1n[11], gfint_2n[11]);
  NOR3 I2578 (internal_0n[481], gfint_3n[11], gfint_4n[11], gfint_5n[11]);
  NOR3 I2579 (internal_0n[482], gfint_6n[11], gfint_7n[11], gfint_8n[11]);
  NAND3 I2580 (ofint_0n[11], internal_0n[480], internal_0n[481], internal_0n[482]);
  NOR3 I2581 (internal_0n[483], gfint_0n[12], gfint_1n[12], gfint_2n[12]);
  NOR3 I2582 (internal_0n[484], gfint_3n[12], gfint_4n[12], gfint_5n[12]);
  NOR3 I2583 (internal_0n[485], gfint_6n[12], gfint_7n[12], gfint_8n[12]);
  NAND3 I2584 (ofint_0n[12], internal_0n[483], internal_0n[484], internal_0n[485]);
  NOR3 I2585 (internal_0n[486], gfint_0n[13], gfint_1n[13], gfint_2n[13]);
  NOR3 I2586 (internal_0n[487], gfint_3n[13], gfint_4n[13], gfint_5n[13]);
  NOR3 I2587 (internal_0n[488], gfint_6n[13], gfint_7n[13], gfint_8n[13]);
  NAND3 I2588 (ofint_0n[13], internal_0n[486], internal_0n[487], internal_0n[488]);
  NOR3 I2589 (internal_0n[489], gfint_0n[14], gfint_1n[14], gfint_2n[14]);
  NOR3 I2590 (internal_0n[490], gfint_3n[14], gfint_4n[14], gfint_5n[14]);
  NOR3 I2591 (internal_0n[491], gfint_6n[14], gfint_7n[14], gfint_8n[14]);
  NAND3 I2592 (ofint_0n[14], internal_0n[489], internal_0n[490], internal_0n[491]);
  NOR3 I2593 (internal_0n[492], gfint_0n[15], gfint_1n[15], gfint_2n[15]);
  NOR3 I2594 (internal_0n[493], gfint_3n[15], gfint_4n[15], gfint_5n[15]);
  NOR3 I2595 (internal_0n[494], gfint_6n[15], gfint_7n[15], gfint_8n[15]);
  NAND3 I2596 (ofint_0n[15], internal_0n[492], internal_0n[493], internal_0n[494]);
  NOR3 I2597 (internal_0n[495], gfint_0n[16], gfint_1n[16], gfint_2n[16]);
  NOR3 I2598 (internal_0n[496], gfint_3n[16], gfint_4n[16], gfint_5n[16]);
  NOR3 I2599 (internal_0n[497], gfint_6n[16], gfint_7n[16], gfint_8n[16]);
  NAND3 I2600 (ofint_0n[16], internal_0n[495], internal_0n[496], internal_0n[497]);
  NOR3 I2601 (internal_0n[498], gfint_0n[17], gfint_1n[17], gfint_2n[17]);
  NOR3 I2602 (internal_0n[499], gfint_3n[17], gfint_4n[17], gfint_5n[17]);
  NOR3 I2603 (internal_0n[500], gfint_6n[17], gfint_7n[17], gfint_8n[17]);
  NAND3 I2604 (ofint_0n[17], internal_0n[498], internal_0n[499], internal_0n[500]);
  NOR3 I2605 (internal_0n[501], gfint_0n[18], gfint_1n[18], gfint_2n[18]);
  NOR3 I2606 (internal_0n[502], gfint_3n[18], gfint_4n[18], gfint_5n[18]);
  NOR3 I2607 (internal_0n[503], gfint_6n[18], gfint_7n[18], gfint_8n[18]);
  NAND3 I2608 (ofint_0n[18], internal_0n[501], internal_0n[502], internal_0n[503]);
  NOR3 I2609 (internal_0n[504], gfint_0n[19], gfint_1n[19], gfint_2n[19]);
  NOR3 I2610 (internal_0n[505], gfint_3n[19], gfint_4n[19], gfint_5n[19]);
  NOR3 I2611 (internal_0n[506], gfint_6n[19], gfint_7n[19], gfint_8n[19]);
  NAND3 I2612 (ofint_0n[19], internal_0n[504], internal_0n[505], internal_0n[506]);
  NOR3 I2613 (internal_0n[507], gfint_0n[20], gfint_1n[20], gfint_2n[20]);
  NOR3 I2614 (internal_0n[508], gfint_3n[20], gfint_4n[20], gfint_5n[20]);
  NOR3 I2615 (internal_0n[509], gfint_6n[20], gfint_7n[20], gfint_8n[20]);
  NAND3 I2616 (ofint_0n[20], internal_0n[507], internal_0n[508], internal_0n[509]);
  NOR3 I2617 (internal_0n[510], gfint_0n[21], gfint_1n[21], gfint_2n[21]);
  NOR3 I2618 (internal_0n[511], gfint_3n[21], gfint_4n[21], gfint_5n[21]);
  NOR3 I2619 (internal_0n[512], gfint_6n[21], gfint_7n[21], gfint_8n[21]);
  NAND3 I2620 (ofint_0n[21], internal_0n[510], internal_0n[511], internal_0n[512]);
  NOR3 I2621 (internal_0n[513], gfint_0n[22], gfint_1n[22], gfint_2n[22]);
  NOR3 I2622 (internal_0n[514], gfint_3n[22], gfint_4n[22], gfint_5n[22]);
  NOR3 I2623 (internal_0n[515], gfint_6n[22], gfint_7n[22], gfint_8n[22]);
  NAND3 I2624 (ofint_0n[22], internal_0n[513], internal_0n[514], internal_0n[515]);
  NOR3 I2625 (internal_0n[516], gfint_0n[23], gfint_1n[23], gfint_2n[23]);
  NOR3 I2626 (internal_0n[517], gfint_3n[23], gfint_4n[23], gfint_5n[23]);
  NOR3 I2627 (internal_0n[518], gfint_6n[23], gfint_7n[23], gfint_8n[23]);
  NAND3 I2628 (ofint_0n[23], internal_0n[516], internal_0n[517], internal_0n[518]);
  NOR3 I2629 (internal_0n[519], gfint_0n[24], gfint_1n[24], gfint_2n[24]);
  NOR3 I2630 (internal_0n[520], gfint_3n[24], gfint_4n[24], gfint_5n[24]);
  NOR3 I2631 (internal_0n[521], gfint_6n[24], gfint_7n[24], gfint_8n[24]);
  NAND3 I2632 (ofint_0n[24], internal_0n[519], internal_0n[520], internal_0n[521]);
  NOR3 I2633 (internal_0n[522], gfint_0n[25], gfint_1n[25], gfint_2n[25]);
  NOR3 I2634 (internal_0n[523], gfint_3n[25], gfint_4n[25], gfint_5n[25]);
  NOR3 I2635 (internal_0n[524], gfint_6n[25], gfint_7n[25], gfint_8n[25]);
  NAND3 I2636 (ofint_0n[25], internal_0n[522], internal_0n[523], internal_0n[524]);
  NOR3 I2637 (internal_0n[525], gfint_0n[26], gfint_1n[26], gfint_2n[26]);
  NOR3 I2638 (internal_0n[526], gfint_3n[26], gfint_4n[26], gfint_5n[26]);
  NOR3 I2639 (internal_0n[527], gfint_6n[26], gfint_7n[26], gfint_8n[26]);
  NAND3 I2640 (ofint_0n[26], internal_0n[525], internal_0n[526], internal_0n[527]);
  NOR3 I2641 (internal_0n[528], gfint_0n[27], gfint_1n[27], gfint_2n[27]);
  NOR3 I2642 (internal_0n[529], gfint_3n[27], gfint_4n[27], gfint_5n[27]);
  NOR3 I2643 (internal_0n[530], gfint_6n[27], gfint_7n[27], gfint_8n[27]);
  NAND3 I2644 (ofint_0n[27], internal_0n[528], internal_0n[529], internal_0n[530]);
  NOR3 I2645 (internal_0n[531], gfint_0n[28], gfint_1n[28], gfint_2n[28]);
  NOR3 I2646 (internal_0n[532], gfint_3n[28], gfint_4n[28], gfint_5n[28]);
  NOR3 I2647 (internal_0n[533], gfint_6n[28], gfint_7n[28], gfint_8n[28]);
  NAND3 I2648 (ofint_0n[28], internal_0n[531], internal_0n[532], internal_0n[533]);
  NOR3 I2649 (internal_0n[534], gfint_0n[29], gfint_1n[29], gfint_2n[29]);
  NOR3 I2650 (internal_0n[535], gfint_3n[29], gfint_4n[29], gfint_5n[29]);
  NOR3 I2651 (internal_0n[536], gfint_6n[29], gfint_7n[29], gfint_8n[29]);
  NAND3 I2652 (ofint_0n[29], internal_0n[534], internal_0n[535], internal_0n[536]);
  NOR3 I2653 (internal_0n[537], gfint_0n[30], gfint_1n[30], gfint_2n[30]);
  NOR3 I2654 (internal_0n[538], gfint_3n[30], gfint_4n[30], gfint_5n[30]);
  NOR3 I2655 (internal_0n[539], gfint_6n[30], gfint_7n[30], gfint_8n[30]);
  NAND3 I2656 (ofint_0n[30], internal_0n[537], internal_0n[538], internal_0n[539]);
  NOR3 I2657 (internal_0n[540], gfint_0n[31], gfint_1n[31], gfint_2n[31]);
  NOR3 I2658 (internal_0n[541], gfint_3n[31], gfint_4n[31], gfint_5n[31]);
  NOR3 I2659 (internal_0n[542], gfint_6n[31], gfint_7n[31], gfint_8n[31]);
  NAND3 I2660 (ofint_0n[31], internal_0n[540], internal_0n[541], internal_0n[542]);
  NOR3 I2661 (internal_0n[543], gfint_0n[32], gfint_1n[32], gfint_2n[32]);
  NOR3 I2662 (internal_0n[544], gfint_3n[32], gfint_4n[32], gfint_5n[32]);
  NOR3 I2663 (internal_0n[545], gfint_6n[32], gfint_7n[32], gfint_8n[32]);
  NAND3 I2664 (ofint_0n[32], internal_0n[543], internal_0n[544], internal_0n[545]);
  NOR3 I2665 (internal_0n[546], gfint_0n[33], gfint_1n[33], gfint_2n[33]);
  NOR3 I2666 (internal_0n[547], gfint_3n[33], gfint_4n[33], gfint_5n[33]);
  NOR3 I2667 (internal_0n[548], gfint_6n[33], gfint_7n[33], gfint_8n[33]);
  NAND3 I2668 (ofint_0n[33], internal_0n[546], internal_0n[547], internal_0n[548]);
  NOR3 I2669 (internal_0n[549], gfint_0n[34], gfint_1n[34], gfint_2n[34]);
  NOR3 I2670 (internal_0n[550], gfint_3n[34], gfint_4n[34], gfint_5n[34]);
  NOR3 I2671 (internal_0n[551], gfint_6n[34], gfint_7n[34], gfint_8n[34]);
  NAND3 I2672 (ofint_0n[34], internal_0n[549], internal_0n[550], internal_0n[551]);
endmodule

module BrzM_36_2 (
  i_0r0d, i_0r1d, i_0a,
  i_1r0d, i_1r1d, i_1a,
  o_0r0d, o_0r1d, o_0a,
  initialise
);
  input [35:0] i_0r0d;
  input [35:0] i_0r1d;
  output i_0a;
  input [35:0] i_1r0d;
  input [35:0] i_1r1d;
  output i_1a;
  output [35:0] o_0r0d;
  output [35:0] o_0r1d;
  input o_0a;
  input initialise;
  wire [89:0] internal_0n;
  wire [1:0] sel_0n;
  wire [35:0] ofint_0n;
  wire [35:0] otint_0n;
  wire oaint_0n;
  wire [35:0] ifint_0n;
  wire [35:0] ifint_1n;
  wire [35:0] itint_0n;
  wire [35:0] itint_1n;
  wire iaint_0n;
  wire iaint_1n;
  wire [1:0] gate_0n;
  wire [35:0] gfint_0n;
  wire [35:0] gfint_1n;
  wire [35:0] gtint_0n;
  wire [35:0] gtint_1n;
  wire [35:0] complete960_0n;
  wire gate959_0n;
  wire [35:0] complete956_0n;
  wire gate955_0n;
  wire [35:0] complete952_0n;
  wire gate951_0n;
  wire [35:0] complete948_0n;
  wire [35:0] complete947_0n;
  wire selcomp_0n;
  wire selcomp_1n;
  C3 I0 (internal_0n[0], complete960_0n[0], complete960_0n[1], complete960_0n[2]);
  C3 I1 (internal_0n[1], complete960_0n[3], complete960_0n[4], complete960_0n[5]);
  C3 I2 (internal_0n[2], complete960_0n[6], complete960_0n[7], complete960_0n[8]);
  C3 I3 (internal_0n[3], complete960_0n[9], complete960_0n[10], complete960_0n[11]);
  C3 I4 (internal_0n[4], complete960_0n[12], complete960_0n[13], complete960_0n[14]);
  C3 I5 (internal_0n[5], complete960_0n[15], complete960_0n[16], complete960_0n[17]);
  C3 I6 (internal_0n[6], complete960_0n[18], complete960_0n[19], complete960_0n[20]);
  C3 I7 (internal_0n[7], complete960_0n[21], complete960_0n[22], complete960_0n[23]);
  C3 I8 (internal_0n[8], complete960_0n[24], complete960_0n[25], complete960_0n[26]);
  C3 I9 (internal_0n[9], complete960_0n[27], complete960_0n[28], complete960_0n[29]);
  C3 I10 (internal_0n[10], complete960_0n[30], complete960_0n[31], complete960_0n[32]);
  C3 I11 (internal_0n[11], complete960_0n[33], complete960_0n[34], complete960_0n[35]);
  C3 I12 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I13 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I14 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I15 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I16 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I17 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I18 (i_1a, internal_0n[16], internal_0n[17]);
  OR2 I19 (complete960_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I20 (complete960_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I21 (complete960_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I22 (complete960_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I23 (complete960_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I24 (complete960_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I25 (complete960_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I26 (complete960_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I27 (complete960_0n[8], ifint_1n[8], itint_1n[8]);
  OR2 I28 (complete960_0n[9], ifint_1n[9], itint_1n[9]);
  OR2 I29 (complete960_0n[10], ifint_1n[10], itint_1n[10]);
  OR2 I30 (complete960_0n[11], ifint_1n[11], itint_1n[11]);
  OR2 I31 (complete960_0n[12], ifint_1n[12], itint_1n[12]);
  OR2 I32 (complete960_0n[13], ifint_1n[13], itint_1n[13]);
  OR2 I33 (complete960_0n[14], ifint_1n[14], itint_1n[14]);
  OR2 I34 (complete960_0n[15], ifint_1n[15], itint_1n[15]);
  OR2 I35 (complete960_0n[16], ifint_1n[16], itint_1n[16]);
  OR2 I36 (complete960_0n[17], ifint_1n[17], itint_1n[17]);
  OR2 I37 (complete960_0n[18], ifint_1n[18], itint_1n[18]);
  OR2 I38 (complete960_0n[19], ifint_1n[19], itint_1n[19]);
  OR2 I39 (complete960_0n[20], ifint_1n[20], itint_1n[20]);
  OR2 I40 (complete960_0n[21], ifint_1n[21], itint_1n[21]);
  OR2 I41 (complete960_0n[22], ifint_1n[22], itint_1n[22]);
  OR2 I42 (complete960_0n[23], ifint_1n[23], itint_1n[23]);
  OR2 I43 (complete960_0n[24], ifint_1n[24], itint_1n[24]);
  OR2 I44 (complete960_0n[25], ifint_1n[25], itint_1n[25]);
  OR2 I45 (complete960_0n[26], ifint_1n[26], itint_1n[26]);
  OR2 I46 (complete960_0n[27], ifint_1n[27], itint_1n[27]);
  OR2 I47 (complete960_0n[28], ifint_1n[28], itint_1n[28]);
  OR2 I48 (complete960_0n[29], ifint_1n[29], itint_1n[29]);
  OR2 I49 (complete960_0n[30], ifint_1n[30], itint_1n[30]);
  OR2 I50 (complete960_0n[31], ifint_1n[31], itint_1n[31]);
  OR2 I51 (complete960_0n[32], ifint_1n[32], itint_1n[32]);
  OR2 I52 (complete960_0n[33], ifint_1n[33], itint_1n[33]);
  OR2 I53 (complete960_0n[34], ifint_1n[34], itint_1n[34]);
  OR2 I54 (complete960_0n[35], ifint_1n[35], itint_1n[35]);
  INV I55 (gate959_0n, iaint_1n);
  C2RI I56 (itint_1n[0], i_1r1d[0], gate959_0n, initialise);
  C2RI I57 (itint_1n[1], i_1r1d[1], gate959_0n, initialise);
  C2RI I58 (itint_1n[2], i_1r1d[2], gate959_0n, initialise);
  C2RI I59 (itint_1n[3], i_1r1d[3], gate959_0n, initialise);
  C2RI I60 (itint_1n[4], i_1r1d[4], gate959_0n, initialise);
  C2RI I61 (itint_1n[5], i_1r1d[5], gate959_0n, initialise);
  C2RI I62 (itint_1n[6], i_1r1d[6], gate959_0n, initialise);
  C2RI I63 (itint_1n[7], i_1r1d[7], gate959_0n, initialise);
  C2RI I64 (itint_1n[8], i_1r1d[8], gate959_0n, initialise);
  C2RI I65 (itint_1n[9], i_1r1d[9], gate959_0n, initialise);
  C2RI I66 (itint_1n[10], i_1r1d[10], gate959_0n, initialise);
  C2RI I67 (itint_1n[11], i_1r1d[11], gate959_0n, initialise);
  C2RI I68 (itint_1n[12], i_1r1d[12], gate959_0n, initialise);
  C2RI I69 (itint_1n[13], i_1r1d[13], gate959_0n, initialise);
  C2RI I70 (itint_1n[14], i_1r1d[14], gate959_0n, initialise);
  C2RI I71 (itint_1n[15], i_1r1d[15], gate959_0n, initialise);
  C2RI I72 (itint_1n[16], i_1r1d[16], gate959_0n, initialise);
  C2RI I73 (itint_1n[17], i_1r1d[17], gate959_0n, initialise);
  C2RI I74 (itint_1n[18], i_1r1d[18], gate959_0n, initialise);
  C2RI I75 (itint_1n[19], i_1r1d[19], gate959_0n, initialise);
  C2RI I76 (itint_1n[20], i_1r1d[20], gate959_0n, initialise);
  C2RI I77 (itint_1n[21], i_1r1d[21], gate959_0n, initialise);
  C2RI I78 (itint_1n[22], i_1r1d[22], gate959_0n, initialise);
  C2RI I79 (itint_1n[23], i_1r1d[23], gate959_0n, initialise);
  C2RI I80 (itint_1n[24], i_1r1d[24], gate959_0n, initialise);
  C2RI I81 (itint_1n[25], i_1r1d[25], gate959_0n, initialise);
  C2RI I82 (itint_1n[26], i_1r1d[26], gate959_0n, initialise);
  C2RI I83 (itint_1n[27], i_1r1d[27], gate959_0n, initialise);
  C2RI I84 (itint_1n[28], i_1r1d[28], gate959_0n, initialise);
  C2RI I85 (itint_1n[29], i_1r1d[29], gate959_0n, initialise);
  C2RI I86 (itint_1n[30], i_1r1d[30], gate959_0n, initialise);
  C2RI I87 (itint_1n[31], i_1r1d[31], gate959_0n, initialise);
  C2RI I88 (itint_1n[32], i_1r1d[32], gate959_0n, initialise);
  C2RI I89 (itint_1n[33], i_1r1d[33], gate959_0n, initialise);
  C2RI I90 (itint_1n[34], i_1r1d[34], gate959_0n, initialise);
  C2RI I91 (itint_1n[35], i_1r1d[35], gate959_0n, initialise);
  C2RI I92 (ifint_1n[0], i_1r0d[0], gate959_0n, initialise);
  C2RI I93 (ifint_1n[1], i_1r0d[1], gate959_0n, initialise);
  C2RI I94 (ifint_1n[2], i_1r0d[2], gate959_0n, initialise);
  C2RI I95 (ifint_1n[3], i_1r0d[3], gate959_0n, initialise);
  C2RI I96 (ifint_1n[4], i_1r0d[4], gate959_0n, initialise);
  C2RI I97 (ifint_1n[5], i_1r0d[5], gate959_0n, initialise);
  C2RI I98 (ifint_1n[6], i_1r0d[6], gate959_0n, initialise);
  C2RI I99 (ifint_1n[7], i_1r0d[7], gate959_0n, initialise);
  C2RI I100 (ifint_1n[8], i_1r0d[8], gate959_0n, initialise);
  C2RI I101 (ifint_1n[9], i_1r0d[9], gate959_0n, initialise);
  C2RI I102 (ifint_1n[10], i_1r0d[10], gate959_0n, initialise);
  C2RI I103 (ifint_1n[11], i_1r0d[11], gate959_0n, initialise);
  C2RI I104 (ifint_1n[12], i_1r0d[12], gate959_0n, initialise);
  C2RI I105 (ifint_1n[13], i_1r0d[13], gate959_0n, initialise);
  C2RI I106 (ifint_1n[14], i_1r0d[14], gate959_0n, initialise);
  C2RI I107 (ifint_1n[15], i_1r0d[15], gate959_0n, initialise);
  C2RI I108 (ifint_1n[16], i_1r0d[16], gate959_0n, initialise);
  C2RI I109 (ifint_1n[17], i_1r0d[17], gate959_0n, initialise);
  C2RI I110 (ifint_1n[18], i_1r0d[18], gate959_0n, initialise);
  C2RI I111 (ifint_1n[19], i_1r0d[19], gate959_0n, initialise);
  C2RI I112 (ifint_1n[20], i_1r0d[20], gate959_0n, initialise);
  C2RI I113 (ifint_1n[21], i_1r0d[21], gate959_0n, initialise);
  C2RI I114 (ifint_1n[22], i_1r0d[22], gate959_0n, initialise);
  C2RI I115 (ifint_1n[23], i_1r0d[23], gate959_0n, initialise);
  C2RI I116 (ifint_1n[24], i_1r0d[24], gate959_0n, initialise);
  C2RI I117 (ifint_1n[25], i_1r0d[25], gate959_0n, initialise);
  C2RI I118 (ifint_1n[26], i_1r0d[26], gate959_0n, initialise);
  C2RI I119 (ifint_1n[27], i_1r0d[27], gate959_0n, initialise);
  C2RI I120 (ifint_1n[28], i_1r0d[28], gate959_0n, initialise);
  C2RI I121 (ifint_1n[29], i_1r0d[29], gate959_0n, initialise);
  C2RI I122 (ifint_1n[30], i_1r0d[30], gate959_0n, initialise);
  C2RI I123 (ifint_1n[31], i_1r0d[31], gate959_0n, initialise);
  C2RI I124 (ifint_1n[32], i_1r0d[32], gate959_0n, initialise);
  C2RI I125 (ifint_1n[33], i_1r0d[33], gate959_0n, initialise);
  C2RI I126 (ifint_1n[34], i_1r0d[34], gate959_0n, initialise);
  C2RI I127 (ifint_1n[35], i_1r0d[35], gate959_0n, initialise);
  C3 I128 (internal_0n[18], complete956_0n[0], complete956_0n[1], complete956_0n[2]);
  C3 I129 (internal_0n[19], complete956_0n[3], complete956_0n[4], complete956_0n[5]);
  C3 I130 (internal_0n[20], complete956_0n[6], complete956_0n[7], complete956_0n[8]);
  C3 I131 (internal_0n[21], complete956_0n[9], complete956_0n[10], complete956_0n[11]);
  C3 I132 (internal_0n[22], complete956_0n[12], complete956_0n[13], complete956_0n[14]);
  C3 I133 (internal_0n[23], complete956_0n[15], complete956_0n[16], complete956_0n[17]);
  C3 I134 (internal_0n[24], complete956_0n[18], complete956_0n[19], complete956_0n[20]);
  C3 I135 (internal_0n[25], complete956_0n[21], complete956_0n[22], complete956_0n[23]);
  C3 I136 (internal_0n[26], complete956_0n[24], complete956_0n[25], complete956_0n[26]);
  C3 I137 (internal_0n[27], complete956_0n[27], complete956_0n[28], complete956_0n[29]);
  C3 I138 (internal_0n[28], complete956_0n[30], complete956_0n[31], complete956_0n[32]);
  C3 I139 (internal_0n[29], complete956_0n[33], complete956_0n[34], complete956_0n[35]);
  C3 I140 (internal_0n[30], internal_0n[18], internal_0n[19], internal_0n[20]);
  C3 I141 (internal_0n[31], internal_0n[21], internal_0n[22], internal_0n[23]);
  C3 I142 (internal_0n[32], internal_0n[24], internal_0n[25], internal_0n[26]);
  C3 I143 (internal_0n[33], internal_0n[27], internal_0n[28], internal_0n[29]);
  C2 I144 (internal_0n[34], internal_0n[30], internal_0n[31]);
  C2 I145 (internal_0n[35], internal_0n[32], internal_0n[33]);
  C2 I146 (i_0a, internal_0n[34], internal_0n[35]);
  OR2 I147 (complete956_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I148 (complete956_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I149 (complete956_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I150 (complete956_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I151 (complete956_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I152 (complete956_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I153 (complete956_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I154 (complete956_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I155 (complete956_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I156 (complete956_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I157 (complete956_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I158 (complete956_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I159 (complete956_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I160 (complete956_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I161 (complete956_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I162 (complete956_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I163 (complete956_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I164 (complete956_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I165 (complete956_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I166 (complete956_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I167 (complete956_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I168 (complete956_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I169 (complete956_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I170 (complete956_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I171 (complete956_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I172 (complete956_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I173 (complete956_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I174 (complete956_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I175 (complete956_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I176 (complete956_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I177 (complete956_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I178 (complete956_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I179 (complete956_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I180 (complete956_0n[33], ifint_0n[33], itint_0n[33]);
  OR2 I181 (complete956_0n[34], ifint_0n[34], itint_0n[34]);
  OR2 I182 (complete956_0n[35], ifint_0n[35], itint_0n[35]);
  INV I183 (gate955_0n, iaint_0n);
  C2RI I184 (itint_0n[0], i_0r1d[0], gate955_0n, initialise);
  C2RI I185 (itint_0n[1], i_0r1d[1], gate955_0n, initialise);
  C2RI I186 (itint_0n[2], i_0r1d[2], gate955_0n, initialise);
  C2RI I187 (itint_0n[3], i_0r1d[3], gate955_0n, initialise);
  C2RI I188 (itint_0n[4], i_0r1d[4], gate955_0n, initialise);
  C2RI I189 (itint_0n[5], i_0r1d[5], gate955_0n, initialise);
  C2RI I190 (itint_0n[6], i_0r1d[6], gate955_0n, initialise);
  C2RI I191 (itint_0n[7], i_0r1d[7], gate955_0n, initialise);
  C2RI I192 (itint_0n[8], i_0r1d[8], gate955_0n, initialise);
  C2RI I193 (itint_0n[9], i_0r1d[9], gate955_0n, initialise);
  C2RI I194 (itint_0n[10], i_0r1d[10], gate955_0n, initialise);
  C2RI I195 (itint_0n[11], i_0r1d[11], gate955_0n, initialise);
  C2RI I196 (itint_0n[12], i_0r1d[12], gate955_0n, initialise);
  C2RI I197 (itint_0n[13], i_0r1d[13], gate955_0n, initialise);
  C2RI I198 (itint_0n[14], i_0r1d[14], gate955_0n, initialise);
  C2RI I199 (itint_0n[15], i_0r1d[15], gate955_0n, initialise);
  C2RI I200 (itint_0n[16], i_0r1d[16], gate955_0n, initialise);
  C2RI I201 (itint_0n[17], i_0r1d[17], gate955_0n, initialise);
  C2RI I202 (itint_0n[18], i_0r1d[18], gate955_0n, initialise);
  C2RI I203 (itint_0n[19], i_0r1d[19], gate955_0n, initialise);
  C2RI I204 (itint_0n[20], i_0r1d[20], gate955_0n, initialise);
  C2RI I205 (itint_0n[21], i_0r1d[21], gate955_0n, initialise);
  C2RI I206 (itint_0n[22], i_0r1d[22], gate955_0n, initialise);
  C2RI I207 (itint_0n[23], i_0r1d[23], gate955_0n, initialise);
  C2RI I208 (itint_0n[24], i_0r1d[24], gate955_0n, initialise);
  C2RI I209 (itint_0n[25], i_0r1d[25], gate955_0n, initialise);
  C2RI I210 (itint_0n[26], i_0r1d[26], gate955_0n, initialise);
  C2RI I211 (itint_0n[27], i_0r1d[27], gate955_0n, initialise);
  C2RI I212 (itint_0n[28], i_0r1d[28], gate955_0n, initialise);
  C2RI I213 (itint_0n[29], i_0r1d[29], gate955_0n, initialise);
  C2RI I214 (itint_0n[30], i_0r1d[30], gate955_0n, initialise);
  C2RI I215 (itint_0n[31], i_0r1d[31], gate955_0n, initialise);
  C2RI I216 (itint_0n[32], i_0r1d[32], gate955_0n, initialise);
  C2RI I217 (itint_0n[33], i_0r1d[33], gate955_0n, initialise);
  C2RI I218 (itint_0n[34], i_0r1d[34], gate955_0n, initialise);
  C2RI I219 (itint_0n[35], i_0r1d[35], gate955_0n, initialise);
  C2RI I220 (ifint_0n[0], i_0r0d[0], gate955_0n, initialise);
  C2RI I221 (ifint_0n[1], i_0r0d[1], gate955_0n, initialise);
  C2RI I222 (ifint_0n[2], i_0r0d[2], gate955_0n, initialise);
  C2RI I223 (ifint_0n[3], i_0r0d[3], gate955_0n, initialise);
  C2RI I224 (ifint_0n[4], i_0r0d[4], gate955_0n, initialise);
  C2RI I225 (ifint_0n[5], i_0r0d[5], gate955_0n, initialise);
  C2RI I226 (ifint_0n[6], i_0r0d[6], gate955_0n, initialise);
  C2RI I227 (ifint_0n[7], i_0r0d[7], gate955_0n, initialise);
  C2RI I228 (ifint_0n[8], i_0r0d[8], gate955_0n, initialise);
  C2RI I229 (ifint_0n[9], i_0r0d[9], gate955_0n, initialise);
  C2RI I230 (ifint_0n[10], i_0r0d[10], gate955_0n, initialise);
  C2RI I231 (ifint_0n[11], i_0r0d[11], gate955_0n, initialise);
  C2RI I232 (ifint_0n[12], i_0r0d[12], gate955_0n, initialise);
  C2RI I233 (ifint_0n[13], i_0r0d[13], gate955_0n, initialise);
  C2RI I234 (ifint_0n[14], i_0r0d[14], gate955_0n, initialise);
  C2RI I235 (ifint_0n[15], i_0r0d[15], gate955_0n, initialise);
  C2RI I236 (ifint_0n[16], i_0r0d[16], gate955_0n, initialise);
  C2RI I237 (ifint_0n[17], i_0r0d[17], gate955_0n, initialise);
  C2RI I238 (ifint_0n[18], i_0r0d[18], gate955_0n, initialise);
  C2RI I239 (ifint_0n[19], i_0r0d[19], gate955_0n, initialise);
  C2RI I240 (ifint_0n[20], i_0r0d[20], gate955_0n, initialise);
  C2RI I241 (ifint_0n[21], i_0r0d[21], gate955_0n, initialise);
  C2RI I242 (ifint_0n[22], i_0r0d[22], gate955_0n, initialise);
  C2RI I243 (ifint_0n[23], i_0r0d[23], gate955_0n, initialise);
  C2RI I244 (ifint_0n[24], i_0r0d[24], gate955_0n, initialise);
  C2RI I245 (ifint_0n[25], i_0r0d[25], gate955_0n, initialise);
  C2RI I246 (ifint_0n[26], i_0r0d[26], gate955_0n, initialise);
  C2RI I247 (ifint_0n[27], i_0r0d[27], gate955_0n, initialise);
  C2RI I248 (ifint_0n[28], i_0r0d[28], gate955_0n, initialise);
  C2RI I249 (ifint_0n[29], i_0r0d[29], gate955_0n, initialise);
  C2RI I250 (ifint_0n[30], i_0r0d[30], gate955_0n, initialise);
  C2RI I251 (ifint_0n[31], i_0r0d[31], gate955_0n, initialise);
  C2RI I252 (ifint_0n[32], i_0r0d[32], gate955_0n, initialise);
  C2RI I253 (ifint_0n[33], i_0r0d[33], gate955_0n, initialise);
  C2RI I254 (ifint_0n[34], i_0r0d[34], gate955_0n, initialise);
  C2RI I255 (ifint_0n[35], i_0r0d[35], gate955_0n, initialise);
  C3 I256 (internal_0n[36], complete952_0n[0], complete952_0n[1], complete952_0n[2]);
  C3 I257 (internal_0n[37], complete952_0n[3], complete952_0n[4], complete952_0n[5]);
  C3 I258 (internal_0n[38], complete952_0n[6], complete952_0n[7], complete952_0n[8]);
  C3 I259 (internal_0n[39], complete952_0n[9], complete952_0n[10], complete952_0n[11]);
  C3 I260 (internal_0n[40], complete952_0n[12], complete952_0n[13], complete952_0n[14]);
  C3 I261 (internal_0n[41], complete952_0n[15], complete952_0n[16], complete952_0n[17]);
  C3 I262 (internal_0n[42], complete952_0n[18], complete952_0n[19], complete952_0n[20]);
  C3 I263 (internal_0n[43], complete952_0n[21], complete952_0n[22], complete952_0n[23]);
  C3 I264 (internal_0n[44], complete952_0n[24], complete952_0n[25], complete952_0n[26]);
  C3 I265 (internal_0n[45], complete952_0n[27], complete952_0n[28], complete952_0n[29]);
  C3 I266 (internal_0n[46], complete952_0n[30], complete952_0n[31], complete952_0n[32]);
  C3 I267 (internal_0n[47], complete952_0n[33], complete952_0n[34], complete952_0n[35]);
  C3 I268 (internal_0n[48], internal_0n[36], internal_0n[37], internal_0n[38]);
  C3 I269 (internal_0n[49], internal_0n[39], internal_0n[40], internal_0n[41]);
  C3 I270 (internal_0n[50], internal_0n[42], internal_0n[43], internal_0n[44]);
  C3 I271 (internal_0n[51], internal_0n[45], internal_0n[46], internal_0n[47]);
  C2 I272 (internal_0n[52], internal_0n[48], internal_0n[49]);
  C2 I273 (internal_0n[53], internal_0n[50], internal_0n[51]);
  C2 I274 (oaint_0n, internal_0n[52], internal_0n[53]);
  OR2 I275 (complete952_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I276 (complete952_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I277 (complete952_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I278 (complete952_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I279 (complete952_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I280 (complete952_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I281 (complete952_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I282 (complete952_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I283 (complete952_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I284 (complete952_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I285 (complete952_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I286 (complete952_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I287 (complete952_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I288 (complete952_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I289 (complete952_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I290 (complete952_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I291 (complete952_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I292 (complete952_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I293 (complete952_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I294 (complete952_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I295 (complete952_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I296 (complete952_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I297 (complete952_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I298 (complete952_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I299 (complete952_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I300 (complete952_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I301 (complete952_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I302 (complete952_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I303 (complete952_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I304 (complete952_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I305 (complete952_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I306 (complete952_0n[31], o_0r0d[31], o_0r1d[31]);
  OR2 I307 (complete952_0n[32], o_0r0d[32], o_0r1d[32]);
  OR2 I308 (complete952_0n[33], o_0r0d[33], o_0r1d[33]);
  OR2 I309 (complete952_0n[34], o_0r0d[34], o_0r1d[34]);
  OR2 I310 (complete952_0n[35], o_0r0d[35], o_0r1d[35]);
  INV I311 (gate951_0n, o_0a);
  C2RI I312 (o_0r1d[0], otint_0n[0], gate951_0n, initialise);
  C2RI I313 (o_0r1d[1], otint_0n[1], gate951_0n, initialise);
  C2RI I314 (o_0r1d[2], otint_0n[2], gate951_0n, initialise);
  C2RI I315 (o_0r1d[3], otint_0n[3], gate951_0n, initialise);
  C2RI I316 (o_0r1d[4], otint_0n[4], gate951_0n, initialise);
  C2RI I317 (o_0r1d[5], otint_0n[5], gate951_0n, initialise);
  C2RI I318 (o_0r1d[6], otint_0n[6], gate951_0n, initialise);
  C2RI I319 (o_0r1d[7], otint_0n[7], gate951_0n, initialise);
  C2RI I320 (o_0r1d[8], otint_0n[8], gate951_0n, initialise);
  C2RI I321 (o_0r1d[9], otint_0n[9], gate951_0n, initialise);
  C2RI I322 (o_0r1d[10], otint_0n[10], gate951_0n, initialise);
  C2RI I323 (o_0r1d[11], otint_0n[11], gate951_0n, initialise);
  C2RI I324 (o_0r1d[12], otint_0n[12], gate951_0n, initialise);
  C2RI I325 (o_0r1d[13], otint_0n[13], gate951_0n, initialise);
  C2RI I326 (o_0r1d[14], otint_0n[14], gate951_0n, initialise);
  C2RI I327 (o_0r1d[15], otint_0n[15], gate951_0n, initialise);
  C2RI I328 (o_0r1d[16], otint_0n[16], gate951_0n, initialise);
  C2RI I329 (o_0r1d[17], otint_0n[17], gate951_0n, initialise);
  C2RI I330 (o_0r1d[18], otint_0n[18], gate951_0n, initialise);
  C2RI I331 (o_0r1d[19], otint_0n[19], gate951_0n, initialise);
  C2RI I332 (o_0r1d[20], otint_0n[20], gate951_0n, initialise);
  C2RI I333 (o_0r1d[21], otint_0n[21], gate951_0n, initialise);
  C2RI I334 (o_0r1d[22], otint_0n[22], gate951_0n, initialise);
  C2RI I335 (o_0r1d[23], otint_0n[23], gate951_0n, initialise);
  C2RI I336 (o_0r1d[24], otint_0n[24], gate951_0n, initialise);
  C2RI I337 (o_0r1d[25], otint_0n[25], gate951_0n, initialise);
  C2RI I338 (o_0r1d[26], otint_0n[26], gate951_0n, initialise);
  C2RI I339 (o_0r1d[27], otint_0n[27], gate951_0n, initialise);
  C2RI I340 (o_0r1d[28], otint_0n[28], gate951_0n, initialise);
  C2RI I341 (o_0r1d[29], otint_0n[29], gate951_0n, initialise);
  C2RI I342 (o_0r1d[30], otint_0n[30], gate951_0n, initialise);
  C2RI I343 (o_0r1d[31], otint_0n[31], gate951_0n, initialise);
  C2RI I344 (o_0r1d[32], otint_0n[32], gate951_0n, initialise);
  C2RI I345 (o_0r1d[33], otint_0n[33], gate951_0n, initialise);
  C2RI I346 (o_0r1d[34], otint_0n[34], gate951_0n, initialise);
  C2RI I347 (o_0r1d[35], otint_0n[35], gate951_0n, initialise);
  C2RI I348 (o_0r0d[0], ofint_0n[0], gate951_0n, initialise);
  C2RI I349 (o_0r0d[1], ofint_0n[1], gate951_0n, initialise);
  C2RI I350 (o_0r0d[2], ofint_0n[2], gate951_0n, initialise);
  C2RI I351 (o_0r0d[3], ofint_0n[3], gate951_0n, initialise);
  C2RI I352 (o_0r0d[4], ofint_0n[4], gate951_0n, initialise);
  C2RI I353 (o_0r0d[5], ofint_0n[5], gate951_0n, initialise);
  C2RI I354 (o_0r0d[6], ofint_0n[6], gate951_0n, initialise);
  C2RI I355 (o_0r0d[7], ofint_0n[7], gate951_0n, initialise);
  C2RI I356 (o_0r0d[8], ofint_0n[8], gate951_0n, initialise);
  C2RI I357 (o_0r0d[9], ofint_0n[9], gate951_0n, initialise);
  C2RI I358 (o_0r0d[10], ofint_0n[10], gate951_0n, initialise);
  C2RI I359 (o_0r0d[11], ofint_0n[11], gate951_0n, initialise);
  C2RI I360 (o_0r0d[12], ofint_0n[12], gate951_0n, initialise);
  C2RI I361 (o_0r0d[13], ofint_0n[13], gate951_0n, initialise);
  C2RI I362 (o_0r0d[14], ofint_0n[14], gate951_0n, initialise);
  C2RI I363 (o_0r0d[15], ofint_0n[15], gate951_0n, initialise);
  C2RI I364 (o_0r0d[16], ofint_0n[16], gate951_0n, initialise);
  C2RI I365 (o_0r0d[17], ofint_0n[17], gate951_0n, initialise);
  C2RI I366 (o_0r0d[18], ofint_0n[18], gate951_0n, initialise);
  C2RI I367 (o_0r0d[19], ofint_0n[19], gate951_0n, initialise);
  C2RI I368 (o_0r0d[20], ofint_0n[20], gate951_0n, initialise);
  C2RI I369 (o_0r0d[21], ofint_0n[21], gate951_0n, initialise);
  C2RI I370 (o_0r0d[22], ofint_0n[22], gate951_0n, initialise);
  C2RI I371 (o_0r0d[23], ofint_0n[23], gate951_0n, initialise);
  C2RI I372 (o_0r0d[24], ofint_0n[24], gate951_0n, initialise);
  C2RI I373 (o_0r0d[25], ofint_0n[25], gate951_0n, initialise);
  C2RI I374 (o_0r0d[26], ofint_0n[26], gate951_0n, initialise);
  C2RI I375 (o_0r0d[27], ofint_0n[27], gate951_0n, initialise);
  C2RI I376 (o_0r0d[28], ofint_0n[28], gate951_0n, initialise);
  C2RI I377 (o_0r0d[29], ofint_0n[29], gate951_0n, initialise);
  C2RI I378 (o_0r0d[30], ofint_0n[30], gate951_0n, initialise);
  C2RI I379 (o_0r0d[31], ofint_0n[31], gate951_0n, initialise);
  C2RI I380 (o_0r0d[32], ofint_0n[32], gate951_0n, initialise);
  C2RI I381 (o_0r0d[33], ofint_0n[33], gate951_0n, initialise);
  C2RI I382 (o_0r0d[34], ofint_0n[34], gate951_0n, initialise);
  C2RI I383 (o_0r0d[35], ofint_0n[35], gate951_0n, initialise);
  C2RI I384 (iaint_0n, sel_0n[0], oaint_0n, initialise);
  C2RI I385 (iaint_1n, sel_0n[1], oaint_0n, initialise);
  assign gate_0n[0] = sel_0n[0];
  assign gate_0n[1] = sel_0n[1];
  assign sel_0n[0] = selcomp_0n;
  assign sel_0n[1] = selcomp_1n;
  C3 I390 (internal_0n[54], complete948_0n[0], complete948_0n[1], complete948_0n[2]);
  C3 I391 (internal_0n[55], complete948_0n[3], complete948_0n[4], complete948_0n[5]);
  C3 I392 (internal_0n[56], complete948_0n[6], complete948_0n[7], complete948_0n[8]);
  C3 I393 (internal_0n[57], complete948_0n[9], complete948_0n[10], complete948_0n[11]);
  C3 I394 (internal_0n[58], complete948_0n[12], complete948_0n[13], complete948_0n[14]);
  C3 I395 (internal_0n[59], complete948_0n[15], complete948_0n[16], complete948_0n[17]);
  C3 I396 (internal_0n[60], complete948_0n[18], complete948_0n[19], complete948_0n[20]);
  C3 I397 (internal_0n[61], complete948_0n[21], complete948_0n[22], complete948_0n[23]);
  C3 I398 (internal_0n[62], complete948_0n[24], complete948_0n[25], complete948_0n[26]);
  C3 I399 (internal_0n[63], complete948_0n[27], complete948_0n[28], complete948_0n[29]);
  C3 I400 (internal_0n[64], complete948_0n[30], complete948_0n[31], complete948_0n[32]);
  C3 I401 (internal_0n[65], complete948_0n[33], complete948_0n[34], complete948_0n[35]);
  C3 I402 (internal_0n[66], internal_0n[54], internal_0n[55], internal_0n[56]);
  C3 I403 (internal_0n[67], internal_0n[57], internal_0n[58], internal_0n[59]);
  C3 I404 (internal_0n[68], internal_0n[60], internal_0n[61], internal_0n[62]);
  C3 I405 (internal_0n[69], internal_0n[63], internal_0n[64], internal_0n[65]);
  C2 I406 (internal_0n[70], internal_0n[66], internal_0n[67]);
  C2 I407 (internal_0n[71], internal_0n[68], internal_0n[69]);
  C2 I408 (selcomp_1n, internal_0n[70], internal_0n[71]);
  OR2 I409 (complete948_0n[0], ifint_1n[0], itint_1n[0]);
  OR2 I410 (complete948_0n[1], ifint_1n[1], itint_1n[1]);
  OR2 I411 (complete948_0n[2], ifint_1n[2], itint_1n[2]);
  OR2 I412 (complete948_0n[3], ifint_1n[3], itint_1n[3]);
  OR2 I413 (complete948_0n[4], ifint_1n[4], itint_1n[4]);
  OR2 I414 (complete948_0n[5], ifint_1n[5], itint_1n[5]);
  OR2 I415 (complete948_0n[6], ifint_1n[6], itint_1n[6]);
  OR2 I416 (complete948_0n[7], ifint_1n[7], itint_1n[7]);
  OR2 I417 (complete948_0n[8], ifint_1n[8], itint_1n[8]);
  OR2 I418 (complete948_0n[9], ifint_1n[9], itint_1n[9]);
  OR2 I419 (complete948_0n[10], ifint_1n[10], itint_1n[10]);
  OR2 I420 (complete948_0n[11], ifint_1n[11], itint_1n[11]);
  OR2 I421 (complete948_0n[12], ifint_1n[12], itint_1n[12]);
  OR2 I422 (complete948_0n[13], ifint_1n[13], itint_1n[13]);
  OR2 I423 (complete948_0n[14], ifint_1n[14], itint_1n[14]);
  OR2 I424 (complete948_0n[15], ifint_1n[15], itint_1n[15]);
  OR2 I425 (complete948_0n[16], ifint_1n[16], itint_1n[16]);
  OR2 I426 (complete948_0n[17], ifint_1n[17], itint_1n[17]);
  OR2 I427 (complete948_0n[18], ifint_1n[18], itint_1n[18]);
  OR2 I428 (complete948_0n[19], ifint_1n[19], itint_1n[19]);
  OR2 I429 (complete948_0n[20], ifint_1n[20], itint_1n[20]);
  OR2 I430 (complete948_0n[21], ifint_1n[21], itint_1n[21]);
  OR2 I431 (complete948_0n[22], ifint_1n[22], itint_1n[22]);
  OR2 I432 (complete948_0n[23], ifint_1n[23], itint_1n[23]);
  OR2 I433 (complete948_0n[24], ifint_1n[24], itint_1n[24]);
  OR2 I434 (complete948_0n[25], ifint_1n[25], itint_1n[25]);
  OR2 I435 (complete948_0n[26], ifint_1n[26], itint_1n[26]);
  OR2 I436 (complete948_0n[27], ifint_1n[27], itint_1n[27]);
  OR2 I437 (complete948_0n[28], ifint_1n[28], itint_1n[28]);
  OR2 I438 (complete948_0n[29], ifint_1n[29], itint_1n[29]);
  OR2 I439 (complete948_0n[30], ifint_1n[30], itint_1n[30]);
  OR2 I440 (complete948_0n[31], ifint_1n[31], itint_1n[31]);
  OR2 I441 (complete948_0n[32], ifint_1n[32], itint_1n[32]);
  OR2 I442 (complete948_0n[33], ifint_1n[33], itint_1n[33]);
  OR2 I443 (complete948_0n[34], ifint_1n[34], itint_1n[34]);
  OR2 I444 (complete948_0n[35], ifint_1n[35], itint_1n[35]);
  C3 I445 (internal_0n[72], complete947_0n[0], complete947_0n[1], complete947_0n[2]);
  C3 I446 (internal_0n[73], complete947_0n[3], complete947_0n[4], complete947_0n[5]);
  C3 I447 (internal_0n[74], complete947_0n[6], complete947_0n[7], complete947_0n[8]);
  C3 I448 (internal_0n[75], complete947_0n[9], complete947_0n[10], complete947_0n[11]);
  C3 I449 (internal_0n[76], complete947_0n[12], complete947_0n[13], complete947_0n[14]);
  C3 I450 (internal_0n[77], complete947_0n[15], complete947_0n[16], complete947_0n[17]);
  C3 I451 (internal_0n[78], complete947_0n[18], complete947_0n[19], complete947_0n[20]);
  C3 I452 (internal_0n[79], complete947_0n[21], complete947_0n[22], complete947_0n[23]);
  C3 I453 (internal_0n[80], complete947_0n[24], complete947_0n[25], complete947_0n[26]);
  C3 I454 (internal_0n[81], complete947_0n[27], complete947_0n[28], complete947_0n[29]);
  C3 I455 (internal_0n[82], complete947_0n[30], complete947_0n[31], complete947_0n[32]);
  C3 I456 (internal_0n[83], complete947_0n[33], complete947_0n[34], complete947_0n[35]);
  C3 I457 (internal_0n[84], internal_0n[72], internal_0n[73], internal_0n[74]);
  C3 I458 (internal_0n[85], internal_0n[75], internal_0n[76], internal_0n[77]);
  C3 I459 (internal_0n[86], internal_0n[78], internal_0n[79], internal_0n[80]);
  C3 I460 (internal_0n[87], internal_0n[81], internal_0n[82], internal_0n[83]);
  C2 I461 (internal_0n[88], internal_0n[84], internal_0n[85]);
  C2 I462 (internal_0n[89], internal_0n[86], internal_0n[87]);
  C2 I463 (selcomp_0n, internal_0n[88], internal_0n[89]);
  OR2 I464 (complete947_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I465 (complete947_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I466 (complete947_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I467 (complete947_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I468 (complete947_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I469 (complete947_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I470 (complete947_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I471 (complete947_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I472 (complete947_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I473 (complete947_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I474 (complete947_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I475 (complete947_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I476 (complete947_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I477 (complete947_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I478 (complete947_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I479 (complete947_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I480 (complete947_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I481 (complete947_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I482 (complete947_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I483 (complete947_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I484 (complete947_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I485 (complete947_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I486 (complete947_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I487 (complete947_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I488 (complete947_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I489 (complete947_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I490 (complete947_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I491 (complete947_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I492 (complete947_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I493 (complete947_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I494 (complete947_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I495 (complete947_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I496 (complete947_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I497 (complete947_0n[33], ifint_0n[33], itint_0n[33]);
  OR2 I498 (complete947_0n[34], ifint_0n[34], itint_0n[34]);
  OR2 I499 (complete947_0n[35], ifint_0n[35], itint_0n[35]);
  AND2 I500 (gfint_0n[0], gate_0n[0], ifint_0n[0]);
  AND2 I501 (gfint_0n[1], gate_0n[0], ifint_0n[1]);
  AND2 I502 (gfint_0n[2], gate_0n[0], ifint_0n[2]);
  AND2 I503 (gfint_0n[3], gate_0n[0], ifint_0n[3]);
  AND2 I504 (gfint_0n[4], gate_0n[0], ifint_0n[4]);
  AND2 I505 (gfint_0n[5], gate_0n[0], ifint_0n[5]);
  AND2 I506 (gfint_0n[6], gate_0n[0], ifint_0n[6]);
  AND2 I507 (gfint_0n[7], gate_0n[0], ifint_0n[7]);
  AND2 I508 (gfint_0n[8], gate_0n[0], ifint_0n[8]);
  AND2 I509 (gfint_0n[9], gate_0n[0], ifint_0n[9]);
  AND2 I510 (gfint_0n[10], gate_0n[0], ifint_0n[10]);
  AND2 I511 (gfint_0n[11], gate_0n[0], ifint_0n[11]);
  AND2 I512 (gfint_0n[12], gate_0n[0], ifint_0n[12]);
  AND2 I513 (gfint_0n[13], gate_0n[0], ifint_0n[13]);
  AND2 I514 (gfint_0n[14], gate_0n[0], ifint_0n[14]);
  AND2 I515 (gfint_0n[15], gate_0n[0], ifint_0n[15]);
  AND2 I516 (gfint_0n[16], gate_0n[0], ifint_0n[16]);
  AND2 I517 (gfint_0n[17], gate_0n[0], ifint_0n[17]);
  AND2 I518 (gfint_0n[18], gate_0n[0], ifint_0n[18]);
  AND2 I519 (gfint_0n[19], gate_0n[0], ifint_0n[19]);
  AND2 I520 (gfint_0n[20], gate_0n[0], ifint_0n[20]);
  AND2 I521 (gfint_0n[21], gate_0n[0], ifint_0n[21]);
  AND2 I522 (gfint_0n[22], gate_0n[0], ifint_0n[22]);
  AND2 I523 (gfint_0n[23], gate_0n[0], ifint_0n[23]);
  AND2 I524 (gfint_0n[24], gate_0n[0], ifint_0n[24]);
  AND2 I525 (gfint_0n[25], gate_0n[0], ifint_0n[25]);
  AND2 I526 (gfint_0n[26], gate_0n[0], ifint_0n[26]);
  AND2 I527 (gfint_0n[27], gate_0n[0], ifint_0n[27]);
  AND2 I528 (gfint_0n[28], gate_0n[0], ifint_0n[28]);
  AND2 I529 (gfint_0n[29], gate_0n[0], ifint_0n[29]);
  AND2 I530 (gfint_0n[30], gate_0n[0], ifint_0n[30]);
  AND2 I531 (gfint_0n[31], gate_0n[0], ifint_0n[31]);
  AND2 I532 (gfint_0n[32], gate_0n[0], ifint_0n[32]);
  AND2 I533 (gfint_0n[33], gate_0n[0], ifint_0n[33]);
  AND2 I534 (gfint_0n[34], gate_0n[0], ifint_0n[34]);
  AND2 I535 (gfint_0n[35], gate_0n[0], ifint_0n[35]);
  AND2 I536 (gfint_1n[0], gate_0n[1], ifint_1n[0]);
  AND2 I537 (gfint_1n[1], gate_0n[1], ifint_1n[1]);
  AND2 I538 (gfint_1n[2], gate_0n[1], ifint_1n[2]);
  AND2 I539 (gfint_1n[3], gate_0n[1], ifint_1n[3]);
  AND2 I540 (gfint_1n[4], gate_0n[1], ifint_1n[4]);
  AND2 I541 (gfint_1n[5], gate_0n[1], ifint_1n[5]);
  AND2 I542 (gfint_1n[6], gate_0n[1], ifint_1n[6]);
  AND2 I543 (gfint_1n[7], gate_0n[1], ifint_1n[7]);
  AND2 I544 (gfint_1n[8], gate_0n[1], ifint_1n[8]);
  AND2 I545 (gfint_1n[9], gate_0n[1], ifint_1n[9]);
  AND2 I546 (gfint_1n[10], gate_0n[1], ifint_1n[10]);
  AND2 I547 (gfint_1n[11], gate_0n[1], ifint_1n[11]);
  AND2 I548 (gfint_1n[12], gate_0n[1], ifint_1n[12]);
  AND2 I549 (gfint_1n[13], gate_0n[1], ifint_1n[13]);
  AND2 I550 (gfint_1n[14], gate_0n[1], ifint_1n[14]);
  AND2 I551 (gfint_1n[15], gate_0n[1], ifint_1n[15]);
  AND2 I552 (gfint_1n[16], gate_0n[1], ifint_1n[16]);
  AND2 I553 (gfint_1n[17], gate_0n[1], ifint_1n[17]);
  AND2 I554 (gfint_1n[18], gate_0n[1], ifint_1n[18]);
  AND2 I555 (gfint_1n[19], gate_0n[1], ifint_1n[19]);
  AND2 I556 (gfint_1n[20], gate_0n[1], ifint_1n[20]);
  AND2 I557 (gfint_1n[21], gate_0n[1], ifint_1n[21]);
  AND2 I558 (gfint_1n[22], gate_0n[1], ifint_1n[22]);
  AND2 I559 (gfint_1n[23], gate_0n[1], ifint_1n[23]);
  AND2 I560 (gfint_1n[24], gate_0n[1], ifint_1n[24]);
  AND2 I561 (gfint_1n[25], gate_0n[1], ifint_1n[25]);
  AND2 I562 (gfint_1n[26], gate_0n[1], ifint_1n[26]);
  AND2 I563 (gfint_1n[27], gate_0n[1], ifint_1n[27]);
  AND2 I564 (gfint_1n[28], gate_0n[1], ifint_1n[28]);
  AND2 I565 (gfint_1n[29], gate_0n[1], ifint_1n[29]);
  AND2 I566 (gfint_1n[30], gate_0n[1], ifint_1n[30]);
  AND2 I567 (gfint_1n[31], gate_0n[1], ifint_1n[31]);
  AND2 I568 (gfint_1n[32], gate_0n[1], ifint_1n[32]);
  AND2 I569 (gfint_1n[33], gate_0n[1], ifint_1n[33]);
  AND2 I570 (gfint_1n[34], gate_0n[1], ifint_1n[34]);
  AND2 I571 (gfint_1n[35], gate_0n[1], ifint_1n[35]);
  AND2 I572 (gtint_0n[0], gate_0n[0], itint_0n[0]);
  AND2 I573 (gtint_0n[1], gate_0n[0], itint_0n[1]);
  AND2 I574 (gtint_0n[2], gate_0n[0], itint_0n[2]);
  AND2 I575 (gtint_0n[3], gate_0n[0], itint_0n[3]);
  AND2 I576 (gtint_0n[4], gate_0n[0], itint_0n[4]);
  AND2 I577 (gtint_0n[5], gate_0n[0], itint_0n[5]);
  AND2 I578 (gtint_0n[6], gate_0n[0], itint_0n[6]);
  AND2 I579 (gtint_0n[7], gate_0n[0], itint_0n[7]);
  AND2 I580 (gtint_0n[8], gate_0n[0], itint_0n[8]);
  AND2 I581 (gtint_0n[9], gate_0n[0], itint_0n[9]);
  AND2 I582 (gtint_0n[10], gate_0n[0], itint_0n[10]);
  AND2 I583 (gtint_0n[11], gate_0n[0], itint_0n[11]);
  AND2 I584 (gtint_0n[12], gate_0n[0], itint_0n[12]);
  AND2 I585 (gtint_0n[13], gate_0n[0], itint_0n[13]);
  AND2 I586 (gtint_0n[14], gate_0n[0], itint_0n[14]);
  AND2 I587 (gtint_0n[15], gate_0n[0], itint_0n[15]);
  AND2 I588 (gtint_0n[16], gate_0n[0], itint_0n[16]);
  AND2 I589 (gtint_0n[17], gate_0n[0], itint_0n[17]);
  AND2 I590 (gtint_0n[18], gate_0n[0], itint_0n[18]);
  AND2 I591 (gtint_0n[19], gate_0n[0], itint_0n[19]);
  AND2 I592 (gtint_0n[20], gate_0n[0], itint_0n[20]);
  AND2 I593 (gtint_0n[21], gate_0n[0], itint_0n[21]);
  AND2 I594 (gtint_0n[22], gate_0n[0], itint_0n[22]);
  AND2 I595 (gtint_0n[23], gate_0n[0], itint_0n[23]);
  AND2 I596 (gtint_0n[24], gate_0n[0], itint_0n[24]);
  AND2 I597 (gtint_0n[25], gate_0n[0], itint_0n[25]);
  AND2 I598 (gtint_0n[26], gate_0n[0], itint_0n[26]);
  AND2 I599 (gtint_0n[27], gate_0n[0], itint_0n[27]);
  AND2 I600 (gtint_0n[28], gate_0n[0], itint_0n[28]);
  AND2 I601 (gtint_0n[29], gate_0n[0], itint_0n[29]);
  AND2 I602 (gtint_0n[30], gate_0n[0], itint_0n[30]);
  AND2 I603 (gtint_0n[31], gate_0n[0], itint_0n[31]);
  AND2 I604 (gtint_0n[32], gate_0n[0], itint_0n[32]);
  AND2 I605 (gtint_0n[33], gate_0n[0], itint_0n[33]);
  AND2 I606 (gtint_0n[34], gate_0n[0], itint_0n[34]);
  AND2 I607 (gtint_0n[35], gate_0n[0], itint_0n[35]);
  AND2 I608 (gtint_1n[0], gate_0n[1], itint_1n[0]);
  AND2 I609 (gtint_1n[1], gate_0n[1], itint_1n[1]);
  AND2 I610 (gtint_1n[2], gate_0n[1], itint_1n[2]);
  AND2 I611 (gtint_1n[3], gate_0n[1], itint_1n[3]);
  AND2 I612 (gtint_1n[4], gate_0n[1], itint_1n[4]);
  AND2 I613 (gtint_1n[5], gate_0n[1], itint_1n[5]);
  AND2 I614 (gtint_1n[6], gate_0n[1], itint_1n[6]);
  AND2 I615 (gtint_1n[7], gate_0n[1], itint_1n[7]);
  AND2 I616 (gtint_1n[8], gate_0n[1], itint_1n[8]);
  AND2 I617 (gtint_1n[9], gate_0n[1], itint_1n[9]);
  AND2 I618 (gtint_1n[10], gate_0n[1], itint_1n[10]);
  AND2 I619 (gtint_1n[11], gate_0n[1], itint_1n[11]);
  AND2 I620 (gtint_1n[12], gate_0n[1], itint_1n[12]);
  AND2 I621 (gtint_1n[13], gate_0n[1], itint_1n[13]);
  AND2 I622 (gtint_1n[14], gate_0n[1], itint_1n[14]);
  AND2 I623 (gtint_1n[15], gate_0n[1], itint_1n[15]);
  AND2 I624 (gtint_1n[16], gate_0n[1], itint_1n[16]);
  AND2 I625 (gtint_1n[17], gate_0n[1], itint_1n[17]);
  AND2 I626 (gtint_1n[18], gate_0n[1], itint_1n[18]);
  AND2 I627 (gtint_1n[19], gate_0n[1], itint_1n[19]);
  AND2 I628 (gtint_1n[20], gate_0n[1], itint_1n[20]);
  AND2 I629 (gtint_1n[21], gate_0n[1], itint_1n[21]);
  AND2 I630 (gtint_1n[22], gate_0n[1], itint_1n[22]);
  AND2 I631 (gtint_1n[23], gate_0n[1], itint_1n[23]);
  AND2 I632 (gtint_1n[24], gate_0n[1], itint_1n[24]);
  AND2 I633 (gtint_1n[25], gate_0n[1], itint_1n[25]);
  AND2 I634 (gtint_1n[26], gate_0n[1], itint_1n[26]);
  AND2 I635 (gtint_1n[27], gate_0n[1], itint_1n[27]);
  AND2 I636 (gtint_1n[28], gate_0n[1], itint_1n[28]);
  AND2 I637 (gtint_1n[29], gate_0n[1], itint_1n[29]);
  AND2 I638 (gtint_1n[30], gate_0n[1], itint_1n[30]);
  AND2 I639 (gtint_1n[31], gate_0n[1], itint_1n[31]);
  AND2 I640 (gtint_1n[32], gate_0n[1], itint_1n[32]);
  AND2 I641 (gtint_1n[33], gate_0n[1], itint_1n[33]);
  AND2 I642 (gtint_1n[34], gate_0n[1], itint_1n[34]);
  AND2 I643 (gtint_1n[35], gate_0n[1], itint_1n[35]);
  OR2 I644 (otint_0n[0], gtint_0n[0], gtint_1n[0]);
  OR2 I645 (otint_0n[1], gtint_0n[1], gtint_1n[1]);
  OR2 I646 (otint_0n[2], gtint_0n[2], gtint_1n[2]);
  OR2 I647 (otint_0n[3], gtint_0n[3], gtint_1n[3]);
  OR2 I648 (otint_0n[4], gtint_0n[4], gtint_1n[4]);
  OR2 I649 (otint_0n[5], gtint_0n[5], gtint_1n[5]);
  OR2 I650 (otint_0n[6], gtint_0n[6], gtint_1n[6]);
  OR2 I651 (otint_0n[7], gtint_0n[7], gtint_1n[7]);
  OR2 I652 (otint_0n[8], gtint_0n[8], gtint_1n[8]);
  OR2 I653 (otint_0n[9], gtint_0n[9], gtint_1n[9]);
  OR2 I654 (otint_0n[10], gtint_0n[10], gtint_1n[10]);
  OR2 I655 (otint_0n[11], gtint_0n[11], gtint_1n[11]);
  OR2 I656 (otint_0n[12], gtint_0n[12], gtint_1n[12]);
  OR2 I657 (otint_0n[13], gtint_0n[13], gtint_1n[13]);
  OR2 I658 (otint_0n[14], gtint_0n[14], gtint_1n[14]);
  OR2 I659 (otint_0n[15], gtint_0n[15], gtint_1n[15]);
  OR2 I660 (otint_0n[16], gtint_0n[16], gtint_1n[16]);
  OR2 I661 (otint_0n[17], gtint_0n[17], gtint_1n[17]);
  OR2 I662 (otint_0n[18], gtint_0n[18], gtint_1n[18]);
  OR2 I663 (otint_0n[19], gtint_0n[19], gtint_1n[19]);
  OR2 I664 (otint_0n[20], gtint_0n[20], gtint_1n[20]);
  OR2 I665 (otint_0n[21], gtint_0n[21], gtint_1n[21]);
  OR2 I666 (otint_0n[22], gtint_0n[22], gtint_1n[22]);
  OR2 I667 (otint_0n[23], gtint_0n[23], gtint_1n[23]);
  OR2 I668 (otint_0n[24], gtint_0n[24], gtint_1n[24]);
  OR2 I669 (otint_0n[25], gtint_0n[25], gtint_1n[25]);
  OR2 I670 (otint_0n[26], gtint_0n[26], gtint_1n[26]);
  OR2 I671 (otint_0n[27], gtint_0n[27], gtint_1n[27]);
  OR2 I672 (otint_0n[28], gtint_0n[28], gtint_1n[28]);
  OR2 I673 (otint_0n[29], gtint_0n[29], gtint_1n[29]);
  OR2 I674 (otint_0n[30], gtint_0n[30], gtint_1n[30]);
  OR2 I675 (otint_0n[31], gtint_0n[31], gtint_1n[31]);
  OR2 I676 (otint_0n[32], gtint_0n[32], gtint_1n[32]);
  OR2 I677 (otint_0n[33], gtint_0n[33], gtint_1n[33]);
  OR2 I678 (otint_0n[34], gtint_0n[34], gtint_1n[34]);
  OR2 I679 (otint_0n[35], gtint_0n[35], gtint_1n[35]);
  OR2 I680 (ofint_0n[0], gfint_0n[0], gfint_1n[0]);
  OR2 I681 (ofint_0n[1], gfint_0n[1], gfint_1n[1]);
  OR2 I682 (ofint_0n[2], gfint_0n[2], gfint_1n[2]);
  OR2 I683 (ofint_0n[3], gfint_0n[3], gfint_1n[3]);
  OR2 I684 (ofint_0n[4], gfint_0n[4], gfint_1n[4]);
  OR2 I685 (ofint_0n[5], gfint_0n[5], gfint_1n[5]);
  OR2 I686 (ofint_0n[6], gfint_0n[6], gfint_1n[6]);
  OR2 I687 (ofint_0n[7], gfint_0n[7], gfint_1n[7]);
  OR2 I688 (ofint_0n[8], gfint_0n[8], gfint_1n[8]);
  OR2 I689 (ofint_0n[9], gfint_0n[9], gfint_1n[9]);
  OR2 I690 (ofint_0n[10], gfint_0n[10], gfint_1n[10]);
  OR2 I691 (ofint_0n[11], gfint_0n[11], gfint_1n[11]);
  OR2 I692 (ofint_0n[12], gfint_0n[12], gfint_1n[12]);
  OR2 I693 (ofint_0n[13], gfint_0n[13], gfint_1n[13]);
  OR2 I694 (ofint_0n[14], gfint_0n[14], gfint_1n[14]);
  OR2 I695 (ofint_0n[15], gfint_0n[15], gfint_1n[15]);
  OR2 I696 (ofint_0n[16], gfint_0n[16], gfint_1n[16]);
  OR2 I697 (ofint_0n[17], gfint_0n[17], gfint_1n[17]);
  OR2 I698 (ofint_0n[18], gfint_0n[18], gfint_1n[18]);
  OR2 I699 (ofint_0n[19], gfint_0n[19], gfint_1n[19]);
  OR2 I700 (ofint_0n[20], gfint_0n[20], gfint_1n[20]);
  OR2 I701 (ofint_0n[21], gfint_0n[21], gfint_1n[21]);
  OR2 I702 (ofint_0n[22], gfint_0n[22], gfint_1n[22]);
  OR2 I703 (ofint_0n[23], gfint_0n[23], gfint_1n[23]);
  OR2 I704 (ofint_0n[24], gfint_0n[24], gfint_1n[24]);
  OR2 I705 (ofint_0n[25], gfint_0n[25], gfint_1n[25]);
  OR2 I706 (ofint_0n[26], gfint_0n[26], gfint_1n[26]);
  OR2 I707 (ofint_0n[27], gfint_0n[27], gfint_1n[27]);
  OR2 I708 (ofint_0n[28], gfint_0n[28], gfint_1n[28]);
  OR2 I709 (ofint_0n[29], gfint_0n[29], gfint_1n[29]);
  OR2 I710 (ofint_0n[30], gfint_0n[30], gfint_1n[30]);
  OR2 I711 (ofint_0n[31], gfint_0n[31], gfint_1n[31]);
  OR2 I712 (ofint_0n[32], gfint_0n[32], gfint_1n[32]);
  OR2 I713 (ofint_0n[33], gfint_0n[33], gfint_1n[33]);
  OR2 I714 (ofint_0n[34], gfint_0n[34], gfint_1n[34]);
  OR2 I715 (ofint_0n[35], gfint_0n[35], gfint_1n[35]);
endmodule

module BrzO_0_1_l23__28_28num_201_200_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output o_0r0d;
  output o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d = gnd;
  assign o_0r0d = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_1_l23__28_28num_201_201_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output o_0r0d;
  output o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r0d = gnd;
  assign o_0r1d = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_2_l23__28_28num_202_200_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [1:0] o_0r0d;
  output [1:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[0] = gnd;
  assign o_0r1d[1] = gnd;
  assign o_0r0d[0] = go_0n;
  assign o_0r0d[1] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_2_l23__28_28num_202_201_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [1:0] o_0r0d;
  output [1:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[1] = gnd;
  assign o_0r0d[1] = go_0n;
  assign o_0r0d[0] = gnd;
  assign o_0r1d[0] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_2_l23__28_28num_202_202_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [1:0] o_0r0d;
  output [1:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[0] = gnd;
  assign o_0r0d[0] = go_0n;
  assign o_0r0d[1] = gnd;
  assign o_0r1d[1] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_3_l23__28_28num_203_201_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [2:0] o_0r0d;
  output [2:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[1] = gnd;
  assign o_0r1d[2] = gnd;
  assign o_0r0d[1] = go_0n;
  assign o_0r0d[2] = go_0n;
  assign o_0r0d[0] = gnd;
  assign o_0r1d[0] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_3_l23__28_28num_203_202_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [2:0] o_0r0d;
  output [2:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[0] = gnd;
  assign o_0r1d[2] = gnd;
  assign o_0r0d[0] = go_0n;
  assign o_0r0d[2] = go_0n;
  assign o_0r0d[1] = gnd;
  assign o_0r1d[1] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_3_l23__28_28num_203_204_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [2:0] o_0r0d;
  output [2:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[0] = gnd;
  assign o_0r1d[1] = gnd;
  assign o_0r0d[0] = go_0n;
  assign o_0r0d[1] = go_0n;
  assign o_0r0d[2] = gnd;
  assign o_0r1d[2] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_9_l23__28_28num_209_201_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [8:0] o_0r0d;
  output [8:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[1] = gnd;
  assign o_0r1d[2] = gnd;
  assign o_0r1d[3] = gnd;
  assign o_0r1d[4] = gnd;
  assign o_0r1d[5] = gnd;
  assign o_0r1d[6] = gnd;
  assign o_0r1d[7] = gnd;
  assign o_0r1d[8] = gnd;
  assign o_0r0d[1] = go_0n;
  assign o_0r0d[2] = go_0n;
  assign o_0r0d[3] = go_0n;
  assign o_0r0d[4] = go_0n;
  assign o_0r0d[5] = go_0n;
  assign o_0r0d[6] = go_0n;
  assign o_0r0d[7] = go_0n;
  assign o_0r0d[8] = go_0n;
  assign o_0r0d[0] = gnd;
  assign o_0r1d[0] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_9_l23__28_28num_209_202_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [8:0] o_0r0d;
  output [8:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[0] = gnd;
  assign o_0r1d[2] = gnd;
  assign o_0r1d[3] = gnd;
  assign o_0r1d[4] = gnd;
  assign o_0r1d[5] = gnd;
  assign o_0r1d[6] = gnd;
  assign o_0r1d[7] = gnd;
  assign o_0r1d[8] = gnd;
  assign o_0r0d[0] = go_0n;
  assign o_0r0d[2] = go_0n;
  assign o_0r0d[3] = go_0n;
  assign o_0r0d[4] = go_0n;
  assign o_0r0d[5] = go_0n;
  assign o_0r0d[6] = go_0n;
  assign o_0r0d[7] = go_0n;
  assign o_0r0d[8] = go_0n;
  assign o_0r0d[1] = gnd;
  assign o_0r1d[1] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_9_l23__28_28num_209_204_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [8:0] o_0r0d;
  output [8:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[0] = gnd;
  assign o_0r1d[1] = gnd;
  assign o_0r1d[3] = gnd;
  assign o_0r1d[4] = gnd;
  assign o_0r1d[5] = gnd;
  assign o_0r1d[6] = gnd;
  assign o_0r1d[7] = gnd;
  assign o_0r1d[8] = gnd;
  assign o_0r0d[0] = go_0n;
  assign o_0r0d[1] = go_0n;
  assign o_0r0d[3] = go_0n;
  assign o_0r0d[4] = go_0n;
  assign o_0r0d[5] = go_0n;
  assign o_0r0d[6] = go_0n;
  assign o_0r0d[7] = go_0n;
  assign o_0r0d[8] = go_0n;
  assign o_0r0d[2] = gnd;
  assign o_0r1d[2] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_9_l23__28_28num_209_208_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [8:0] o_0r0d;
  output [8:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[0] = gnd;
  assign o_0r1d[1] = gnd;
  assign o_0r1d[2] = gnd;
  assign o_0r1d[4] = gnd;
  assign o_0r1d[5] = gnd;
  assign o_0r1d[6] = gnd;
  assign o_0r1d[7] = gnd;
  assign o_0r1d[8] = gnd;
  assign o_0r0d[0] = go_0n;
  assign o_0r0d[1] = go_0n;
  assign o_0r0d[2] = go_0n;
  assign o_0r0d[4] = go_0n;
  assign o_0r0d[5] = go_0n;
  assign o_0r0d[6] = go_0n;
  assign o_0r0d[7] = go_0n;
  assign o_0r0d[8] = go_0n;
  assign o_0r0d[3] = gnd;
  assign o_0r1d[3] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_9_l24__28_28num_209_2016_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [8:0] o_0r0d;
  output [8:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[0] = gnd;
  assign o_0r1d[1] = gnd;
  assign o_0r1d[2] = gnd;
  assign o_0r1d[3] = gnd;
  assign o_0r1d[5] = gnd;
  assign o_0r1d[6] = gnd;
  assign o_0r1d[7] = gnd;
  assign o_0r1d[8] = gnd;
  assign o_0r0d[0] = go_0n;
  assign o_0r0d[1] = go_0n;
  assign o_0r0d[2] = go_0n;
  assign o_0r0d[3] = go_0n;
  assign o_0r0d[5] = go_0n;
  assign o_0r0d[6] = go_0n;
  assign o_0r0d[7] = go_0n;
  assign o_0r0d[8] = go_0n;
  assign o_0r0d[4] = gnd;
  assign o_0r1d[4] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_9_l24__28_28num_209_2032_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [8:0] o_0r0d;
  output [8:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[0] = gnd;
  assign o_0r1d[1] = gnd;
  assign o_0r1d[2] = gnd;
  assign o_0r1d[3] = gnd;
  assign o_0r1d[4] = gnd;
  assign o_0r1d[6] = gnd;
  assign o_0r1d[7] = gnd;
  assign o_0r1d[8] = gnd;
  assign o_0r0d[0] = go_0n;
  assign o_0r0d[1] = go_0n;
  assign o_0r0d[2] = go_0n;
  assign o_0r0d[3] = go_0n;
  assign o_0r0d[4] = go_0n;
  assign o_0r0d[6] = go_0n;
  assign o_0r0d[7] = go_0n;
  assign o_0r0d[8] = go_0n;
  assign o_0r0d[5] = gnd;
  assign o_0r1d[5] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_9_l24__28_28num_209_2064_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [8:0] o_0r0d;
  output [8:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[0] = gnd;
  assign o_0r1d[1] = gnd;
  assign o_0r1d[2] = gnd;
  assign o_0r1d[3] = gnd;
  assign o_0r1d[4] = gnd;
  assign o_0r1d[5] = gnd;
  assign o_0r1d[7] = gnd;
  assign o_0r1d[8] = gnd;
  assign o_0r0d[0] = go_0n;
  assign o_0r0d[1] = go_0n;
  assign o_0r0d[2] = go_0n;
  assign o_0r0d[3] = go_0n;
  assign o_0r0d[4] = go_0n;
  assign o_0r0d[5] = go_0n;
  assign o_0r0d[7] = go_0n;
  assign o_0r0d[8] = go_0n;
  assign o_0r0d[6] = gnd;
  assign o_0r1d[6] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_9_l25__28_28num_209_20128_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [8:0] o_0r0d;
  output [8:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[0] = gnd;
  assign o_0r1d[1] = gnd;
  assign o_0r1d[2] = gnd;
  assign o_0r1d[3] = gnd;
  assign o_0r1d[4] = gnd;
  assign o_0r1d[5] = gnd;
  assign o_0r1d[6] = gnd;
  assign o_0r1d[8] = gnd;
  assign o_0r0d[0] = go_0n;
  assign o_0r0d[1] = go_0n;
  assign o_0r0d[2] = go_0n;
  assign o_0r0d[3] = go_0n;
  assign o_0r0d[4] = go_0n;
  assign o_0r0d[5] = go_0n;
  assign o_0r0d[6] = go_0n;
  assign o_0r0d[8] = go_0n;
  assign o_0r0d[7] = gnd;
  assign o_0r1d[7] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_9_l25__28_28num_209_20256_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [8:0] o_0r0d;
  output [8:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[0] = gnd;
  assign o_0r1d[1] = gnd;
  assign o_0r1d[2] = gnd;
  assign o_0r1d[3] = gnd;
  assign o_0r1d[4] = gnd;
  assign o_0r1d[5] = gnd;
  assign o_0r1d[6] = gnd;
  assign o_0r1d[7] = gnd;
  assign o_0r0d[0] = go_0n;
  assign o_0r0d[1] = go_0n;
  assign o_0r0d[2] = go_0n;
  assign o_0r0d[3] = go_0n;
  assign o_0r0d[4] = go_0n;
  assign o_0r0d[5] = go_0n;
  assign o_0r0d[6] = go_0n;
  assign o_0r0d[7] = go_0n;
  assign o_0r0d[8] = gnd;
  assign o_0r1d[8] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_10_l26__28_28num_2010_20256_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [9:0] o_0r0d;
  output [9:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[0] = gnd;
  assign o_0r1d[1] = gnd;
  assign o_0r1d[2] = gnd;
  assign o_0r1d[3] = gnd;
  assign o_0r1d[4] = gnd;
  assign o_0r1d[5] = gnd;
  assign o_0r1d[6] = gnd;
  assign o_0r1d[7] = gnd;
  assign o_0r1d[9] = gnd;
  assign o_0r0d[0] = go_0n;
  assign o_0r0d[1] = go_0n;
  assign o_0r0d[2] = go_0n;
  assign o_0r0d[3] = go_0n;
  assign o_0r0d[4] = go_0n;
  assign o_0r0d[5] = go_0n;
  assign o_0r0d[6] = go_0n;
  assign o_0r0d[7] = go_0n;
  assign o_0r0d[9] = go_0n;
  assign o_0r0d[8] = gnd;
  assign o_0r1d[8] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_32_l24__28_28num_2032_200_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [31:0] o_0r0d;
  output [31:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[0] = gnd;
  assign o_0r1d[1] = gnd;
  assign o_0r1d[2] = gnd;
  assign o_0r1d[3] = gnd;
  assign o_0r1d[4] = gnd;
  assign o_0r1d[5] = gnd;
  assign o_0r1d[6] = gnd;
  assign o_0r1d[7] = gnd;
  assign o_0r1d[8] = gnd;
  assign o_0r1d[9] = gnd;
  assign o_0r1d[10] = gnd;
  assign o_0r1d[11] = gnd;
  assign o_0r1d[12] = gnd;
  assign o_0r1d[13] = gnd;
  assign o_0r1d[14] = gnd;
  assign o_0r1d[15] = gnd;
  assign o_0r1d[16] = gnd;
  assign o_0r1d[17] = gnd;
  assign o_0r1d[18] = gnd;
  assign o_0r1d[19] = gnd;
  assign o_0r1d[20] = gnd;
  assign o_0r1d[21] = gnd;
  assign o_0r1d[22] = gnd;
  assign o_0r1d[23] = gnd;
  assign o_0r1d[24] = gnd;
  assign o_0r1d[25] = gnd;
  assign o_0r1d[26] = gnd;
  assign o_0r1d[27] = gnd;
  assign o_0r1d[28] = gnd;
  assign o_0r1d[29] = gnd;
  assign o_0r1d[30] = gnd;
  assign o_0r1d[31] = gnd;
  assign o_0r0d[0] = go_0n;
  assign o_0r0d[1] = go_0n;
  assign o_0r0d[2] = go_0n;
  assign o_0r0d[3] = go_0n;
  assign o_0r0d[4] = go_0n;
  assign o_0r0d[5] = go_0n;
  assign o_0r0d[6] = go_0n;
  assign o_0r0d[7] = go_0n;
  assign o_0r0d[8] = go_0n;
  assign o_0r0d[9] = go_0n;
  assign o_0r0d[10] = go_0n;
  assign o_0r0d[11] = go_0n;
  assign o_0r0d[12] = go_0n;
  assign o_0r0d[13] = go_0n;
  assign o_0r0d[14] = go_0n;
  assign o_0r0d[15] = go_0n;
  assign o_0r0d[16] = go_0n;
  assign o_0r0d[17] = go_0n;
  assign o_0r0d[18] = go_0n;
  assign o_0r0d[19] = go_0n;
  assign o_0r0d[20] = go_0n;
  assign o_0r0d[21] = go_0n;
  assign o_0r0d[22] = go_0n;
  assign o_0r0d[23] = go_0n;
  assign o_0r0d[24] = go_0n;
  assign o_0r0d[25] = go_0n;
  assign o_0r0d[26] = go_0n;
  assign o_0r0d[27] = go_0n;
  assign o_0r0d[28] = go_0n;
  assign o_0r0d[29] = go_0n;
  assign o_0r0d[30] = go_0n;
  assign o_0r0d[31] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_35_l24__28_28num_2035_200_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [34:0] o_0r0d;
  output [34:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[0] = gnd;
  assign o_0r1d[1] = gnd;
  assign o_0r1d[2] = gnd;
  assign o_0r1d[3] = gnd;
  assign o_0r1d[4] = gnd;
  assign o_0r1d[5] = gnd;
  assign o_0r1d[6] = gnd;
  assign o_0r1d[7] = gnd;
  assign o_0r1d[8] = gnd;
  assign o_0r1d[9] = gnd;
  assign o_0r1d[10] = gnd;
  assign o_0r1d[11] = gnd;
  assign o_0r1d[12] = gnd;
  assign o_0r1d[13] = gnd;
  assign o_0r1d[14] = gnd;
  assign o_0r1d[15] = gnd;
  assign o_0r1d[16] = gnd;
  assign o_0r1d[17] = gnd;
  assign o_0r1d[18] = gnd;
  assign o_0r1d[19] = gnd;
  assign o_0r1d[20] = gnd;
  assign o_0r1d[21] = gnd;
  assign o_0r1d[22] = gnd;
  assign o_0r1d[23] = gnd;
  assign o_0r1d[24] = gnd;
  assign o_0r1d[25] = gnd;
  assign o_0r1d[26] = gnd;
  assign o_0r1d[27] = gnd;
  assign o_0r1d[28] = gnd;
  assign o_0r1d[29] = gnd;
  assign o_0r1d[30] = gnd;
  assign o_0r1d[31] = gnd;
  assign o_0r1d[32] = gnd;
  assign o_0r1d[33] = gnd;
  assign o_0r1d[34] = gnd;
  assign o_0r0d[0] = go_0n;
  assign o_0r0d[1] = go_0n;
  assign o_0r0d[2] = go_0n;
  assign o_0r0d[3] = go_0n;
  assign o_0r0d[4] = go_0n;
  assign o_0r0d[5] = go_0n;
  assign o_0r0d[6] = go_0n;
  assign o_0r0d[7] = go_0n;
  assign o_0r0d[8] = go_0n;
  assign o_0r0d[9] = go_0n;
  assign o_0r0d[10] = go_0n;
  assign o_0r0d[11] = go_0n;
  assign o_0r0d[12] = go_0n;
  assign o_0r0d[13] = go_0n;
  assign o_0r0d[14] = go_0n;
  assign o_0r0d[15] = go_0n;
  assign o_0r0d[16] = go_0n;
  assign o_0r0d[17] = go_0n;
  assign o_0r0d[18] = go_0n;
  assign o_0r0d[19] = go_0n;
  assign o_0r0d[20] = go_0n;
  assign o_0r0d[21] = go_0n;
  assign o_0r0d[22] = go_0n;
  assign o_0r0d[23] = go_0n;
  assign o_0r0d[24] = go_0n;
  assign o_0r0d[25] = go_0n;
  assign o_0r0d[26] = go_0n;
  assign o_0r0d[27] = go_0n;
  assign o_0r0d[28] = go_0n;
  assign o_0r0d[29] = go_0n;
  assign o_0r0d[30] = go_0n;
  assign o_0r0d[31] = go_0n;
  assign o_0r0d[32] = go_0n;
  assign o_0r0d[33] = go_0n;
  assign o_0r0d[34] = go_0n;
  assign go_0n = i_0r;
endmodule

module BrzO_0_36_l24__28_28num_2036_200_29_29 (
  i_0r, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input i_0r;
  output i_0a;
  output [35:0] o_0r0d;
  output [35:0] o_0r1d;
  input o_0a;
  wire go_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[0] = gnd;
  assign o_0r1d[1] = gnd;
  assign o_0r1d[2] = gnd;
  assign o_0r1d[3] = gnd;
  assign o_0r1d[4] = gnd;
  assign o_0r1d[5] = gnd;
  assign o_0r1d[6] = gnd;
  assign o_0r1d[7] = gnd;
  assign o_0r1d[8] = gnd;
  assign o_0r1d[9] = gnd;
  assign o_0r1d[10] = gnd;
  assign o_0r1d[11] = gnd;
  assign o_0r1d[12] = gnd;
  assign o_0r1d[13] = gnd;
  assign o_0r1d[14] = gnd;
  assign o_0r1d[15] = gnd;
  assign o_0r1d[16] = gnd;
  assign o_0r1d[17] = gnd;
  assign o_0r1d[18] = gnd;
  assign o_0r1d[19] = gnd;
  assign o_0r1d[20] = gnd;
  assign o_0r1d[21] = gnd;
  assign o_0r1d[22] = gnd;
  assign o_0r1d[23] = gnd;
  assign o_0r1d[24] = gnd;
  assign o_0r1d[25] = gnd;
  assign o_0r1d[26] = gnd;
  assign o_0r1d[27] = gnd;
  assign o_0r1d[28] = gnd;
  assign o_0r1d[29] = gnd;
  assign o_0r1d[30] = gnd;
  assign o_0r1d[31] = gnd;
  assign o_0r1d[32] = gnd;
  assign o_0r1d[33] = gnd;
  assign o_0r1d[34] = gnd;
  assign o_0r1d[35] = gnd;
  assign o_0r0d[0] = go_0n;
  assign o_0r0d[1] = go_0n;
  assign o_0r0d[2] = go_0n;
  assign o_0r0d[3] = go_0n;
  assign o_0r0d[4] = go_0n;
  assign o_0r0d[5] = go_0n;
  assign o_0r0d[6] = go_0n;
  assign o_0r0d[7] = go_0n;
  assign o_0r0d[8] = go_0n;
  assign o_0r0d[9] = go_0n;
  assign o_0r0d[10] = go_0n;
  assign o_0r0d[11] = go_0n;
  assign o_0r0d[12] = go_0n;
  assign o_0r0d[13] = go_0n;
  assign o_0r0d[14] = go_0n;
  assign o_0r0d[15] = go_0n;
  assign o_0r0d[16] = go_0n;
  assign o_0r0d[17] = go_0n;
  assign o_0r0d[18] = go_0n;
  assign o_0r0d[19] = go_0n;
  assign o_0r0d[20] = go_0n;
  assign o_0r0d[21] = go_0n;
  assign o_0r0d[22] = go_0n;
  assign o_0r0d[23] = go_0n;
  assign o_0r0d[24] = go_0n;
  assign o_0r0d[25] = go_0n;
  assign o_0r0d[26] = go_0n;
  assign o_0r0d[27] = go_0n;
  assign o_0r0d[28] = go_0n;
  assign o_0r0d[29] = go_0n;
  assign o_0r0d[30] = go_0n;
  assign o_0r0d[31] = go_0n;
  assign o_0r0d[32] = go_0n;
  assign o_0r0d[33] = go_0n;
  assign o_0r0d[34] = go_0n;
  assign o_0r0d[35] = go_0n;
  assign go_0n = i_0r;
endmodule

module DRAND2 (
  i0_0,
  i0_1,
  i1_0,
  i1_1,
  q_0,
  q_1
);
  input i0_0;
  input i0_1;
  input i1_0;
  input i1_1;
  output q_0;
  output q_1;
  wire n0_0n;
  wire n1_0n;
  wire n2_0n;
  OR3 I0 (q_0, n0_0n, n1_0n, n2_0n);
  C2 I1 (n0_0n, i0_0, i1_0);
  C2 I2 (n1_0n, i0_0, i1_1);
  C2 I3 (n2_0n, i0_1, i1_0);
  C2 I4 (q_1, i0_1, i1_1);
endmodule

module BrzO_2_1_l119__28_28app_201_20_280_200_201_m47m (
  i_0r0d, i_0r1d, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input [1:0] i_0r0d;
  input [1:0] i_0r1d;
  output i_0a;
  output o_0r0d;
  output o_0r1d;
  input o_0a;
  wire termf_0n;
  wire termf_1n;
  wire termt_0n;
  wire termt_1n;
  assign i_0a = o_0a;
  DRAND2 I1 (termf_0n, termt_0n, termf_1n, termt_1n, o_0r0d, o_0r1d);
  assign termt_1n = i_0r1d[1];
  assign termf_1n = i_0r0d[1];
  assign termt_0n = i_0r1d[0];
  assign termf_0n = i_0r0d[0];
endmodule

module BrzO_4_35_l91__28_28app_2031_20_280_203_20_m48m (
  i_0r0d, i_0r1d, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input [3:0] i_0r0d;
  input [3:0] i_0r1d;
  output i_0a;
  output [34:0] o_0r0d;
  output [34:0] o_0r1d;
  input o_0a;
  wire [30:0] termf_0n;
  wire [30:0] termt_0n;
  assign i_0a = o_0a;
  assign o_0r1d[4] = termt_0n[0];
  assign o_0r1d[5] = termt_0n[1];
  assign o_0r1d[6] = termt_0n[2];
  assign o_0r1d[7] = termt_0n[3];
  assign o_0r1d[8] = termt_0n[4];
  assign o_0r1d[9] = termt_0n[5];
  assign o_0r1d[10] = termt_0n[6];
  assign o_0r1d[11] = termt_0n[7];
  assign o_0r1d[12] = termt_0n[8];
  assign o_0r1d[13] = termt_0n[9];
  assign o_0r1d[14] = termt_0n[10];
  assign o_0r1d[15] = termt_0n[11];
  assign o_0r1d[16] = termt_0n[12];
  assign o_0r1d[17] = termt_0n[13];
  assign o_0r1d[18] = termt_0n[14];
  assign o_0r1d[19] = termt_0n[15];
  assign o_0r1d[20] = termt_0n[16];
  assign o_0r1d[21] = termt_0n[17];
  assign o_0r1d[22] = termt_0n[18];
  assign o_0r1d[23] = termt_0n[19];
  assign o_0r1d[24] = termt_0n[20];
  assign o_0r1d[25] = termt_0n[21];
  assign o_0r1d[26] = termt_0n[22];
  assign o_0r1d[27] = termt_0n[23];
  assign o_0r1d[28] = termt_0n[24];
  assign o_0r1d[29] = termt_0n[25];
  assign o_0r1d[30] = termt_0n[26];
  assign o_0r1d[31] = termt_0n[27];
  assign o_0r1d[32] = termt_0n[28];
  assign o_0r1d[33] = termt_0n[29];
  assign o_0r1d[34] = termt_0n[30];
  assign o_0r0d[4] = termf_0n[0];
  assign o_0r0d[5] = termf_0n[1];
  assign o_0r0d[6] = termf_0n[2];
  assign o_0r0d[7] = termf_0n[3];
  assign o_0r0d[8] = termf_0n[4];
  assign o_0r0d[9] = termf_0n[5];
  assign o_0r0d[10] = termf_0n[6];
  assign o_0r0d[11] = termf_0n[7];
  assign o_0r0d[12] = termf_0n[8];
  assign o_0r0d[13] = termf_0n[9];
  assign o_0r0d[14] = termf_0n[10];
  assign o_0r0d[15] = termf_0n[11];
  assign o_0r0d[16] = termf_0n[12];
  assign o_0r0d[17] = termf_0n[13];
  assign o_0r0d[18] = termf_0n[14];
  assign o_0r0d[19] = termf_0n[15];
  assign o_0r0d[20] = termf_0n[16];
  assign o_0r0d[21] = termf_0n[17];
  assign o_0r0d[22] = termf_0n[18];
  assign o_0r0d[23] = termf_0n[19];
  assign o_0r0d[24] = termf_0n[20];
  assign o_0r0d[25] = termf_0n[21];
  assign o_0r0d[26] = termf_0n[22];
  assign o_0r0d[27] = termf_0n[23];
  assign o_0r0d[28] = termf_0n[24];
  assign o_0r0d[29] = termf_0n[25];
  assign o_0r0d[30] = termf_0n[26];
  assign o_0r0d[31] = termf_0n[27];
  assign o_0r0d[32] = termf_0n[28];
  assign o_0r0d[33] = termf_0n[29];
  assign o_0r0d[34] = termf_0n[30];
  assign o_0r1d[0] = i_0r1d[0];
  assign o_0r1d[1] = i_0r1d[1];
  assign o_0r1d[2] = i_0r1d[2];
  assign o_0r1d[3] = i_0r1d[3];
  assign o_0r0d[0] = i_0r0d[0];
  assign o_0r0d[1] = i_0r0d[1];
  assign o_0r0d[2] = i_0r0d[2];
  assign o_0r0d[3] = i_0r0d[3];
  assign termt_0n[30] = i_0r1d[3];
  assign termf_0n[30] = i_0r0d[3];
  assign termt_0n[29] = i_0r1d[3];
  assign termf_0n[29] = i_0r0d[3];
  assign termt_0n[28] = i_0r1d[3];
  assign termf_0n[28] = i_0r0d[3];
  assign termt_0n[27] = i_0r1d[3];
  assign termf_0n[27] = i_0r0d[3];
  assign termt_0n[26] = i_0r1d[3];
  assign termf_0n[26] = i_0r0d[3];
  assign termt_0n[25] = i_0r1d[3];
  assign termf_0n[25] = i_0r0d[3];
  assign termt_0n[24] = i_0r1d[3];
  assign termf_0n[24] = i_0r0d[3];
  assign termt_0n[23] = i_0r1d[3];
  assign termf_0n[23] = i_0r0d[3];
  assign termt_0n[22] = i_0r1d[3];
  assign termf_0n[22] = i_0r0d[3];
  assign termt_0n[21] = i_0r1d[3];
  assign termf_0n[21] = i_0r0d[3];
  assign termt_0n[20] = i_0r1d[3];
  assign termf_0n[20] = i_0r0d[3];
  assign termt_0n[19] = i_0r1d[3];
  assign termf_0n[19] = i_0r0d[3];
  assign termt_0n[18] = i_0r1d[3];
  assign termf_0n[18] = i_0r0d[3];
  assign termt_0n[17] = i_0r1d[3];
  assign termf_0n[17] = i_0r0d[3];
  assign termt_0n[16] = i_0r1d[3];
  assign termf_0n[16] = i_0r0d[3];
  assign termt_0n[15] = i_0r1d[3];
  assign termf_0n[15] = i_0r0d[3];
  assign termt_0n[14] = i_0r1d[3];
  assign termf_0n[14] = i_0r0d[3];
  assign termt_0n[13] = i_0r1d[3];
  assign termf_0n[13] = i_0r0d[3];
  assign termt_0n[12] = i_0r1d[3];
  assign termf_0n[12] = i_0r0d[3];
  assign termt_0n[11] = i_0r1d[3];
  assign termf_0n[11] = i_0r0d[3];
  assign termt_0n[10] = i_0r1d[3];
  assign termf_0n[10] = i_0r0d[3];
  assign termt_0n[9] = i_0r1d[3];
  assign termf_0n[9] = i_0r0d[3];
  assign termt_0n[8] = i_0r1d[3];
  assign termf_0n[8] = i_0r0d[3];
  assign termt_0n[7] = i_0r1d[3];
  assign termf_0n[7] = i_0r0d[3];
  assign termt_0n[6] = i_0r1d[3];
  assign termf_0n[6] = i_0r0d[3];
  assign termt_0n[5] = i_0r1d[3];
  assign termf_0n[5] = i_0r0d[3];
  assign termt_0n[4] = i_0r1d[3];
  assign termf_0n[4] = i_0r0d[3];
  assign termt_0n[3] = i_0r1d[3];
  assign termf_0n[3] = i_0r0d[3];
  assign termt_0n[2] = i_0r1d[3];
  assign termf_0n[2] = i_0r0d[3];
  assign termt_0n[1] = i_0r1d[3];
  assign termf_0n[1] = i_0r0d[3];
  assign termt_0n[0] = i_0r1d[3];
  assign termf_0n[0] = i_0r0d[3];
endmodule

module BrzO_9_10_l75__28_28num_201_200_29_20_28ap_m49m (
  i_0r0d, i_0r1d, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input [8:0] i_0r0d;
  input [8:0] i_0r1d;
  output i_0a;
  output [9:0] o_0r0d;
  output [9:0] o_0r1d;
  input o_0a;
  wire go_0n;
  wire termf_0n;
  wire termt_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[9] = termt_0n;
  assign o_0r0d[9] = termf_0n;
  assign o_0r1d[0] = i_0r1d[0];
  assign o_0r1d[1] = i_0r1d[1];
  assign o_0r1d[2] = i_0r1d[2];
  assign o_0r1d[3] = i_0r1d[3];
  assign o_0r1d[4] = i_0r1d[4];
  assign o_0r1d[5] = i_0r1d[5];
  assign o_0r1d[6] = i_0r1d[6];
  assign o_0r1d[7] = i_0r1d[7];
  assign o_0r1d[8] = i_0r1d[8];
  assign o_0r0d[0] = i_0r0d[0];
  assign o_0r0d[1] = i_0r0d[1];
  assign o_0r0d[2] = i_0r0d[2];
  assign o_0r0d[3] = i_0r0d[3];
  assign o_0r0d[4] = i_0r0d[4];
  assign o_0r0d[5] = i_0r0d[5];
  assign o_0r0d[6] = i_0r0d[6];
  assign o_0r0d[7] = i_0r0d[7];
  assign o_0r0d[8] = i_0r0d[8];
  assign termt_0n = gnd;
  assign termf_0n = go_0n;
  OR2 I23 (go_0n, i_0r0d[0], i_0r1d[0]);
endmodule

module BrzO_32_35_l91__28_28app_203_20_280_2031_2_m50m (
  i_0r0d, i_0r1d, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input [31:0] i_0r0d;
  input [31:0] i_0r1d;
  output i_0a;
  output [34:0] o_0r0d;
  output [34:0] o_0r1d;
  input o_0a;
  wire [2:0] termf_0n;
  wire [2:0] termt_0n;
  assign i_0a = o_0a;
  assign o_0r1d[32] = termt_0n[0];
  assign o_0r1d[33] = termt_0n[1];
  assign o_0r1d[34] = termt_0n[2];
  assign o_0r0d[32] = termf_0n[0];
  assign o_0r0d[33] = termf_0n[1];
  assign o_0r0d[34] = termf_0n[2];
  assign o_0r1d[0] = i_0r1d[0];
  assign o_0r1d[1] = i_0r1d[1];
  assign o_0r1d[2] = i_0r1d[2];
  assign o_0r1d[3] = i_0r1d[3];
  assign o_0r1d[4] = i_0r1d[4];
  assign o_0r1d[5] = i_0r1d[5];
  assign o_0r1d[6] = i_0r1d[6];
  assign o_0r1d[7] = i_0r1d[7];
  assign o_0r1d[8] = i_0r1d[8];
  assign o_0r1d[9] = i_0r1d[9];
  assign o_0r1d[10] = i_0r1d[10];
  assign o_0r1d[11] = i_0r1d[11];
  assign o_0r1d[12] = i_0r1d[12];
  assign o_0r1d[13] = i_0r1d[13];
  assign o_0r1d[14] = i_0r1d[14];
  assign o_0r1d[15] = i_0r1d[15];
  assign o_0r1d[16] = i_0r1d[16];
  assign o_0r1d[17] = i_0r1d[17];
  assign o_0r1d[18] = i_0r1d[18];
  assign o_0r1d[19] = i_0r1d[19];
  assign o_0r1d[20] = i_0r1d[20];
  assign o_0r1d[21] = i_0r1d[21];
  assign o_0r1d[22] = i_0r1d[22];
  assign o_0r1d[23] = i_0r1d[23];
  assign o_0r1d[24] = i_0r1d[24];
  assign o_0r1d[25] = i_0r1d[25];
  assign o_0r1d[26] = i_0r1d[26];
  assign o_0r1d[27] = i_0r1d[27];
  assign o_0r1d[28] = i_0r1d[28];
  assign o_0r1d[29] = i_0r1d[29];
  assign o_0r1d[30] = i_0r1d[30];
  assign o_0r1d[31] = i_0r1d[31];
  assign o_0r0d[0] = i_0r0d[0];
  assign o_0r0d[1] = i_0r0d[1];
  assign o_0r0d[2] = i_0r0d[2];
  assign o_0r0d[3] = i_0r0d[3];
  assign o_0r0d[4] = i_0r0d[4];
  assign o_0r0d[5] = i_0r0d[5];
  assign o_0r0d[6] = i_0r0d[6];
  assign o_0r0d[7] = i_0r0d[7];
  assign o_0r0d[8] = i_0r0d[8];
  assign o_0r0d[9] = i_0r0d[9];
  assign o_0r0d[10] = i_0r0d[10];
  assign o_0r0d[11] = i_0r0d[11];
  assign o_0r0d[12] = i_0r0d[12];
  assign o_0r0d[13] = i_0r0d[13];
  assign o_0r0d[14] = i_0r0d[14];
  assign o_0r0d[15] = i_0r0d[15];
  assign o_0r0d[16] = i_0r0d[16];
  assign o_0r0d[17] = i_0r0d[17];
  assign o_0r0d[18] = i_0r0d[18];
  assign o_0r0d[19] = i_0r0d[19];
  assign o_0r0d[20] = i_0r0d[20];
  assign o_0r0d[21] = i_0r0d[21];
  assign o_0r0d[22] = i_0r0d[22];
  assign o_0r0d[23] = i_0r0d[23];
  assign o_0r0d[24] = i_0r0d[24];
  assign o_0r0d[25] = i_0r0d[25];
  assign o_0r0d[26] = i_0r0d[26];
  assign o_0r0d[27] = i_0r0d[27];
  assign o_0r0d[28] = i_0r0d[28];
  assign o_0r0d[29] = i_0r0d[29];
  assign o_0r0d[30] = i_0r0d[30];
  assign o_0r0d[31] = i_0r0d[31];
  assign termt_0n[2] = i_0r1d[31];
  assign termf_0n[2] = i_0r0d[31];
  assign termt_0n[1] = i_0r1d[31];
  assign termf_0n[1] = i_0r0d[31];
  assign termt_0n[0] = i_0r1d[31];
  assign termf_0n[0] = i_0r0d[31];
endmodule

module BrzO_32_35_l76__28_28num_203_200_29_20_28a_m51m (
  i_0r0d, i_0r1d, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input [31:0] i_0r0d;
  input [31:0] i_0r1d;
  output i_0a;
  output [34:0] o_0r0d;
  output [34:0] o_0r1d;
  input o_0a;
  wire go_0n;
  wire [2:0] termf_0n;
  wire [2:0] termt_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[32] = termt_0n[0];
  assign o_0r1d[33] = termt_0n[1];
  assign o_0r1d[34] = termt_0n[2];
  assign o_0r0d[32] = termf_0n[0];
  assign o_0r0d[33] = termf_0n[1];
  assign o_0r0d[34] = termf_0n[2];
  assign o_0r1d[0] = i_0r1d[0];
  assign o_0r1d[1] = i_0r1d[1];
  assign o_0r1d[2] = i_0r1d[2];
  assign o_0r1d[3] = i_0r1d[3];
  assign o_0r1d[4] = i_0r1d[4];
  assign o_0r1d[5] = i_0r1d[5];
  assign o_0r1d[6] = i_0r1d[6];
  assign o_0r1d[7] = i_0r1d[7];
  assign o_0r1d[8] = i_0r1d[8];
  assign o_0r1d[9] = i_0r1d[9];
  assign o_0r1d[10] = i_0r1d[10];
  assign o_0r1d[11] = i_0r1d[11];
  assign o_0r1d[12] = i_0r1d[12];
  assign o_0r1d[13] = i_0r1d[13];
  assign o_0r1d[14] = i_0r1d[14];
  assign o_0r1d[15] = i_0r1d[15];
  assign o_0r1d[16] = i_0r1d[16];
  assign o_0r1d[17] = i_0r1d[17];
  assign o_0r1d[18] = i_0r1d[18];
  assign o_0r1d[19] = i_0r1d[19];
  assign o_0r1d[20] = i_0r1d[20];
  assign o_0r1d[21] = i_0r1d[21];
  assign o_0r1d[22] = i_0r1d[22];
  assign o_0r1d[23] = i_0r1d[23];
  assign o_0r1d[24] = i_0r1d[24];
  assign o_0r1d[25] = i_0r1d[25];
  assign o_0r1d[26] = i_0r1d[26];
  assign o_0r1d[27] = i_0r1d[27];
  assign o_0r1d[28] = i_0r1d[28];
  assign o_0r1d[29] = i_0r1d[29];
  assign o_0r1d[30] = i_0r1d[30];
  assign o_0r1d[31] = i_0r1d[31];
  assign o_0r0d[0] = i_0r0d[0];
  assign o_0r0d[1] = i_0r0d[1];
  assign o_0r0d[2] = i_0r0d[2];
  assign o_0r0d[3] = i_0r0d[3];
  assign o_0r0d[4] = i_0r0d[4];
  assign o_0r0d[5] = i_0r0d[5];
  assign o_0r0d[6] = i_0r0d[6];
  assign o_0r0d[7] = i_0r0d[7];
  assign o_0r0d[8] = i_0r0d[8];
  assign o_0r0d[9] = i_0r0d[9];
  assign o_0r0d[10] = i_0r0d[10];
  assign o_0r0d[11] = i_0r0d[11];
  assign o_0r0d[12] = i_0r0d[12];
  assign o_0r0d[13] = i_0r0d[13];
  assign o_0r0d[14] = i_0r0d[14];
  assign o_0r0d[15] = i_0r0d[15];
  assign o_0r0d[16] = i_0r0d[16];
  assign o_0r0d[17] = i_0r0d[17];
  assign o_0r0d[18] = i_0r0d[18];
  assign o_0r0d[19] = i_0r0d[19];
  assign o_0r0d[20] = i_0r0d[20];
  assign o_0r0d[21] = i_0r0d[21];
  assign o_0r0d[22] = i_0r0d[22];
  assign o_0r0d[23] = i_0r0d[23];
  assign o_0r0d[24] = i_0r0d[24];
  assign o_0r0d[25] = i_0r0d[25];
  assign o_0r0d[26] = i_0r0d[26];
  assign o_0r0d[27] = i_0r0d[27];
  assign o_0r0d[28] = i_0r0d[28];
  assign o_0r0d[29] = i_0r0d[29];
  assign o_0r0d[30] = i_0r0d[30];
  assign o_0r0d[31] = i_0r0d[31];
  assign termt_0n[0] = gnd;
  assign termt_0n[1] = gnd;
  assign termt_0n[2] = gnd;
  assign termf_0n[0] = go_0n;
  assign termf_0n[1] = go_0n;
  assign termf_0n[2] = go_0n;
  OR2 I77 (go_0n, i_0r0d[0], i_0r1d[0]);
endmodule

module DRXOR2 (
  i0_0,
  i0_1,
  i1_0,
  i1_1,
  q_0,
  q_1
);
  input i0_0;
  input i0_1;
  input i1_0;
  input i1_1;
  output q_0;
  output q_1;
  wire n0_0n;
  wire n1_0n;
  wire n2_0n;
  wire n3_0n;
  OR2 I0 (q_0, n0_0n, n3_0n);
  C2 I1 (n3_0n, i0_1, i1_1);
  C2 I2 (n0_0n, i0_0, i1_0);
  OR2 I3 (q_1, n1_0n, n2_0n);
  C2 I4 (n1_0n, i0_0, i1_1);
  C2 I5 (n2_0n, i0_1, i1_0);
endmodule

module BrzO_33_1_l196__28_28app_201_20_280_200_20_m52m (
  i_0r0d, i_0r1d, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input [32:0] i_0r0d;
  input [32:0] i_0r1d;
  output i_0a;
  output o_0r0d;
  output o_0r1d;
  input o_0a;
  wire go_0n;
  wire [31:0] termf_0n;
  wire termf_1n;
  wire [30:0] termf_2n;
  wire [31:0] termf_3n;
  wire [31:0] termt_0n;
  wire termt_1n;
  wire [30:0] termt_2n;
  wire [31:0] termt_3n;
  wire [1:0] drr968__1_0n;
  wire [1:0] drr967__0_0n;
  wire [1:0] drr970__1_0n;
  wire [1:0] drr969__0_0n;
  wire [1:0] drr966__1_0n;
  wire [1:0] drr965__0_0n;
  wire [1:0] drr974__1_0n;
  wire [1:0] drr973__0_0n;
  wire [1:0] drr976__1_0n;
  wire [1:0] drr975__0_0n;
  wire [1:0] drr972__1_0n;
  wire [1:0] drr971__0_0n;
  wire [1:0] drr964__1_0n;
  wire [1:0] drr963__0_0n;
  wire [1:0] drr982__1_0n;
  wire [1:0] drr981__0_0n;
  wire [1:0] drr984__1_0n;
  wire [1:0] drr983__0_0n;
  wire [1:0] drr980__1_0n;
  wire [1:0] drr979__0_0n;
  wire [1:0] drr988__1_0n;
  wire [1:0] drr987__0_0n;
  wire [1:0] drr990__1_0n;
  wire [1:0] drr989__0_0n;
  wire [1:0] drr986__1_0n;
  wire [1:0] drr985__0_0n;
  wire [1:0] drr978__1_0n;
  wire [1:0] drr977__0_0n;
  wire [1:0] drr962__1_0n;
  wire [1:0] drr961__0_0n;
  wire [31:0] eqf5_0n;
  wire [31:0] eqt5_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  DRAND2 I1 (drr961__0_0n[0], drr962__1_0n[0], drr961__0_0n[1], drr962__1_0n[1], o_0r0d, o_0r1d);
  DRAND2 I2 (drr963__0_0n[0], drr964__1_0n[0], drr963__0_0n[1], drr964__1_0n[1], drr961__0_0n[1], drr962__1_0n[1]);
  DRAND2 I3 (drr965__0_0n[0], drr966__1_0n[0], drr965__0_0n[1], drr966__1_0n[1], drr963__0_0n[1], drr964__1_0n[1]);
  DRAND2 I4 (drr967__0_0n[0], drr968__1_0n[0], drr967__0_0n[1], drr968__1_0n[1], drr965__0_0n[1], drr966__1_0n[1]);
  DRAND2 I5 (eqt5_0n[30], eqf5_0n[30], eqt5_0n[31], eqf5_0n[31], drr967__0_0n[1], drr968__1_0n[1]);
  DRAND2 I6 (eqt5_0n[28], eqf5_0n[28], eqt5_0n[29], eqf5_0n[29], drr967__0_0n[0], drr968__1_0n[0]);
  DRAND2 I7 (drr969__0_0n[0], drr970__1_0n[0], drr969__0_0n[1], drr970__1_0n[1], drr965__0_0n[0], drr966__1_0n[0]);
  DRAND2 I8 (eqt5_0n[26], eqf5_0n[26], eqt5_0n[27], eqf5_0n[27], drr969__0_0n[1], drr970__1_0n[1]);
  DRAND2 I9 (eqt5_0n[24], eqf5_0n[24], eqt5_0n[25], eqf5_0n[25], drr969__0_0n[0], drr970__1_0n[0]);
  DRAND2 I10 (drr971__0_0n[0], drr972__1_0n[0], drr971__0_0n[1], drr972__1_0n[1], drr963__0_0n[0], drr964__1_0n[0]);
  DRAND2 I11 (drr973__0_0n[0], drr974__1_0n[0], drr973__0_0n[1], drr974__1_0n[1], drr971__0_0n[1], drr972__1_0n[1]);
  DRAND2 I12 (eqt5_0n[22], eqf5_0n[22], eqt5_0n[23], eqf5_0n[23], drr973__0_0n[1], drr974__1_0n[1]);
  DRAND2 I13 (eqt5_0n[20], eqf5_0n[20], eqt5_0n[21], eqf5_0n[21], drr973__0_0n[0], drr974__1_0n[0]);
  DRAND2 I14 (drr975__0_0n[0], drr976__1_0n[0], drr975__0_0n[1], drr976__1_0n[1], drr971__0_0n[0], drr972__1_0n[0]);
  DRAND2 I15 (eqt5_0n[18], eqf5_0n[18], eqt5_0n[19], eqf5_0n[19], drr975__0_0n[1], drr976__1_0n[1]);
  DRAND2 I16 (eqt5_0n[16], eqf5_0n[16], eqt5_0n[17], eqf5_0n[17], drr975__0_0n[0], drr976__1_0n[0]);
  DRAND2 I17 (drr977__0_0n[0], drr978__1_0n[0], drr977__0_0n[1], drr978__1_0n[1], drr961__0_0n[0], drr962__1_0n[0]);
  DRAND2 I18 (drr979__0_0n[0], drr980__1_0n[0], drr979__0_0n[1], drr980__1_0n[1], drr977__0_0n[1], drr978__1_0n[1]);
  DRAND2 I19 (drr981__0_0n[0], drr982__1_0n[0], drr981__0_0n[1], drr982__1_0n[1], drr979__0_0n[1], drr980__1_0n[1]);
  DRAND2 I20 (eqt5_0n[14], eqf5_0n[14], eqt5_0n[15], eqf5_0n[15], drr981__0_0n[1], drr982__1_0n[1]);
  DRAND2 I21 (eqt5_0n[12], eqf5_0n[12], eqt5_0n[13], eqf5_0n[13], drr981__0_0n[0], drr982__1_0n[0]);
  DRAND2 I22 (drr983__0_0n[0], drr984__1_0n[0], drr983__0_0n[1], drr984__1_0n[1], drr979__0_0n[0], drr980__1_0n[0]);
  DRAND2 I23 (eqt5_0n[10], eqf5_0n[10], eqt5_0n[11], eqf5_0n[11], drr983__0_0n[1], drr984__1_0n[1]);
  DRAND2 I24 (eqt5_0n[8], eqf5_0n[8], eqt5_0n[9], eqf5_0n[9], drr983__0_0n[0], drr984__1_0n[0]);
  DRAND2 I25 (drr985__0_0n[0], drr986__1_0n[0], drr985__0_0n[1], drr986__1_0n[1], drr977__0_0n[0], drr978__1_0n[0]);
  DRAND2 I26 (drr987__0_0n[0], drr988__1_0n[0], drr987__0_0n[1], drr988__1_0n[1], drr985__0_0n[1], drr986__1_0n[1]);
  DRAND2 I27 (eqt5_0n[6], eqf5_0n[6], eqt5_0n[7], eqf5_0n[7], drr987__0_0n[1], drr988__1_0n[1]);
  DRAND2 I28 (eqt5_0n[4], eqf5_0n[4], eqt5_0n[5], eqf5_0n[5], drr987__0_0n[0], drr988__1_0n[0]);
  DRAND2 I29 (drr989__0_0n[0], drr990__1_0n[0], drr989__0_0n[1], drr990__1_0n[1], drr985__0_0n[0], drr986__1_0n[0]);
  DRAND2 I30 (eqt5_0n[2], eqf5_0n[2], eqt5_0n[3], eqf5_0n[3], drr989__0_0n[1], drr990__1_0n[1]);
  DRAND2 I31 (eqt5_0n[0], eqf5_0n[0], eqt5_0n[1], eqf5_0n[1], drr989__0_0n[0], drr990__1_0n[0]);
  DRXOR2 I32 (termf_0n[0], termt_0n[0], termf_3n[0], termt_3n[0], eqf5_0n[0], eqt5_0n[0]);
  DRXOR2 I33 (termf_0n[1], termt_0n[1], termf_3n[1], termt_3n[1], eqf5_0n[1], eqt5_0n[1]);
  DRXOR2 I34 (termf_0n[2], termt_0n[2], termf_3n[2], termt_3n[2], eqf5_0n[2], eqt5_0n[2]);
  DRXOR2 I35 (termf_0n[3], termt_0n[3], termf_3n[3], termt_3n[3], eqf5_0n[3], eqt5_0n[3]);
  DRXOR2 I36 (termf_0n[4], termt_0n[4], termf_3n[4], termt_3n[4], eqf5_0n[4], eqt5_0n[4]);
  DRXOR2 I37 (termf_0n[5], termt_0n[5], termf_3n[5], termt_3n[5], eqf5_0n[5], eqt5_0n[5]);
  DRXOR2 I38 (termf_0n[6], termt_0n[6], termf_3n[6], termt_3n[6], eqf5_0n[6], eqt5_0n[6]);
  DRXOR2 I39 (termf_0n[7], termt_0n[7], termf_3n[7], termt_3n[7], eqf5_0n[7], eqt5_0n[7]);
  DRXOR2 I40 (termf_0n[8], termt_0n[8], termf_3n[8], termt_3n[8], eqf5_0n[8], eqt5_0n[8]);
  DRXOR2 I41 (termf_0n[9], termt_0n[9], termf_3n[9], termt_3n[9], eqf5_0n[9], eqt5_0n[9]);
  DRXOR2 I42 (termf_0n[10], termt_0n[10], termf_3n[10], termt_3n[10], eqf5_0n[10], eqt5_0n[10]);
  DRXOR2 I43 (termf_0n[11], termt_0n[11], termf_3n[11], termt_3n[11], eqf5_0n[11], eqt5_0n[11]);
  DRXOR2 I44 (termf_0n[12], termt_0n[12], termf_3n[12], termt_3n[12], eqf5_0n[12], eqt5_0n[12]);
  DRXOR2 I45 (termf_0n[13], termt_0n[13], termf_3n[13], termt_3n[13], eqf5_0n[13], eqt5_0n[13]);
  DRXOR2 I46 (termf_0n[14], termt_0n[14], termf_3n[14], termt_3n[14], eqf5_0n[14], eqt5_0n[14]);
  DRXOR2 I47 (termf_0n[15], termt_0n[15], termf_3n[15], termt_3n[15], eqf5_0n[15], eqt5_0n[15]);
  DRXOR2 I48 (termf_0n[16], termt_0n[16], termf_3n[16], termt_3n[16], eqf5_0n[16], eqt5_0n[16]);
  DRXOR2 I49 (termf_0n[17], termt_0n[17], termf_3n[17], termt_3n[17], eqf5_0n[17], eqt5_0n[17]);
  DRXOR2 I50 (termf_0n[18], termt_0n[18], termf_3n[18], termt_3n[18], eqf5_0n[18], eqt5_0n[18]);
  DRXOR2 I51 (termf_0n[19], termt_0n[19], termf_3n[19], termt_3n[19], eqf5_0n[19], eqt5_0n[19]);
  DRXOR2 I52 (termf_0n[20], termt_0n[20], termf_3n[20], termt_3n[20], eqf5_0n[20], eqt5_0n[20]);
  DRXOR2 I53 (termf_0n[21], termt_0n[21], termf_3n[21], termt_3n[21], eqf5_0n[21], eqt5_0n[21]);
  DRXOR2 I54 (termf_0n[22], termt_0n[22], termf_3n[22], termt_3n[22], eqf5_0n[22], eqt5_0n[22]);
  DRXOR2 I55 (termf_0n[23], termt_0n[23], termf_3n[23], termt_3n[23], eqf5_0n[23], eqt5_0n[23]);
  DRXOR2 I56 (termf_0n[24], termt_0n[24], termf_3n[24], termt_3n[24], eqf5_0n[24], eqt5_0n[24]);
  DRXOR2 I57 (termf_0n[25], termt_0n[25], termf_3n[25], termt_3n[25], eqf5_0n[25], eqt5_0n[25]);
  DRXOR2 I58 (termf_0n[26], termt_0n[26], termf_3n[26], termt_3n[26], eqf5_0n[26], eqt5_0n[26]);
  DRXOR2 I59 (termf_0n[27], termt_0n[27], termf_3n[27], termt_3n[27], eqf5_0n[27], eqt5_0n[27]);
  DRXOR2 I60 (termf_0n[28], termt_0n[28], termf_3n[28], termt_3n[28], eqf5_0n[28], eqt5_0n[28]);
  DRXOR2 I61 (termf_0n[29], termt_0n[29], termf_3n[29], termt_3n[29], eqf5_0n[29], eqt5_0n[29]);
  DRXOR2 I62 (termf_0n[30], termt_0n[30], termf_3n[30], termt_3n[30], eqf5_0n[30], eqt5_0n[30]);
  DRXOR2 I63 (termf_0n[31], termt_0n[31], termf_3n[31], termt_3n[31], eqf5_0n[31], eqt5_0n[31]);
  assign termt_3n[1] = termt_2n[0];
  assign termt_3n[2] = termt_2n[1];
  assign termt_3n[3] = termt_2n[2];
  assign termt_3n[4] = termt_2n[3];
  assign termt_3n[5] = termt_2n[4];
  assign termt_3n[6] = termt_2n[5];
  assign termt_3n[7] = termt_2n[6];
  assign termt_3n[8] = termt_2n[7];
  assign termt_3n[9] = termt_2n[8];
  assign termt_3n[10] = termt_2n[9];
  assign termt_3n[11] = termt_2n[10];
  assign termt_3n[12] = termt_2n[11];
  assign termt_3n[13] = termt_2n[12];
  assign termt_3n[14] = termt_2n[13];
  assign termt_3n[15] = termt_2n[14];
  assign termt_3n[16] = termt_2n[15];
  assign termt_3n[17] = termt_2n[16];
  assign termt_3n[18] = termt_2n[17];
  assign termt_3n[19] = termt_2n[18];
  assign termt_3n[20] = termt_2n[19];
  assign termt_3n[21] = termt_2n[20];
  assign termt_3n[22] = termt_2n[21];
  assign termt_3n[23] = termt_2n[22];
  assign termt_3n[24] = termt_2n[23];
  assign termt_3n[25] = termt_2n[24];
  assign termt_3n[26] = termt_2n[25];
  assign termt_3n[27] = termt_2n[26];
  assign termt_3n[28] = termt_2n[27];
  assign termt_3n[29] = termt_2n[28];
  assign termt_3n[30] = termt_2n[29];
  assign termt_3n[31] = termt_2n[30];
  assign termf_3n[1] = termf_2n[0];
  assign termf_3n[2] = termf_2n[1];
  assign termf_3n[3] = termf_2n[2];
  assign termf_3n[4] = termf_2n[3];
  assign termf_3n[5] = termf_2n[4];
  assign termf_3n[6] = termf_2n[5];
  assign termf_3n[7] = termf_2n[6];
  assign termf_3n[8] = termf_2n[7];
  assign termf_3n[9] = termf_2n[8];
  assign termf_3n[10] = termf_2n[9];
  assign termf_3n[11] = termf_2n[10];
  assign termf_3n[12] = termf_2n[11];
  assign termf_3n[13] = termf_2n[12];
  assign termf_3n[14] = termf_2n[13];
  assign termf_3n[15] = termf_2n[14];
  assign termf_3n[16] = termf_2n[15];
  assign termf_3n[17] = termf_2n[16];
  assign termf_3n[18] = termf_2n[17];
  assign termf_3n[19] = termf_2n[18];
  assign termf_3n[20] = termf_2n[19];
  assign termf_3n[21] = termf_2n[20];
  assign termf_3n[22] = termf_2n[21];
  assign termf_3n[23] = termf_2n[22];
  assign termf_3n[24] = termf_2n[23];
  assign termf_3n[25] = termf_2n[24];
  assign termf_3n[26] = termf_2n[25];
  assign termf_3n[27] = termf_2n[26];
  assign termf_3n[28] = termf_2n[27];
  assign termf_3n[29] = termf_2n[28];
  assign termf_3n[30] = termf_2n[29];
  assign termf_3n[31] = termf_2n[30];
  assign termt_3n[0] = termt_1n;
  assign termf_3n[0] = termf_1n;
  assign termt_2n[0] = gnd;
  assign termt_2n[1] = gnd;
  assign termt_2n[2] = gnd;
  assign termt_2n[3] = gnd;
  assign termt_2n[4] = gnd;
  assign termt_2n[5] = gnd;
  assign termt_2n[6] = gnd;
  assign termt_2n[7] = gnd;
  assign termt_2n[8] = gnd;
  assign termt_2n[9] = gnd;
  assign termt_2n[10] = gnd;
  assign termt_2n[11] = gnd;
  assign termt_2n[12] = gnd;
  assign termt_2n[13] = gnd;
  assign termt_2n[14] = gnd;
  assign termt_2n[15] = gnd;
  assign termt_2n[16] = gnd;
  assign termt_2n[17] = gnd;
  assign termt_2n[18] = gnd;
  assign termt_2n[19] = gnd;
  assign termt_2n[20] = gnd;
  assign termt_2n[21] = gnd;
  assign termt_2n[22] = gnd;
  assign termt_2n[23] = gnd;
  assign termt_2n[24] = gnd;
  assign termt_2n[25] = gnd;
  assign termt_2n[26] = gnd;
  assign termt_2n[27] = gnd;
  assign termt_2n[28] = gnd;
  assign termt_2n[29] = gnd;
  assign termt_2n[30] = gnd;
  assign termf_2n[0] = go_0n;
  assign termf_2n[1] = go_0n;
  assign termf_2n[2] = go_0n;
  assign termf_2n[3] = go_0n;
  assign termf_2n[4] = go_0n;
  assign termf_2n[5] = go_0n;
  assign termf_2n[6] = go_0n;
  assign termf_2n[7] = go_0n;
  assign termf_2n[8] = go_0n;
  assign termf_2n[9] = go_0n;
  assign termf_2n[10] = go_0n;
  assign termf_2n[11] = go_0n;
  assign termf_2n[12] = go_0n;
  assign termf_2n[13] = go_0n;
  assign termf_2n[14] = go_0n;
  assign termf_2n[15] = go_0n;
  assign termf_2n[16] = go_0n;
  assign termf_2n[17] = go_0n;
  assign termf_2n[18] = go_0n;
  assign termf_2n[19] = go_0n;
  assign termf_2n[20] = go_0n;
  assign termf_2n[21] = go_0n;
  assign termf_2n[22] = go_0n;
  assign termf_2n[23] = go_0n;
  assign termf_2n[24] = go_0n;
  assign termf_2n[25] = go_0n;
  assign termf_2n[26] = go_0n;
  assign termf_2n[27] = go_0n;
  assign termf_2n[28] = go_0n;
  assign termf_2n[29] = go_0n;
  assign termf_2n[30] = go_0n;
  assign termt_1n = i_0r1d[32];
  assign termf_1n = i_0r0d[32];
  assign termt_0n[0] = i_0r1d[0];
  assign termt_0n[1] = i_0r1d[1];
  assign termt_0n[2] = i_0r1d[2];
  assign termt_0n[3] = i_0r1d[3];
  assign termt_0n[4] = i_0r1d[4];
  assign termt_0n[5] = i_0r1d[5];
  assign termt_0n[6] = i_0r1d[6];
  assign termt_0n[7] = i_0r1d[7];
  assign termt_0n[8] = i_0r1d[8];
  assign termt_0n[9] = i_0r1d[9];
  assign termt_0n[10] = i_0r1d[10];
  assign termt_0n[11] = i_0r1d[11];
  assign termt_0n[12] = i_0r1d[12];
  assign termt_0n[13] = i_0r1d[13];
  assign termt_0n[14] = i_0r1d[14];
  assign termt_0n[15] = i_0r1d[15];
  assign termt_0n[16] = i_0r1d[16];
  assign termt_0n[17] = i_0r1d[17];
  assign termt_0n[18] = i_0r1d[18];
  assign termt_0n[19] = i_0r1d[19];
  assign termt_0n[20] = i_0r1d[20];
  assign termt_0n[21] = i_0r1d[21];
  assign termt_0n[22] = i_0r1d[22];
  assign termt_0n[23] = i_0r1d[23];
  assign termt_0n[24] = i_0r1d[24];
  assign termt_0n[25] = i_0r1d[25];
  assign termt_0n[26] = i_0r1d[26];
  assign termt_0n[27] = i_0r1d[27];
  assign termt_0n[28] = i_0r1d[28];
  assign termt_0n[29] = i_0r1d[29];
  assign termt_0n[30] = i_0r1d[30];
  assign termt_0n[31] = i_0r1d[31];
  assign termf_0n[0] = i_0r0d[0];
  assign termf_0n[1] = i_0r0d[1];
  assign termf_0n[2] = i_0r0d[2];
  assign termf_0n[3] = i_0r0d[3];
  assign termf_0n[4] = i_0r0d[4];
  assign termf_0n[5] = i_0r0d[5];
  assign termf_0n[6] = i_0r0d[6];
  assign termf_0n[7] = i_0r0d[7];
  assign termf_0n[8] = i_0r0d[8];
  assign termf_0n[9] = i_0r0d[9];
  assign termf_0n[10] = i_0r0d[10];
  assign termf_0n[11] = i_0r0d[11];
  assign termf_0n[12] = i_0r0d[12];
  assign termf_0n[13] = i_0r0d[13];
  assign termf_0n[14] = i_0r0d[14];
  assign termf_0n[15] = i_0r0d[15];
  assign termf_0n[16] = i_0r0d[16];
  assign termf_0n[17] = i_0r0d[17];
  assign termf_0n[18] = i_0r0d[18];
  assign termf_0n[19] = i_0r0d[19];
  assign termf_0n[20] = i_0r0d[20];
  assign termf_0n[21] = i_0r0d[21];
  assign termf_0n[22] = i_0r0d[22];
  assign termf_0n[23] = i_0r0d[23];
  assign termf_0n[24] = i_0r0d[24];
  assign termf_0n[25] = i_0r0d[25];
  assign termf_0n[26] = i_0r0d[26];
  assign termf_0n[27] = i_0r0d[27];
  assign termf_0n[28] = i_0r0d[28];
  assign termf_0n[29] = i_0r0d[29];
  assign termf_0n[30] = i_0r0d[30];
  assign termf_0n[31] = i_0r0d[31];
  OR2 I256 (go_0n, i_0r0d[0], i_0r1d[0]);
endmodule

module BrzO_33_36_l91__28_28app_203_20_280_2032_2_m53m (
  i_0r0d, i_0r1d, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input [32:0] i_0r0d;
  input [32:0] i_0r1d;
  output i_0a;
  output [35:0] o_0r0d;
  output [35:0] o_0r1d;
  input o_0a;
  wire [2:0] termf_0n;
  wire [2:0] termt_0n;
  assign i_0a = o_0a;
  assign o_0r1d[33] = termt_0n[0];
  assign o_0r1d[34] = termt_0n[1];
  assign o_0r1d[35] = termt_0n[2];
  assign o_0r0d[33] = termf_0n[0];
  assign o_0r0d[34] = termf_0n[1];
  assign o_0r0d[35] = termf_0n[2];
  assign o_0r1d[0] = i_0r1d[0];
  assign o_0r1d[1] = i_0r1d[1];
  assign o_0r1d[2] = i_0r1d[2];
  assign o_0r1d[3] = i_0r1d[3];
  assign o_0r1d[4] = i_0r1d[4];
  assign o_0r1d[5] = i_0r1d[5];
  assign o_0r1d[6] = i_0r1d[6];
  assign o_0r1d[7] = i_0r1d[7];
  assign o_0r1d[8] = i_0r1d[8];
  assign o_0r1d[9] = i_0r1d[9];
  assign o_0r1d[10] = i_0r1d[10];
  assign o_0r1d[11] = i_0r1d[11];
  assign o_0r1d[12] = i_0r1d[12];
  assign o_0r1d[13] = i_0r1d[13];
  assign o_0r1d[14] = i_0r1d[14];
  assign o_0r1d[15] = i_0r1d[15];
  assign o_0r1d[16] = i_0r1d[16];
  assign o_0r1d[17] = i_0r1d[17];
  assign o_0r1d[18] = i_0r1d[18];
  assign o_0r1d[19] = i_0r1d[19];
  assign o_0r1d[20] = i_0r1d[20];
  assign o_0r1d[21] = i_0r1d[21];
  assign o_0r1d[22] = i_0r1d[22];
  assign o_0r1d[23] = i_0r1d[23];
  assign o_0r1d[24] = i_0r1d[24];
  assign o_0r1d[25] = i_0r1d[25];
  assign o_0r1d[26] = i_0r1d[26];
  assign o_0r1d[27] = i_0r1d[27];
  assign o_0r1d[28] = i_0r1d[28];
  assign o_0r1d[29] = i_0r1d[29];
  assign o_0r1d[30] = i_0r1d[30];
  assign o_0r1d[31] = i_0r1d[31];
  assign o_0r1d[32] = i_0r1d[32];
  assign o_0r0d[0] = i_0r0d[0];
  assign o_0r0d[1] = i_0r0d[1];
  assign o_0r0d[2] = i_0r0d[2];
  assign o_0r0d[3] = i_0r0d[3];
  assign o_0r0d[4] = i_0r0d[4];
  assign o_0r0d[5] = i_0r0d[5];
  assign o_0r0d[6] = i_0r0d[6];
  assign o_0r0d[7] = i_0r0d[7];
  assign o_0r0d[8] = i_0r0d[8];
  assign o_0r0d[9] = i_0r0d[9];
  assign o_0r0d[10] = i_0r0d[10];
  assign o_0r0d[11] = i_0r0d[11];
  assign o_0r0d[12] = i_0r0d[12];
  assign o_0r0d[13] = i_0r0d[13];
  assign o_0r0d[14] = i_0r0d[14];
  assign o_0r0d[15] = i_0r0d[15];
  assign o_0r0d[16] = i_0r0d[16];
  assign o_0r0d[17] = i_0r0d[17];
  assign o_0r0d[18] = i_0r0d[18];
  assign o_0r0d[19] = i_0r0d[19];
  assign o_0r0d[20] = i_0r0d[20];
  assign o_0r0d[21] = i_0r0d[21];
  assign o_0r0d[22] = i_0r0d[22];
  assign o_0r0d[23] = i_0r0d[23];
  assign o_0r0d[24] = i_0r0d[24];
  assign o_0r0d[25] = i_0r0d[25];
  assign o_0r0d[26] = i_0r0d[26];
  assign o_0r0d[27] = i_0r0d[27];
  assign o_0r0d[28] = i_0r0d[28];
  assign o_0r0d[29] = i_0r0d[29];
  assign o_0r0d[30] = i_0r0d[30];
  assign o_0r0d[31] = i_0r0d[31];
  assign o_0r0d[32] = i_0r0d[32];
  assign termt_0n[2] = i_0r1d[32];
  assign termf_0n[2] = i_0r0d[32];
  assign termt_0n[1] = i_0r1d[32];
  assign termf_0n[1] = i_0r0d[32];
  assign termt_0n[0] = i_0r1d[32];
  assign termf_0n[0] = i_0r0d[32];
endmodule

module BrzO_33_36_l76__28_28num_203_200_29_20_28a_m54m (
  i_0r0d, i_0r1d, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input [32:0] i_0r0d;
  input [32:0] i_0r1d;
  output i_0a;
  output [35:0] o_0r0d;
  output [35:0] o_0r1d;
  input o_0a;
  wire go_0n;
  wire [2:0] termf_0n;
  wire [2:0] termt_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[33] = termt_0n[0];
  assign o_0r1d[34] = termt_0n[1];
  assign o_0r1d[35] = termt_0n[2];
  assign o_0r0d[33] = termf_0n[0];
  assign o_0r0d[34] = termf_0n[1];
  assign o_0r0d[35] = termf_0n[2];
  assign o_0r1d[0] = i_0r1d[0];
  assign o_0r1d[1] = i_0r1d[1];
  assign o_0r1d[2] = i_0r1d[2];
  assign o_0r1d[3] = i_0r1d[3];
  assign o_0r1d[4] = i_0r1d[4];
  assign o_0r1d[5] = i_0r1d[5];
  assign o_0r1d[6] = i_0r1d[6];
  assign o_0r1d[7] = i_0r1d[7];
  assign o_0r1d[8] = i_0r1d[8];
  assign o_0r1d[9] = i_0r1d[9];
  assign o_0r1d[10] = i_0r1d[10];
  assign o_0r1d[11] = i_0r1d[11];
  assign o_0r1d[12] = i_0r1d[12];
  assign o_0r1d[13] = i_0r1d[13];
  assign o_0r1d[14] = i_0r1d[14];
  assign o_0r1d[15] = i_0r1d[15];
  assign o_0r1d[16] = i_0r1d[16];
  assign o_0r1d[17] = i_0r1d[17];
  assign o_0r1d[18] = i_0r1d[18];
  assign o_0r1d[19] = i_0r1d[19];
  assign o_0r1d[20] = i_0r1d[20];
  assign o_0r1d[21] = i_0r1d[21];
  assign o_0r1d[22] = i_0r1d[22];
  assign o_0r1d[23] = i_0r1d[23];
  assign o_0r1d[24] = i_0r1d[24];
  assign o_0r1d[25] = i_0r1d[25];
  assign o_0r1d[26] = i_0r1d[26];
  assign o_0r1d[27] = i_0r1d[27];
  assign o_0r1d[28] = i_0r1d[28];
  assign o_0r1d[29] = i_0r1d[29];
  assign o_0r1d[30] = i_0r1d[30];
  assign o_0r1d[31] = i_0r1d[31];
  assign o_0r1d[32] = i_0r1d[32];
  assign o_0r0d[0] = i_0r0d[0];
  assign o_0r0d[1] = i_0r0d[1];
  assign o_0r0d[2] = i_0r0d[2];
  assign o_0r0d[3] = i_0r0d[3];
  assign o_0r0d[4] = i_0r0d[4];
  assign o_0r0d[5] = i_0r0d[5];
  assign o_0r0d[6] = i_0r0d[6];
  assign o_0r0d[7] = i_0r0d[7];
  assign o_0r0d[8] = i_0r0d[8];
  assign o_0r0d[9] = i_0r0d[9];
  assign o_0r0d[10] = i_0r0d[10];
  assign o_0r0d[11] = i_0r0d[11];
  assign o_0r0d[12] = i_0r0d[12];
  assign o_0r0d[13] = i_0r0d[13];
  assign o_0r0d[14] = i_0r0d[14];
  assign o_0r0d[15] = i_0r0d[15];
  assign o_0r0d[16] = i_0r0d[16];
  assign o_0r0d[17] = i_0r0d[17];
  assign o_0r0d[18] = i_0r0d[18];
  assign o_0r0d[19] = i_0r0d[19];
  assign o_0r0d[20] = i_0r0d[20];
  assign o_0r0d[21] = i_0r0d[21];
  assign o_0r0d[22] = i_0r0d[22];
  assign o_0r0d[23] = i_0r0d[23];
  assign o_0r0d[24] = i_0r0d[24];
  assign o_0r0d[25] = i_0r0d[25];
  assign o_0r0d[26] = i_0r0d[26];
  assign o_0r0d[27] = i_0r0d[27];
  assign o_0r0d[28] = i_0r0d[28];
  assign o_0r0d[29] = i_0r0d[29];
  assign o_0r0d[30] = i_0r0d[30];
  assign o_0r0d[31] = i_0r0d[31];
  assign o_0r0d[32] = i_0r0d[32];
  assign termt_0n[0] = gnd;
  assign termt_0n[1] = gnd;
  assign termt_0n[2] = gnd;
  assign termf_0n[0] = go_0n;
  assign termf_0n[1] = go_0n;
  assign termf_0n[2] = go_0n;
  OR2 I79 (go_0n, i_0r0d[0], i_0r1d[0]);
endmodule

module BrzO_35_35_l34__28_28not_20_280_200_2035_2_m55m (
  i_0r0d, i_0r1d, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input [34:0] i_0r0d;
  input [34:0] i_0r1d;
  output i_0a;
  output [34:0] o_0r0d;
  output [34:0] o_0r1d;
  input o_0a;
  assign i_0a = o_0a;
  assign o_0r0d[0] = i_0r1d[0];
  assign o_0r0d[1] = i_0r1d[1];
  assign o_0r0d[2] = i_0r1d[2];
  assign o_0r0d[3] = i_0r1d[3];
  assign o_0r0d[4] = i_0r1d[4];
  assign o_0r0d[5] = i_0r1d[5];
  assign o_0r0d[6] = i_0r1d[6];
  assign o_0r0d[7] = i_0r1d[7];
  assign o_0r0d[8] = i_0r1d[8];
  assign o_0r0d[9] = i_0r1d[9];
  assign o_0r0d[10] = i_0r1d[10];
  assign o_0r0d[11] = i_0r1d[11];
  assign o_0r0d[12] = i_0r1d[12];
  assign o_0r0d[13] = i_0r1d[13];
  assign o_0r0d[14] = i_0r1d[14];
  assign o_0r0d[15] = i_0r1d[15];
  assign o_0r0d[16] = i_0r1d[16];
  assign o_0r0d[17] = i_0r1d[17];
  assign o_0r0d[18] = i_0r1d[18];
  assign o_0r0d[19] = i_0r1d[19];
  assign o_0r0d[20] = i_0r1d[20];
  assign o_0r0d[21] = i_0r1d[21];
  assign o_0r0d[22] = i_0r1d[22];
  assign o_0r0d[23] = i_0r1d[23];
  assign o_0r0d[24] = i_0r1d[24];
  assign o_0r0d[25] = i_0r1d[25];
  assign o_0r0d[26] = i_0r1d[26];
  assign o_0r0d[27] = i_0r1d[27];
  assign o_0r0d[28] = i_0r1d[28];
  assign o_0r0d[29] = i_0r1d[29];
  assign o_0r0d[30] = i_0r1d[30];
  assign o_0r0d[31] = i_0r1d[31];
  assign o_0r0d[32] = i_0r1d[32];
  assign o_0r0d[33] = i_0r1d[33];
  assign o_0r0d[34] = i_0r1d[34];
  assign o_0r1d[0] = i_0r0d[0];
  assign o_0r1d[1] = i_0r0d[1];
  assign o_0r1d[2] = i_0r0d[2];
  assign o_0r1d[3] = i_0r0d[3];
  assign o_0r1d[4] = i_0r0d[4];
  assign o_0r1d[5] = i_0r0d[5];
  assign o_0r1d[6] = i_0r0d[6];
  assign o_0r1d[7] = i_0r0d[7];
  assign o_0r1d[8] = i_0r0d[8];
  assign o_0r1d[9] = i_0r0d[9];
  assign o_0r1d[10] = i_0r0d[10];
  assign o_0r1d[11] = i_0r0d[11];
  assign o_0r1d[12] = i_0r0d[12];
  assign o_0r1d[13] = i_0r0d[13];
  assign o_0r1d[14] = i_0r0d[14];
  assign o_0r1d[15] = i_0r0d[15];
  assign o_0r1d[16] = i_0r0d[16];
  assign o_0r1d[17] = i_0r0d[17];
  assign o_0r1d[18] = i_0r0d[18];
  assign o_0r1d[19] = i_0r0d[19];
  assign o_0r1d[20] = i_0r0d[20];
  assign o_0r1d[21] = i_0r0d[21];
  assign o_0r1d[22] = i_0r0d[22];
  assign o_0r1d[23] = i_0r0d[23];
  assign o_0r1d[24] = i_0r0d[24];
  assign o_0r1d[25] = i_0r0d[25];
  assign o_0r1d[26] = i_0r0d[26];
  assign o_0r1d[27] = i_0r0d[27];
  assign o_0r1d[28] = i_0r0d[28];
  assign o_0r1d[29] = i_0r0d[29];
  assign o_0r1d[30] = i_0r0d[30];
  assign o_0r1d[31] = i_0r0d[31];
  assign o_0r1d[32] = i_0r0d[32];
  assign o_0r1d[33] = i_0r0d[33];
  assign o_0r1d[34] = i_0r0d[34];
endmodule

module BrzO_35_36_l76__28_28num_201_200_29_20_28a_m56m (
  i_0r0d, i_0r1d, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input [34:0] i_0r0d;
  input [34:0] i_0r1d;
  output i_0a;
  output [35:0] o_0r0d;
  output [35:0] o_0r1d;
  input o_0a;
  wire go_0n;
  wire termf_0n;
  wire termt_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  assign o_0r1d[35] = termt_0n;
  assign o_0r0d[35] = termf_0n;
  assign o_0r1d[0] = i_0r1d[0];
  assign o_0r1d[1] = i_0r1d[1];
  assign o_0r1d[2] = i_0r1d[2];
  assign o_0r1d[3] = i_0r1d[3];
  assign o_0r1d[4] = i_0r1d[4];
  assign o_0r1d[5] = i_0r1d[5];
  assign o_0r1d[6] = i_0r1d[6];
  assign o_0r1d[7] = i_0r1d[7];
  assign o_0r1d[8] = i_0r1d[8];
  assign o_0r1d[9] = i_0r1d[9];
  assign o_0r1d[10] = i_0r1d[10];
  assign o_0r1d[11] = i_0r1d[11];
  assign o_0r1d[12] = i_0r1d[12];
  assign o_0r1d[13] = i_0r1d[13];
  assign o_0r1d[14] = i_0r1d[14];
  assign o_0r1d[15] = i_0r1d[15];
  assign o_0r1d[16] = i_0r1d[16];
  assign o_0r1d[17] = i_0r1d[17];
  assign o_0r1d[18] = i_0r1d[18];
  assign o_0r1d[19] = i_0r1d[19];
  assign o_0r1d[20] = i_0r1d[20];
  assign o_0r1d[21] = i_0r1d[21];
  assign o_0r1d[22] = i_0r1d[22];
  assign o_0r1d[23] = i_0r1d[23];
  assign o_0r1d[24] = i_0r1d[24];
  assign o_0r1d[25] = i_0r1d[25];
  assign o_0r1d[26] = i_0r1d[26];
  assign o_0r1d[27] = i_0r1d[27];
  assign o_0r1d[28] = i_0r1d[28];
  assign o_0r1d[29] = i_0r1d[29];
  assign o_0r1d[30] = i_0r1d[30];
  assign o_0r1d[31] = i_0r1d[31];
  assign o_0r1d[32] = i_0r1d[32];
  assign o_0r1d[33] = i_0r1d[33];
  assign o_0r1d[34] = i_0r1d[34];
  assign o_0r0d[0] = i_0r0d[0];
  assign o_0r0d[1] = i_0r0d[1];
  assign o_0r0d[2] = i_0r0d[2];
  assign o_0r0d[3] = i_0r0d[3];
  assign o_0r0d[4] = i_0r0d[4];
  assign o_0r0d[5] = i_0r0d[5];
  assign o_0r0d[6] = i_0r0d[6];
  assign o_0r0d[7] = i_0r0d[7];
  assign o_0r0d[8] = i_0r0d[8];
  assign o_0r0d[9] = i_0r0d[9];
  assign o_0r0d[10] = i_0r0d[10];
  assign o_0r0d[11] = i_0r0d[11];
  assign o_0r0d[12] = i_0r0d[12];
  assign o_0r0d[13] = i_0r0d[13];
  assign o_0r0d[14] = i_0r0d[14];
  assign o_0r0d[15] = i_0r0d[15];
  assign o_0r0d[16] = i_0r0d[16];
  assign o_0r0d[17] = i_0r0d[17];
  assign o_0r0d[18] = i_0r0d[18];
  assign o_0r0d[19] = i_0r0d[19];
  assign o_0r0d[20] = i_0r0d[20];
  assign o_0r0d[21] = i_0r0d[21];
  assign o_0r0d[22] = i_0r0d[22];
  assign o_0r0d[23] = i_0r0d[23];
  assign o_0r0d[24] = i_0r0d[24];
  assign o_0r0d[25] = i_0r0d[25];
  assign o_0r0d[26] = i_0r0d[26];
  assign o_0r0d[27] = i_0r0d[27];
  assign o_0r0d[28] = i_0r0d[28];
  assign o_0r0d[29] = i_0r0d[29];
  assign o_0r0d[30] = i_0r0d[30];
  assign o_0r0d[31] = i_0r0d[31];
  assign o_0r0d[32] = i_0r0d[32];
  assign o_0r0d[33] = i_0r0d[33];
  assign o_0r0d[34] = i_0r0d[34];
  assign termt_0n = gnd;
  assign termf_0n = go_0n;
  OR2 I75 (go_0n, i_0r0d[0], i_0r1d[0]);
endmodule

module AO222 (
  q,
  i0,
  i1,
  i2,
  i3,
  i4,
  i5
);
  output q;
  input i0;
  input i1;
  input i2;
  input i3;
  input i4;
  input i5;
  wire [2:0] int_0n;
  OR3 I0 (q, int_0n[0], int_0n[1], int_0n[2]);
  AND2 I1 (int_0n[2], i4, i5);
  AND2 I2 (int_0n[1], i2, i3);
  AND2 I3 (int_0n[0], i0, i1);
endmodule

module DRFA (
  a0,
  a1,
  b0,
  b1,
  ci0,
  ci1,
  co0,
  co1,
  sum0,
  sum1
);
  input a0;
  input a1;
  input b0;
  input b1;
  input ci0;
  input ci1;
  output co0;
  output co1;
  output sum0;
  output sum1;
  wire [7:0] internal_0n;
  wire [7:0] minterm_0n;
  AO222 I0 (co0, a0, b0, a0, ci0, b0, ci0);
  AO222 I1 (co1, a1, b1, a1, ci1, b1, ci1);
  NAND2 I2 (sum0, internal_0n[4], internal_0n[5]);
  NOR2 I3 (internal_0n[5], minterm_0n[5], minterm_0n[6]);
  NOR2 I4 (internal_0n[4], minterm_0n[0], minterm_0n[3]);
  NAND2 I5 (sum1, internal_0n[6], internal_0n[7]);
  NOR2 I6 (internal_0n[7], minterm_0n[4], minterm_0n[7]);
  NOR2 I7 (internal_0n[6], minterm_0n[1], minterm_0n[2]);
  C3 I8 (minterm_0n[7], a1, b1, ci1);
  C3 I9 (minterm_0n[6], a1, b1, ci0);
  C3 I10 (minterm_0n[5], a1, b0, ci1);
  C3 I11 (minterm_0n[4], a1, b0, ci0);
  C3 I12 (minterm_0n[3], a0, b1, ci1);
  C3 I13 (minterm_0n[2], a0, b1, ci0);
  C3 I14 (minterm_0n[1], a0, b0, ci1);
  C3 I15 (minterm_0n[0], a0, b0, ci0);
endmodule

module AO21 (
  q,
  i0,
  i1,
  i2
);
  output q;
  input i0;
  input i1;
  input i2;
  wire int_0n;
  OR2 I0 (q, i2, int_0n);
  AND2 I1 (int_0n, i0, i1);
endmodule

module DRHA (
  a_0,
  a_1,
  b_0,
  b_1,
  co_0,
  co_1,
  sum_0,
  sum_1
);
  input a_0;
  input a_1;
  input b_0;
  input b_1;
  output co_0;
  output co_1;
  output sum_0;
  output sum_1;
  wire n0_0n;
  wire n1_0n;
  wire n2_0n;
  wire n3_0n;
  AND2 I0 (co_1, a_1, b_1);
  AO21 I1 (co_0, a_1, b_0, a_0);
  OR2 I2 (sum_1, n1_0n, n2_0n);
  OR2 I3 (sum_0, n0_0n, n3_0n);
  C2 I4 (n3_0n, a_1, b_1);
  C2 I5 (n2_0n, a_1, b_0);
  C2 I6 (n1_0n, a_0, b_1);
  C2 I7 (n0_0n, a_0, b_0);
endmodule

module BrzO_66_34_l270__28_28app_201_20_280_200_2_m57m (
  i_0r0d, i_0r1d, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input [65:0] i_0r0d;
  input [65:0] i_0r1d;
  output i_0a;
  output [33:0] o_0r0d;
  output [33:0] o_0r1d;
  input o_0a;
  wire go_0n;
  wire [32:0] termf_0n;
  wire [32:0] termf_1n;
  wire termf_2n;
  wire [33:0] termf_3n;
  wire termf_4n;
  wire [33:0] termf_5n;
  wire [32:0] termt_0n;
  wire [32:0] termt_1n;
  wire termt_2n;
  wire [33:0] termt_3n;
  wire termt_4n;
  wire [33:0] termt_5n;
  wire [33:0] carryt7_0n;
  wire [33:0] carryf7_0n;
  supply0 gnd;
  assign i_0a = o_0a;
  DRFA I1 (termf_3n[1], termt_3n[1], termf_5n[1], termt_5n[1], carryf7_0n[0], carryt7_0n[0], carryf7_0n[1], carryt7_0n[1], o_0r0d[1], o_0r1d[1]);
  DRFA I2 (termf_3n[2], termt_3n[2], termf_5n[2], termt_5n[2], carryf7_0n[1], carryt7_0n[1], carryf7_0n[2], carryt7_0n[2], o_0r0d[2], o_0r1d[2]);
  DRFA I3 (termf_3n[3], termt_3n[3], termf_5n[3], termt_5n[3], carryf7_0n[2], carryt7_0n[2], carryf7_0n[3], carryt7_0n[3], o_0r0d[3], o_0r1d[3]);
  DRFA I4 (termf_3n[4], termt_3n[4], termf_5n[4], termt_5n[4], carryf7_0n[3], carryt7_0n[3], carryf7_0n[4], carryt7_0n[4], o_0r0d[4], o_0r1d[4]);
  DRFA I5 (termf_3n[5], termt_3n[5], termf_5n[5], termt_5n[5], carryf7_0n[4], carryt7_0n[4], carryf7_0n[5], carryt7_0n[5], o_0r0d[5], o_0r1d[5]);
  DRFA I6 (termf_3n[6], termt_3n[6], termf_5n[6], termt_5n[6], carryf7_0n[5], carryt7_0n[5], carryf7_0n[6], carryt7_0n[6], o_0r0d[6], o_0r1d[6]);
  DRFA I7 (termf_3n[7], termt_3n[7], termf_5n[7], termt_5n[7], carryf7_0n[6], carryt7_0n[6], carryf7_0n[7], carryt7_0n[7], o_0r0d[7], o_0r1d[7]);
  DRFA I8 (termf_3n[8], termt_3n[8], termf_5n[8], termt_5n[8], carryf7_0n[7], carryt7_0n[7], carryf7_0n[8], carryt7_0n[8], o_0r0d[8], o_0r1d[8]);
  DRFA I9 (termf_3n[9], termt_3n[9], termf_5n[9], termt_5n[9], carryf7_0n[8], carryt7_0n[8], carryf7_0n[9], carryt7_0n[9], o_0r0d[9], o_0r1d[9]);
  DRFA I10 (termf_3n[10], termt_3n[10], termf_5n[10], termt_5n[10], carryf7_0n[9], carryt7_0n[9], carryf7_0n[10], carryt7_0n[10], o_0r0d[10], o_0r1d[10]);
  DRFA I11 (termf_3n[11], termt_3n[11], termf_5n[11], termt_5n[11], carryf7_0n[10], carryt7_0n[10], carryf7_0n[11], carryt7_0n[11], o_0r0d[11], o_0r1d[11]);
  DRFA I12 (termf_3n[12], termt_3n[12], termf_5n[12], termt_5n[12], carryf7_0n[11], carryt7_0n[11], carryf7_0n[12], carryt7_0n[12], o_0r0d[12], o_0r1d[12]);
  DRFA I13 (termf_3n[13], termt_3n[13], termf_5n[13], termt_5n[13], carryf7_0n[12], carryt7_0n[12], carryf7_0n[13], carryt7_0n[13], o_0r0d[13], o_0r1d[13]);
  DRFA I14 (termf_3n[14], termt_3n[14], termf_5n[14], termt_5n[14], carryf7_0n[13], carryt7_0n[13], carryf7_0n[14], carryt7_0n[14], o_0r0d[14], o_0r1d[14]);
  DRFA I15 (termf_3n[15], termt_3n[15], termf_5n[15], termt_5n[15], carryf7_0n[14], carryt7_0n[14], carryf7_0n[15], carryt7_0n[15], o_0r0d[15], o_0r1d[15]);
  DRFA I16 (termf_3n[16], termt_3n[16], termf_5n[16], termt_5n[16], carryf7_0n[15], carryt7_0n[15], carryf7_0n[16], carryt7_0n[16], o_0r0d[16], o_0r1d[16]);
  DRFA I17 (termf_3n[17], termt_3n[17], termf_5n[17], termt_5n[17], carryf7_0n[16], carryt7_0n[16], carryf7_0n[17], carryt7_0n[17], o_0r0d[17], o_0r1d[17]);
  DRFA I18 (termf_3n[18], termt_3n[18], termf_5n[18], termt_5n[18], carryf7_0n[17], carryt7_0n[17], carryf7_0n[18], carryt7_0n[18], o_0r0d[18], o_0r1d[18]);
  DRFA I19 (termf_3n[19], termt_3n[19], termf_5n[19], termt_5n[19], carryf7_0n[18], carryt7_0n[18], carryf7_0n[19], carryt7_0n[19], o_0r0d[19], o_0r1d[19]);
  DRFA I20 (termf_3n[20], termt_3n[20], termf_5n[20], termt_5n[20], carryf7_0n[19], carryt7_0n[19], carryf7_0n[20], carryt7_0n[20], o_0r0d[20], o_0r1d[20]);
  DRFA I21 (termf_3n[21], termt_3n[21], termf_5n[21], termt_5n[21], carryf7_0n[20], carryt7_0n[20], carryf7_0n[21], carryt7_0n[21], o_0r0d[21], o_0r1d[21]);
  DRFA I22 (termf_3n[22], termt_3n[22], termf_5n[22], termt_5n[22], carryf7_0n[21], carryt7_0n[21], carryf7_0n[22], carryt7_0n[22], o_0r0d[22], o_0r1d[22]);
  DRFA I23 (termf_3n[23], termt_3n[23], termf_5n[23], termt_5n[23], carryf7_0n[22], carryt7_0n[22], carryf7_0n[23], carryt7_0n[23], o_0r0d[23], o_0r1d[23]);
  DRFA I24 (termf_3n[24], termt_3n[24], termf_5n[24], termt_5n[24], carryf7_0n[23], carryt7_0n[23], carryf7_0n[24], carryt7_0n[24], o_0r0d[24], o_0r1d[24]);
  DRFA I25 (termf_3n[25], termt_3n[25], termf_5n[25], termt_5n[25], carryf7_0n[24], carryt7_0n[24], carryf7_0n[25], carryt7_0n[25], o_0r0d[25], o_0r1d[25]);
  DRFA I26 (termf_3n[26], termt_3n[26], termf_5n[26], termt_5n[26], carryf7_0n[25], carryt7_0n[25], carryf7_0n[26], carryt7_0n[26], o_0r0d[26], o_0r1d[26]);
  DRFA I27 (termf_3n[27], termt_3n[27], termf_5n[27], termt_5n[27], carryf7_0n[26], carryt7_0n[26], carryf7_0n[27], carryt7_0n[27], o_0r0d[27], o_0r1d[27]);
  DRFA I28 (termf_3n[28], termt_3n[28], termf_5n[28], termt_5n[28], carryf7_0n[27], carryt7_0n[27], carryf7_0n[28], carryt7_0n[28], o_0r0d[28], o_0r1d[28]);
  DRFA I29 (termf_3n[29], termt_3n[29], termf_5n[29], termt_5n[29], carryf7_0n[28], carryt7_0n[28], carryf7_0n[29], carryt7_0n[29], o_0r0d[29], o_0r1d[29]);
  DRFA I30 (termf_3n[30], termt_3n[30], termf_5n[30], termt_5n[30], carryf7_0n[29], carryt7_0n[29], carryf7_0n[30], carryt7_0n[30], o_0r0d[30], o_0r1d[30]);
  DRFA I31 (termf_3n[31], termt_3n[31], termf_5n[31], termt_5n[31], carryf7_0n[30], carryt7_0n[30], carryf7_0n[31], carryt7_0n[31], o_0r0d[31], o_0r1d[31]);
  DRFA I32 (termf_3n[32], termt_3n[32], termf_5n[32], termt_5n[32], carryf7_0n[31], carryt7_0n[31], carryf7_0n[32], carryt7_0n[32], o_0r0d[32], o_0r1d[32]);
  DRFA I33 (termf_3n[33], termt_3n[33], termf_5n[33], termt_5n[33], carryf7_0n[32], carryt7_0n[32], carryf7_0n[33], carryt7_0n[33], o_0r0d[33], o_0r1d[33]);
  DRHA I34 (termf_3n[0], termt_3n[0], termf_5n[0], termt_5n[0], carryf7_0n[0], carryt7_0n[0], o_0r0d[0], o_0r1d[0]);
  assign termt_5n[33] = termt_4n;
  assign termf_5n[33] = termf_4n;
  assign termt_5n[0] = termt_1n[0];
  assign termt_5n[1] = termt_1n[1];
  assign termt_5n[2] = termt_1n[2];
  assign termt_5n[3] = termt_1n[3];
  assign termt_5n[4] = termt_1n[4];
  assign termt_5n[5] = termt_1n[5];
  assign termt_5n[6] = termt_1n[6];
  assign termt_5n[7] = termt_1n[7];
  assign termt_5n[8] = termt_1n[8];
  assign termt_5n[9] = termt_1n[9];
  assign termt_5n[10] = termt_1n[10];
  assign termt_5n[11] = termt_1n[11];
  assign termt_5n[12] = termt_1n[12];
  assign termt_5n[13] = termt_1n[13];
  assign termt_5n[14] = termt_1n[14];
  assign termt_5n[15] = termt_1n[15];
  assign termt_5n[16] = termt_1n[16];
  assign termt_5n[17] = termt_1n[17];
  assign termt_5n[18] = termt_1n[18];
  assign termt_5n[19] = termt_1n[19];
  assign termt_5n[20] = termt_1n[20];
  assign termt_5n[21] = termt_1n[21];
  assign termt_5n[22] = termt_1n[22];
  assign termt_5n[23] = termt_1n[23];
  assign termt_5n[24] = termt_1n[24];
  assign termt_5n[25] = termt_1n[25];
  assign termt_5n[26] = termt_1n[26];
  assign termt_5n[27] = termt_1n[27];
  assign termt_5n[28] = termt_1n[28];
  assign termt_5n[29] = termt_1n[29];
  assign termt_5n[30] = termt_1n[30];
  assign termt_5n[31] = termt_1n[31];
  assign termt_5n[32] = termt_1n[32];
  assign termf_5n[0] = termf_1n[0];
  assign termf_5n[1] = termf_1n[1];
  assign termf_5n[2] = termf_1n[2];
  assign termf_5n[3] = termf_1n[3];
  assign termf_5n[4] = termf_1n[4];
  assign termf_5n[5] = termf_1n[5];
  assign termf_5n[6] = termf_1n[6];
  assign termf_5n[7] = termf_1n[7];
  assign termf_5n[8] = termf_1n[8];
  assign termf_5n[9] = termf_1n[9];
  assign termf_5n[10] = termf_1n[10];
  assign termf_5n[11] = termf_1n[11];
  assign termf_5n[12] = termf_1n[12];
  assign termf_5n[13] = termf_1n[13];
  assign termf_5n[14] = termf_1n[14];
  assign termf_5n[15] = termf_1n[15];
  assign termf_5n[16] = termf_1n[16];
  assign termf_5n[17] = termf_1n[17];
  assign termf_5n[18] = termf_1n[18];
  assign termf_5n[19] = termf_1n[19];
  assign termf_5n[20] = termf_1n[20];
  assign termf_5n[21] = termf_1n[21];
  assign termf_5n[22] = termf_1n[22];
  assign termf_5n[23] = termf_1n[23];
  assign termf_5n[24] = termf_1n[24];
  assign termf_5n[25] = termf_1n[25];
  assign termf_5n[26] = termf_1n[26];
  assign termf_5n[27] = termf_1n[27];
  assign termf_5n[28] = termf_1n[28];
  assign termf_5n[29] = termf_1n[29];
  assign termf_5n[30] = termf_1n[30];
  assign termf_5n[31] = termf_1n[31];
  assign termf_5n[32] = termf_1n[32];
  assign termt_4n = gnd;
  assign termf_4n = go_0n;
  assign termt_3n[33] = termt_2n;
  assign termf_3n[33] = termf_2n;
  assign termt_3n[0] = termt_0n[0];
  assign termt_3n[1] = termt_0n[1];
  assign termt_3n[2] = termt_0n[2];
  assign termt_3n[3] = termt_0n[3];
  assign termt_3n[4] = termt_0n[4];
  assign termt_3n[5] = termt_0n[5];
  assign termt_3n[6] = termt_0n[6];
  assign termt_3n[7] = termt_0n[7];
  assign termt_3n[8] = termt_0n[8];
  assign termt_3n[9] = termt_0n[9];
  assign termt_3n[10] = termt_0n[10];
  assign termt_3n[11] = termt_0n[11];
  assign termt_3n[12] = termt_0n[12];
  assign termt_3n[13] = termt_0n[13];
  assign termt_3n[14] = termt_0n[14];
  assign termt_3n[15] = termt_0n[15];
  assign termt_3n[16] = termt_0n[16];
  assign termt_3n[17] = termt_0n[17];
  assign termt_3n[18] = termt_0n[18];
  assign termt_3n[19] = termt_0n[19];
  assign termt_3n[20] = termt_0n[20];
  assign termt_3n[21] = termt_0n[21];
  assign termt_3n[22] = termt_0n[22];
  assign termt_3n[23] = termt_0n[23];
  assign termt_3n[24] = termt_0n[24];
  assign termt_3n[25] = termt_0n[25];
  assign termt_3n[26] = termt_0n[26];
  assign termt_3n[27] = termt_0n[27];
  assign termt_3n[28] = termt_0n[28];
  assign termt_3n[29] = termt_0n[29];
  assign termt_3n[30] = termt_0n[30];
  assign termt_3n[31] = termt_0n[31];
  assign termt_3n[32] = termt_0n[32];
  assign termf_3n[0] = termf_0n[0];
  assign termf_3n[1] = termf_0n[1];
  assign termf_3n[2] = termf_0n[2];
  assign termf_3n[3] = termf_0n[3];
  assign termf_3n[4] = termf_0n[4];
  assign termf_3n[5] = termf_0n[5];
  assign termf_3n[6] = termf_0n[6];
  assign termf_3n[7] = termf_0n[7];
  assign termf_3n[8] = termf_0n[8];
  assign termf_3n[9] = termf_0n[9];
  assign termf_3n[10] = termf_0n[10];
  assign termf_3n[11] = termf_0n[11];
  assign termf_3n[12] = termf_0n[12];
  assign termf_3n[13] = termf_0n[13];
  assign termf_3n[14] = termf_0n[14];
  assign termf_3n[15] = termf_0n[15];
  assign termf_3n[16] = termf_0n[16];
  assign termf_3n[17] = termf_0n[17];
  assign termf_3n[18] = termf_0n[18];
  assign termf_3n[19] = termf_0n[19];
  assign termf_3n[20] = termf_0n[20];
  assign termf_3n[21] = termf_0n[21];
  assign termf_3n[22] = termf_0n[22];
  assign termf_3n[23] = termf_0n[23];
  assign termf_3n[24] = termf_0n[24];
  assign termf_3n[25] = termf_0n[25];
  assign termf_3n[26] = termf_0n[26];
  assign termf_3n[27] = termf_0n[27];
  assign termf_3n[28] = termf_0n[28];
  assign termf_3n[29] = termf_0n[29];
  assign termf_3n[30] = termf_0n[30];
  assign termf_3n[31] = termf_0n[31];
  assign termf_3n[32] = termf_0n[32];
  assign termt_2n = gnd;
  assign termf_2n = go_0n;
  assign termt_1n[0] = i_0r1d[33];
  assign termt_1n[1] = i_0r1d[34];
  assign termt_1n[2] = i_0r1d[35];
  assign termt_1n[3] = i_0r1d[36];
  assign termt_1n[4] = i_0r1d[37];
  assign termt_1n[5] = i_0r1d[38];
  assign termt_1n[6] = i_0r1d[39];
  assign termt_1n[7] = i_0r1d[40];
  assign termt_1n[8] = i_0r1d[41];
  assign termt_1n[9] = i_0r1d[42];
  assign termt_1n[10] = i_0r1d[43];
  assign termt_1n[11] = i_0r1d[44];
  assign termt_1n[12] = i_0r1d[45];
  assign termt_1n[13] = i_0r1d[46];
  assign termt_1n[14] = i_0r1d[47];
  assign termt_1n[15] = i_0r1d[48];
  assign termt_1n[16] = i_0r1d[49];
  assign termt_1n[17] = i_0r1d[50];
  assign termt_1n[18] = i_0r1d[51];
  assign termt_1n[19] = i_0r1d[52];
  assign termt_1n[20] = i_0r1d[53];
  assign termt_1n[21] = i_0r1d[54];
  assign termt_1n[22] = i_0r1d[55];
  assign termt_1n[23] = i_0r1d[56];
  assign termt_1n[24] = i_0r1d[57];
  assign termt_1n[25] = i_0r1d[58];
  assign termt_1n[26] = i_0r1d[59];
  assign termt_1n[27] = i_0r1d[60];
  assign termt_1n[28] = i_0r1d[61];
  assign termt_1n[29] = i_0r1d[62];
  assign termt_1n[30] = i_0r1d[63];
  assign termt_1n[31] = i_0r1d[64];
  assign termt_1n[32] = i_0r1d[65];
  assign termf_1n[0] = i_0r0d[33];
  assign termf_1n[1] = i_0r0d[34];
  assign termf_1n[2] = i_0r0d[35];
  assign termf_1n[3] = i_0r0d[36];
  assign termf_1n[4] = i_0r0d[37];
  assign termf_1n[5] = i_0r0d[38];
  assign termf_1n[6] = i_0r0d[39];
  assign termf_1n[7] = i_0r0d[40];
  assign termf_1n[8] = i_0r0d[41];
  assign termf_1n[9] = i_0r0d[42];
  assign termf_1n[10] = i_0r0d[43];
  assign termf_1n[11] = i_0r0d[44];
  assign termf_1n[12] = i_0r0d[45];
  assign termf_1n[13] = i_0r0d[46];
  assign termf_1n[14] = i_0r0d[47];
  assign termf_1n[15] = i_0r0d[48];
  assign termf_1n[16] = i_0r0d[49];
  assign termf_1n[17] = i_0r0d[50];
  assign termf_1n[18] = i_0r0d[51];
  assign termf_1n[19] = i_0r0d[52];
  assign termf_1n[20] = i_0r0d[53];
  assign termf_1n[21] = i_0r0d[54];
  assign termf_1n[22] = i_0r0d[55];
  assign termf_1n[23] = i_0r0d[56];
  assign termf_1n[24] = i_0r0d[57];
  assign termf_1n[25] = i_0r0d[58];
  assign termf_1n[26] = i_0r0d[59];
  assign termf_1n[27] = i_0r0d[60];
  assign termf_1n[28] = i_0r0d[61];
  assign termf_1n[29] = i_0r0d[62];
  assign termf_1n[30] = i_0r0d[63];
  assign termf_1n[31] = i_0r0d[64];
  assign termf_1n[32] = i_0r0d[65];
  assign termt_0n[0] = i_0r1d[0];
  assign termt_0n[1] = i_0r1d[1];
  assign termt_0n[2] = i_0r1d[2];
  assign termt_0n[3] = i_0r1d[3];
  assign termt_0n[4] = i_0r1d[4];
  assign termt_0n[5] = i_0r1d[5];
  assign termt_0n[6] = i_0r1d[6];
  assign termt_0n[7] = i_0r1d[7];
  assign termt_0n[8] = i_0r1d[8];
  assign termt_0n[9] = i_0r1d[9];
  assign termt_0n[10] = i_0r1d[10];
  assign termt_0n[11] = i_0r1d[11];
  assign termt_0n[12] = i_0r1d[12];
  assign termt_0n[13] = i_0r1d[13];
  assign termt_0n[14] = i_0r1d[14];
  assign termt_0n[15] = i_0r1d[15];
  assign termt_0n[16] = i_0r1d[16];
  assign termt_0n[17] = i_0r1d[17];
  assign termt_0n[18] = i_0r1d[18];
  assign termt_0n[19] = i_0r1d[19];
  assign termt_0n[20] = i_0r1d[20];
  assign termt_0n[21] = i_0r1d[21];
  assign termt_0n[22] = i_0r1d[22];
  assign termt_0n[23] = i_0r1d[23];
  assign termt_0n[24] = i_0r1d[24];
  assign termt_0n[25] = i_0r1d[25];
  assign termt_0n[26] = i_0r1d[26];
  assign termt_0n[27] = i_0r1d[27];
  assign termt_0n[28] = i_0r1d[28];
  assign termt_0n[29] = i_0r1d[29];
  assign termt_0n[30] = i_0r1d[30];
  assign termt_0n[31] = i_0r1d[31];
  assign termt_0n[32] = i_0r1d[32];
  assign termf_0n[0] = i_0r0d[0];
  assign termf_0n[1] = i_0r0d[1];
  assign termf_0n[2] = i_0r0d[2];
  assign termf_0n[3] = i_0r0d[3];
  assign termf_0n[4] = i_0r0d[4];
  assign termf_0n[5] = i_0r0d[5];
  assign termf_0n[6] = i_0r0d[6];
  assign termf_0n[7] = i_0r0d[7];
  assign termf_0n[8] = i_0r0d[8];
  assign termf_0n[9] = i_0r0d[9];
  assign termf_0n[10] = i_0r0d[10];
  assign termf_0n[11] = i_0r0d[11];
  assign termf_0n[12] = i_0r0d[12];
  assign termf_0n[13] = i_0r0d[13];
  assign termf_0n[14] = i_0r0d[14];
  assign termf_0n[15] = i_0r0d[15];
  assign termf_0n[16] = i_0r0d[16];
  assign termf_0n[17] = i_0r0d[17];
  assign termf_0n[18] = i_0r0d[18];
  assign termf_0n[19] = i_0r0d[19];
  assign termf_0n[20] = i_0r0d[20];
  assign termf_0n[21] = i_0r0d[21];
  assign termf_0n[22] = i_0r0d[22];
  assign termf_0n[23] = i_0r0d[23];
  assign termf_0n[24] = i_0r0d[24];
  assign termf_0n[25] = i_0r0d[25];
  assign termf_0n[26] = i_0r0d[26];
  assign termf_0n[27] = i_0r0d[27];
  assign termf_0n[28] = i_0r0d[28];
  assign termf_0n[29] = i_0r0d[29];
  assign termf_0n[30] = i_0r0d[30];
  assign termf_0n[31] = i_0r0d[31];
  assign termf_0n[32] = i_0r0d[32];
  OR2 I307 (go_0n, i_0r0d[0], i_0r1d[0]);
endmodule

module BrzO_70_35_l124__28_28app_201_20_280_200_2_m58m (
  i_0r0d, i_0r1d, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input [69:0] i_0r0d;
  input [69:0] i_0r1d;
  output i_0a;
  output [34:0] o_0r0d;
  output [34:0] o_0r1d;
  input o_0a;
  wire [34:0] termf_0n;
  wire [34:0] termf_1n;
  wire [34:0] termt_0n;
  wire [34:0] termt_1n;
  assign i_0a = o_0a;
  DRAND2 I1 (termf_0n[0], termt_0n[0], termf_1n[0], termt_1n[0], o_0r0d[0], o_0r1d[0]);
  DRAND2 I2 (termf_0n[1], termt_0n[1], termf_1n[1], termt_1n[1], o_0r0d[1], o_0r1d[1]);
  DRAND2 I3 (termf_0n[2], termt_0n[2], termf_1n[2], termt_1n[2], o_0r0d[2], o_0r1d[2]);
  DRAND2 I4 (termf_0n[3], termt_0n[3], termf_1n[3], termt_1n[3], o_0r0d[3], o_0r1d[3]);
  DRAND2 I5 (termf_0n[4], termt_0n[4], termf_1n[4], termt_1n[4], o_0r0d[4], o_0r1d[4]);
  DRAND2 I6 (termf_0n[5], termt_0n[5], termf_1n[5], termt_1n[5], o_0r0d[5], o_0r1d[5]);
  DRAND2 I7 (termf_0n[6], termt_0n[6], termf_1n[6], termt_1n[6], o_0r0d[6], o_0r1d[6]);
  DRAND2 I8 (termf_0n[7], termt_0n[7], termf_1n[7], termt_1n[7], o_0r0d[7], o_0r1d[7]);
  DRAND2 I9 (termf_0n[8], termt_0n[8], termf_1n[8], termt_1n[8], o_0r0d[8], o_0r1d[8]);
  DRAND2 I10 (termf_0n[9], termt_0n[9], termf_1n[9], termt_1n[9], o_0r0d[9], o_0r1d[9]);
  DRAND2 I11 (termf_0n[10], termt_0n[10], termf_1n[10], termt_1n[10], o_0r0d[10], o_0r1d[10]);
  DRAND2 I12 (termf_0n[11], termt_0n[11], termf_1n[11], termt_1n[11], o_0r0d[11], o_0r1d[11]);
  DRAND2 I13 (termf_0n[12], termt_0n[12], termf_1n[12], termt_1n[12], o_0r0d[12], o_0r1d[12]);
  DRAND2 I14 (termf_0n[13], termt_0n[13], termf_1n[13], termt_1n[13], o_0r0d[13], o_0r1d[13]);
  DRAND2 I15 (termf_0n[14], termt_0n[14], termf_1n[14], termt_1n[14], o_0r0d[14], o_0r1d[14]);
  DRAND2 I16 (termf_0n[15], termt_0n[15], termf_1n[15], termt_1n[15], o_0r0d[15], o_0r1d[15]);
  DRAND2 I17 (termf_0n[16], termt_0n[16], termf_1n[16], termt_1n[16], o_0r0d[16], o_0r1d[16]);
  DRAND2 I18 (termf_0n[17], termt_0n[17], termf_1n[17], termt_1n[17], o_0r0d[17], o_0r1d[17]);
  DRAND2 I19 (termf_0n[18], termt_0n[18], termf_1n[18], termt_1n[18], o_0r0d[18], o_0r1d[18]);
  DRAND2 I20 (termf_0n[19], termt_0n[19], termf_1n[19], termt_1n[19], o_0r0d[19], o_0r1d[19]);
  DRAND2 I21 (termf_0n[20], termt_0n[20], termf_1n[20], termt_1n[20], o_0r0d[20], o_0r1d[20]);
  DRAND2 I22 (termf_0n[21], termt_0n[21], termf_1n[21], termt_1n[21], o_0r0d[21], o_0r1d[21]);
  DRAND2 I23 (termf_0n[22], termt_0n[22], termf_1n[22], termt_1n[22], o_0r0d[22], o_0r1d[22]);
  DRAND2 I24 (termf_0n[23], termt_0n[23], termf_1n[23], termt_1n[23], o_0r0d[23], o_0r1d[23]);
  DRAND2 I25 (termf_0n[24], termt_0n[24], termf_1n[24], termt_1n[24], o_0r0d[24], o_0r1d[24]);
  DRAND2 I26 (termf_0n[25], termt_0n[25], termf_1n[25], termt_1n[25], o_0r0d[25], o_0r1d[25]);
  DRAND2 I27 (termf_0n[26], termt_0n[26], termf_1n[26], termt_1n[26], o_0r0d[26], o_0r1d[26]);
  DRAND2 I28 (termf_0n[27], termt_0n[27], termf_1n[27], termt_1n[27], o_0r0d[27], o_0r1d[27]);
  DRAND2 I29 (termf_0n[28], termt_0n[28], termf_1n[28], termt_1n[28], o_0r0d[28], o_0r1d[28]);
  DRAND2 I30 (termf_0n[29], termt_0n[29], termf_1n[29], termt_1n[29], o_0r0d[29], o_0r1d[29]);
  DRAND2 I31 (termf_0n[30], termt_0n[30], termf_1n[30], termt_1n[30], o_0r0d[30], o_0r1d[30]);
  DRAND2 I32 (termf_0n[31], termt_0n[31], termf_1n[31], termt_1n[31], o_0r0d[31], o_0r1d[31]);
  DRAND2 I33 (termf_0n[32], termt_0n[32], termf_1n[32], termt_1n[32], o_0r0d[32], o_0r1d[32]);
  DRAND2 I34 (termf_0n[33], termt_0n[33], termf_1n[33], termt_1n[33], o_0r0d[33], o_0r1d[33]);
  DRAND2 I35 (termf_0n[34], termt_0n[34], termf_1n[34], termt_1n[34], o_0r0d[34], o_0r1d[34]);
  assign termt_1n[0] = i_0r1d[35];
  assign termt_1n[1] = i_0r1d[36];
  assign termt_1n[2] = i_0r1d[37];
  assign termt_1n[3] = i_0r1d[38];
  assign termt_1n[4] = i_0r1d[39];
  assign termt_1n[5] = i_0r1d[40];
  assign termt_1n[6] = i_0r1d[41];
  assign termt_1n[7] = i_0r1d[42];
  assign termt_1n[8] = i_0r1d[43];
  assign termt_1n[9] = i_0r1d[44];
  assign termt_1n[10] = i_0r1d[45];
  assign termt_1n[11] = i_0r1d[46];
  assign termt_1n[12] = i_0r1d[47];
  assign termt_1n[13] = i_0r1d[48];
  assign termt_1n[14] = i_0r1d[49];
  assign termt_1n[15] = i_0r1d[50];
  assign termt_1n[16] = i_0r1d[51];
  assign termt_1n[17] = i_0r1d[52];
  assign termt_1n[18] = i_0r1d[53];
  assign termt_1n[19] = i_0r1d[54];
  assign termt_1n[20] = i_0r1d[55];
  assign termt_1n[21] = i_0r1d[56];
  assign termt_1n[22] = i_0r1d[57];
  assign termt_1n[23] = i_0r1d[58];
  assign termt_1n[24] = i_0r1d[59];
  assign termt_1n[25] = i_0r1d[60];
  assign termt_1n[26] = i_0r1d[61];
  assign termt_1n[27] = i_0r1d[62];
  assign termt_1n[28] = i_0r1d[63];
  assign termt_1n[29] = i_0r1d[64];
  assign termt_1n[30] = i_0r1d[65];
  assign termt_1n[31] = i_0r1d[66];
  assign termt_1n[32] = i_0r1d[67];
  assign termt_1n[33] = i_0r1d[68];
  assign termt_1n[34] = i_0r1d[69];
  assign termf_1n[0] = i_0r0d[35];
  assign termf_1n[1] = i_0r0d[36];
  assign termf_1n[2] = i_0r0d[37];
  assign termf_1n[3] = i_0r0d[38];
  assign termf_1n[4] = i_0r0d[39];
  assign termf_1n[5] = i_0r0d[40];
  assign termf_1n[6] = i_0r0d[41];
  assign termf_1n[7] = i_0r0d[42];
  assign termf_1n[8] = i_0r0d[43];
  assign termf_1n[9] = i_0r0d[44];
  assign termf_1n[10] = i_0r0d[45];
  assign termf_1n[11] = i_0r0d[46];
  assign termf_1n[12] = i_0r0d[47];
  assign termf_1n[13] = i_0r0d[48];
  assign termf_1n[14] = i_0r0d[49];
  assign termf_1n[15] = i_0r0d[50];
  assign termf_1n[16] = i_0r0d[51];
  assign termf_1n[17] = i_0r0d[52];
  assign termf_1n[18] = i_0r0d[53];
  assign termf_1n[19] = i_0r0d[54];
  assign termf_1n[20] = i_0r0d[55];
  assign termf_1n[21] = i_0r0d[56];
  assign termf_1n[22] = i_0r0d[57];
  assign termf_1n[23] = i_0r0d[58];
  assign termf_1n[24] = i_0r0d[59];
  assign termf_1n[25] = i_0r0d[60];
  assign termf_1n[26] = i_0r0d[61];
  assign termf_1n[27] = i_0r0d[62];
  assign termf_1n[28] = i_0r0d[63];
  assign termf_1n[29] = i_0r0d[64];
  assign termf_1n[30] = i_0r0d[65];
  assign termf_1n[31] = i_0r0d[66];
  assign termf_1n[32] = i_0r0d[67];
  assign termf_1n[33] = i_0r0d[68];
  assign termf_1n[34] = i_0r0d[69];
  assign termt_0n[0] = i_0r1d[0];
  assign termt_0n[1] = i_0r1d[1];
  assign termt_0n[2] = i_0r1d[2];
  assign termt_0n[3] = i_0r1d[3];
  assign termt_0n[4] = i_0r1d[4];
  assign termt_0n[5] = i_0r1d[5];
  assign termt_0n[6] = i_0r1d[6];
  assign termt_0n[7] = i_0r1d[7];
  assign termt_0n[8] = i_0r1d[8];
  assign termt_0n[9] = i_0r1d[9];
  assign termt_0n[10] = i_0r1d[10];
  assign termt_0n[11] = i_0r1d[11];
  assign termt_0n[12] = i_0r1d[12];
  assign termt_0n[13] = i_0r1d[13];
  assign termt_0n[14] = i_0r1d[14];
  assign termt_0n[15] = i_0r1d[15];
  assign termt_0n[16] = i_0r1d[16];
  assign termt_0n[17] = i_0r1d[17];
  assign termt_0n[18] = i_0r1d[18];
  assign termt_0n[19] = i_0r1d[19];
  assign termt_0n[20] = i_0r1d[20];
  assign termt_0n[21] = i_0r1d[21];
  assign termt_0n[22] = i_0r1d[22];
  assign termt_0n[23] = i_0r1d[23];
  assign termt_0n[24] = i_0r1d[24];
  assign termt_0n[25] = i_0r1d[25];
  assign termt_0n[26] = i_0r1d[26];
  assign termt_0n[27] = i_0r1d[27];
  assign termt_0n[28] = i_0r1d[28];
  assign termt_0n[29] = i_0r1d[29];
  assign termt_0n[30] = i_0r1d[30];
  assign termt_0n[31] = i_0r1d[31];
  assign termt_0n[32] = i_0r1d[32];
  assign termt_0n[33] = i_0r1d[33];
  assign termt_0n[34] = i_0r1d[34];
  assign termf_0n[0] = i_0r0d[0];
  assign termf_0n[1] = i_0r0d[1];
  assign termf_0n[2] = i_0r0d[2];
  assign termf_0n[3] = i_0r0d[3];
  assign termf_0n[4] = i_0r0d[4];
  assign termf_0n[5] = i_0r0d[5];
  assign termf_0n[6] = i_0r0d[6];
  assign termf_0n[7] = i_0r0d[7];
  assign termf_0n[8] = i_0r0d[8];
  assign termf_0n[9] = i_0r0d[9];
  assign termf_0n[10] = i_0r0d[10];
  assign termf_0n[11] = i_0r0d[11];
  assign termf_0n[12] = i_0r0d[12];
  assign termf_0n[13] = i_0r0d[13];
  assign termf_0n[14] = i_0r0d[14];
  assign termf_0n[15] = i_0r0d[15];
  assign termf_0n[16] = i_0r0d[16];
  assign termf_0n[17] = i_0r0d[17];
  assign termf_0n[18] = i_0r0d[18];
  assign termf_0n[19] = i_0r0d[19];
  assign termf_0n[20] = i_0r0d[20];
  assign termf_0n[21] = i_0r0d[21];
  assign termf_0n[22] = i_0r0d[22];
  assign termf_0n[23] = i_0r0d[23];
  assign termf_0n[24] = i_0r0d[24];
  assign termf_0n[25] = i_0r0d[25];
  assign termf_0n[26] = i_0r0d[26];
  assign termf_0n[27] = i_0r0d[27];
  assign termf_0n[28] = i_0r0d[28];
  assign termf_0n[29] = i_0r0d[29];
  assign termf_0n[30] = i_0r0d[30];
  assign termf_0n[31] = i_0r0d[31];
  assign termf_0n[32] = i_0r0d[32];
  assign termf_0n[33] = i_0r0d[33];
  assign termf_0n[34] = i_0r0d[34];
endmodule

module DROR2 (
  i0_0,
  i0_1,
  i1_0,
  i1_1,
  q_0,
  q_1
);
  input i0_0;
  input i0_1;
  input i1_0;
  input i1_1;
  output q_0;
  output q_1;
  wire n0_0n;
  wire n1_0n;
  wire n2_0n;
  C2 I0 (q_0, i0_0, i1_0);
  OR3 I1 (q_1, n0_0n, n1_0n, n2_0n);
  C2 I2 (n2_0n, i0_1, i1_1);
  C2 I3 (n1_0n, i0_1, i1_0);
  C2 I4 (n0_0n, i0_0, i1_1);
endmodule

module BrzO_70_35_l123__28_28app_201_20_280_200_2_m59m (
  i_0r0d, i_0r1d, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input [69:0] i_0r0d;
  input [69:0] i_0r1d;
  output i_0a;
  output [34:0] o_0r0d;
  output [34:0] o_0r1d;
  input o_0a;
  wire [34:0] termf_0n;
  wire [34:0] termf_1n;
  wire [34:0] termt_0n;
  wire [34:0] termt_1n;
  assign i_0a = o_0a;
  DROR2 I1 (termf_0n[0], termt_0n[0], termf_1n[0], termt_1n[0], o_0r0d[0], o_0r1d[0]);
  DROR2 I2 (termf_0n[1], termt_0n[1], termf_1n[1], termt_1n[1], o_0r0d[1], o_0r1d[1]);
  DROR2 I3 (termf_0n[2], termt_0n[2], termf_1n[2], termt_1n[2], o_0r0d[2], o_0r1d[2]);
  DROR2 I4 (termf_0n[3], termt_0n[3], termf_1n[3], termt_1n[3], o_0r0d[3], o_0r1d[3]);
  DROR2 I5 (termf_0n[4], termt_0n[4], termf_1n[4], termt_1n[4], o_0r0d[4], o_0r1d[4]);
  DROR2 I6 (termf_0n[5], termt_0n[5], termf_1n[5], termt_1n[5], o_0r0d[5], o_0r1d[5]);
  DROR2 I7 (termf_0n[6], termt_0n[6], termf_1n[6], termt_1n[6], o_0r0d[6], o_0r1d[6]);
  DROR2 I8 (termf_0n[7], termt_0n[7], termf_1n[7], termt_1n[7], o_0r0d[7], o_0r1d[7]);
  DROR2 I9 (termf_0n[8], termt_0n[8], termf_1n[8], termt_1n[8], o_0r0d[8], o_0r1d[8]);
  DROR2 I10 (termf_0n[9], termt_0n[9], termf_1n[9], termt_1n[9], o_0r0d[9], o_0r1d[9]);
  DROR2 I11 (termf_0n[10], termt_0n[10], termf_1n[10], termt_1n[10], o_0r0d[10], o_0r1d[10]);
  DROR2 I12 (termf_0n[11], termt_0n[11], termf_1n[11], termt_1n[11], o_0r0d[11], o_0r1d[11]);
  DROR2 I13 (termf_0n[12], termt_0n[12], termf_1n[12], termt_1n[12], o_0r0d[12], o_0r1d[12]);
  DROR2 I14 (termf_0n[13], termt_0n[13], termf_1n[13], termt_1n[13], o_0r0d[13], o_0r1d[13]);
  DROR2 I15 (termf_0n[14], termt_0n[14], termf_1n[14], termt_1n[14], o_0r0d[14], o_0r1d[14]);
  DROR2 I16 (termf_0n[15], termt_0n[15], termf_1n[15], termt_1n[15], o_0r0d[15], o_0r1d[15]);
  DROR2 I17 (termf_0n[16], termt_0n[16], termf_1n[16], termt_1n[16], o_0r0d[16], o_0r1d[16]);
  DROR2 I18 (termf_0n[17], termt_0n[17], termf_1n[17], termt_1n[17], o_0r0d[17], o_0r1d[17]);
  DROR2 I19 (termf_0n[18], termt_0n[18], termf_1n[18], termt_1n[18], o_0r0d[18], o_0r1d[18]);
  DROR2 I20 (termf_0n[19], termt_0n[19], termf_1n[19], termt_1n[19], o_0r0d[19], o_0r1d[19]);
  DROR2 I21 (termf_0n[20], termt_0n[20], termf_1n[20], termt_1n[20], o_0r0d[20], o_0r1d[20]);
  DROR2 I22 (termf_0n[21], termt_0n[21], termf_1n[21], termt_1n[21], o_0r0d[21], o_0r1d[21]);
  DROR2 I23 (termf_0n[22], termt_0n[22], termf_1n[22], termt_1n[22], o_0r0d[22], o_0r1d[22]);
  DROR2 I24 (termf_0n[23], termt_0n[23], termf_1n[23], termt_1n[23], o_0r0d[23], o_0r1d[23]);
  DROR2 I25 (termf_0n[24], termt_0n[24], termf_1n[24], termt_1n[24], o_0r0d[24], o_0r1d[24]);
  DROR2 I26 (termf_0n[25], termt_0n[25], termf_1n[25], termt_1n[25], o_0r0d[25], o_0r1d[25]);
  DROR2 I27 (termf_0n[26], termt_0n[26], termf_1n[26], termt_1n[26], o_0r0d[26], o_0r1d[26]);
  DROR2 I28 (termf_0n[27], termt_0n[27], termf_1n[27], termt_1n[27], o_0r0d[27], o_0r1d[27]);
  DROR2 I29 (termf_0n[28], termt_0n[28], termf_1n[28], termt_1n[28], o_0r0d[28], o_0r1d[28]);
  DROR2 I30 (termf_0n[29], termt_0n[29], termf_1n[29], termt_1n[29], o_0r0d[29], o_0r1d[29]);
  DROR2 I31 (termf_0n[30], termt_0n[30], termf_1n[30], termt_1n[30], o_0r0d[30], o_0r1d[30]);
  DROR2 I32 (termf_0n[31], termt_0n[31], termf_1n[31], termt_1n[31], o_0r0d[31], o_0r1d[31]);
  DROR2 I33 (termf_0n[32], termt_0n[32], termf_1n[32], termt_1n[32], o_0r0d[32], o_0r1d[32]);
  DROR2 I34 (termf_0n[33], termt_0n[33], termf_1n[33], termt_1n[33], o_0r0d[33], o_0r1d[33]);
  DROR2 I35 (termf_0n[34], termt_0n[34], termf_1n[34], termt_1n[34], o_0r0d[34], o_0r1d[34]);
  assign termt_1n[0] = i_0r1d[35];
  assign termt_1n[1] = i_0r1d[36];
  assign termt_1n[2] = i_0r1d[37];
  assign termt_1n[3] = i_0r1d[38];
  assign termt_1n[4] = i_0r1d[39];
  assign termt_1n[5] = i_0r1d[40];
  assign termt_1n[6] = i_0r1d[41];
  assign termt_1n[7] = i_0r1d[42];
  assign termt_1n[8] = i_0r1d[43];
  assign termt_1n[9] = i_0r1d[44];
  assign termt_1n[10] = i_0r1d[45];
  assign termt_1n[11] = i_0r1d[46];
  assign termt_1n[12] = i_0r1d[47];
  assign termt_1n[13] = i_0r1d[48];
  assign termt_1n[14] = i_0r1d[49];
  assign termt_1n[15] = i_0r1d[50];
  assign termt_1n[16] = i_0r1d[51];
  assign termt_1n[17] = i_0r1d[52];
  assign termt_1n[18] = i_0r1d[53];
  assign termt_1n[19] = i_0r1d[54];
  assign termt_1n[20] = i_0r1d[55];
  assign termt_1n[21] = i_0r1d[56];
  assign termt_1n[22] = i_0r1d[57];
  assign termt_1n[23] = i_0r1d[58];
  assign termt_1n[24] = i_0r1d[59];
  assign termt_1n[25] = i_0r1d[60];
  assign termt_1n[26] = i_0r1d[61];
  assign termt_1n[27] = i_0r1d[62];
  assign termt_1n[28] = i_0r1d[63];
  assign termt_1n[29] = i_0r1d[64];
  assign termt_1n[30] = i_0r1d[65];
  assign termt_1n[31] = i_0r1d[66];
  assign termt_1n[32] = i_0r1d[67];
  assign termt_1n[33] = i_0r1d[68];
  assign termt_1n[34] = i_0r1d[69];
  assign termf_1n[0] = i_0r0d[35];
  assign termf_1n[1] = i_0r0d[36];
  assign termf_1n[2] = i_0r0d[37];
  assign termf_1n[3] = i_0r0d[38];
  assign termf_1n[4] = i_0r0d[39];
  assign termf_1n[5] = i_0r0d[40];
  assign termf_1n[6] = i_0r0d[41];
  assign termf_1n[7] = i_0r0d[42];
  assign termf_1n[8] = i_0r0d[43];
  assign termf_1n[9] = i_0r0d[44];
  assign termf_1n[10] = i_0r0d[45];
  assign termf_1n[11] = i_0r0d[46];
  assign termf_1n[12] = i_0r0d[47];
  assign termf_1n[13] = i_0r0d[48];
  assign termf_1n[14] = i_0r0d[49];
  assign termf_1n[15] = i_0r0d[50];
  assign termf_1n[16] = i_0r0d[51];
  assign termf_1n[17] = i_0r0d[52];
  assign termf_1n[18] = i_0r0d[53];
  assign termf_1n[19] = i_0r0d[54];
  assign termf_1n[20] = i_0r0d[55];
  assign termf_1n[21] = i_0r0d[56];
  assign termf_1n[22] = i_0r0d[57];
  assign termf_1n[23] = i_0r0d[58];
  assign termf_1n[24] = i_0r0d[59];
  assign termf_1n[25] = i_0r0d[60];
  assign termf_1n[26] = i_0r0d[61];
  assign termf_1n[27] = i_0r0d[62];
  assign termf_1n[28] = i_0r0d[63];
  assign termf_1n[29] = i_0r0d[64];
  assign termf_1n[30] = i_0r0d[65];
  assign termf_1n[31] = i_0r0d[66];
  assign termf_1n[32] = i_0r0d[67];
  assign termf_1n[33] = i_0r0d[68];
  assign termf_1n[34] = i_0r0d[69];
  assign termt_0n[0] = i_0r1d[0];
  assign termt_0n[1] = i_0r1d[1];
  assign termt_0n[2] = i_0r1d[2];
  assign termt_0n[3] = i_0r1d[3];
  assign termt_0n[4] = i_0r1d[4];
  assign termt_0n[5] = i_0r1d[5];
  assign termt_0n[6] = i_0r1d[6];
  assign termt_0n[7] = i_0r1d[7];
  assign termt_0n[8] = i_0r1d[8];
  assign termt_0n[9] = i_0r1d[9];
  assign termt_0n[10] = i_0r1d[10];
  assign termt_0n[11] = i_0r1d[11];
  assign termt_0n[12] = i_0r1d[12];
  assign termt_0n[13] = i_0r1d[13];
  assign termt_0n[14] = i_0r1d[14];
  assign termt_0n[15] = i_0r1d[15];
  assign termt_0n[16] = i_0r1d[16];
  assign termt_0n[17] = i_0r1d[17];
  assign termt_0n[18] = i_0r1d[18];
  assign termt_0n[19] = i_0r1d[19];
  assign termt_0n[20] = i_0r1d[20];
  assign termt_0n[21] = i_0r1d[21];
  assign termt_0n[22] = i_0r1d[22];
  assign termt_0n[23] = i_0r1d[23];
  assign termt_0n[24] = i_0r1d[24];
  assign termt_0n[25] = i_0r1d[25];
  assign termt_0n[26] = i_0r1d[26];
  assign termt_0n[27] = i_0r1d[27];
  assign termt_0n[28] = i_0r1d[28];
  assign termt_0n[29] = i_0r1d[29];
  assign termt_0n[30] = i_0r1d[30];
  assign termt_0n[31] = i_0r1d[31];
  assign termt_0n[32] = i_0r1d[32];
  assign termt_0n[33] = i_0r1d[33];
  assign termt_0n[34] = i_0r1d[34];
  assign termf_0n[0] = i_0r0d[0];
  assign termf_0n[1] = i_0r0d[1];
  assign termf_0n[2] = i_0r0d[2];
  assign termf_0n[3] = i_0r0d[3];
  assign termf_0n[4] = i_0r0d[4];
  assign termf_0n[5] = i_0r0d[5];
  assign termf_0n[6] = i_0r0d[6];
  assign termf_0n[7] = i_0r0d[7];
  assign termf_0n[8] = i_0r0d[8];
  assign termf_0n[9] = i_0r0d[9];
  assign termf_0n[10] = i_0r0d[10];
  assign termf_0n[11] = i_0r0d[11];
  assign termf_0n[12] = i_0r0d[12];
  assign termf_0n[13] = i_0r0d[13];
  assign termf_0n[14] = i_0r0d[14];
  assign termf_0n[15] = i_0r0d[15];
  assign termf_0n[16] = i_0r0d[16];
  assign termf_0n[17] = i_0r0d[17];
  assign termf_0n[18] = i_0r0d[18];
  assign termf_0n[19] = i_0r0d[19];
  assign termf_0n[20] = i_0r0d[20];
  assign termf_0n[21] = i_0r0d[21];
  assign termf_0n[22] = i_0r0d[22];
  assign termf_0n[23] = i_0r0d[23];
  assign termf_0n[24] = i_0r0d[24];
  assign termf_0n[25] = i_0r0d[25];
  assign termf_0n[26] = i_0r0d[26];
  assign termf_0n[27] = i_0r0d[27];
  assign termf_0n[28] = i_0r0d[28];
  assign termf_0n[29] = i_0r0d[29];
  assign termf_0n[30] = i_0r0d[30];
  assign termf_0n[31] = i_0r0d[31];
  assign termf_0n[32] = i_0r0d[32];
  assign termf_0n[33] = i_0r0d[33];
  assign termf_0n[34] = i_0r0d[34];
endmodule

module BrzO_70_35_l124__28_28app_201_20_280_200_2_m60m (
  i_0r0d, i_0r1d, i_0a,
  o_0r0d, o_0r1d, o_0a
);
  input [69:0] i_0r0d;
  input [69:0] i_0r1d;
  output i_0a;
  output [34:0] o_0r0d;
  output [34:0] o_0r1d;
  input o_0a;
  wire [34:0] termf_0n;
  wire [34:0] termf_1n;
  wire [34:0] termt_0n;
  wire [34:0] termt_1n;
  assign i_0a = o_0a;
  DRXOR2 I1 (termf_0n[0], termt_0n[0], termf_1n[0], termt_1n[0], o_0r0d[0], o_0r1d[0]);
  DRXOR2 I2 (termf_0n[1], termt_0n[1], termf_1n[1], termt_1n[1], o_0r0d[1], o_0r1d[1]);
  DRXOR2 I3 (termf_0n[2], termt_0n[2], termf_1n[2], termt_1n[2], o_0r0d[2], o_0r1d[2]);
  DRXOR2 I4 (termf_0n[3], termt_0n[3], termf_1n[3], termt_1n[3], o_0r0d[3], o_0r1d[3]);
  DRXOR2 I5 (termf_0n[4], termt_0n[4], termf_1n[4], termt_1n[4], o_0r0d[4], o_0r1d[4]);
  DRXOR2 I6 (termf_0n[5], termt_0n[5], termf_1n[5], termt_1n[5], o_0r0d[5], o_0r1d[5]);
  DRXOR2 I7 (termf_0n[6], termt_0n[6], termf_1n[6], termt_1n[6], o_0r0d[6], o_0r1d[6]);
  DRXOR2 I8 (termf_0n[7], termt_0n[7], termf_1n[7], termt_1n[7], o_0r0d[7], o_0r1d[7]);
  DRXOR2 I9 (termf_0n[8], termt_0n[8], termf_1n[8], termt_1n[8], o_0r0d[8], o_0r1d[8]);
  DRXOR2 I10 (termf_0n[9], termt_0n[9], termf_1n[9], termt_1n[9], o_0r0d[9], o_0r1d[9]);
  DRXOR2 I11 (termf_0n[10], termt_0n[10], termf_1n[10], termt_1n[10], o_0r0d[10], o_0r1d[10]);
  DRXOR2 I12 (termf_0n[11], termt_0n[11], termf_1n[11], termt_1n[11], o_0r0d[11], o_0r1d[11]);
  DRXOR2 I13 (termf_0n[12], termt_0n[12], termf_1n[12], termt_1n[12], o_0r0d[12], o_0r1d[12]);
  DRXOR2 I14 (termf_0n[13], termt_0n[13], termf_1n[13], termt_1n[13], o_0r0d[13], o_0r1d[13]);
  DRXOR2 I15 (termf_0n[14], termt_0n[14], termf_1n[14], termt_1n[14], o_0r0d[14], o_0r1d[14]);
  DRXOR2 I16 (termf_0n[15], termt_0n[15], termf_1n[15], termt_1n[15], o_0r0d[15], o_0r1d[15]);
  DRXOR2 I17 (termf_0n[16], termt_0n[16], termf_1n[16], termt_1n[16], o_0r0d[16], o_0r1d[16]);
  DRXOR2 I18 (termf_0n[17], termt_0n[17], termf_1n[17], termt_1n[17], o_0r0d[17], o_0r1d[17]);
  DRXOR2 I19 (termf_0n[18], termt_0n[18], termf_1n[18], termt_1n[18], o_0r0d[18], o_0r1d[18]);
  DRXOR2 I20 (termf_0n[19], termt_0n[19], termf_1n[19], termt_1n[19], o_0r0d[19], o_0r1d[19]);
  DRXOR2 I21 (termf_0n[20], termt_0n[20], termf_1n[20], termt_1n[20], o_0r0d[20], o_0r1d[20]);
  DRXOR2 I22 (termf_0n[21], termt_0n[21], termf_1n[21], termt_1n[21], o_0r0d[21], o_0r1d[21]);
  DRXOR2 I23 (termf_0n[22], termt_0n[22], termf_1n[22], termt_1n[22], o_0r0d[22], o_0r1d[22]);
  DRXOR2 I24 (termf_0n[23], termt_0n[23], termf_1n[23], termt_1n[23], o_0r0d[23], o_0r1d[23]);
  DRXOR2 I25 (termf_0n[24], termt_0n[24], termf_1n[24], termt_1n[24], o_0r0d[24], o_0r1d[24]);
  DRXOR2 I26 (termf_0n[25], termt_0n[25], termf_1n[25], termt_1n[25], o_0r0d[25], o_0r1d[25]);
  DRXOR2 I27 (termf_0n[26], termt_0n[26], termf_1n[26], termt_1n[26], o_0r0d[26], o_0r1d[26]);
  DRXOR2 I28 (termf_0n[27], termt_0n[27], termf_1n[27], termt_1n[27], o_0r0d[27], o_0r1d[27]);
  DRXOR2 I29 (termf_0n[28], termt_0n[28], termf_1n[28], termt_1n[28], o_0r0d[28], o_0r1d[28]);
  DRXOR2 I30 (termf_0n[29], termt_0n[29], termf_1n[29], termt_1n[29], o_0r0d[29], o_0r1d[29]);
  DRXOR2 I31 (termf_0n[30], termt_0n[30], termf_1n[30], termt_1n[30], o_0r0d[30], o_0r1d[30]);
  DRXOR2 I32 (termf_0n[31], termt_0n[31], termf_1n[31], termt_1n[31], o_0r0d[31], o_0r1d[31]);
  DRXOR2 I33 (termf_0n[32], termt_0n[32], termf_1n[32], termt_1n[32], o_0r0d[32], o_0r1d[32]);
  DRXOR2 I34 (termf_0n[33], termt_0n[33], termf_1n[33], termt_1n[33], o_0r0d[33], o_0r1d[33]);
  DRXOR2 I35 (termf_0n[34], termt_0n[34], termf_1n[34], termt_1n[34], o_0r0d[34], o_0r1d[34]);
  assign termt_1n[0] = i_0r1d[35];
  assign termt_1n[1] = i_0r1d[36];
  assign termt_1n[2] = i_0r1d[37];
  assign termt_1n[3] = i_0r1d[38];
  assign termt_1n[4] = i_0r1d[39];
  assign termt_1n[5] = i_0r1d[40];
  assign termt_1n[6] = i_0r1d[41];
  assign termt_1n[7] = i_0r1d[42];
  assign termt_1n[8] = i_0r1d[43];
  assign termt_1n[9] = i_0r1d[44];
  assign termt_1n[10] = i_0r1d[45];
  assign termt_1n[11] = i_0r1d[46];
  assign termt_1n[12] = i_0r1d[47];
  assign termt_1n[13] = i_0r1d[48];
  assign termt_1n[14] = i_0r1d[49];
  assign termt_1n[15] = i_0r1d[50];
  assign termt_1n[16] = i_0r1d[51];
  assign termt_1n[17] = i_0r1d[52];
  assign termt_1n[18] = i_0r1d[53];
  assign termt_1n[19] = i_0r1d[54];
  assign termt_1n[20] = i_0r1d[55];
  assign termt_1n[21] = i_0r1d[56];
  assign termt_1n[22] = i_0r1d[57];
  assign termt_1n[23] = i_0r1d[58];
  assign termt_1n[24] = i_0r1d[59];
  assign termt_1n[25] = i_0r1d[60];
  assign termt_1n[26] = i_0r1d[61];
  assign termt_1n[27] = i_0r1d[62];
  assign termt_1n[28] = i_0r1d[63];
  assign termt_1n[29] = i_0r1d[64];
  assign termt_1n[30] = i_0r1d[65];
  assign termt_1n[31] = i_0r1d[66];
  assign termt_1n[32] = i_0r1d[67];
  assign termt_1n[33] = i_0r1d[68];
  assign termt_1n[34] = i_0r1d[69];
  assign termf_1n[0] = i_0r0d[35];
  assign termf_1n[1] = i_0r0d[36];
  assign termf_1n[2] = i_0r0d[37];
  assign termf_1n[3] = i_0r0d[38];
  assign termf_1n[4] = i_0r0d[39];
  assign termf_1n[5] = i_0r0d[40];
  assign termf_1n[6] = i_0r0d[41];
  assign termf_1n[7] = i_0r0d[42];
  assign termf_1n[8] = i_0r0d[43];
  assign termf_1n[9] = i_0r0d[44];
  assign termf_1n[10] = i_0r0d[45];
  assign termf_1n[11] = i_0r0d[46];
  assign termf_1n[12] = i_0r0d[47];
  assign termf_1n[13] = i_0r0d[48];
  assign termf_1n[14] = i_0r0d[49];
  assign termf_1n[15] = i_0r0d[50];
  assign termf_1n[16] = i_0r0d[51];
  assign termf_1n[17] = i_0r0d[52];
  assign termf_1n[18] = i_0r0d[53];
  assign termf_1n[19] = i_0r0d[54];
  assign termf_1n[20] = i_0r0d[55];
  assign termf_1n[21] = i_0r0d[56];
  assign termf_1n[22] = i_0r0d[57];
  assign termf_1n[23] = i_0r0d[58];
  assign termf_1n[24] = i_0r0d[59];
  assign termf_1n[25] = i_0r0d[60];
  assign termf_1n[26] = i_0r0d[61];
  assign termf_1n[27] = i_0r0d[62];
  assign termf_1n[28] = i_0r0d[63];
  assign termf_1n[29] = i_0r0d[64];
  assign termf_1n[30] = i_0r0d[65];
  assign termf_1n[31] = i_0r0d[66];
  assign termf_1n[32] = i_0r0d[67];
  assign termf_1n[33] = i_0r0d[68];
  assign termf_1n[34] = i_0r0d[69];
  assign termt_0n[0] = i_0r1d[0];
  assign termt_0n[1] = i_0r1d[1];
  assign termt_0n[2] = i_0r1d[2];
  assign termt_0n[3] = i_0r1d[3];
  assign termt_0n[4] = i_0r1d[4];
  assign termt_0n[5] = i_0r1d[5];
  assign termt_0n[6] = i_0r1d[6];
  assign termt_0n[7] = i_0r1d[7];
  assign termt_0n[8] = i_0r1d[8];
  assign termt_0n[9] = i_0r1d[9];
  assign termt_0n[10] = i_0r1d[10];
  assign termt_0n[11] = i_0r1d[11];
  assign termt_0n[12] = i_0r1d[12];
  assign termt_0n[13] = i_0r1d[13];
  assign termt_0n[14] = i_0r1d[14];
  assign termt_0n[15] = i_0r1d[15];
  assign termt_0n[16] = i_0r1d[16];
  assign termt_0n[17] = i_0r1d[17];
  assign termt_0n[18] = i_0r1d[18];
  assign termt_0n[19] = i_0r1d[19];
  assign termt_0n[20] = i_0r1d[20];
  assign termt_0n[21] = i_0r1d[21];
  assign termt_0n[22] = i_0r1d[22];
  assign termt_0n[23] = i_0r1d[23];
  assign termt_0n[24] = i_0r1d[24];
  assign termt_0n[25] = i_0r1d[25];
  assign termt_0n[26] = i_0r1d[26];
  assign termt_0n[27] = i_0r1d[27];
  assign termt_0n[28] = i_0r1d[28];
  assign termt_0n[29] = i_0r1d[29];
  assign termt_0n[30] = i_0r1d[30];
  assign termt_0n[31] = i_0r1d[31];
  assign termt_0n[32] = i_0r1d[32];
  assign termt_0n[33] = i_0r1d[33];
  assign termt_0n[34] = i_0r1d[34];
  assign termf_0n[0] = i_0r0d[0];
  assign termf_0n[1] = i_0r0d[1];
  assign termf_0n[2] = i_0r0d[2];
  assign termf_0n[3] = i_0r0d[3];
  assign termf_0n[4] = i_0r0d[4];
  assign termf_0n[5] = i_0r0d[5];
  assign termf_0n[6] = i_0r0d[6];
  assign termf_0n[7] = i_0r0d[7];
  assign termf_0n[8] = i_0r0d[8];
  assign termf_0n[9] = i_0r0d[9];
  assign termf_0n[10] = i_0r0d[10];
  assign termf_0n[11] = i_0r0d[11];
  assign termf_0n[12] = i_0r0d[12];
  assign termf_0n[13] = i_0r0d[13];
  assign termf_0n[14] = i_0r0d[14];
  assign termf_0n[15] = i_0r0d[15];
  assign termf_0n[16] = i_0r0d[16];
  assign termf_0n[17] = i_0r0d[17];
  assign termf_0n[18] = i_0r0d[18];
  assign termf_0n[19] = i_0r0d[19];
  assign termf_0n[20] = i_0r0d[20];
  assign termf_0n[21] = i_0r0d[21];
  assign termf_0n[22] = i_0r0d[22];
  assign termf_0n[23] = i_0r0d[23];
  assign termf_0n[24] = i_0r0d[24];
  assign termf_0n[25] = i_0r0d[25];
  assign termf_0n[26] = i_0r0d[26];
  assign termf_0n[27] = i_0r0d[27];
  assign termf_0n[28] = i_0r0d[28];
  assign termf_0n[29] = i_0r0d[29];
  assign termf_0n[30] = i_0r0d[30];
  assign termf_0n[31] = i_0r0d[31];
  assign termf_0n[32] = i_0r0d[32];
  assign termf_0n[33] = i_0r0d[33];
  assign termf_0n[34] = i_0r0d[34];
endmodule

module BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m (
  i_0r0d, i_0r1d, i_0a,
  o_0r, o_0a,
  o_1r, o_1a,
  initialise
);
  input i_0r0d;
  input i_0r1d;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input initialise;
  wire icomplete_0n;
  wire sel_0n;
  wire sel_1n;
  wire matchi_0n;
  wire matchi_1n;
  wire ifint_0n;
  wire itint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire ofint_1n;
  wire oaint_0n;
  wire oaint_1n;
  wire oack_0n;
  wire gate1001_0n;
  wire gate998_0n;
  wire complete995_0n;
  wire gate994_0n;
  wire complete991_0n;
  C2 I0 (iaint_0n, oack_0n, icomplete_0n);
  OR2 I1 (oack_0n, oaint_0n, oaint_1n);
  assign oaint_1n = o_1r;
  INV I3 (gate1001_0n, o_1a);
  C2RI I4 (o_1r, ofint_1n, gate1001_0n, initialise);
  assign oaint_0n = o_0r;
  INV I6 (gate998_0n, o_0a);
  C2RI I7 (o_0r, ofint_0n, gate998_0n, initialise);
  assign i_0a = complete995_0n;
  OR2 I9 (complete995_0n, ifint_0n, itint_0n);
  INV I10 (gate994_0n, iaint_0n);
  C2RI I11 (itint_0n, i_0r1d, gate994_0n, initialise);
  C2RI I12 (ifint_0n, i_0r0d, gate994_0n, initialise);
  assign ofint_1n = sel_1n;
  assign ofint_0n = sel_0n;
  assign icomplete_0n = complete991_0n;
  OR2 I16 (complete991_0n, ifint_0n, itint_0n);
  assign matchi_1n = itint_0n;
  assign sel_1n = matchi_1n;
  assign matchi_0n = ifint_0n;
  assign sel_0n = matchi_0n;
endmodule

module BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m (
  i_0r0d, i_0r1d, i_0a,
  o_0r, o_0a,
  o_1r, o_1a,
  initialise
);
  input [1:0] i_0r0d;
  input [1:0] i_0r1d;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input initialise;
  wire icomplete_0n;
  wire sel_0n;
  wire sel_1n;
  wire matchi_0n;
  wire matchi_1n;
  wire [1:0] ifint_0n;
  wire [1:0] itint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire ofint_1n;
  wire oaint_0n;
  wire oaint_1n;
  wire oack_0n;
  wire gate1012_0n;
  wire gate1009_0n;
  wire [1:0] complete1006_0n;
  wire gate1005_0n;
  wire [1:0] complete1002_0n;
  C2 I0 (iaint_0n, oack_0n, icomplete_0n);
  OR2 I1 (oack_0n, oaint_0n, oaint_1n);
  assign oaint_1n = o_1r;
  INV I3 (gate1012_0n, o_1a);
  C2RI I4 (o_1r, ofint_1n, gate1012_0n, initialise);
  assign oaint_0n = o_0r;
  INV I6 (gate1009_0n, o_0a);
  C2RI I7 (o_0r, ofint_0n, gate1009_0n, initialise);
  C2 I8 (i_0a, complete1006_0n[0], complete1006_0n[1]);
  OR2 I9 (complete1006_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I10 (complete1006_0n[1], ifint_0n[1], itint_0n[1]);
  INV I11 (gate1005_0n, iaint_0n);
  C2RI I12 (itint_0n[0], i_0r1d[0], gate1005_0n, initialise);
  C2RI I13 (itint_0n[1], i_0r1d[1], gate1005_0n, initialise);
  C2RI I14 (ifint_0n[0], i_0r0d[0], gate1005_0n, initialise);
  C2RI I15 (ifint_0n[1], i_0r0d[1], gate1005_0n, initialise);
  assign ofint_1n = sel_1n;
  assign ofint_0n = sel_0n;
  C2 I18 (icomplete_0n, complete1002_0n[0], complete1002_0n[1]);
  OR2 I19 (complete1002_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I20 (complete1002_0n[1], ifint_0n[1], itint_0n[1]);
  C2 I21 (matchi_1n, ifint_0n[0], itint_0n[1]);
  assign sel_1n = matchi_1n;
  C2 I23 (matchi_0n, ifint_0n[1], itint_0n[0]);
  assign sel_0n = matchi_0n;
endmodule

module BrzS_3_l11__280_203_29_l137__28_28_28_280__m63m (
  i_0r0d, i_0r1d, i_0a,
  o_0r, o_0a,
  o_1r, o_1a,
  initialise
);
  input [2:0] i_0r0d;
  input [2:0] i_0r1d;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input initialise;
  wire icomplete_0n;
  wire sel_0n;
  wire sel_1n;
  wire [1:0] matchi_0n;
  wire [2:0] matchi_1n;
  wire [2:0] ifint_0n;
  wire [2:0] itint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire ofint_1n;
  wire oaint_0n;
  wire oaint_1n;
  wire oack_0n;
  wire gate1023_0n;
  wire gate1020_0n;
  wire [2:0] complete1017_0n;
  wire gate1016_0n;
  wire [2:0] complete1013_0n;
  C2 I0 (iaint_0n, oack_0n, icomplete_0n);
  OR2 I1 (oack_0n, oaint_0n, oaint_1n);
  assign oaint_1n = o_1r;
  INV I3 (gate1023_0n, o_1a);
  C2RI I4 (o_1r, ofint_1n, gate1023_0n, initialise);
  assign oaint_0n = o_0r;
  INV I6 (gate1020_0n, o_0a);
  C2RI I7 (o_0r, ofint_0n, gate1020_0n, initialise);
  C3 I8 (i_0a, complete1017_0n[0], complete1017_0n[1], complete1017_0n[2]);
  OR2 I9 (complete1017_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I10 (complete1017_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I11 (complete1017_0n[2], ifint_0n[2], itint_0n[2]);
  INV I12 (gate1016_0n, iaint_0n);
  C2RI I13 (itint_0n[0], i_0r1d[0], gate1016_0n, initialise);
  C2RI I14 (itint_0n[1], i_0r1d[1], gate1016_0n, initialise);
  C2RI I15 (itint_0n[2], i_0r1d[2], gate1016_0n, initialise);
  C2RI I16 (ifint_0n[0], i_0r0d[0], gate1016_0n, initialise);
  C2RI I17 (ifint_0n[1], i_0r0d[1], gate1016_0n, initialise);
  C2RI I18 (ifint_0n[2], i_0r0d[2], gate1016_0n, initialise);
  assign ofint_1n = sel_1n;
  assign ofint_0n = sel_0n;
  C3 I21 (icomplete_0n, complete1013_0n[0], complete1013_0n[1], complete1013_0n[2]);
  OR2 I22 (complete1013_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I23 (complete1013_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I24 (complete1013_0n[2], ifint_0n[2], itint_0n[2]);
  C3 I25 (matchi_1n[2], itint_0n[2], itint_0n[1], itint_0n[0]);
  C3 I26 (matchi_1n[1], ifint_0n[1], itint_0n[2], itint_0n[0]);
  C3 I27 (matchi_1n[0], ifint_0n[2], ifint_0n[1], itint_0n[0]);
  OR3 I28 (sel_1n, matchi_1n[0], matchi_1n[1], matchi_1n[2]);
  C3 I29 (matchi_0n[1], ifint_0n[2], itint_0n[1], itint_0n[0]);
  assign matchi_0n[0] = ifint_0n[0];
  OR2 I31 (sel_0n, matchi_0n[0], matchi_0n[1]);
endmodule

module BrzS_3_l11__280_203_29_l141__28_28_28_281__m64m (
  i_0r0d, i_0r1d, i_0a,
  o_0r, o_0a,
  o_1r, o_1a,
  o_2r, o_2a,
  initialise
);
  input [2:0] i_0r0d;
  input [2:0] i_0r1d;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  input initialise;
  wire icomplete_0n;
  wire sel_0n;
  wire sel_1n;
  wire sel_2n;
  wire matchi_0n;
  wire matchi_1n;
  wire matchi_2n;
  wire [2:0] ifint_0n;
  wire [2:0] itint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire ofint_1n;
  wire ofint_2n;
  wire oaint_0n;
  wire oaint_1n;
  wire oaint_2n;
  wire oack_0n;
  wire gate1037_0n;
  wire gate1034_0n;
  wire gate1031_0n;
  wire [2:0] complete1028_0n;
  wire gate1027_0n;
  wire [2:0] complete1024_0n;
  C2 I0 (iaint_0n, oack_0n, icomplete_0n);
  OR3 I1 (oack_0n, oaint_0n, oaint_1n, oaint_2n);
  assign oaint_2n = o_2r;
  INV I3 (gate1037_0n, o_2a);
  C2RI I4 (o_2r, ofint_2n, gate1037_0n, initialise);
  assign oaint_1n = o_1r;
  INV I6 (gate1034_0n, o_1a);
  C2RI I7 (o_1r, ofint_1n, gate1034_0n, initialise);
  assign oaint_0n = o_0r;
  INV I9 (gate1031_0n, o_0a);
  C2RI I10 (o_0r, ofint_0n, gate1031_0n, initialise);
  C3 I11 (i_0a, complete1028_0n[0], complete1028_0n[1], complete1028_0n[2]);
  OR2 I12 (complete1028_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I13 (complete1028_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I14 (complete1028_0n[2], ifint_0n[2], itint_0n[2]);
  INV I15 (gate1027_0n, iaint_0n);
  C2RI I16 (itint_0n[0], i_0r1d[0], gate1027_0n, initialise);
  C2RI I17 (itint_0n[1], i_0r1d[1], gate1027_0n, initialise);
  C2RI I18 (itint_0n[2], i_0r1d[2], gate1027_0n, initialise);
  C2RI I19 (ifint_0n[0], i_0r0d[0], gate1027_0n, initialise);
  C2RI I20 (ifint_0n[1], i_0r0d[1], gate1027_0n, initialise);
  C2RI I21 (ifint_0n[2], i_0r0d[2], gate1027_0n, initialise);
  assign ofint_2n = sel_2n;
  assign ofint_1n = sel_1n;
  assign ofint_0n = sel_0n;
  C3 I25 (icomplete_0n, complete1024_0n[0], complete1024_0n[1], complete1024_0n[2]);
  OR2 I26 (complete1024_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I27 (complete1024_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I28 (complete1024_0n[2], ifint_0n[2], itint_0n[2]);
  C3 I29 (matchi_2n, ifint_0n[1], ifint_0n[0], itint_0n[2]);
  assign sel_2n = matchi_2n;
  C3 I31 (matchi_1n, ifint_0n[2], ifint_0n[0], itint_0n[1]);
  assign sel_1n = matchi_1n;
  C3 I33 (matchi_0n, ifint_0n[2], ifint_0n[1], itint_0n[0]);
  assign sel_0n = matchi_0n;
endmodule

module BrzS_3_l11__280_203_29_l151__28_28_28_281__m65m (
  i_0r0d, i_0r1d, i_0a,
  o_0r, o_0a,
  o_1r, o_1a,
  initialise
);
  input [2:0] i_0r0d;
  input [2:0] i_0r1d;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input initialise;
  wire icomplete_0n;
  wire sel_0n;
  wire sel_1n;
  wire [2:0] matchi_0n;
  wire [2:0] matchi_1n;
  wire [2:0] ifint_0n;
  wire [2:0] itint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire ofint_1n;
  wire oaint_0n;
  wire oaint_1n;
  wire oack_0n;
  wire gate1048_0n;
  wire gate1045_0n;
  wire [2:0] complete1042_0n;
  wire gate1041_0n;
  wire [2:0] complete1038_0n;
  C2 I0 (iaint_0n, oack_0n, icomplete_0n);
  OR2 I1 (oack_0n, oaint_0n, oaint_1n);
  assign oaint_1n = o_1r;
  INV I3 (gate1048_0n, o_1a);
  C2RI I4 (o_1r, ofint_1n, gate1048_0n, initialise);
  assign oaint_0n = o_0r;
  INV I6 (gate1045_0n, o_0a);
  C2RI I7 (o_0r, ofint_0n, gate1045_0n, initialise);
  C3 I8 (i_0a, complete1042_0n[0], complete1042_0n[1], complete1042_0n[2]);
  OR2 I9 (complete1042_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I10 (complete1042_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I11 (complete1042_0n[2], ifint_0n[2], itint_0n[2]);
  INV I12 (gate1041_0n, iaint_0n);
  C2RI I13 (itint_0n[0], i_0r1d[0], gate1041_0n, initialise);
  C2RI I14 (itint_0n[1], i_0r1d[1], gate1041_0n, initialise);
  C2RI I15 (itint_0n[2], i_0r1d[2], gate1041_0n, initialise);
  C2RI I16 (ifint_0n[0], i_0r0d[0], gate1041_0n, initialise);
  C2RI I17 (ifint_0n[1], i_0r0d[1], gate1041_0n, initialise);
  C2RI I18 (ifint_0n[2], i_0r0d[2], gate1041_0n, initialise);
  assign ofint_1n = sel_1n;
  assign ofint_0n = sel_0n;
  C3 I21 (icomplete_0n, complete1038_0n[0], complete1038_0n[1], complete1038_0n[2]);
  OR2 I22 (complete1038_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I23 (complete1038_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I24 (complete1038_0n[2], ifint_0n[2], itint_0n[2]);
  C3 I25 (matchi_1n[2], ifint_0n[1], itint_0n[2], itint_0n[0]);
  C3 I26 (matchi_1n[1], ifint_0n[1], ifint_0n[0], itint_0n[2]);
  C3 I27 (matchi_1n[0], ifint_0n[2], ifint_0n[1], ifint_0n[0]);
  OR3 I28 (sel_1n, matchi_1n[0], matchi_1n[1], matchi_1n[2]);
  C2 I29 (matchi_0n[2], itint_0n[1], itint_0n[0]);
  C2 I30 (matchi_0n[1], ifint_0n[0], itint_0n[1]);
  C3 I31 (matchi_0n[0], ifint_0n[2], ifint_0n[1], itint_0n[0]);
  OR3 I32 (sel_0n, matchi_0n[0], matchi_0n[1], matchi_0n[2]);
endmodule

module BrzS_4_l11__280_204_29_l521__28_28_28_280__m66m (
  i_0r0d, i_0r1d, i_0a,
  o_0r, o_0a,
  o_1r, o_1a,
  o_2r, o_2a,
  o_3r, o_3a,
  o_4r, o_4a,
  o_5r, o_5a,
  o_6r, o_6a,
  o_7r, o_7a,
  o_8r, o_8a,
  initialise
);
  input [3:0] i_0r0d;
  input [3:0] i_0r1d;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  output o_7r;
  input o_7a;
  output o_8r;
  input o_8a;
  input initialise;
  wire [38:0] internal_0n;
  wire icomplete_0n;
  wire sel_0n;
  wire sel_1n;
  wire sel_2n;
  wire sel_3n;
  wire sel_4n;
  wire sel_5n;
  wire sel_6n;
  wire sel_7n;
  wire sel_8n;
  wire [1:0] matchi_0n;
  wire [1:0] matchi_1n;
  wire [1:0] matchi_2n;
  wire [1:0] matchi_3n;
  wire matchi_4n;
  wire matchi_5n;
  wire [1:0] matchi_6n;
  wire [1:0] matchi_7n;
  wire [1:0] matchi_8n;
  wire [3:0] ifint_0n;
  wire [3:0] itint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire ofint_1n;
  wire ofint_2n;
  wire ofint_3n;
  wire ofint_4n;
  wire ofint_5n;
  wire ofint_6n;
  wire ofint_7n;
  wire ofint_8n;
  wire oaint_0n;
  wire oaint_1n;
  wire oaint_2n;
  wire oaint_3n;
  wire oaint_4n;
  wire oaint_5n;
  wire oaint_6n;
  wire oaint_7n;
  wire oaint_8n;
  wire oack_0n;
  wire gate1080_0n;
  wire gate1077_0n;
  wire gate1074_0n;
  wire gate1071_0n;
  wire gate1068_0n;
  wire gate1065_0n;
  wire gate1062_0n;
  wire gate1059_0n;
  wire gate1056_0n;
  wire [3:0] complete1053_0n;
  wire gate1052_0n;
  wire [3:0] complete1049_0n;
  C2 I0 (iaint_0n, oack_0n, icomplete_0n);
  NOR3 I1 (internal_0n[0], oaint_0n, oaint_1n, oaint_2n);
  NOR3 I2 (internal_0n[1], oaint_3n, oaint_4n, oaint_5n);
  NOR3 I3 (internal_0n[2], oaint_6n, oaint_7n, oaint_8n);
  NAND3 I4 (oack_0n, internal_0n[0], internal_0n[1], internal_0n[2]);
  assign oaint_8n = o_8r;
  INV I6 (gate1080_0n, o_8a);
  C2RI I7 (o_8r, ofint_8n, gate1080_0n, initialise);
  assign oaint_7n = o_7r;
  INV I9 (gate1077_0n, o_7a);
  C2RI I10 (o_7r, ofint_7n, gate1077_0n, initialise);
  assign oaint_6n = o_6r;
  INV I12 (gate1074_0n, o_6a);
  C2RI I13 (o_6r, ofint_6n, gate1074_0n, initialise);
  assign oaint_5n = o_5r;
  INV I15 (gate1071_0n, o_5a);
  C2RI I16 (o_5r, ofint_5n, gate1071_0n, initialise);
  assign oaint_4n = o_4r;
  INV I18 (gate1068_0n, o_4a);
  C2RI I19 (o_4r, ofint_4n, gate1068_0n, initialise);
  assign oaint_3n = o_3r;
  INV I21 (gate1065_0n, o_3a);
  C2RI I22 (o_3r, ofint_3n, gate1065_0n, initialise);
  assign oaint_2n = o_2r;
  INV I24 (gate1062_0n, o_2a);
  C2RI I25 (o_2r, ofint_2n, gate1062_0n, initialise);
  assign oaint_1n = o_1r;
  INV I27 (gate1059_0n, o_1a);
  C2RI I28 (o_1r, ofint_1n, gate1059_0n, initialise);
  assign oaint_0n = o_0r;
  INV I30 (gate1056_0n, o_0a);
  C2RI I31 (o_0r, ofint_0n, gate1056_0n, initialise);
  C2 I32 (internal_0n[3], complete1053_0n[0], complete1053_0n[1]);
  C2 I33 (internal_0n[4], complete1053_0n[2], complete1053_0n[3]);
  C2 I34 (i_0a, internal_0n[3], internal_0n[4]);
  OR2 I35 (complete1053_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I36 (complete1053_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I37 (complete1053_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I38 (complete1053_0n[3], ifint_0n[3], itint_0n[3]);
  INV I39 (gate1052_0n, iaint_0n);
  C2RI I40 (itint_0n[0], i_0r1d[0], gate1052_0n, initialise);
  C2RI I41 (itint_0n[1], i_0r1d[1], gate1052_0n, initialise);
  C2RI I42 (itint_0n[2], i_0r1d[2], gate1052_0n, initialise);
  C2RI I43 (itint_0n[3], i_0r1d[3], gate1052_0n, initialise);
  C2RI I44 (ifint_0n[0], i_0r0d[0], gate1052_0n, initialise);
  C2RI I45 (ifint_0n[1], i_0r0d[1], gate1052_0n, initialise);
  C2RI I46 (ifint_0n[2], i_0r0d[2], gate1052_0n, initialise);
  C2RI I47 (ifint_0n[3], i_0r0d[3], gate1052_0n, initialise);
  assign ofint_8n = sel_8n;
  assign ofint_7n = sel_7n;
  assign ofint_6n = sel_6n;
  assign ofint_5n = sel_5n;
  assign ofint_4n = sel_4n;
  assign ofint_3n = sel_3n;
  assign ofint_2n = sel_2n;
  assign ofint_1n = sel_1n;
  assign ofint_0n = sel_0n;
  C2 I57 (internal_0n[5], complete1049_0n[0], complete1049_0n[1]);
  C2 I58 (internal_0n[6], complete1049_0n[2], complete1049_0n[3]);
  C2 I59 (icomplete_0n, internal_0n[5], internal_0n[6]);
  OR2 I60 (complete1049_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I61 (complete1049_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I62 (complete1049_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I63 (complete1049_0n[3], ifint_0n[3], itint_0n[3]);
  C2 I64 (internal_0n[7], ifint_0n[0], itint_0n[3]);
  C2 I65 (internal_0n[8], itint_0n[2], itint_0n[1]);
  C2 I66 (matchi_8n[1], internal_0n[7], internal_0n[8]);
  C2 I67 (internal_0n[9], ifint_0n[1], itint_0n[3]);
  C2 I68 (internal_0n[10], itint_0n[2], itint_0n[0]);
  C2 I69 (matchi_8n[0], internal_0n[9], internal_0n[10]);
  OR2 I70 (sel_8n, matchi_8n[0], matchi_8n[1]);
  C2 I71 (internal_0n[11], ifint_0n[1], ifint_0n[0]);
  C2 I72 (internal_0n[12], itint_0n[3], itint_0n[2]);
  C2 I73 (matchi_7n[1], internal_0n[11], internal_0n[12]);
  C2 I74 (internal_0n[13], ifint_0n[2], itint_0n[3]);
  C2 I75 (internal_0n[14], itint_0n[1], itint_0n[0]);
  C2 I76 (matchi_7n[0], internal_0n[13], internal_0n[14]);
  OR2 I77 (sel_7n, matchi_7n[0], matchi_7n[1]);
  C2 I78 (internal_0n[15], ifint_0n[2], ifint_0n[0]);
  C2 I79 (internal_0n[16], itint_0n[3], itint_0n[1]);
  C2 I80 (matchi_6n[1], internal_0n[15], internal_0n[16]);
  C2 I81 (internal_0n[17], ifint_0n[2], ifint_0n[1]);
  C2 I82 (internal_0n[18], itint_0n[3], itint_0n[0]);
  C2 I83 (matchi_6n[0], internal_0n[17], internal_0n[18]);
  OR2 I84 (sel_6n, matchi_6n[0], matchi_6n[1]);
  C2 I85 (internal_0n[19], ifint_0n[2], ifint_0n[1]);
  C2 I86 (internal_0n[20], ifint_0n[0], itint_0n[3]);
  C2 I87 (matchi_5n, internal_0n[19], internal_0n[20]);
  assign sel_5n = matchi_5n;
  C2 I89 (internal_0n[21], ifint_0n[3], itint_0n[2]);
  C2 I90 (internal_0n[22], itint_0n[1], itint_0n[0]);
  C2 I91 (matchi_4n, internal_0n[21], internal_0n[22]);
  assign sel_4n = matchi_4n;
  C2 I93 (internal_0n[23], ifint_0n[3], ifint_0n[0]);
  C2 I94 (internal_0n[24], itint_0n[2], itint_0n[1]);
  C2 I95 (matchi_3n[1], internal_0n[23], internal_0n[24]);
  C2 I96 (internal_0n[25], ifint_0n[3], ifint_0n[1]);
  C2 I97 (internal_0n[26], itint_0n[2], itint_0n[0]);
  C2 I98 (matchi_3n[0], internal_0n[25], internal_0n[26]);
  OR2 I99 (sel_3n, matchi_3n[0], matchi_3n[1]);
  C2 I100 (internal_0n[27], ifint_0n[3], ifint_0n[1]);
  C2 I101 (internal_0n[28], ifint_0n[0], itint_0n[2]);
  C2 I102 (matchi_2n[1], internal_0n[27], internal_0n[28]);
  C2 I103 (internal_0n[29], ifint_0n[3], ifint_0n[2]);
  C2 I104 (internal_0n[30], itint_0n[1], itint_0n[0]);
  C2 I105 (matchi_2n[0], internal_0n[29], internal_0n[30]);
  OR2 I106 (sel_2n, matchi_2n[0], matchi_2n[1]);
  C2 I107 (internal_0n[31], ifint_0n[3], ifint_0n[2]);
  C2 I108 (internal_0n[32], ifint_0n[0], itint_0n[1]);
  C2 I109 (matchi_1n[1], internal_0n[31], internal_0n[32]);
  C2 I110 (internal_0n[33], ifint_0n[3], ifint_0n[2]);
  C2 I111 (internal_0n[34], ifint_0n[1], itint_0n[0]);
  C2 I112 (matchi_1n[0], internal_0n[33], internal_0n[34]);
  OR2 I113 (sel_1n, matchi_1n[0], matchi_1n[1]);
  C2 I114 (internal_0n[35], itint_0n[3], itint_0n[2]);
  C2 I115 (internal_0n[36], itint_0n[1], itint_0n[0]);
  C2 I116 (matchi_0n[1], internal_0n[35], internal_0n[36]);
  C2 I117 (internal_0n[37], ifint_0n[3], ifint_0n[2]);
  C2 I118 (internal_0n[38], ifint_0n[1], ifint_0n[0]);
  C2 I119 (matchi_0n[0], internal_0n[37], internal_0n[38]);
  OR2 I120 (sel_0n, matchi_0n[0], matchi_0n[1]);
endmodule

module BrzS_4_l11__281_203_29_l141__28_28_28_281__m67m (
  i_0r0d, i_0r1d, i_0a,
  o_0r0d, o_0r1d, o_0a,
  o_1r0d, o_1r1d, o_1a,
  o_2r0d, o_2r1d, o_2a,
  initialise
);
  input [3:0] i_0r0d;
  input [3:0] i_0r1d;
  output i_0a;
  output o_0r0d;
  output o_0r1d;
  input o_0a;
  output o_1r0d;
  output o_1r1d;
  input o_1a;
  output o_2r0d;
  output o_2r1d;
  input o_2a;
  input initialise;
  wire [3:0] internal_0n;
  wire icomplete_0n;
  wire sel_0n;
  wire sel_1n;
  wire sel_2n;
  wire matchi_0n;
  wire matchi_1n;
  wire matchi_2n;
  wire [3:0] ifint_0n;
  wire [3:0] itint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire ofint_1n;
  wire ofint_2n;
  wire otint_0n;
  wire otint_1n;
  wire otint_2n;
  wire oaint_0n;
  wire oaint_1n;
  wire oaint_2n;
  wire oack_0n;
  wire complete1097_0n;
  wire gate1096_0n;
  wire complete1093_0n;
  wire gate1092_0n;
  wire complete1089_0n;
  wire gate1088_0n;
  wire [3:0] complete1085_0n;
  wire gate1084_0n;
  wire [3:0] complete1081_0n;
  C2 I0 (iaint_0n, oack_0n, icomplete_0n);
  OR3 I1 (oack_0n, oaint_0n, oaint_1n, oaint_2n);
  assign oaint_2n = complete1097_0n;
  OR2 I3 (complete1097_0n, o_2r0d, o_2r1d);
  INV I4 (gate1096_0n, o_2a);
  C2RI I5 (o_2r1d, otint_2n, gate1096_0n, initialise);
  C2RI I6 (o_2r0d, ofint_2n, gate1096_0n, initialise);
  assign oaint_1n = complete1093_0n;
  OR2 I8 (complete1093_0n, o_1r0d, o_1r1d);
  INV I9 (gate1092_0n, o_1a);
  C2RI I10 (o_1r1d, otint_1n, gate1092_0n, initialise);
  C2RI I11 (o_1r0d, ofint_1n, gate1092_0n, initialise);
  assign oaint_0n = complete1089_0n;
  OR2 I13 (complete1089_0n, o_0r0d, o_0r1d);
  INV I14 (gate1088_0n, o_0a);
  C2RI I15 (o_0r1d, otint_0n, gate1088_0n, initialise);
  C2RI I16 (o_0r0d, ofint_0n, gate1088_0n, initialise);
  C2 I17 (internal_0n[0], complete1085_0n[0], complete1085_0n[1]);
  C2 I18 (internal_0n[1], complete1085_0n[2], complete1085_0n[3]);
  C2 I19 (i_0a, internal_0n[0], internal_0n[1]);
  OR2 I20 (complete1085_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I21 (complete1085_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I22 (complete1085_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I23 (complete1085_0n[3], ifint_0n[3], itint_0n[3]);
  INV I24 (gate1084_0n, iaint_0n);
  C2RI I25 (itint_0n[0], i_0r1d[0], gate1084_0n, initialise);
  C2RI I26 (itint_0n[1], i_0r1d[1], gate1084_0n, initialise);
  C2RI I27 (itint_0n[2], i_0r1d[2], gate1084_0n, initialise);
  C2RI I28 (itint_0n[3], i_0r1d[3], gate1084_0n, initialise);
  C2RI I29 (ifint_0n[0], i_0r0d[0], gate1084_0n, initialise);
  C2RI I30 (ifint_0n[1], i_0r0d[1], gate1084_0n, initialise);
  C2RI I31 (ifint_0n[2], i_0r0d[2], gate1084_0n, initialise);
  C2RI I32 (ifint_0n[3], i_0r0d[3], gate1084_0n, initialise);
  C2 I33 (otint_2n, sel_2n, itint_0n[0]);
  C2 I34 (otint_1n, sel_1n, itint_0n[0]);
  C2 I35 (otint_0n, sel_0n, itint_0n[0]);
  C2 I36 (ofint_2n, sel_2n, ifint_0n[0]);
  C2 I37 (ofint_1n, sel_1n, ifint_0n[0]);
  C2 I38 (ofint_0n, sel_0n, ifint_0n[0]);
  C2 I39 (internal_0n[2], complete1081_0n[0], complete1081_0n[1]);
  C2 I40 (internal_0n[3], complete1081_0n[2], complete1081_0n[3]);
  C2 I41 (icomplete_0n, internal_0n[2], internal_0n[3]);
  OR2 I42 (complete1081_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I43 (complete1081_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I44 (complete1081_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I45 (complete1081_0n[3], ifint_0n[3], itint_0n[3]);
  C3 I46 (matchi_2n, ifint_0n[2], ifint_0n[1], itint_0n[3]);
  assign sel_2n = matchi_2n;
  C3 I48 (matchi_1n, ifint_0n[3], ifint_0n[1], itint_0n[2]);
  assign sel_1n = matchi_1n;
  C3 I50 (matchi_0n, ifint_0n[3], ifint_0n[2], itint_0n[1]);
  assign sel_0n = matchi_0n;
endmodule

module BrzS_9_l11__280_209_29_l424__28_28_28_281__m68m (
  i_0r0d, i_0r1d, i_0a,
  o_0r, o_0a,
  o_1r, o_1a,
  o_2r, o_2a,
  o_3r, o_3a,
  o_4r, o_4a,
  o_5r, o_5a,
  o_6r, o_6a,
  o_7r, o_7a,
  o_8r, o_8a,
  initialise
);
  input [8:0] i_0r0d;
  input [8:0] i_0r1d;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  output o_7r;
  input o_7a;
  output o_8r;
  input o_8a;
  input initialise;
  wire [35:0] internal_0n;
  wire icomplete_0n;
  wire sel_0n;
  wire sel_1n;
  wire sel_2n;
  wire sel_3n;
  wire sel_4n;
  wire sel_5n;
  wire sel_6n;
  wire sel_7n;
  wire sel_8n;
  wire matchi_0n;
  wire matchi_1n;
  wire matchi_2n;
  wire matchi_3n;
  wire matchi_4n;
  wire matchi_5n;
  wire matchi_6n;
  wire matchi_7n;
  wire matchi_8n;
  wire [8:0] ifint_0n;
  wire [8:0] itint_0n;
  wire iaint_0n;
  wire ofint_0n;
  wire ofint_1n;
  wire ofint_2n;
  wire ofint_3n;
  wire ofint_4n;
  wire ofint_5n;
  wire ofint_6n;
  wire ofint_7n;
  wire ofint_8n;
  wire oaint_0n;
  wire oaint_1n;
  wire oaint_2n;
  wire oaint_3n;
  wire oaint_4n;
  wire oaint_5n;
  wire oaint_6n;
  wire oaint_7n;
  wire oaint_8n;
  wire oack_0n;
  wire gate1129_0n;
  wire gate1126_0n;
  wire gate1123_0n;
  wire gate1120_0n;
  wire gate1117_0n;
  wire gate1114_0n;
  wire gate1111_0n;
  wire gate1108_0n;
  wire gate1105_0n;
  wire [8:0] complete1102_0n;
  wire gate1101_0n;
  wire [8:0] complete1098_0n;
  C2 I0 (iaint_0n, oack_0n, icomplete_0n);
  NOR3 I1 (internal_0n[0], oaint_0n, oaint_1n, oaint_2n);
  NOR3 I2 (internal_0n[1], oaint_3n, oaint_4n, oaint_5n);
  NOR3 I3 (internal_0n[2], oaint_6n, oaint_7n, oaint_8n);
  NAND3 I4 (oack_0n, internal_0n[0], internal_0n[1], internal_0n[2]);
  assign oaint_8n = o_8r;
  INV I6 (gate1129_0n, o_8a);
  C2RI I7 (o_8r, ofint_8n, gate1129_0n, initialise);
  assign oaint_7n = o_7r;
  INV I9 (gate1126_0n, o_7a);
  C2RI I10 (o_7r, ofint_7n, gate1126_0n, initialise);
  assign oaint_6n = o_6r;
  INV I12 (gate1123_0n, o_6a);
  C2RI I13 (o_6r, ofint_6n, gate1123_0n, initialise);
  assign oaint_5n = o_5r;
  INV I15 (gate1120_0n, o_5a);
  C2RI I16 (o_5r, ofint_5n, gate1120_0n, initialise);
  assign oaint_4n = o_4r;
  INV I18 (gate1117_0n, o_4a);
  C2RI I19 (o_4r, ofint_4n, gate1117_0n, initialise);
  assign oaint_3n = o_3r;
  INV I21 (gate1114_0n, o_3a);
  C2RI I22 (o_3r, ofint_3n, gate1114_0n, initialise);
  assign oaint_2n = o_2r;
  INV I24 (gate1111_0n, o_2a);
  C2RI I25 (o_2r, ofint_2n, gate1111_0n, initialise);
  assign oaint_1n = o_1r;
  INV I27 (gate1108_0n, o_1a);
  C2RI I28 (o_1r, ofint_1n, gate1108_0n, initialise);
  assign oaint_0n = o_0r;
  INV I30 (gate1105_0n, o_0a);
  C2RI I31 (o_0r, ofint_0n, gate1105_0n, initialise);
  C3 I32 (internal_0n[3], complete1102_0n[0], complete1102_0n[1], complete1102_0n[2]);
  C3 I33 (internal_0n[4], complete1102_0n[3], complete1102_0n[4], complete1102_0n[5]);
  C3 I34 (internal_0n[5], complete1102_0n[6], complete1102_0n[7], complete1102_0n[8]);
  C3 I35 (i_0a, internal_0n[3], internal_0n[4], internal_0n[5]);
  OR2 I36 (complete1102_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I37 (complete1102_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I38 (complete1102_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I39 (complete1102_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I40 (complete1102_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I41 (complete1102_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I42 (complete1102_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I43 (complete1102_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I44 (complete1102_0n[8], ifint_0n[8], itint_0n[8]);
  INV I45 (gate1101_0n, iaint_0n);
  C2RI I46 (itint_0n[0], i_0r1d[0], gate1101_0n, initialise);
  C2RI I47 (itint_0n[1], i_0r1d[1], gate1101_0n, initialise);
  C2RI I48 (itint_0n[2], i_0r1d[2], gate1101_0n, initialise);
  C2RI I49 (itint_0n[3], i_0r1d[3], gate1101_0n, initialise);
  C2RI I50 (itint_0n[4], i_0r1d[4], gate1101_0n, initialise);
  C2RI I51 (itint_0n[5], i_0r1d[5], gate1101_0n, initialise);
  C2RI I52 (itint_0n[6], i_0r1d[6], gate1101_0n, initialise);
  C2RI I53 (itint_0n[7], i_0r1d[7], gate1101_0n, initialise);
  C2RI I54 (itint_0n[8], i_0r1d[8], gate1101_0n, initialise);
  C2RI I55 (ifint_0n[0], i_0r0d[0], gate1101_0n, initialise);
  C2RI I56 (ifint_0n[1], i_0r0d[1], gate1101_0n, initialise);
  C2RI I57 (ifint_0n[2], i_0r0d[2], gate1101_0n, initialise);
  C2RI I58 (ifint_0n[3], i_0r0d[3], gate1101_0n, initialise);
  C2RI I59 (ifint_0n[4], i_0r0d[4], gate1101_0n, initialise);
  C2RI I60 (ifint_0n[5], i_0r0d[5], gate1101_0n, initialise);
  C2RI I61 (ifint_0n[6], i_0r0d[6], gate1101_0n, initialise);
  C2RI I62 (ifint_0n[7], i_0r0d[7], gate1101_0n, initialise);
  C2RI I63 (ifint_0n[8], i_0r0d[8], gate1101_0n, initialise);
  assign ofint_8n = sel_8n;
  assign ofint_7n = sel_7n;
  assign ofint_6n = sel_6n;
  assign ofint_5n = sel_5n;
  assign ofint_4n = sel_4n;
  assign ofint_3n = sel_3n;
  assign ofint_2n = sel_2n;
  assign ofint_1n = sel_1n;
  assign ofint_0n = sel_0n;
  C3 I73 (internal_0n[6], complete1098_0n[0], complete1098_0n[1], complete1098_0n[2]);
  C3 I74 (internal_0n[7], complete1098_0n[3], complete1098_0n[4], complete1098_0n[5]);
  C3 I75 (internal_0n[8], complete1098_0n[6], complete1098_0n[7], complete1098_0n[8]);
  C3 I76 (icomplete_0n, internal_0n[6], internal_0n[7], internal_0n[8]);
  OR2 I77 (complete1098_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I78 (complete1098_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I79 (complete1098_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I80 (complete1098_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I81 (complete1098_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I82 (complete1098_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I83 (complete1098_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I84 (complete1098_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I85 (complete1098_0n[8], ifint_0n[8], itint_0n[8]);
  C3 I86 (internal_0n[9], ifint_0n[7], ifint_0n[6], ifint_0n[5]);
  C3 I87 (internal_0n[10], ifint_0n[4], ifint_0n[3], ifint_0n[2]);
  C3 I88 (internal_0n[11], ifint_0n[1], ifint_0n[0], itint_0n[8]);
  C3 I89 (matchi_8n, internal_0n[9], internal_0n[10], internal_0n[11]);
  assign sel_8n = matchi_8n;
  C3 I91 (internal_0n[12], ifint_0n[8], ifint_0n[6], ifint_0n[5]);
  C3 I92 (internal_0n[13], ifint_0n[4], ifint_0n[3], ifint_0n[2]);
  C3 I93 (internal_0n[14], ifint_0n[1], ifint_0n[0], itint_0n[7]);
  C3 I94 (matchi_7n, internal_0n[12], internal_0n[13], internal_0n[14]);
  assign sel_7n = matchi_7n;
  C3 I96 (internal_0n[15], ifint_0n[8], ifint_0n[7], ifint_0n[5]);
  C3 I97 (internal_0n[16], ifint_0n[4], ifint_0n[3], ifint_0n[2]);
  C3 I98 (internal_0n[17], ifint_0n[1], ifint_0n[0], itint_0n[6]);
  C3 I99 (matchi_6n, internal_0n[15], internal_0n[16], internal_0n[17]);
  assign sel_6n = matchi_6n;
  C3 I101 (internal_0n[18], ifint_0n[8], ifint_0n[7], ifint_0n[6]);
  C3 I102 (internal_0n[19], ifint_0n[4], ifint_0n[3], ifint_0n[2]);
  C3 I103 (internal_0n[20], ifint_0n[1], ifint_0n[0], itint_0n[5]);
  C3 I104 (matchi_5n, internal_0n[18], internal_0n[19], internal_0n[20]);
  assign sel_5n = matchi_5n;
  C3 I106 (internal_0n[21], ifint_0n[8], ifint_0n[7], ifint_0n[6]);
  C3 I107 (internal_0n[22], ifint_0n[5], ifint_0n[3], ifint_0n[2]);
  C3 I108 (internal_0n[23], ifint_0n[1], ifint_0n[0], itint_0n[4]);
  C3 I109 (matchi_4n, internal_0n[21], internal_0n[22], internal_0n[23]);
  assign sel_4n = matchi_4n;
  C3 I111 (internal_0n[24], ifint_0n[8], ifint_0n[7], ifint_0n[6]);
  C3 I112 (internal_0n[25], ifint_0n[5], ifint_0n[4], ifint_0n[2]);
  C3 I113 (internal_0n[26], ifint_0n[1], ifint_0n[0], itint_0n[3]);
  C3 I114 (matchi_3n, internal_0n[24], internal_0n[25], internal_0n[26]);
  assign sel_3n = matchi_3n;
  C3 I116 (internal_0n[27], ifint_0n[8], ifint_0n[7], ifint_0n[6]);
  C3 I117 (internal_0n[28], ifint_0n[5], ifint_0n[4], ifint_0n[3]);
  C3 I118 (internal_0n[29], ifint_0n[1], ifint_0n[0], itint_0n[2]);
  C3 I119 (matchi_2n, internal_0n[27], internal_0n[28], internal_0n[29]);
  assign sel_2n = matchi_2n;
  C3 I121 (internal_0n[30], ifint_0n[8], ifint_0n[7], ifint_0n[6]);
  C3 I122 (internal_0n[31], ifint_0n[5], ifint_0n[4], ifint_0n[3]);
  C3 I123 (internal_0n[32], ifint_0n[2], ifint_0n[0], itint_0n[1]);
  C3 I124 (matchi_1n, internal_0n[30], internal_0n[31], internal_0n[32]);
  assign sel_1n = matchi_1n;
  C3 I126 (internal_0n[33], ifint_0n[8], ifint_0n[7], ifint_0n[6]);
  C3 I127 (internal_0n[34], ifint_0n[5], ifint_0n[4], ifint_0n[3]);
  C3 I128 (internal_0n[35], ifint_0n[2], ifint_0n[1], itint_0n[0]);
  C3 I129 (matchi_0n, internal_0n[33], internal_0n[34], internal_0n[35]);
  assign sel_0n = matchi_0n;
endmodule

module BrzS_34_l12__2832_202_29_l97__28_28_28_281_m69m (
  i_0r0d, i_0r1d, i_0a,
  o_0r0d, o_0r1d, o_0a,
  o_1r0d, o_1r1d, o_1a,
  initialise
);
  input [33:0] i_0r0d;
  input [33:0] i_0r1d;
  output i_0a;
  output [31:0] o_0r0d;
  output [31:0] o_0r1d;
  input o_0a;
  output [31:0] o_1r0d;
  output [31:0] o_1r1d;
  input o_1a;
  input initialise;
  wire [69:0] internal_0n;
  wire icomplete_0n;
  wire sel_0n;
  wire sel_1n;
  wire matchi_0n;
  wire matchi_1n;
  wire [33:0] ifint_0n;
  wire [33:0] itint_0n;
  wire iaint_0n;
  wire [31:0] ofint_0n;
  wire [31:0] ofint_1n;
  wire [31:0] otint_0n;
  wire [31:0] otint_1n;
  wire oaint_0n;
  wire oaint_1n;
  wire oack_0n;
  wire [31:0] complete1142_0n;
  wire gate1141_0n;
  wire [31:0] complete1138_0n;
  wire gate1137_0n;
  wire [33:0] complete1134_0n;
  wire gate1133_0n;
  wire [33:0] complete1130_0n;
  C2 I0 (iaint_0n, oack_0n, icomplete_0n);
  OR2 I1 (oack_0n, oaint_0n, oaint_1n);
  C3 I2 (internal_0n[0], complete1142_0n[0], complete1142_0n[1], complete1142_0n[2]);
  C3 I3 (internal_0n[1], complete1142_0n[3], complete1142_0n[4], complete1142_0n[5]);
  C3 I4 (internal_0n[2], complete1142_0n[6], complete1142_0n[7], complete1142_0n[8]);
  C3 I5 (internal_0n[3], complete1142_0n[9], complete1142_0n[10], complete1142_0n[11]);
  C3 I6 (internal_0n[4], complete1142_0n[12], complete1142_0n[13], complete1142_0n[14]);
  C3 I7 (internal_0n[5], complete1142_0n[15], complete1142_0n[16], complete1142_0n[17]);
  C3 I8 (internal_0n[6], complete1142_0n[18], complete1142_0n[19], complete1142_0n[20]);
  C3 I9 (internal_0n[7], complete1142_0n[21], complete1142_0n[22], complete1142_0n[23]);
  C3 I10 (internal_0n[8], complete1142_0n[24], complete1142_0n[25], complete1142_0n[26]);
  C3 I11 (internal_0n[9], complete1142_0n[27], complete1142_0n[28], complete1142_0n[29]);
  C2 I12 (internal_0n[10], complete1142_0n[30], complete1142_0n[31]);
  C3 I13 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I14 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I15 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I16 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I17 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I18 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I19 (oaint_1n, internal_0n[15], internal_0n[16]);
  OR2 I20 (complete1142_0n[0], o_1r0d[0], o_1r1d[0]);
  OR2 I21 (complete1142_0n[1], o_1r0d[1], o_1r1d[1]);
  OR2 I22 (complete1142_0n[2], o_1r0d[2], o_1r1d[2]);
  OR2 I23 (complete1142_0n[3], o_1r0d[3], o_1r1d[3]);
  OR2 I24 (complete1142_0n[4], o_1r0d[4], o_1r1d[4]);
  OR2 I25 (complete1142_0n[5], o_1r0d[5], o_1r1d[5]);
  OR2 I26 (complete1142_0n[6], o_1r0d[6], o_1r1d[6]);
  OR2 I27 (complete1142_0n[7], o_1r0d[7], o_1r1d[7]);
  OR2 I28 (complete1142_0n[8], o_1r0d[8], o_1r1d[8]);
  OR2 I29 (complete1142_0n[9], o_1r0d[9], o_1r1d[9]);
  OR2 I30 (complete1142_0n[10], o_1r0d[10], o_1r1d[10]);
  OR2 I31 (complete1142_0n[11], o_1r0d[11], o_1r1d[11]);
  OR2 I32 (complete1142_0n[12], o_1r0d[12], o_1r1d[12]);
  OR2 I33 (complete1142_0n[13], o_1r0d[13], o_1r1d[13]);
  OR2 I34 (complete1142_0n[14], o_1r0d[14], o_1r1d[14]);
  OR2 I35 (complete1142_0n[15], o_1r0d[15], o_1r1d[15]);
  OR2 I36 (complete1142_0n[16], o_1r0d[16], o_1r1d[16]);
  OR2 I37 (complete1142_0n[17], o_1r0d[17], o_1r1d[17]);
  OR2 I38 (complete1142_0n[18], o_1r0d[18], o_1r1d[18]);
  OR2 I39 (complete1142_0n[19], o_1r0d[19], o_1r1d[19]);
  OR2 I40 (complete1142_0n[20], o_1r0d[20], o_1r1d[20]);
  OR2 I41 (complete1142_0n[21], o_1r0d[21], o_1r1d[21]);
  OR2 I42 (complete1142_0n[22], o_1r0d[22], o_1r1d[22]);
  OR2 I43 (complete1142_0n[23], o_1r0d[23], o_1r1d[23]);
  OR2 I44 (complete1142_0n[24], o_1r0d[24], o_1r1d[24]);
  OR2 I45 (complete1142_0n[25], o_1r0d[25], o_1r1d[25]);
  OR2 I46 (complete1142_0n[26], o_1r0d[26], o_1r1d[26]);
  OR2 I47 (complete1142_0n[27], o_1r0d[27], o_1r1d[27]);
  OR2 I48 (complete1142_0n[28], o_1r0d[28], o_1r1d[28]);
  OR2 I49 (complete1142_0n[29], o_1r0d[29], o_1r1d[29]);
  OR2 I50 (complete1142_0n[30], o_1r0d[30], o_1r1d[30]);
  OR2 I51 (complete1142_0n[31], o_1r0d[31], o_1r1d[31]);
  INV I52 (gate1141_0n, o_1a);
  C2RI I53 (o_1r1d[0], otint_1n[0], gate1141_0n, initialise);
  C2RI I54 (o_1r1d[1], otint_1n[1], gate1141_0n, initialise);
  C2RI I55 (o_1r1d[2], otint_1n[2], gate1141_0n, initialise);
  C2RI I56 (o_1r1d[3], otint_1n[3], gate1141_0n, initialise);
  C2RI I57 (o_1r1d[4], otint_1n[4], gate1141_0n, initialise);
  C2RI I58 (o_1r1d[5], otint_1n[5], gate1141_0n, initialise);
  C2RI I59 (o_1r1d[6], otint_1n[6], gate1141_0n, initialise);
  C2RI I60 (o_1r1d[7], otint_1n[7], gate1141_0n, initialise);
  C2RI I61 (o_1r1d[8], otint_1n[8], gate1141_0n, initialise);
  C2RI I62 (o_1r1d[9], otint_1n[9], gate1141_0n, initialise);
  C2RI I63 (o_1r1d[10], otint_1n[10], gate1141_0n, initialise);
  C2RI I64 (o_1r1d[11], otint_1n[11], gate1141_0n, initialise);
  C2RI I65 (o_1r1d[12], otint_1n[12], gate1141_0n, initialise);
  C2RI I66 (o_1r1d[13], otint_1n[13], gate1141_0n, initialise);
  C2RI I67 (o_1r1d[14], otint_1n[14], gate1141_0n, initialise);
  C2RI I68 (o_1r1d[15], otint_1n[15], gate1141_0n, initialise);
  C2RI I69 (o_1r1d[16], otint_1n[16], gate1141_0n, initialise);
  C2RI I70 (o_1r1d[17], otint_1n[17], gate1141_0n, initialise);
  C2RI I71 (o_1r1d[18], otint_1n[18], gate1141_0n, initialise);
  C2RI I72 (o_1r1d[19], otint_1n[19], gate1141_0n, initialise);
  C2RI I73 (o_1r1d[20], otint_1n[20], gate1141_0n, initialise);
  C2RI I74 (o_1r1d[21], otint_1n[21], gate1141_0n, initialise);
  C2RI I75 (o_1r1d[22], otint_1n[22], gate1141_0n, initialise);
  C2RI I76 (o_1r1d[23], otint_1n[23], gate1141_0n, initialise);
  C2RI I77 (o_1r1d[24], otint_1n[24], gate1141_0n, initialise);
  C2RI I78 (o_1r1d[25], otint_1n[25], gate1141_0n, initialise);
  C2RI I79 (o_1r1d[26], otint_1n[26], gate1141_0n, initialise);
  C2RI I80 (o_1r1d[27], otint_1n[27], gate1141_0n, initialise);
  C2RI I81 (o_1r1d[28], otint_1n[28], gate1141_0n, initialise);
  C2RI I82 (o_1r1d[29], otint_1n[29], gate1141_0n, initialise);
  C2RI I83 (o_1r1d[30], otint_1n[30], gate1141_0n, initialise);
  C2RI I84 (o_1r1d[31], otint_1n[31], gate1141_0n, initialise);
  C2RI I85 (o_1r0d[0], ofint_1n[0], gate1141_0n, initialise);
  C2RI I86 (o_1r0d[1], ofint_1n[1], gate1141_0n, initialise);
  C2RI I87 (o_1r0d[2], ofint_1n[2], gate1141_0n, initialise);
  C2RI I88 (o_1r0d[3], ofint_1n[3], gate1141_0n, initialise);
  C2RI I89 (o_1r0d[4], ofint_1n[4], gate1141_0n, initialise);
  C2RI I90 (o_1r0d[5], ofint_1n[5], gate1141_0n, initialise);
  C2RI I91 (o_1r0d[6], ofint_1n[6], gate1141_0n, initialise);
  C2RI I92 (o_1r0d[7], ofint_1n[7], gate1141_0n, initialise);
  C2RI I93 (o_1r0d[8], ofint_1n[8], gate1141_0n, initialise);
  C2RI I94 (o_1r0d[9], ofint_1n[9], gate1141_0n, initialise);
  C2RI I95 (o_1r0d[10], ofint_1n[10], gate1141_0n, initialise);
  C2RI I96 (o_1r0d[11], ofint_1n[11], gate1141_0n, initialise);
  C2RI I97 (o_1r0d[12], ofint_1n[12], gate1141_0n, initialise);
  C2RI I98 (o_1r0d[13], ofint_1n[13], gate1141_0n, initialise);
  C2RI I99 (o_1r0d[14], ofint_1n[14], gate1141_0n, initialise);
  C2RI I100 (o_1r0d[15], ofint_1n[15], gate1141_0n, initialise);
  C2RI I101 (o_1r0d[16], ofint_1n[16], gate1141_0n, initialise);
  C2RI I102 (o_1r0d[17], ofint_1n[17], gate1141_0n, initialise);
  C2RI I103 (o_1r0d[18], ofint_1n[18], gate1141_0n, initialise);
  C2RI I104 (o_1r0d[19], ofint_1n[19], gate1141_0n, initialise);
  C2RI I105 (o_1r0d[20], ofint_1n[20], gate1141_0n, initialise);
  C2RI I106 (o_1r0d[21], ofint_1n[21], gate1141_0n, initialise);
  C2RI I107 (o_1r0d[22], ofint_1n[22], gate1141_0n, initialise);
  C2RI I108 (o_1r0d[23], ofint_1n[23], gate1141_0n, initialise);
  C2RI I109 (o_1r0d[24], ofint_1n[24], gate1141_0n, initialise);
  C2RI I110 (o_1r0d[25], ofint_1n[25], gate1141_0n, initialise);
  C2RI I111 (o_1r0d[26], ofint_1n[26], gate1141_0n, initialise);
  C2RI I112 (o_1r0d[27], ofint_1n[27], gate1141_0n, initialise);
  C2RI I113 (o_1r0d[28], ofint_1n[28], gate1141_0n, initialise);
  C2RI I114 (o_1r0d[29], ofint_1n[29], gate1141_0n, initialise);
  C2RI I115 (o_1r0d[30], ofint_1n[30], gate1141_0n, initialise);
  C2RI I116 (o_1r0d[31], ofint_1n[31], gate1141_0n, initialise);
  C3 I117 (internal_0n[17], complete1138_0n[0], complete1138_0n[1], complete1138_0n[2]);
  C3 I118 (internal_0n[18], complete1138_0n[3], complete1138_0n[4], complete1138_0n[5]);
  C3 I119 (internal_0n[19], complete1138_0n[6], complete1138_0n[7], complete1138_0n[8]);
  C3 I120 (internal_0n[20], complete1138_0n[9], complete1138_0n[10], complete1138_0n[11]);
  C3 I121 (internal_0n[21], complete1138_0n[12], complete1138_0n[13], complete1138_0n[14]);
  C3 I122 (internal_0n[22], complete1138_0n[15], complete1138_0n[16], complete1138_0n[17]);
  C3 I123 (internal_0n[23], complete1138_0n[18], complete1138_0n[19], complete1138_0n[20]);
  C3 I124 (internal_0n[24], complete1138_0n[21], complete1138_0n[22], complete1138_0n[23]);
  C3 I125 (internal_0n[25], complete1138_0n[24], complete1138_0n[25], complete1138_0n[26]);
  C3 I126 (internal_0n[26], complete1138_0n[27], complete1138_0n[28], complete1138_0n[29]);
  C2 I127 (internal_0n[27], complete1138_0n[30], complete1138_0n[31]);
  C3 I128 (internal_0n[28], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I129 (internal_0n[29], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I130 (internal_0n[30], internal_0n[23], internal_0n[24], internal_0n[25]);
  C2 I131 (internal_0n[31], internal_0n[26], internal_0n[27]);
  C2 I132 (internal_0n[32], internal_0n[28], internal_0n[29]);
  C2 I133 (internal_0n[33], internal_0n[30], internal_0n[31]);
  C2 I134 (oaint_0n, internal_0n[32], internal_0n[33]);
  OR2 I135 (complete1138_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I136 (complete1138_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I137 (complete1138_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I138 (complete1138_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I139 (complete1138_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I140 (complete1138_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I141 (complete1138_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I142 (complete1138_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I143 (complete1138_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I144 (complete1138_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I145 (complete1138_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I146 (complete1138_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I147 (complete1138_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I148 (complete1138_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I149 (complete1138_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I150 (complete1138_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I151 (complete1138_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I152 (complete1138_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I153 (complete1138_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I154 (complete1138_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I155 (complete1138_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I156 (complete1138_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I157 (complete1138_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I158 (complete1138_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I159 (complete1138_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I160 (complete1138_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I161 (complete1138_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I162 (complete1138_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I163 (complete1138_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I164 (complete1138_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I165 (complete1138_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I166 (complete1138_0n[31], o_0r0d[31], o_0r1d[31]);
  INV I167 (gate1137_0n, o_0a);
  C2RI I168 (o_0r1d[0], otint_0n[0], gate1137_0n, initialise);
  C2RI I169 (o_0r1d[1], otint_0n[1], gate1137_0n, initialise);
  C2RI I170 (o_0r1d[2], otint_0n[2], gate1137_0n, initialise);
  C2RI I171 (o_0r1d[3], otint_0n[3], gate1137_0n, initialise);
  C2RI I172 (o_0r1d[4], otint_0n[4], gate1137_0n, initialise);
  C2RI I173 (o_0r1d[5], otint_0n[5], gate1137_0n, initialise);
  C2RI I174 (o_0r1d[6], otint_0n[6], gate1137_0n, initialise);
  C2RI I175 (o_0r1d[7], otint_0n[7], gate1137_0n, initialise);
  C2RI I176 (o_0r1d[8], otint_0n[8], gate1137_0n, initialise);
  C2RI I177 (o_0r1d[9], otint_0n[9], gate1137_0n, initialise);
  C2RI I178 (o_0r1d[10], otint_0n[10], gate1137_0n, initialise);
  C2RI I179 (o_0r1d[11], otint_0n[11], gate1137_0n, initialise);
  C2RI I180 (o_0r1d[12], otint_0n[12], gate1137_0n, initialise);
  C2RI I181 (o_0r1d[13], otint_0n[13], gate1137_0n, initialise);
  C2RI I182 (o_0r1d[14], otint_0n[14], gate1137_0n, initialise);
  C2RI I183 (o_0r1d[15], otint_0n[15], gate1137_0n, initialise);
  C2RI I184 (o_0r1d[16], otint_0n[16], gate1137_0n, initialise);
  C2RI I185 (o_0r1d[17], otint_0n[17], gate1137_0n, initialise);
  C2RI I186 (o_0r1d[18], otint_0n[18], gate1137_0n, initialise);
  C2RI I187 (o_0r1d[19], otint_0n[19], gate1137_0n, initialise);
  C2RI I188 (o_0r1d[20], otint_0n[20], gate1137_0n, initialise);
  C2RI I189 (o_0r1d[21], otint_0n[21], gate1137_0n, initialise);
  C2RI I190 (o_0r1d[22], otint_0n[22], gate1137_0n, initialise);
  C2RI I191 (o_0r1d[23], otint_0n[23], gate1137_0n, initialise);
  C2RI I192 (o_0r1d[24], otint_0n[24], gate1137_0n, initialise);
  C2RI I193 (o_0r1d[25], otint_0n[25], gate1137_0n, initialise);
  C2RI I194 (o_0r1d[26], otint_0n[26], gate1137_0n, initialise);
  C2RI I195 (o_0r1d[27], otint_0n[27], gate1137_0n, initialise);
  C2RI I196 (o_0r1d[28], otint_0n[28], gate1137_0n, initialise);
  C2RI I197 (o_0r1d[29], otint_0n[29], gate1137_0n, initialise);
  C2RI I198 (o_0r1d[30], otint_0n[30], gate1137_0n, initialise);
  C2RI I199 (o_0r1d[31], otint_0n[31], gate1137_0n, initialise);
  C2RI I200 (o_0r0d[0], ofint_0n[0], gate1137_0n, initialise);
  C2RI I201 (o_0r0d[1], ofint_0n[1], gate1137_0n, initialise);
  C2RI I202 (o_0r0d[2], ofint_0n[2], gate1137_0n, initialise);
  C2RI I203 (o_0r0d[3], ofint_0n[3], gate1137_0n, initialise);
  C2RI I204 (o_0r0d[4], ofint_0n[4], gate1137_0n, initialise);
  C2RI I205 (o_0r0d[5], ofint_0n[5], gate1137_0n, initialise);
  C2RI I206 (o_0r0d[6], ofint_0n[6], gate1137_0n, initialise);
  C2RI I207 (o_0r0d[7], ofint_0n[7], gate1137_0n, initialise);
  C2RI I208 (o_0r0d[8], ofint_0n[8], gate1137_0n, initialise);
  C2RI I209 (o_0r0d[9], ofint_0n[9], gate1137_0n, initialise);
  C2RI I210 (o_0r0d[10], ofint_0n[10], gate1137_0n, initialise);
  C2RI I211 (o_0r0d[11], ofint_0n[11], gate1137_0n, initialise);
  C2RI I212 (o_0r0d[12], ofint_0n[12], gate1137_0n, initialise);
  C2RI I213 (o_0r0d[13], ofint_0n[13], gate1137_0n, initialise);
  C2RI I214 (o_0r0d[14], ofint_0n[14], gate1137_0n, initialise);
  C2RI I215 (o_0r0d[15], ofint_0n[15], gate1137_0n, initialise);
  C2RI I216 (o_0r0d[16], ofint_0n[16], gate1137_0n, initialise);
  C2RI I217 (o_0r0d[17], ofint_0n[17], gate1137_0n, initialise);
  C2RI I218 (o_0r0d[18], ofint_0n[18], gate1137_0n, initialise);
  C2RI I219 (o_0r0d[19], ofint_0n[19], gate1137_0n, initialise);
  C2RI I220 (o_0r0d[20], ofint_0n[20], gate1137_0n, initialise);
  C2RI I221 (o_0r0d[21], ofint_0n[21], gate1137_0n, initialise);
  C2RI I222 (o_0r0d[22], ofint_0n[22], gate1137_0n, initialise);
  C2RI I223 (o_0r0d[23], ofint_0n[23], gate1137_0n, initialise);
  C2RI I224 (o_0r0d[24], ofint_0n[24], gate1137_0n, initialise);
  C2RI I225 (o_0r0d[25], ofint_0n[25], gate1137_0n, initialise);
  C2RI I226 (o_0r0d[26], ofint_0n[26], gate1137_0n, initialise);
  C2RI I227 (o_0r0d[27], ofint_0n[27], gate1137_0n, initialise);
  C2RI I228 (o_0r0d[28], ofint_0n[28], gate1137_0n, initialise);
  C2RI I229 (o_0r0d[29], ofint_0n[29], gate1137_0n, initialise);
  C2RI I230 (o_0r0d[30], ofint_0n[30], gate1137_0n, initialise);
  C2RI I231 (o_0r0d[31], ofint_0n[31], gate1137_0n, initialise);
  C3 I232 (internal_0n[34], complete1134_0n[0], complete1134_0n[1], complete1134_0n[2]);
  C3 I233 (internal_0n[35], complete1134_0n[3], complete1134_0n[4], complete1134_0n[5]);
  C3 I234 (internal_0n[36], complete1134_0n[6], complete1134_0n[7], complete1134_0n[8]);
  C3 I235 (internal_0n[37], complete1134_0n[9], complete1134_0n[10], complete1134_0n[11]);
  C3 I236 (internal_0n[38], complete1134_0n[12], complete1134_0n[13], complete1134_0n[14]);
  C3 I237 (internal_0n[39], complete1134_0n[15], complete1134_0n[16], complete1134_0n[17]);
  C3 I238 (internal_0n[40], complete1134_0n[18], complete1134_0n[19], complete1134_0n[20]);
  C3 I239 (internal_0n[41], complete1134_0n[21], complete1134_0n[22], complete1134_0n[23]);
  C3 I240 (internal_0n[42], complete1134_0n[24], complete1134_0n[25], complete1134_0n[26]);
  C3 I241 (internal_0n[43], complete1134_0n[27], complete1134_0n[28], complete1134_0n[29]);
  C2 I242 (internal_0n[44], complete1134_0n[30], complete1134_0n[31]);
  C2 I243 (internal_0n[45], complete1134_0n[32], complete1134_0n[33]);
  C3 I244 (internal_0n[46], internal_0n[34], internal_0n[35], internal_0n[36]);
  C3 I245 (internal_0n[47], internal_0n[37], internal_0n[38], internal_0n[39]);
  C3 I246 (internal_0n[48], internal_0n[40], internal_0n[41], internal_0n[42]);
  C3 I247 (internal_0n[49], internal_0n[43], internal_0n[44], internal_0n[45]);
  C2 I248 (internal_0n[50], internal_0n[46], internal_0n[47]);
  C2 I249 (internal_0n[51], internal_0n[48], internal_0n[49]);
  C2 I250 (i_0a, internal_0n[50], internal_0n[51]);
  OR2 I251 (complete1134_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I252 (complete1134_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I253 (complete1134_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I254 (complete1134_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I255 (complete1134_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I256 (complete1134_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I257 (complete1134_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I258 (complete1134_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I259 (complete1134_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I260 (complete1134_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I261 (complete1134_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I262 (complete1134_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I263 (complete1134_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I264 (complete1134_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I265 (complete1134_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I266 (complete1134_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I267 (complete1134_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I268 (complete1134_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I269 (complete1134_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I270 (complete1134_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I271 (complete1134_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I272 (complete1134_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I273 (complete1134_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I274 (complete1134_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I275 (complete1134_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I276 (complete1134_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I277 (complete1134_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I278 (complete1134_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I279 (complete1134_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I280 (complete1134_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I281 (complete1134_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I282 (complete1134_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I283 (complete1134_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I284 (complete1134_0n[33], ifint_0n[33], itint_0n[33]);
  INV I285 (gate1133_0n, iaint_0n);
  C2RI I286 (itint_0n[0], i_0r1d[0], gate1133_0n, initialise);
  C2RI I287 (itint_0n[1], i_0r1d[1], gate1133_0n, initialise);
  C2RI I288 (itint_0n[2], i_0r1d[2], gate1133_0n, initialise);
  C2RI I289 (itint_0n[3], i_0r1d[3], gate1133_0n, initialise);
  C2RI I290 (itint_0n[4], i_0r1d[4], gate1133_0n, initialise);
  C2RI I291 (itint_0n[5], i_0r1d[5], gate1133_0n, initialise);
  C2RI I292 (itint_0n[6], i_0r1d[6], gate1133_0n, initialise);
  C2RI I293 (itint_0n[7], i_0r1d[7], gate1133_0n, initialise);
  C2RI I294 (itint_0n[8], i_0r1d[8], gate1133_0n, initialise);
  C2RI I295 (itint_0n[9], i_0r1d[9], gate1133_0n, initialise);
  C2RI I296 (itint_0n[10], i_0r1d[10], gate1133_0n, initialise);
  C2RI I297 (itint_0n[11], i_0r1d[11], gate1133_0n, initialise);
  C2RI I298 (itint_0n[12], i_0r1d[12], gate1133_0n, initialise);
  C2RI I299 (itint_0n[13], i_0r1d[13], gate1133_0n, initialise);
  C2RI I300 (itint_0n[14], i_0r1d[14], gate1133_0n, initialise);
  C2RI I301 (itint_0n[15], i_0r1d[15], gate1133_0n, initialise);
  C2RI I302 (itint_0n[16], i_0r1d[16], gate1133_0n, initialise);
  C2RI I303 (itint_0n[17], i_0r1d[17], gate1133_0n, initialise);
  C2RI I304 (itint_0n[18], i_0r1d[18], gate1133_0n, initialise);
  C2RI I305 (itint_0n[19], i_0r1d[19], gate1133_0n, initialise);
  C2RI I306 (itint_0n[20], i_0r1d[20], gate1133_0n, initialise);
  C2RI I307 (itint_0n[21], i_0r1d[21], gate1133_0n, initialise);
  C2RI I308 (itint_0n[22], i_0r1d[22], gate1133_0n, initialise);
  C2RI I309 (itint_0n[23], i_0r1d[23], gate1133_0n, initialise);
  C2RI I310 (itint_0n[24], i_0r1d[24], gate1133_0n, initialise);
  C2RI I311 (itint_0n[25], i_0r1d[25], gate1133_0n, initialise);
  C2RI I312 (itint_0n[26], i_0r1d[26], gate1133_0n, initialise);
  C2RI I313 (itint_0n[27], i_0r1d[27], gate1133_0n, initialise);
  C2RI I314 (itint_0n[28], i_0r1d[28], gate1133_0n, initialise);
  C2RI I315 (itint_0n[29], i_0r1d[29], gate1133_0n, initialise);
  C2RI I316 (itint_0n[30], i_0r1d[30], gate1133_0n, initialise);
  C2RI I317 (itint_0n[31], i_0r1d[31], gate1133_0n, initialise);
  C2RI I318 (itint_0n[32], i_0r1d[32], gate1133_0n, initialise);
  C2RI I319 (itint_0n[33], i_0r1d[33], gate1133_0n, initialise);
  C2RI I320 (ifint_0n[0], i_0r0d[0], gate1133_0n, initialise);
  C2RI I321 (ifint_0n[1], i_0r0d[1], gate1133_0n, initialise);
  C2RI I322 (ifint_0n[2], i_0r0d[2], gate1133_0n, initialise);
  C2RI I323 (ifint_0n[3], i_0r0d[3], gate1133_0n, initialise);
  C2RI I324 (ifint_0n[4], i_0r0d[4], gate1133_0n, initialise);
  C2RI I325 (ifint_0n[5], i_0r0d[5], gate1133_0n, initialise);
  C2RI I326 (ifint_0n[6], i_0r0d[6], gate1133_0n, initialise);
  C2RI I327 (ifint_0n[7], i_0r0d[7], gate1133_0n, initialise);
  C2RI I328 (ifint_0n[8], i_0r0d[8], gate1133_0n, initialise);
  C2RI I329 (ifint_0n[9], i_0r0d[9], gate1133_0n, initialise);
  C2RI I330 (ifint_0n[10], i_0r0d[10], gate1133_0n, initialise);
  C2RI I331 (ifint_0n[11], i_0r0d[11], gate1133_0n, initialise);
  C2RI I332 (ifint_0n[12], i_0r0d[12], gate1133_0n, initialise);
  C2RI I333 (ifint_0n[13], i_0r0d[13], gate1133_0n, initialise);
  C2RI I334 (ifint_0n[14], i_0r0d[14], gate1133_0n, initialise);
  C2RI I335 (ifint_0n[15], i_0r0d[15], gate1133_0n, initialise);
  C2RI I336 (ifint_0n[16], i_0r0d[16], gate1133_0n, initialise);
  C2RI I337 (ifint_0n[17], i_0r0d[17], gate1133_0n, initialise);
  C2RI I338 (ifint_0n[18], i_0r0d[18], gate1133_0n, initialise);
  C2RI I339 (ifint_0n[19], i_0r0d[19], gate1133_0n, initialise);
  C2RI I340 (ifint_0n[20], i_0r0d[20], gate1133_0n, initialise);
  C2RI I341 (ifint_0n[21], i_0r0d[21], gate1133_0n, initialise);
  C2RI I342 (ifint_0n[22], i_0r0d[22], gate1133_0n, initialise);
  C2RI I343 (ifint_0n[23], i_0r0d[23], gate1133_0n, initialise);
  C2RI I344 (ifint_0n[24], i_0r0d[24], gate1133_0n, initialise);
  C2RI I345 (ifint_0n[25], i_0r0d[25], gate1133_0n, initialise);
  C2RI I346 (ifint_0n[26], i_0r0d[26], gate1133_0n, initialise);
  C2RI I347 (ifint_0n[27], i_0r0d[27], gate1133_0n, initialise);
  C2RI I348 (ifint_0n[28], i_0r0d[28], gate1133_0n, initialise);
  C2RI I349 (ifint_0n[29], i_0r0d[29], gate1133_0n, initialise);
  C2RI I350 (ifint_0n[30], i_0r0d[30], gate1133_0n, initialise);
  C2RI I351 (ifint_0n[31], i_0r0d[31], gate1133_0n, initialise);
  C2RI I352 (ifint_0n[32], i_0r0d[32], gate1133_0n, initialise);
  C2RI I353 (ifint_0n[33], i_0r0d[33], gate1133_0n, initialise);
  C2 I354 (otint_1n[0], sel_1n, itint_0n[0]);
  C2 I355 (otint_1n[1], sel_1n, itint_0n[1]);
  C2 I356 (otint_1n[2], sel_1n, itint_0n[2]);
  C2 I357 (otint_1n[3], sel_1n, itint_0n[3]);
  C2 I358 (otint_1n[4], sel_1n, itint_0n[4]);
  C2 I359 (otint_1n[5], sel_1n, itint_0n[5]);
  C2 I360 (otint_1n[6], sel_1n, itint_0n[6]);
  C2 I361 (otint_1n[7], sel_1n, itint_0n[7]);
  C2 I362 (otint_1n[8], sel_1n, itint_0n[8]);
  C2 I363 (otint_1n[9], sel_1n, itint_0n[9]);
  C2 I364 (otint_1n[10], sel_1n, itint_0n[10]);
  C2 I365 (otint_1n[11], sel_1n, itint_0n[11]);
  C2 I366 (otint_1n[12], sel_1n, itint_0n[12]);
  C2 I367 (otint_1n[13], sel_1n, itint_0n[13]);
  C2 I368 (otint_1n[14], sel_1n, itint_0n[14]);
  C2 I369 (otint_1n[15], sel_1n, itint_0n[15]);
  C2 I370 (otint_1n[16], sel_1n, itint_0n[16]);
  C2 I371 (otint_1n[17], sel_1n, itint_0n[17]);
  C2 I372 (otint_1n[18], sel_1n, itint_0n[18]);
  C2 I373 (otint_1n[19], sel_1n, itint_0n[19]);
  C2 I374 (otint_1n[20], sel_1n, itint_0n[20]);
  C2 I375 (otint_1n[21], sel_1n, itint_0n[21]);
  C2 I376 (otint_1n[22], sel_1n, itint_0n[22]);
  C2 I377 (otint_1n[23], sel_1n, itint_0n[23]);
  C2 I378 (otint_1n[24], sel_1n, itint_0n[24]);
  C2 I379 (otint_1n[25], sel_1n, itint_0n[25]);
  C2 I380 (otint_1n[26], sel_1n, itint_0n[26]);
  C2 I381 (otint_1n[27], sel_1n, itint_0n[27]);
  C2 I382 (otint_1n[28], sel_1n, itint_0n[28]);
  C2 I383 (otint_1n[29], sel_1n, itint_0n[29]);
  C2 I384 (otint_1n[30], sel_1n, itint_0n[30]);
  C2 I385 (otint_1n[31], sel_1n, itint_0n[31]);
  C2 I386 (otint_0n[0], sel_0n, itint_0n[0]);
  C2 I387 (otint_0n[1], sel_0n, itint_0n[1]);
  C2 I388 (otint_0n[2], sel_0n, itint_0n[2]);
  C2 I389 (otint_0n[3], sel_0n, itint_0n[3]);
  C2 I390 (otint_0n[4], sel_0n, itint_0n[4]);
  C2 I391 (otint_0n[5], sel_0n, itint_0n[5]);
  C2 I392 (otint_0n[6], sel_0n, itint_0n[6]);
  C2 I393 (otint_0n[7], sel_0n, itint_0n[7]);
  C2 I394 (otint_0n[8], sel_0n, itint_0n[8]);
  C2 I395 (otint_0n[9], sel_0n, itint_0n[9]);
  C2 I396 (otint_0n[10], sel_0n, itint_0n[10]);
  C2 I397 (otint_0n[11], sel_0n, itint_0n[11]);
  C2 I398 (otint_0n[12], sel_0n, itint_0n[12]);
  C2 I399 (otint_0n[13], sel_0n, itint_0n[13]);
  C2 I400 (otint_0n[14], sel_0n, itint_0n[14]);
  C2 I401 (otint_0n[15], sel_0n, itint_0n[15]);
  C2 I402 (otint_0n[16], sel_0n, itint_0n[16]);
  C2 I403 (otint_0n[17], sel_0n, itint_0n[17]);
  C2 I404 (otint_0n[18], sel_0n, itint_0n[18]);
  C2 I405 (otint_0n[19], sel_0n, itint_0n[19]);
  C2 I406 (otint_0n[20], sel_0n, itint_0n[20]);
  C2 I407 (otint_0n[21], sel_0n, itint_0n[21]);
  C2 I408 (otint_0n[22], sel_0n, itint_0n[22]);
  C2 I409 (otint_0n[23], sel_0n, itint_0n[23]);
  C2 I410 (otint_0n[24], sel_0n, itint_0n[24]);
  C2 I411 (otint_0n[25], sel_0n, itint_0n[25]);
  C2 I412 (otint_0n[26], sel_0n, itint_0n[26]);
  C2 I413 (otint_0n[27], sel_0n, itint_0n[27]);
  C2 I414 (otint_0n[28], sel_0n, itint_0n[28]);
  C2 I415 (otint_0n[29], sel_0n, itint_0n[29]);
  C2 I416 (otint_0n[30], sel_0n, itint_0n[30]);
  C2 I417 (otint_0n[31], sel_0n, itint_0n[31]);
  C2 I418 (ofint_1n[0], sel_1n, ifint_0n[0]);
  C2 I419 (ofint_1n[1], sel_1n, ifint_0n[1]);
  C2 I420 (ofint_1n[2], sel_1n, ifint_0n[2]);
  C2 I421 (ofint_1n[3], sel_1n, ifint_0n[3]);
  C2 I422 (ofint_1n[4], sel_1n, ifint_0n[4]);
  C2 I423 (ofint_1n[5], sel_1n, ifint_0n[5]);
  C2 I424 (ofint_1n[6], sel_1n, ifint_0n[6]);
  C2 I425 (ofint_1n[7], sel_1n, ifint_0n[7]);
  C2 I426 (ofint_1n[8], sel_1n, ifint_0n[8]);
  C2 I427 (ofint_1n[9], sel_1n, ifint_0n[9]);
  C2 I428 (ofint_1n[10], sel_1n, ifint_0n[10]);
  C2 I429 (ofint_1n[11], sel_1n, ifint_0n[11]);
  C2 I430 (ofint_1n[12], sel_1n, ifint_0n[12]);
  C2 I431 (ofint_1n[13], sel_1n, ifint_0n[13]);
  C2 I432 (ofint_1n[14], sel_1n, ifint_0n[14]);
  C2 I433 (ofint_1n[15], sel_1n, ifint_0n[15]);
  C2 I434 (ofint_1n[16], sel_1n, ifint_0n[16]);
  C2 I435 (ofint_1n[17], sel_1n, ifint_0n[17]);
  C2 I436 (ofint_1n[18], sel_1n, ifint_0n[18]);
  C2 I437 (ofint_1n[19], sel_1n, ifint_0n[19]);
  C2 I438 (ofint_1n[20], sel_1n, ifint_0n[20]);
  C2 I439 (ofint_1n[21], sel_1n, ifint_0n[21]);
  C2 I440 (ofint_1n[22], sel_1n, ifint_0n[22]);
  C2 I441 (ofint_1n[23], sel_1n, ifint_0n[23]);
  C2 I442 (ofint_1n[24], sel_1n, ifint_0n[24]);
  C2 I443 (ofint_1n[25], sel_1n, ifint_0n[25]);
  C2 I444 (ofint_1n[26], sel_1n, ifint_0n[26]);
  C2 I445 (ofint_1n[27], sel_1n, ifint_0n[27]);
  C2 I446 (ofint_1n[28], sel_1n, ifint_0n[28]);
  C2 I447 (ofint_1n[29], sel_1n, ifint_0n[29]);
  C2 I448 (ofint_1n[30], sel_1n, ifint_0n[30]);
  C2 I449 (ofint_1n[31], sel_1n, ifint_0n[31]);
  C2 I450 (ofint_0n[0], sel_0n, ifint_0n[0]);
  C2 I451 (ofint_0n[1], sel_0n, ifint_0n[1]);
  C2 I452 (ofint_0n[2], sel_0n, ifint_0n[2]);
  C2 I453 (ofint_0n[3], sel_0n, ifint_0n[3]);
  C2 I454 (ofint_0n[4], sel_0n, ifint_0n[4]);
  C2 I455 (ofint_0n[5], sel_0n, ifint_0n[5]);
  C2 I456 (ofint_0n[6], sel_0n, ifint_0n[6]);
  C2 I457 (ofint_0n[7], sel_0n, ifint_0n[7]);
  C2 I458 (ofint_0n[8], sel_0n, ifint_0n[8]);
  C2 I459 (ofint_0n[9], sel_0n, ifint_0n[9]);
  C2 I460 (ofint_0n[10], sel_0n, ifint_0n[10]);
  C2 I461 (ofint_0n[11], sel_0n, ifint_0n[11]);
  C2 I462 (ofint_0n[12], sel_0n, ifint_0n[12]);
  C2 I463 (ofint_0n[13], sel_0n, ifint_0n[13]);
  C2 I464 (ofint_0n[14], sel_0n, ifint_0n[14]);
  C2 I465 (ofint_0n[15], sel_0n, ifint_0n[15]);
  C2 I466 (ofint_0n[16], sel_0n, ifint_0n[16]);
  C2 I467 (ofint_0n[17], sel_0n, ifint_0n[17]);
  C2 I468 (ofint_0n[18], sel_0n, ifint_0n[18]);
  C2 I469 (ofint_0n[19], sel_0n, ifint_0n[19]);
  C2 I470 (ofint_0n[20], sel_0n, ifint_0n[20]);
  C2 I471 (ofint_0n[21], sel_0n, ifint_0n[21]);
  C2 I472 (ofint_0n[22], sel_0n, ifint_0n[22]);
  C2 I473 (ofint_0n[23], sel_0n, ifint_0n[23]);
  C2 I474 (ofint_0n[24], sel_0n, ifint_0n[24]);
  C2 I475 (ofint_0n[25], sel_0n, ifint_0n[25]);
  C2 I476 (ofint_0n[26], sel_0n, ifint_0n[26]);
  C2 I477 (ofint_0n[27], sel_0n, ifint_0n[27]);
  C2 I478 (ofint_0n[28], sel_0n, ifint_0n[28]);
  C2 I479 (ofint_0n[29], sel_0n, ifint_0n[29]);
  C2 I480 (ofint_0n[30], sel_0n, ifint_0n[30]);
  C2 I481 (ofint_0n[31], sel_0n, ifint_0n[31]);
  C3 I482 (internal_0n[52], complete1130_0n[0], complete1130_0n[1], complete1130_0n[2]);
  C3 I483 (internal_0n[53], complete1130_0n[3], complete1130_0n[4], complete1130_0n[5]);
  C3 I484 (internal_0n[54], complete1130_0n[6], complete1130_0n[7], complete1130_0n[8]);
  C3 I485 (internal_0n[55], complete1130_0n[9], complete1130_0n[10], complete1130_0n[11]);
  C3 I486 (internal_0n[56], complete1130_0n[12], complete1130_0n[13], complete1130_0n[14]);
  C3 I487 (internal_0n[57], complete1130_0n[15], complete1130_0n[16], complete1130_0n[17]);
  C3 I488 (internal_0n[58], complete1130_0n[18], complete1130_0n[19], complete1130_0n[20]);
  C3 I489 (internal_0n[59], complete1130_0n[21], complete1130_0n[22], complete1130_0n[23]);
  C3 I490 (internal_0n[60], complete1130_0n[24], complete1130_0n[25], complete1130_0n[26]);
  C3 I491 (internal_0n[61], complete1130_0n[27], complete1130_0n[28], complete1130_0n[29]);
  C2 I492 (internal_0n[62], complete1130_0n[30], complete1130_0n[31]);
  C2 I493 (internal_0n[63], complete1130_0n[32], complete1130_0n[33]);
  C3 I494 (internal_0n[64], internal_0n[52], internal_0n[53], internal_0n[54]);
  C3 I495 (internal_0n[65], internal_0n[55], internal_0n[56], internal_0n[57]);
  C3 I496 (internal_0n[66], internal_0n[58], internal_0n[59], internal_0n[60]);
  C3 I497 (internal_0n[67], internal_0n[61], internal_0n[62], internal_0n[63]);
  C2 I498 (internal_0n[68], internal_0n[64], internal_0n[65]);
  C2 I499 (internal_0n[69], internal_0n[66], internal_0n[67]);
  C2 I500 (icomplete_0n, internal_0n[68], internal_0n[69]);
  OR2 I501 (complete1130_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I502 (complete1130_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I503 (complete1130_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I504 (complete1130_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I505 (complete1130_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I506 (complete1130_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I507 (complete1130_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I508 (complete1130_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I509 (complete1130_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I510 (complete1130_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I511 (complete1130_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I512 (complete1130_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I513 (complete1130_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I514 (complete1130_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I515 (complete1130_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I516 (complete1130_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I517 (complete1130_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I518 (complete1130_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I519 (complete1130_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I520 (complete1130_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I521 (complete1130_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I522 (complete1130_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I523 (complete1130_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I524 (complete1130_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I525 (complete1130_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I526 (complete1130_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I527 (complete1130_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I528 (complete1130_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I529 (complete1130_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I530 (complete1130_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I531 (complete1130_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I532 (complete1130_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I533 (complete1130_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I534 (complete1130_0n[33], ifint_0n[33], itint_0n[33]);
  C2 I535 (matchi_1n, ifint_0n[32], itint_0n[33]);
  assign sel_1n = matchi_1n;
  C2 I537 (matchi_0n, ifint_0n[33], itint_0n[32]);
  assign sel_0n = matchi_0n;
endmodule

module BrzS_35_l12__2832_203_29_l144__28_28_28_28_m70m (
  i_0r0d, i_0r1d, i_0a,
  o_0r0d, o_0r1d, o_0a,
  o_1r0d, o_1r1d, o_1a,
  o_2r0d, o_2r1d, o_2a,
  initialise
);
  input [34:0] i_0r0d;
  input [34:0] i_0r1d;
  output i_0a;
  output [31:0] o_0r0d;
  output [31:0] o_0r1d;
  input o_0a;
  output [31:0] o_1r0d;
  output [31:0] o_1r1d;
  input o_1a;
  output [31:0] o_2r0d;
  output [31:0] o_2r1d;
  input o_2a;
  input initialise;
  wire [86:0] internal_0n;
  wire icomplete_0n;
  wire sel_0n;
  wire sel_1n;
  wire sel_2n;
  wire matchi_0n;
  wire matchi_1n;
  wire matchi_2n;
  wire [34:0] ifint_0n;
  wire [34:0] itint_0n;
  wire iaint_0n;
  wire [31:0] ofint_0n;
  wire [31:0] ofint_1n;
  wire [31:0] ofint_2n;
  wire [31:0] otint_0n;
  wire [31:0] otint_1n;
  wire [31:0] otint_2n;
  wire oaint_0n;
  wire oaint_1n;
  wire oaint_2n;
  wire oack_0n;
  wire [31:0] complete1159_0n;
  wire gate1158_0n;
  wire [31:0] complete1155_0n;
  wire gate1154_0n;
  wire [31:0] complete1151_0n;
  wire gate1150_0n;
  wire [34:0] complete1147_0n;
  wire gate1146_0n;
  wire [34:0] complete1143_0n;
  C2 I0 (iaint_0n, oack_0n, icomplete_0n);
  OR3 I1 (oack_0n, oaint_0n, oaint_1n, oaint_2n);
  C3 I2 (internal_0n[0], complete1159_0n[0], complete1159_0n[1], complete1159_0n[2]);
  C3 I3 (internal_0n[1], complete1159_0n[3], complete1159_0n[4], complete1159_0n[5]);
  C3 I4 (internal_0n[2], complete1159_0n[6], complete1159_0n[7], complete1159_0n[8]);
  C3 I5 (internal_0n[3], complete1159_0n[9], complete1159_0n[10], complete1159_0n[11]);
  C3 I6 (internal_0n[4], complete1159_0n[12], complete1159_0n[13], complete1159_0n[14]);
  C3 I7 (internal_0n[5], complete1159_0n[15], complete1159_0n[16], complete1159_0n[17]);
  C3 I8 (internal_0n[6], complete1159_0n[18], complete1159_0n[19], complete1159_0n[20]);
  C3 I9 (internal_0n[7], complete1159_0n[21], complete1159_0n[22], complete1159_0n[23]);
  C3 I10 (internal_0n[8], complete1159_0n[24], complete1159_0n[25], complete1159_0n[26]);
  C3 I11 (internal_0n[9], complete1159_0n[27], complete1159_0n[28], complete1159_0n[29]);
  C2 I12 (internal_0n[10], complete1159_0n[30], complete1159_0n[31]);
  C3 I13 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I14 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I15 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I16 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I17 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I18 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I19 (oaint_2n, internal_0n[15], internal_0n[16]);
  OR2 I20 (complete1159_0n[0], o_2r0d[0], o_2r1d[0]);
  OR2 I21 (complete1159_0n[1], o_2r0d[1], o_2r1d[1]);
  OR2 I22 (complete1159_0n[2], o_2r0d[2], o_2r1d[2]);
  OR2 I23 (complete1159_0n[3], o_2r0d[3], o_2r1d[3]);
  OR2 I24 (complete1159_0n[4], o_2r0d[4], o_2r1d[4]);
  OR2 I25 (complete1159_0n[5], o_2r0d[5], o_2r1d[5]);
  OR2 I26 (complete1159_0n[6], o_2r0d[6], o_2r1d[6]);
  OR2 I27 (complete1159_0n[7], o_2r0d[7], o_2r1d[7]);
  OR2 I28 (complete1159_0n[8], o_2r0d[8], o_2r1d[8]);
  OR2 I29 (complete1159_0n[9], o_2r0d[9], o_2r1d[9]);
  OR2 I30 (complete1159_0n[10], o_2r0d[10], o_2r1d[10]);
  OR2 I31 (complete1159_0n[11], o_2r0d[11], o_2r1d[11]);
  OR2 I32 (complete1159_0n[12], o_2r0d[12], o_2r1d[12]);
  OR2 I33 (complete1159_0n[13], o_2r0d[13], o_2r1d[13]);
  OR2 I34 (complete1159_0n[14], o_2r0d[14], o_2r1d[14]);
  OR2 I35 (complete1159_0n[15], o_2r0d[15], o_2r1d[15]);
  OR2 I36 (complete1159_0n[16], o_2r0d[16], o_2r1d[16]);
  OR2 I37 (complete1159_0n[17], o_2r0d[17], o_2r1d[17]);
  OR2 I38 (complete1159_0n[18], o_2r0d[18], o_2r1d[18]);
  OR2 I39 (complete1159_0n[19], o_2r0d[19], o_2r1d[19]);
  OR2 I40 (complete1159_0n[20], o_2r0d[20], o_2r1d[20]);
  OR2 I41 (complete1159_0n[21], o_2r0d[21], o_2r1d[21]);
  OR2 I42 (complete1159_0n[22], o_2r0d[22], o_2r1d[22]);
  OR2 I43 (complete1159_0n[23], o_2r0d[23], o_2r1d[23]);
  OR2 I44 (complete1159_0n[24], o_2r0d[24], o_2r1d[24]);
  OR2 I45 (complete1159_0n[25], o_2r0d[25], o_2r1d[25]);
  OR2 I46 (complete1159_0n[26], o_2r0d[26], o_2r1d[26]);
  OR2 I47 (complete1159_0n[27], o_2r0d[27], o_2r1d[27]);
  OR2 I48 (complete1159_0n[28], o_2r0d[28], o_2r1d[28]);
  OR2 I49 (complete1159_0n[29], o_2r0d[29], o_2r1d[29]);
  OR2 I50 (complete1159_0n[30], o_2r0d[30], o_2r1d[30]);
  OR2 I51 (complete1159_0n[31], o_2r0d[31], o_2r1d[31]);
  INV I52 (gate1158_0n, o_2a);
  C2RI I53 (o_2r1d[0], otint_2n[0], gate1158_0n, initialise);
  C2RI I54 (o_2r1d[1], otint_2n[1], gate1158_0n, initialise);
  C2RI I55 (o_2r1d[2], otint_2n[2], gate1158_0n, initialise);
  C2RI I56 (o_2r1d[3], otint_2n[3], gate1158_0n, initialise);
  C2RI I57 (o_2r1d[4], otint_2n[4], gate1158_0n, initialise);
  C2RI I58 (o_2r1d[5], otint_2n[5], gate1158_0n, initialise);
  C2RI I59 (o_2r1d[6], otint_2n[6], gate1158_0n, initialise);
  C2RI I60 (o_2r1d[7], otint_2n[7], gate1158_0n, initialise);
  C2RI I61 (o_2r1d[8], otint_2n[8], gate1158_0n, initialise);
  C2RI I62 (o_2r1d[9], otint_2n[9], gate1158_0n, initialise);
  C2RI I63 (o_2r1d[10], otint_2n[10], gate1158_0n, initialise);
  C2RI I64 (o_2r1d[11], otint_2n[11], gate1158_0n, initialise);
  C2RI I65 (o_2r1d[12], otint_2n[12], gate1158_0n, initialise);
  C2RI I66 (o_2r1d[13], otint_2n[13], gate1158_0n, initialise);
  C2RI I67 (o_2r1d[14], otint_2n[14], gate1158_0n, initialise);
  C2RI I68 (o_2r1d[15], otint_2n[15], gate1158_0n, initialise);
  C2RI I69 (o_2r1d[16], otint_2n[16], gate1158_0n, initialise);
  C2RI I70 (o_2r1d[17], otint_2n[17], gate1158_0n, initialise);
  C2RI I71 (o_2r1d[18], otint_2n[18], gate1158_0n, initialise);
  C2RI I72 (o_2r1d[19], otint_2n[19], gate1158_0n, initialise);
  C2RI I73 (o_2r1d[20], otint_2n[20], gate1158_0n, initialise);
  C2RI I74 (o_2r1d[21], otint_2n[21], gate1158_0n, initialise);
  C2RI I75 (o_2r1d[22], otint_2n[22], gate1158_0n, initialise);
  C2RI I76 (o_2r1d[23], otint_2n[23], gate1158_0n, initialise);
  C2RI I77 (o_2r1d[24], otint_2n[24], gate1158_0n, initialise);
  C2RI I78 (o_2r1d[25], otint_2n[25], gate1158_0n, initialise);
  C2RI I79 (o_2r1d[26], otint_2n[26], gate1158_0n, initialise);
  C2RI I80 (o_2r1d[27], otint_2n[27], gate1158_0n, initialise);
  C2RI I81 (o_2r1d[28], otint_2n[28], gate1158_0n, initialise);
  C2RI I82 (o_2r1d[29], otint_2n[29], gate1158_0n, initialise);
  C2RI I83 (o_2r1d[30], otint_2n[30], gate1158_0n, initialise);
  C2RI I84 (o_2r1d[31], otint_2n[31], gate1158_0n, initialise);
  C2RI I85 (o_2r0d[0], ofint_2n[0], gate1158_0n, initialise);
  C2RI I86 (o_2r0d[1], ofint_2n[1], gate1158_0n, initialise);
  C2RI I87 (o_2r0d[2], ofint_2n[2], gate1158_0n, initialise);
  C2RI I88 (o_2r0d[3], ofint_2n[3], gate1158_0n, initialise);
  C2RI I89 (o_2r0d[4], ofint_2n[4], gate1158_0n, initialise);
  C2RI I90 (o_2r0d[5], ofint_2n[5], gate1158_0n, initialise);
  C2RI I91 (o_2r0d[6], ofint_2n[6], gate1158_0n, initialise);
  C2RI I92 (o_2r0d[7], ofint_2n[7], gate1158_0n, initialise);
  C2RI I93 (o_2r0d[8], ofint_2n[8], gate1158_0n, initialise);
  C2RI I94 (o_2r0d[9], ofint_2n[9], gate1158_0n, initialise);
  C2RI I95 (o_2r0d[10], ofint_2n[10], gate1158_0n, initialise);
  C2RI I96 (o_2r0d[11], ofint_2n[11], gate1158_0n, initialise);
  C2RI I97 (o_2r0d[12], ofint_2n[12], gate1158_0n, initialise);
  C2RI I98 (o_2r0d[13], ofint_2n[13], gate1158_0n, initialise);
  C2RI I99 (o_2r0d[14], ofint_2n[14], gate1158_0n, initialise);
  C2RI I100 (o_2r0d[15], ofint_2n[15], gate1158_0n, initialise);
  C2RI I101 (o_2r0d[16], ofint_2n[16], gate1158_0n, initialise);
  C2RI I102 (o_2r0d[17], ofint_2n[17], gate1158_0n, initialise);
  C2RI I103 (o_2r0d[18], ofint_2n[18], gate1158_0n, initialise);
  C2RI I104 (o_2r0d[19], ofint_2n[19], gate1158_0n, initialise);
  C2RI I105 (o_2r0d[20], ofint_2n[20], gate1158_0n, initialise);
  C2RI I106 (o_2r0d[21], ofint_2n[21], gate1158_0n, initialise);
  C2RI I107 (o_2r0d[22], ofint_2n[22], gate1158_0n, initialise);
  C2RI I108 (o_2r0d[23], ofint_2n[23], gate1158_0n, initialise);
  C2RI I109 (o_2r0d[24], ofint_2n[24], gate1158_0n, initialise);
  C2RI I110 (o_2r0d[25], ofint_2n[25], gate1158_0n, initialise);
  C2RI I111 (o_2r0d[26], ofint_2n[26], gate1158_0n, initialise);
  C2RI I112 (o_2r0d[27], ofint_2n[27], gate1158_0n, initialise);
  C2RI I113 (o_2r0d[28], ofint_2n[28], gate1158_0n, initialise);
  C2RI I114 (o_2r0d[29], ofint_2n[29], gate1158_0n, initialise);
  C2RI I115 (o_2r0d[30], ofint_2n[30], gate1158_0n, initialise);
  C2RI I116 (o_2r0d[31], ofint_2n[31], gate1158_0n, initialise);
  C3 I117 (internal_0n[17], complete1155_0n[0], complete1155_0n[1], complete1155_0n[2]);
  C3 I118 (internal_0n[18], complete1155_0n[3], complete1155_0n[4], complete1155_0n[5]);
  C3 I119 (internal_0n[19], complete1155_0n[6], complete1155_0n[7], complete1155_0n[8]);
  C3 I120 (internal_0n[20], complete1155_0n[9], complete1155_0n[10], complete1155_0n[11]);
  C3 I121 (internal_0n[21], complete1155_0n[12], complete1155_0n[13], complete1155_0n[14]);
  C3 I122 (internal_0n[22], complete1155_0n[15], complete1155_0n[16], complete1155_0n[17]);
  C3 I123 (internal_0n[23], complete1155_0n[18], complete1155_0n[19], complete1155_0n[20]);
  C3 I124 (internal_0n[24], complete1155_0n[21], complete1155_0n[22], complete1155_0n[23]);
  C3 I125 (internal_0n[25], complete1155_0n[24], complete1155_0n[25], complete1155_0n[26]);
  C3 I126 (internal_0n[26], complete1155_0n[27], complete1155_0n[28], complete1155_0n[29]);
  C2 I127 (internal_0n[27], complete1155_0n[30], complete1155_0n[31]);
  C3 I128 (internal_0n[28], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I129 (internal_0n[29], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I130 (internal_0n[30], internal_0n[23], internal_0n[24], internal_0n[25]);
  C2 I131 (internal_0n[31], internal_0n[26], internal_0n[27]);
  C2 I132 (internal_0n[32], internal_0n[28], internal_0n[29]);
  C2 I133 (internal_0n[33], internal_0n[30], internal_0n[31]);
  C2 I134 (oaint_1n, internal_0n[32], internal_0n[33]);
  OR2 I135 (complete1155_0n[0], o_1r0d[0], o_1r1d[0]);
  OR2 I136 (complete1155_0n[1], o_1r0d[1], o_1r1d[1]);
  OR2 I137 (complete1155_0n[2], o_1r0d[2], o_1r1d[2]);
  OR2 I138 (complete1155_0n[3], o_1r0d[3], o_1r1d[3]);
  OR2 I139 (complete1155_0n[4], o_1r0d[4], o_1r1d[4]);
  OR2 I140 (complete1155_0n[5], o_1r0d[5], o_1r1d[5]);
  OR2 I141 (complete1155_0n[6], o_1r0d[6], o_1r1d[6]);
  OR2 I142 (complete1155_0n[7], o_1r0d[7], o_1r1d[7]);
  OR2 I143 (complete1155_0n[8], o_1r0d[8], o_1r1d[8]);
  OR2 I144 (complete1155_0n[9], o_1r0d[9], o_1r1d[9]);
  OR2 I145 (complete1155_0n[10], o_1r0d[10], o_1r1d[10]);
  OR2 I146 (complete1155_0n[11], o_1r0d[11], o_1r1d[11]);
  OR2 I147 (complete1155_0n[12], o_1r0d[12], o_1r1d[12]);
  OR2 I148 (complete1155_0n[13], o_1r0d[13], o_1r1d[13]);
  OR2 I149 (complete1155_0n[14], o_1r0d[14], o_1r1d[14]);
  OR2 I150 (complete1155_0n[15], o_1r0d[15], o_1r1d[15]);
  OR2 I151 (complete1155_0n[16], o_1r0d[16], o_1r1d[16]);
  OR2 I152 (complete1155_0n[17], o_1r0d[17], o_1r1d[17]);
  OR2 I153 (complete1155_0n[18], o_1r0d[18], o_1r1d[18]);
  OR2 I154 (complete1155_0n[19], o_1r0d[19], o_1r1d[19]);
  OR2 I155 (complete1155_0n[20], o_1r0d[20], o_1r1d[20]);
  OR2 I156 (complete1155_0n[21], o_1r0d[21], o_1r1d[21]);
  OR2 I157 (complete1155_0n[22], o_1r0d[22], o_1r1d[22]);
  OR2 I158 (complete1155_0n[23], o_1r0d[23], o_1r1d[23]);
  OR2 I159 (complete1155_0n[24], o_1r0d[24], o_1r1d[24]);
  OR2 I160 (complete1155_0n[25], o_1r0d[25], o_1r1d[25]);
  OR2 I161 (complete1155_0n[26], o_1r0d[26], o_1r1d[26]);
  OR2 I162 (complete1155_0n[27], o_1r0d[27], o_1r1d[27]);
  OR2 I163 (complete1155_0n[28], o_1r0d[28], o_1r1d[28]);
  OR2 I164 (complete1155_0n[29], o_1r0d[29], o_1r1d[29]);
  OR2 I165 (complete1155_0n[30], o_1r0d[30], o_1r1d[30]);
  OR2 I166 (complete1155_0n[31], o_1r0d[31], o_1r1d[31]);
  INV I167 (gate1154_0n, o_1a);
  C2RI I168 (o_1r1d[0], otint_1n[0], gate1154_0n, initialise);
  C2RI I169 (o_1r1d[1], otint_1n[1], gate1154_0n, initialise);
  C2RI I170 (o_1r1d[2], otint_1n[2], gate1154_0n, initialise);
  C2RI I171 (o_1r1d[3], otint_1n[3], gate1154_0n, initialise);
  C2RI I172 (o_1r1d[4], otint_1n[4], gate1154_0n, initialise);
  C2RI I173 (o_1r1d[5], otint_1n[5], gate1154_0n, initialise);
  C2RI I174 (o_1r1d[6], otint_1n[6], gate1154_0n, initialise);
  C2RI I175 (o_1r1d[7], otint_1n[7], gate1154_0n, initialise);
  C2RI I176 (o_1r1d[8], otint_1n[8], gate1154_0n, initialise);
  C2RI I177 (o_1r1d[9], otint_1n[9], gate1154_0n, initialise);
  C2RI I178 (o_1r1d[10], otint_1n[10], gate1154_0n, initialise);
  C2RI I179 (o_1r1d[11], otint_1n[11], gate1154_0n, initialise);
  C2RI I180 (o_1r1d[12], otint_1n[12], gate1154_0n, initialise);
  C2RI I181 (o_1r1d[13], otint_1n[13], gate1154_0n, initialise);
  C2RI I182 (o_1r1d[14], otint_1n[14], gate1154_0n, initialise);
  C2RI I183 (o_1r1d[15], otint_1n[15], gate1154_0n, initialise);
  C2RI I184 (o_1r1d[16], otint_1n[16], gate1154_0n, initialise);
  C2RI I185 (o_1r1d[17], otint_1n[17], gate1154_0n, initialise);
  C2RI I186 (o_1r1d[18], otint_1n[18], gate1154_0n, initialise);
  C2RI I187 (o_1r1d[19], otint_1n[19], gate1154_0n, initialise);
  C2RI I188 (o_1r1d[20], otint_1n[20], gate1154_0n, initialise);
  C2RI I189 (o_1r1d[21], otint_1n[21], gate1154_0n, initialise);
  C2RI I190 (o_1r1d[22], otint_1n[22], gate1154_0n, initialise);
  C2RI I191 (o_1r1d[23], otint_1n[23], gate1154_0n, initialise);
  C2RI I192 (o_1r1d[24], otint_1n[24], gate1154_0n, initialise);
  C2RI I193 (o_1r1d[25], otint_1n[25], gate1154_0n, initialise);
  C2RI I194 (o_1r1d[26], otint_1n[26], gate1154_0n, initialise);
  C2RI I195 (o_1r1d[27], otint_1n[27], gate1154_0n, initialise);
  C2RI I196 (o_1r1d[28], otint_1n[28], gate1154_0n, initialise);
  C2RI I197 (o_1r1d[29], otint_1n[29], gate1154_0n, initialise);
  C2RI I198 (o_1r1d[30], otint_1n[30], gate1154_0n, initialise);
  C2RI I199 (o_1r1d[31], otint_1n[31], gate1154_0n, initialise);
  C2RI I200 (o_1r0d[0], ofint_1n[0], gate1154_0n, initialise);
  C2RI I201 (o_1r0d[1], ofint_1n[1], gate1154_0n, initialise);
  C2RI I202 (o_1r0d[2], ofint_1n[2], gate1154_0n, initialise);
  C2RI I203 (o_1r0d[3], ofint_1n[3], gate1154_0n, initialise);
  C2RI I204 (o_1r0d[4], ofint_1n[4], gate1154_0n, initialise);
  C2RI I205 (o_1r0d[5], ofint_1n[5], gate1154_0n, initialise);
  C2RI I206 (o_1r0d[6], ofint_1n[6], gate1154_0n, initialise);
  C2RI I207 (o_1r0d[7], ofint_1n[7], gate1154_0n, initialise);
  C2RI I208 (o_1r0d[8], ofint_1n[8], gate1154_0n, initialise);
  C2RI I209 (o_1r0d[9], ofint_1n[9], gate1154_0n, initialise);
  C2RI I210 (o_1r0d[10], ofint_1n[10], gate1154_0n, initialise);
  C2RI I211 (o_1r0d[11], ofint_1n[11], gate1154_0n, initialise);
  C2RI I212 (o_1r0d[12], ofint_1n[12], gate1154_0n, initialise);
  C2RI I213 (o_1r0d[13], ofint_1n[13], gate1154_0n, initialise);
  C2RI I214 (o_1r0d[14], ofint_1n[14], gate1154_0n, initialise);
  C2RI I215 (o_1r0d[15], ofint_1n[15], gate1154_0n, initialise);
  C2RI I216 (o_1r0d[16], ofint_1n[16], gate1154_0n, initialise);
  C2RI I217 (o_1r0d[17], ofint_1n[17], gate1154_0n, initialise);
  C2RI I218 (o_1r0d[18], ofint_1n[18], gate1154_0n, initialise);
  C2RI I219 (o_1r0d[19], ofint_1n[19], gate1154_0n, initialise);
  C2RI I220 (o_1r0d[20], ofint_1n[20], gate1154_0n, initialise);
  C2RI I221 (o_1r0d[21], ofint_1n[21], gate1154_0n, initialise);
  C2RI I222 (o_1r0d[22], ofint_1n[22], gate1154_0n, initialise);
  C2RI I223 (o_1r0d[23], ofint_1n[23], gate1154_0n, initialise);
  C2RI I224 (o_1r0d[24], ofint_1n[24], gate1154_0n, initialise);
  C2RI I225 (o_1r0d[25], ofint_1n[25], gate1154_0n, initialise);
  C2RI I226 (o_1r0d[26], ofint_1n[26], gate1154_0n, initialise);
  C2RI I227 (o_1r0d[27], ofint_1n[27], gate1154_0n, initialise);
  C2RI I228 (o_1r0d[28], ofint_1n[28], gate1154_0n, initialise);
  C2RI I229 (o_1r0d[29], ofint_1n[29], gate1154_0n, initialise);
  C2RI I230 (o_1r0d[30], ofint_1n[30], gate1154_0n, initialise);
  C2RI I231 (o_1r0d[31], ofint_1n[31], gate1154_0n, initialise);
  C3 I232 (internal_0n[34], complete1151_0n[0], complete1151_0n[1], complete1151_0n[2]);
  C3 I233 (internal_0n[35], complete1151_0n[3], complete1151_0n[4], complete1151_0n[5]);
  C3 I234 (internal_0n[36], complete1151_0n[6], complete1151_0n[7], complete1151_0n[8]);
  C3 I235 (internal_0n[37], complete1151_0n[9], complete1151_0n[10], complete1151_0n[11]);
  C3 I236 (internal_0n[38], complete1151_0n[12], complete1151_0n[13], complete1151_0n[14]);
  C3 I237 (internal_0n[39], complete1151_0n[15], complete1151_0n[16], complete1151_0n[17]);
  C3 I238 (internal_0n[40], complete1151_0n[18], complete1151_0n[19], complete1151_0n[20]);
  C3 I239 (internal_0n[41], complete1151_0n[21], complete1151_0n[22], complete1151_0n[23]);
  C3 I240 (internal_0n[42], complete1151_0n[24], complete1151_0n[25], complete1151_0n[26]);
  C3 I241 (internal_0n[43], complete1151_0n[27], complete1151_0n[28], complete1151_0n[29]);
  C2 I242 (internal_0n[44], complete1151_0n[30], complete1151_0n[31]);
  C3 I243 (internal_0n[45], internal_0n[34], internal_0n[35], internal_0n[36]);
  C3 I244 (internal_0n[46], internal_0n[37], internal_0n[38], internal_0n[39]);
  C3 I245 (internal_0n[47], internal_0n[40], internal_0n[41], internal_0n[42]);
  C2 I246 (internal_0n[48], internal_0n[43], internal_0n[44]);
  C2 I247 (internal_0n[49], internal_0n[45], internal_0n[46]);
  C2 I248 (internal_0n[50], internal_0n[47], internal_0n[48]);
  C2 I249 (oaint_0n, internal_0n[49], internal_0n[50]);
  OR2 I250 (complete1151_0n[0], o_0r0d[0], o_0r1d[0]);
  OR2 I251 (complete1151_0n[1], o_0r0d[1], o_0r1d[1]);
  OR2 I252 (complete1151_0n[2], o_0r0d[2], o_0r1d[2]);
  OR2 I253 (complete1151_0n[3], o_0r0d[3], o_0r1d[3]);
  OR2 I254 (complete1151_0n[4], o_0r0d[4], o_0r1d[4]);
  OR2 I255 (complete1151_0n[5], o_0r0d[5], o_0r1d[5]);
  OR2 I256 (complete1151_0n[6], o_0r0d[6], o_0r1d[6]);
  OR2 I257 (complete1151_0n[7], o_0r0d[7], o_0r1d[7]);
  OR2 I258 (complete1151_0n[8], o_0r0d[8], o_0r1d[8]);
  OR2 I259 (complete1151_0n[9], o_0r0d[9], o_0r1d[9]);
  OR2 I260 (complete1151_0n[10], o_0r0d[10], o_0r1d[10]);
  OR2 I261 (complete1151_0n[11], o_0r0d[11], o_0r1d[11]);
  OR2 I262 (complete1151_0n[12], o_0r0d[12], o_0r1d[12]);
  OR2 I263 (complete1151_0n[13], o_0r0d[13], o_0r1d[13]);
  OR2 I264 (complete1151_0n[14], o_0r0d[14], o_0r1d[14]);
  OR2 I265 (complete1151_0n[15], o_0r0d[15], o_0r1d[15]);
  OR2 I266 (complete1151_0n[16], o_0r0d[16], o_0r1d[16]);
  OR2 I267 (complete1151_0n[17], o_0r0d[17], o_0r1d[17]);
  OR2 I268 (complete1151_0n[18], o_0r0d[18], o_0r1d[18]);
  OR2 I269 (complete1151_0n[19], o_0r0d[19], o_0r1d[19]);
  OR2 I270 (complete1151_0n[20], o_0r0d[20], o_0r1d[20]);
  OR2 I271 (complete1151_0n[21], o_0r0d[21], o_0r1d[21]);
  OR2 I272 (complete1151_0n[22], o_0r0d[22], o_0r1d[22]);
  OR2 I273 (complete1151_0n[23], o_0r0d[23], o_0r1d[23]);
  OR2 I274 (complete1151_0n[24], o_0r0d[24], o_0r1d[24]);
  OR2 I275 (complete1151_0n[25], o_0r0d[25], o_0r1d[25]);
  OR2 I276 (complete1151_0n[26], o_0r0d[26], o_0r1d[26]);
  OR2 I277 (complete1151_0n[27], o_0r0d[27], o_0r1d[27]);
  OR2 I278 (complete1151_0n[28], o_0r0d[28], o_0r1d[28]);
  OR2 I279 (complete1151_0n[29], o_0r0d[29], o_0r1d[29]);
  OR2 I280 (complete1151_0n[30], o_0r0d[30], o_0r1d[30]);
  OR2 I281 (complete1151_0n[31], o_0r0d[31], o_0r1d[31]);
  INV I282 (gate1150_0n, o_0a);
  C2RI I283 (o_0r1d[0], otint_0n[0], gate1150_0n, initialise);
  C2RI I284 (o_0r1d[1], otint_0n[1], gate1150_0n, initialise);
  C2RI I285 (o_0r1d[2], otint_0n[2], gate1150_0n, initialise);
  C2RI I286 (o_0r1d[3], otint_0n[3], gate1150_0n, initialise);
  C2RI I287 (o_0r1d[4], otint_0n[4], gate1150_0n, initialise);
  C2RI I288 (o_0r1d[5], otint_0n[5], gate1150_0n, initialise);
  C2RI I289 (o_0r1d[6], otint_0n[6], gate1150_0n, initialise);
  C2RI I290 (o_0r1d[7], otint_0n[7], gate1150_0n, initialise);
  C2RI I291 (o_0r1d[8], otint_0n[8], gate1150_0n, initialise);
  C2RI I292 (o_0r1d[9], otint_0n[9], gate1150_0n, initialise);
  C2RI I293 (o_0r1d[10], otint_0n[10], gate1150_0n, initialise);
  C2RI I294 (o_0r1d[11], otint_0n[11], gate1150_0n, initialise);
  C2RI I295 (o_0r1d[12], otint_0n[12], gate1150_0n, initialise);
  C2RI I296 (o_0r1d[13], otint_0n[13], gate1150_0n, initialise);
  C2RI I297 (o_0r1d[14], otint_0n[14], gate1150_0n, initialise);
  C2RI I298 (o_0r1d[15], otint_0n[15], gate1150_0n, initialise);
  C2RI I299 (o_0r1d[16], otint_0n[16], gate1150_0n, initialise);
  C2RI I300 (o_0r1d[17], otint_0n[17], gate1150_0n, initialise);
  C2RI I301 (o_0r1d[18], otint_0n[18], gate1150_0n, initialise);
  C2RI I302 (o_0r1d[19], otint_0n[19], gate1150_0n, initialise);
  C2RI I303 (o_0r1d[20], otint_0n[20], gate1150_0n, initialise);
  C2RI I304 (o_0r1d[21], otint_0n[21], gate1150_0n, initialise);
  C2RI I305 (o_0r1d[22], otint_0n[22], gate1150_0n, initialise);
  C2RI I306 (o_0r1d[23], otint_0n[23], gate1150_0n, initialise);
  C2RI I307 (o_0r1d[24], otint_0n[24], gate1150_0n, initialise);
  C2RI I308 (o_0r1d[25], otint_0n[25], gate1150_0n, initialise);
  C2RI I309 (o_0r1d[26], otint_0n[26], gate1150_0n, initialise);
  C2RI I310 (o_0r1d[27], otint_0n[27], gate1150_0n, initialise);
  C2RI I311 (o_0r1d[28], otint_0n[28], gate1150_0n, initialise);
  C2RI I312 (o_0r1d[29], otint_0n[29], gate1150_0n, initialise);
  C2RI I313 (o_0r1d[30], otint_0n[30], gate1150_0n, initialise);
  C2RI I314 (o_0r1d[31], otint_0n[31], gate1150_0n, initialise);
  C2RI I315 (o_0r0d[0], ofint_0n[0], gate1150_0n, initialise);
  C2RI I316 (o_0r0d[1], ofint_0n[1], gate1150_0n, initialise);
  C2RI I317 (o_0r0d[2], ofint_0n[2], gate1150_0n, initialise);
  C2RI I318 (o_0r0d[3], ofint_0n[3], gate1150_0n, initialise);
  C2RI I319 (o_0r0d[4], ofint_0n[4], gate1150_0n, initialise);
  C2RI I320 (o_0r0d[5], ofint_0n[5], gate1150_0n, initialise);
  C2RI I321 (o_0r0d[6], ofint_0n[6], gate1150_0n, initialise);
  C2RI I322 (o_0r0d[7], ofint_0n[7], gate1150_0n, initialise);
  C2RI I323 (o_0r0d[8], ofint_0n[8], gate1150_0n, initialise);
  C2RI I324 (o_0r0d[9], ofint_0n[9], gate1150_0n, initialise);
  C2RI I325 (o_0r0d[10], ofint_0n[10], gate1150_0n, initialise);
  C2RI I326 (o_0r0d[11], ofint_0n[11], gate1150_0n, initialise);
  C2RI I327 (o_0r0d[12], ofint_0n[12], gate1150_0n, initialise);
  C2RI I328 (o_0r0d[13], ofint_0n[13], gate1150_0n, initialise);
  C2RI I329 (o_0r0d[14], ofint_0n[14], gate1150_0n, initialise);
  C2RI I330 (o_0r0d[15], ofint_0n[15], gate1150_0n, initialise);
  C2RI I331 (o_0r0d[16], ofint_0n[16], gate1150_0n, initialise);
  C2RI I332 (o_0r0d[17], ofint_0n[17], gate1150_0n, initialise);
  C2RI I333 (o_0r0d[18], ofint_0n[18], gate1150_0n, initialise);
  C2RI I334 (o_0r0d[19], ofint_0n[19], gate1150_0n, initialise);
  C2RI I335 (o_0r0d[20], ofint_0n[20], gate1150_0n, initialise);
  C2RI I336 (o_0r0d[21], ofint_0n[21], gate1150_0n, initialise);
  C2RI I337 (o_0r0d[22], ofint_0n[22], gate1150_0n, initialise);
  C2RI I338 (o_0r0d[23], ofint_0n[23], gate1150_0n, initialise);
  C2RI I339 (o_0r0d[24], ofint_0n[24], gate1150_0n, initialise);
  C2RI I340 (o_0r0d[25], ofint_0n[25], gate1150_0n, initialise);
  C2RI I341 (o_0r0d[26], ofint_0n[26], gate1150_0n, initialise);
  C2RI I342 (o_0r0d[27], ofint_0n[27], gate1150_0n, initialise);
  C2RI I343 (o_0r0d[28], ofint_0n[28], gate1150_0n, initialise);
  C2RI I344 (o_0r0d[29], ofint_0n[29], gate1150_0n, initialise);
  C2RI I345 (o_0r0d[30], ofint_0n[30], gate1150_0n, initialise);
  C2RI I346 (o_0r0d[31], ofint_0n[31], gate1150_0n, initialise);
  C3 I347 (internal_0n[51], complete1147_0n[0], complete1147_0n[1], complete1147_0n[2]);
  C3 I348 (internal_0n[52], complete1147_0n[3], complete1147_0n[4], complete1147_0n[5]);
  C3 I349 (internal_0n[53], complete1147_0n[6], complete1147_0n[7], complete1147_0n[8]);
  C3 I350 (internal_0n[54], complete1147_0n[9], complete1147_0n[10], complete1147_0n[11]);
  C3 I351 (internal_0n[55], complete1147_0n[12], complete1147_0n[13], complete1147_0n[14]);
  C3 I352 (internal_0n[56], complete1147_0n[15], complete1147_0n[16], complete1147_0n[17]);
  C3 I353 (internal_0n[57], complete1147_0n[18], complete1147_0n[19], complete1147_0n[20]);
  C3 I354 (internal_0n[58], complete1147_0n[21], complete1147_0n[22], complete1147_0n[23]);
  C3 I355 (internal_0n[59], complete1147_0n[24], complete1147_0n[25], complete1147_0n[26]);
  C3 I356 (internal_0n[60], complete1147_0n[27], complete1147_0n[28], complete1147_0n[29]);
  C3 I357 (internal_0n[61], complete1147_0n[30], complete1147_0n[31], complete1147_0n[32]);
  C2 I358 (internal_0n[62], complete1147_0n[33], complete1147_0n[34]);
  C3 I359 (internal_0n[63], internal_0n[51], internal_0n[52], internal_0n[53]);
  C3 I360 (internal_0n[64], internal_0n[54], internal_0n[55], internal_0n[56]);
  C3 I361 (internal_0n[65], internal_0n[57], internal_0n[58], internal_0n[59]);
  C3 I362 (internal_0n[66], internal_0n[60], internal_0n[61], internal_0n[62]);
  C2 I363 (internal_0n[67], internal_0n[63], internal_0n[64]);
  C2 I364 (internal_0n[68], internal_0n[65], internal_0n[66]);
  C2 I365 (i_0a, internal_0n[67], internal_0n[68]);
  OR2 I366 (complete1147_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I367 (complete1147_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I368 (complete1147_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I369 (complete1147_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I370 (complete1147_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I371 (complete1147_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I372 (complete1147_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I373 (complete1147_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I374 (complete1147_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I375 (complete1147_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I376 (complete1147_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I377 (complete1147_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I378 (complete1147_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I379 (complete1147_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I380 (complete1147_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I381 (complete1147_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I382 (complete1147_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I383 (complete1147_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I384 (complete1147_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I385 (complete1147_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I386 (complete1147_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I387 (complete1147_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I388 (complete1147_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I389 (complete1147_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I390 (complete1147_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I391 (complete1147_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I392 (complete1147_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I393 (complete1147_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I394 (complete1147_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I395 (complete1147_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I396 (complete1147_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I397 (complete1147_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I398 (complete1147_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I399 (complete1147_0n[33], ifint_0n[33], itint_0n[33]);
  OR2 I400 (complete1147_0n[34], ifint_0n[34], itint_0n[34]);
  INV I401 (gate1146_0n, iaint_0n);
  C2RI I402 (itint_0n[0], i_0r1d[0], gate1146_0n, initialise);
  C2RI I403 (itint_0n[1], i_0r1d[1], gate1146_0n, initialise);
  C2RI I404 (itint_0n[2], i_0r1d[2], gate1146_0n, initialise);
  C2RI I405 (itint_0n[3], i_0r1d[3], gate1146_0n, initialise);
  C2RI I406 (itint_0n[4], i_0r1d[4], gate1146_0n, initialise);
  C2RI I407 (itint_0n[5], i_0r1d[5], gate1146_0n, initialise);
  C2RI I408 (itint_0n[6], i_0r1d[6], gate1146_0n, initialise);
  C2RI I409 (itint_0n[7], i_0r1d[7], gate1146_0n, initialise);
  C2RI I410 (itint_0n[8], i_0r1d[8], gate1146_0n, initialise);
  C2RI I411 (itint_0n[9], i_0r1d[9], gate1146_0n, initialise);
  C2RI I412 (itint_0n[10], i_0r1d[10], gate1146_0n, initialise);
  C2RI I413 (itint_0n[11], i_0r1d[11], gate1146_0n, initialise);
  C2RI I414 (itint_0n[12], i_0r1d[12], gate1146_0n, initialise);
  C2RI I415 (itint_0n[13], i_0r1d[13], gate1146_0n, initialise);
  C2RI I416 (itint_0n[14], i_0r1d[14], gate1146_0n, initialise);
  C2RI I417 (itint_0n[15], i_0r1d[15], gate1146_0n, initialise);
  C2RI I418 (itint_0n[16], i_0r1d[16], gate1146_0n, initialise);
  C2RI I419 (itint_0n[17], i_0r1d[17], gate1146_0n, initialise);
  C2RI I420 (itint_0n[18], i_0r1d[18], gate1146_0n, initialise);
  C2RI I421 (itint_0n[19], i_0r1d[19], gate1146_0n, initialise);
  C2RI I422 (itint_0n[20], i_0r1d[20], gate1146_0n, initialise);
  C2RI I423 (itint_0n[21], i_0r1d[21], gate1146_0n, initialise);
  C2RI I424 (itint_0n[22], i_0r1d[22], gate1146_0n, initialise);
  C2RI I425 (itint_0n[23], i_0r1d[23], gate1146_0n, initialise);
  C2RI I426 (itint_0n[24], i_0r1d[24], gate1146_0n, initialise);
  C2RI I427 (itint_0n[25], i_0r1d[25], gate1146_0n, initialise);
  C2RI I428 (itint_0n[26], i_0r1d[26], gate1146_0n, initialise);
  C2RI I429 (itint_0n[27], i_0r1d[27], gate1146_0n, initialise);
  C2RI I430 (itint_0n[28], i_0r1d[28], gate1146_0n, initialise);
  C2RI I431 (itint_0n[29], i_0r1d[29], gate1146_0n, initialise);
  C2RI I432 (itint_0n[30], i_0r1d[30], gate1146_0n, initialise);
  C2RI I433 (itint_0n[31], i_0r1d[31], gate1146_0n, initialise);
  C2RI I434 (itint_0n[32], i_0r1d[32], gate1146_0n, initialise);
  C2RI I435 (itint_0n[33], i_0r1d[33], gate1146_0n, initialise);
  C2RI I436 (itint_0n[34], i_0r1d[34], gate1146_0n, initialise);
  C2RI I437 (ifint_0n[0], i_0r0d[0], gate1146_0n, initialise);
  C2RI I438 (ifint_0n[1], i_0r0d[1], gate1146_0n, initialise);
  C2RI I439 (ifint_0n[2], i_0r0d[2], gate1146_0n, initialise);
  C2RI I440 (ifint_0n[3], i_0r0d[3], gate1146_0n, initialise);
  C2RI I441 (ifint_0n[4], i_0r0d[4], gate1146_0n, initialise);
  C2RI I442 (ifint_0n[5], i_0r0d[5], gate1146_0n, initialise);
  C2RI I443 (ifint_0n[6], i_0r0d[6], gate1146_0n, initialise);
  C2RI I444 (ifint_0n[7], i_0r0d[7], gate1146_0n, initialise);
  C2RI I445 (ifint_0n[8], i_0r0d[8], gate1146_0n, initialise);
  C2RI I446 (ifint_0n[9], i_0r0d[9], gate1146_0n, initialise);
  C2RI I447 (ifint_0n[10], i_0r0d[10], gate1146_0n, initialise);
  C2RI I448 (ifint_0n[11], i_0r0d[11], gate1146_0n, initialise);
  C2RI I449 (ifint_0n[12], i_0r0d[12], gate1146_0n, initialise);
  C2RI I450 (ifint_0n[13], i_0r0d[13], gate1146_0n, initialise);
  C2RI I451 (ifint_0n[14], i_0r0d[14], gate1146_0n, initialise);
  C2RI I452 (ifint_0n[15], i_0r0d[15], gate1146_0n, initialise);
  C2RI I453 (ifint_0n[16], i_0r0d[16], gate1146_0n, initialise);
  C2RI I454 (ifint_0n[17], i_0r0d[17], gate1146_0n, initialise);
  C2RI I455 (ifint_0n[18], i_0r0d[18], gate1146_0n, initialise);
  C2RI I456 (ifint_0n[19], i_0r0d[19], gate1146_0n, initialise);
  C2RI I457 (ifint_0n[20], i_0r0d[20], gate1146_0n, initialise);
  C2RI I458 (ifint_0n[21], i_0r0d[21], gate1146_0n, initialise);
  C2RI I459 (ifint_0n[22], i_0r0d[22], gate1146_0n, initialise);
  C2RI I460 (ifint_0n[23], i_0r0d[23], gate1146_0n, initialise);
  C2RI I461 (ifint_0n[24], i_0r0d[24], gate1146_0n, initialise);
  C2RI I462 (ifint_0n[25], i_0r0d[25], gate1146_0n, initialise);
  C2RI I463 (ifint_0n[26], i_0r0d[26], gate1146_0n, initialise);
  C2RI I464 (ifint_0n[27], i_0r0d[27], gate1146_0n, initialise);
  C2RI I465 (ifint_0n[28], i_0r0d[28], gate1146_0n, initialise);
  C2RI I466 (ifint_0n[29], i_0r0d[29], gate1146_0n, initialise);
  C2RI I467 (ifint_0n[30], i_0r0d[30], gate1146_0n, initialise);
  C2RI I468 (ifint_0n[31], i_0r0d[31], gate1146_0n, initialise);
  C2RI I469 (ifint_0n[32], i_0r0d[32], gate1146_0n, initialise);
  C2RI I470 (ifint_0n[33], i_0r0d[33], gate1146_0n, initialise);
  C2RI I471 (ifint_0n[34], i_0r0d[34], gate1146_0n, initialise);
  C2 I472 (otint_2n[0], sel_2n, itint_0n[0]);
  C2 I473 (otint_2n[1], sel_2n, itint_0n[1]);
  C2 I474 (otint_2n[2], sel_2n, itint_0n[2]);
  C2 I475 (otint_2n[3], sel_2n, itint_0n[3]);
  C2 I476 (otint_2n[4], sel_2n, itint_0n[4]);
  C2 I477 (otint_2n[5], sel_2n, itint_0n[5]);
  C2 I478 (otint_2n[6], sel_2n, itint_0n[6]);
  C2 I479 (otint_2n[7], sel_2n, itint_0n[7]);
  C2 I480 (otint_2n[8], sel_2n, itint_0n[8]);
  C2 I481 (otint_2n[9], sel_2n, itint_0n[9]);
  C2 I482 (otint_2n[10], sel_2n, itint_0n[10]);
  C2 I483 (otint_2n[11], sel_2n, itint_0n[11]);
  C2 I484 (otint_2n[12], sel_2n, itint_0n[12]);
  C2 I485 (otint_2n[13], sel_2n, itint_0n[13]);
  C2 I486 (otint_2n[14], sel_2n, itint_0n[14]);
  C2 I487 (otint_2n[15], sel_2n, itint_0n[15]);
  C2 I488 (otint_2n[16], sel_2n, itint_0n[16]);
  C2 I489 (otint_2n[17], sel_2n, itint_0n[17]);
  C2 I490 (otint_2n[18], sel_2n, itint_0n[18]);
  C2 I491 (otint_2n[19], sel_2n, itint_0n[19]);
  C2 I492 (otint_2n[20], sel_2n, itint_0n[20]);
  C2 I493 (otint_2n[21], sel_2n, itint_0n[21]);
  C2 I494 (otint_2n[22], sel_2n, itint_0n[22]);
  C2 I495 (otint_2n[23], sel_2n, itint_0n[23]);
  C2 I496 (otint_2n[24], sel_2n, itint_0n[24]);
  C2 I497 (otint_2n[25], sel_2n, itint_0n[25]);
  C2 I498 (otint_2n[26], sel_2n, itint_0n[26]);
  C2 I499 (otint_2n[27], sel_2n, itint_0n[27]);
  C2 I500 (otint_2n[28], sel_2n, itint_0n[28]);
  C2 I501 (otint_2n[29], sel_2n, itint_0n[29]);
  C2 I502 (otint_2n[30], sel_2n, itint_0n[30]);
  C2 I503 (otint_2n[31], sel_2n, itint_0n[31]);
  C2 I504 (otint_1n[0], sel_1n, itint_0n[0]);
  C2 I505 (otint_1n[1], sel_1n, itint_0n[1]);
  C2 I506 (otint_1n[2], sel_1n, itint_0n[2]);
  C2 I507 (otint_1n[3], sel_1n, itint_0n[3]);
  C2 I508 (otint_1n[4], sel_1n, itint_0n[4]);
  C2 I509 (otint_1n[5], sel_1n, itint_0n[5]);
  C2 I510 (otint_1n[6], sel_1n, itint_0n[6]);
  C2 I511 (otint_1n[7], sel_1n, itint_0n[7]);
  C2 I512 (otint_1n[8], sel_1n, itint_0n[8]);
  C2 I513 (otint_1n[9], sel_1n, itint_0n[9]);
  C2 I514 (otint_1n[10], sel_1n, itint_0n[10]);
  C2 I515 (otint_1n[11], sel_1n, itint_0n[11]);
  C2 I516 (otint_1n[12], sel_1n, itint_0n[12]);
  C2 I517 (otint_1n[13], sel_1n, itint_0n[13]);
  C2 I518 (otint_1n[14], sel_1n, itint_0n[14]);
  C2 I519 (otint_1n[15], sel_1n, itint_0n[15]);
  C2 I520 (otint_1n[16], sel_1n, itint_0n[16]);
  C2 I521 (otint_1n[17], sel_1n, itint_0n[17]);
  C2 I522 (otint_1n[18], sel_1n, itint_0n[18]);
  C2 I523 (otint_1n[19], sel_1n, itint_0n[19]);
  C2 I524 (otint_1n[20], sel_1n, itint_0n[20]);
  C2 I525 (otint_1n[21], sel_1n, itint_0n[21]);
  C2 I526 (otint_1n[22], sel_1n, itint_0n[22]);
  C2 I527 (otint_1n[23], sel_1n, itint_0n[23]);
  C2 I528 (otint_1n[24], sel_1n, itint_0n[24]);
  C2 I529 (otint_1n[25], sel_1n, itint_0n[25]);
  C2 I530 (otint_1n[26], sel_1n, itint_0n[26]);
  C2 I531 (otint_1n[27], sel_1n, itint_0n[27]);
  C2 I532 (otint_1n[28], sel_1n, itint_0n[28]);
  C2 I533 (otint_1n[29], sel_1n, itint_0n[29]);
  C2 I534 (otint_1n[30], sel_1n, itint_0n[30]);
  C2 I535 (otint_1n[31], sel_1n, itint_0n[31]);
  C2 I536 (otint_0n[0], sel_0n, itint_0n[0]);
  C2 I537 (otint_0n[1], sel_0n, itint_0n[1]);
  C2 I538 (otint_0n[2], sel_0n, itint_0n[2]);
  C2 I539 (otint_0n[3], sel_0n, itint_0n[3]);
  C2 I540 (otint_0n[4], sel_0n, itint_0n[4]);
  C2 I541 (otint_0n[5], sel_0n, itint_0n[5]);
  C2 I542 (otint_0n[6], sel_0n, itint_0n[6]);
  C2 I543 (otint_0n[7], sel_0n, itint_0n[7]);
  C2 I544 (otint_0n[8], sel_0n, itint_0n[8]);
  C2 I545 (otint_0n[9], sel_0n, itint_0n[9]);
  C2 I546 (otint_0n[10], sel_0n, itint_0n[10]);
  C2 I547 (otint_0n[11], sel_0n, itint_0n[11]);
  C2 I548 (otint_0n[12], sel_0n, itint_0n[12]);
  C2 I549 (otint_0n[13], sel_0n, itint_0n[13]);
  C2 I550 (otint_0n[14], sel_0n, itint_0n[14]);
  C2 I551 (otint_0n[15], sel_0n, itint_0n[15]);
  C2 I552 (otint_0n[16], sel_0n, itint_0n[16]);
  C2 I553 (otint_0n[17], sel_0n, itint_0n[17]);
  C2 I554 (otint_0n[18], sel_0n, itint_0n[18]);
  C2 I555 (otint_0n[19], sel_0n, itint_0n[19]);
  C2 I556 (otint_0n[20], sel_0n, itint_0n[20]);
  C2 I557 (otint_0n[21], sel_0n, itint_0n[21]);
  C2 I558 (otint_0n[22], sel_0n, itint_0n[22]);
  C2 I559 (otint_0n[23], sel_0n, itint_0n[23]);
  C2 I560 (otint_0n[24], sel_0n, itint_0n[24]);
  C2 I561 (otint_0n[25], sel_0n, itint_0n[25]);
  C2 I562 (otint_0n[26], sel_0n, itint_0n[26]);
  C2 I563 (otint_0n[27], sel_0n, itint_0n[27]);
  C2 I564 (otint_0n[28], sel_0n, itint_0n[28]);
  C2 I565 (otint_0n[29], sel_0n, itint_0n[29]);
  C2 I566 (otint_0n[30], sel_0n, itint_0n[30]);
  C2 I567 (otint_0n[31], sel_0n, itint_0n[31]);
  C2 I568 (ofint_2n[0], sel_2n, ifint_0n[0]);
  C2 I569 (ofint_2n[1], sel_2n, ifint_0n[1]);
  C2 I570 (ofint_2n[2], sel_2n, ifint_0n[2]);
  C2 I571 (ofint_2n[3], sel_2n, ifint_0n[3]);
  C2 I572 (ofint_2n[4], sel_2n, ifint_0n[4]);
  C2 I573 (ofint_2n[5], sel_2n, ifint_0n[5]);
  C2 I574 (ofint_2n[6], sel_2n, ifint_0n[6]);
  C2 I575 (ofint_2n[7], sel_2n, ifint_0n[7]);
  C2 I576 (ofint_2n[8], sel_2n, ifint_0n[8]);
  C2 I577 (ofint_2n[9], sel_2n, ifint_0n[9]);
  C2 I578 (ofint_2n[10], sel_2n, ifint_0n[10]);
  C2 I579 (ofint_2n[11], sel_2n, ifint_0n[11]);
  C2 I580 (ofint_2n[12], sel_2n, ifint_0n[12]);
  C2 I581 (ofint_2n[13], sel_2n, ifint_0n[13]);
  C2 I582 (ofint_2n[14], sel_2n, ifint_0n[14]);
  C2 I583 (ofint_2n[15], sel_2n, ifint_0n[15]);
  C2 I584 (ofint_2n[16], sel_2n, ifint_0n[16]);
  C2 I585 (ofint_2n[17], sel_2n, ifint_0n[17]);
  C2 I586 (ofint_2n[18], sel_2n, ifint_0n[18]);
  C2 I587 (ofint_2n[19], sel_2n, ifint_0n[19]);
  C2 I588 (ofint_2n[20], sel_2n, ifint_0n[20]);
  C2 I589 (ofint_2n[21], sel_2n, ifint_0n[21]);
  C2 I590 (ofint_2n[22], sel_2n, ifint_0n[22]);
  C2 I591 (ofint_2n[23], sel_2n, ifint_0n[23]);
  C2 I592 (ofint_2n[24], sel_2n, ifint_0n[24]);
  C2 I593 (ofint_2n[25], sel_2n, ifint_0n[25]);
  C2 I594 (ofint_2n[26], sel_2n, ifint_0n[26]);
  C2 I595 (ofint_2n[27], sel_2n, ifint_0n[27]);
  C2 I596 (ofint_2n[28], sel_2n, ifint_0n[28]);
  C2 I597 (ofint_2n[29], sel_2n, ifint_0n[29]);
  C2 I598 (ofint_2n[30], sel_2n, ifint_0n[30]);
  C2 I599 (ofint_2n[31], sel_2n, ifint_0n[31]);
  C2 I600 (ofint_1n[0], sel_1n, ifint_0n[0]);
  C2 I601 (ofint_1n[1], sel_1n, ifint_0n[1]);
  C2 I602 (ofint_1n[2], sel_1n, ifint_0n[2]);
  C2 I603 (ofint_1n[3], sel_1n, ifint_0n[3]);
  C2 I604 (ofint_1n[4], sel_1n, ifint_0n[4]);
  C2 I605 (ofint_1n[5], sel_1n, ifint_0n[5]);
  C2 I606 (ofint_1n[6], sel_1n, ifint_0n[6]);
  C2 I607 (ofint_1n[7], sel_1n, ifint_0n[7]);
  C2 I608 (ofint_1n[8], sel_1n, ifint_0n[8]);
  C2 I609 (ofint_1n[9], sel_1n, ifint_0n[9]);
  C2 I610 (ofint_1n[10], sel_1n, ifint_0n[10]);
  C2 I611 (ofint_1n[11], sel_1n, ifint_0n[11]);
  C2 I612 (ofint_1n[12], sel_1n, ifint_0n[12]);
  C2 I613 (ofint_1n[13], sel_1n, ifint_0n[13]);
  C2 I614 (ofint_1n[14], sel_1n, ifint_0n[14]);
  C2 I615 (ofint_1n[15], sel_1n, ifint_0n[15]);
  C2 I616 (ofint_1n[16], sel_1n, ifint_0n[16]);
  C2 I617 (ofint_1n[17], sel_1n, ifint_0n[17]);
  C2 I618 (ofint_1n[18], sel_1n, ifint_0n[18]);
  C2 I619 (ofint_1n[19], sel_1n, ifint_0n[19]);
  C2 I620 (ofint_1n[20], sel_1n, ifint_0n[20]);
  C2 I621 (ofint_1n[21], sel_1n, ifint_0n[21]);
  C2 I622 (ofint_1n[22], sel_1n, ifint_0n[22]);
  C2 I623 (ofint_1n[23], sel_1n, ifint_0n[23]);
  C2 I624 (ofint_1n[24], sel_1n, ifint_0n[24]);
  C2 I625 (ofint_1n[25], sel_1n, ifint_0n[25]);
  C2 I626 (ofint_1n[26], sel_1n, ifint_0n[26]);
  C2 I627 (ofint_1n[27], sel_1n, ifint_0n[27]);
  C2 I628 (ofint_1n[28], sel_1n, ifint_0n[28]);
  C2 I629 (ofint_1n[29], sel_1n, ifint_0n[29]);
  C2 I630 (ofint_1n[30], sel_1n, ifint_0n[30]);
  C2 I631 (ofint_1n[31], sel_1n, ifint_0n[31]);
  C2 I632 (ofint_0n[0], sel_0n, ifint_0n[0]);
  C2 I633 (ofint_0n[1], sel_0n, ifint_0n[1]);
  C2 I634 (ofint_0n[2], sel_0n, ifint_0n[2]);
  C2 I635 (ofint_0n[3], sel_0n, ifint_0n[3]);
  C2 I636 (ofint_0n[4], sel_0n, ifint_0n[4]);
  C2 I637 (ofint_0n[5], sel_0n, ifint_0n[5]);
  C2 I638 (ofint_0n[6], sel_0n, ifint_0n[6]);
  C2 I639 (ofint_0n[7], sel_0n, ifint_0n[7]);
  C2 I640 (ofint_0n[8], sel_0n, ifint_0n[8]);
  C2 I641 (ofint_0n[9], sel_0n, ifint_0n[9]);
  C2 I642 (ofint_0n[10], sel_0n, ifint_0n[10]);
  C2 I643 (ofint_0n[11], sel_0n, ifint_0n[11]);
  C2 I644 (ofint_0n[12], sel_0n, ifint_0n[12]);
  C2 I645 (ofint_0n[13], sel_0n, ifint_0n[13]);
  C2 I646 (ofint_0n[14], sel_0n, ifint_0n[14]);
  C2 I647 (ofint_0n[15], sel_0n, ifint_0n[15]);
  C2 I648 (ofint_0n[16], sel_0n, ifint_0n[16]);
  C2 I649 (ofint_0n[17], sel_0n, ifint_0n[17]);
  C2 I650 (ofint_0n[18], sel_0n, ifint_0n[18]);
  C2 I651 (ofint_0n[19], sel_0n, ifint_0n[19]);
  C2 I652 (ofint_0n[20], sel_0n, ifint_0n[20]);
  C2 I653 (ofint_0n[21], sel_0n, ifint_0n[21]);
  C2 I654 (ofint_0n[22], sel_0n, ifint_0n[22]);
  C2 I655 (ofint_0n[23], sel_0n, ifint_0n[23]);
  C2 I656 (ofint_0n[24], sel_0n, ifint_0n[24]);
  C2 I657 (ofint_0n[25], sel_0n, ifint_0n[25]);
  C2 I658 (ofint_0n[26], sel_0n, ifint_0n[26]);
  C2 I659 (ofint_0n[27], sel_0n, ifint_0n[27]);
  C2 I660 (ofint_0n[28], sel_0n, ifint_0n[28]);
  C2 I661 (ofint_0n[29], sel_0n, ifint_0n[29]);
  C2 I662 (ofint_0n[30], sel_0n, ifint_0n[30]);
  C2 I663 (ofint_0n[31], sel_0n, ifint_0n[31]);
  C3 I664 (internal_0n[69], complete1143_0n[0], complete1143_0n[1], complete1143_0n[2]);
  C3 I665 (internal_0n[70], complete1143_0n[3], complete1143_0n[4], complete1143_0n[5]);
  C3 I666 (internal_0n[71], complete1143_0n[6], complete1143_0n[7], complete1143_0n[8]);
  C3 I667 (internal_0n[72], complete1143_0n[9], complete1143_0n[10], complete1143_0n[11]);
  C3 I668 (internal_0n[73], complete1143_0n[12], complete1143_0n[13], complete1143_0n[14]);
  C3 I669 (internal_0n[74], complete1143_0n[15], complete1143_0n[16], complete1143_0n[17]);
  C3 I670 (internal_0n[75], complete1143_0n[18], complete1143_0n[19], complete1143_0n[20]);
  C3 I671 (internal_0n[76], complete1143_0n[21], complete1143_0n[22], complete1143_0n[23]);
  C3 I672 (internal_0n[77], complete1143_0n[24], complete1143_0n[25], complete1143_0n[26]);
  C3 I673 (internal_0n[78], complete1143_0n[27], complete1143_0n[28], complete1143_0n[29]);
  C3 I674 (internal_0n[79], complete1143_0n[30], complete1143_0n[31], complete1143_0n[32]);
  C2 I675 (internal_0n[80], complete1143_0n[33], complete1143_0n[34]);
  C3 I676 (internal_0n[81], internal_0n[69], internal_0n[70], internal_0n[71]);
  C3 I677 (internal_0n[82], internal_0n[72], internal_0n[73], internal_0n[74]);
  C3 I678 (internal_0n[83], internal_0n[75], internal_0n[76], internal_0n[77]);
  C3 I679 (internal_0n[84], internal_0n[78], internal_0n[79], internal_0n[80]);
  C2 I680 (internal_0n[85], internal_0n[81], internal_0n[82]);
  C2 I681 (internal_0n[86], internal_0n[83], internal_0n[84]);
  C2 I682 (icomplete_0n, internal_0n[85], internal_0n[86]);
  OR2 I683 (complete1143_0n[0], ifint_0n[0], itint_0n[0]);
  OR2 I684 (complete1143_0n[1], ifint_0n[1], itint_0n[1]);
  OR2 I685 (complete1143_0n[2], ifint_0n[2], itint_0n[2]);
  OR2 I686 (complete1143_0n[3], ifint_0n[3], itint_0n[3]);
  OR2 I687 (complete1143_0n[4], ifint_0n[4], itint_0n[4]);
  OR2 I688 (complete1143_0n[5], ifint_0n[5], itint_0n[5]);
  OR2 I689 (complete1143_0n[6], ifint_0n[6], itint_0n[6]);
  OR2 I690 (complete1143_0n[7], ifint_0n[7], itint_0n[7]);
  OR2 I691 (complete1143_0n[8], ifint_0n[8], itint_0n[8]);
  OR2 I692 (complete1143_0n[9], ifint_0n[9], itint_0n[9]);
  OR2 I693 (complete1143_0n[10], ifint_0n[10], itint_0n[10]);
  OR2 I694 (complete1143_0n[11], ifint_0n[11], itint_0n[11]);
  OR2 I695 (complete1143_0n[12], ifint_0n[12], itint_0n[12]);
  OR2 I696 (complete1143_0n[13], ifint_0n[13], itint_0n[13]);
  OR2 I697 (complete1143_0n[14], ifint_0n[14], itint_0n[14]);
  OR2 I698 (complete1143_0n[15], ifint_0n[15], itint_0n[15]);
  OR2 I699 (complete1143_0n[16], ifint_0n[16], itint_0n[16]);
  OR2 I700 (complete1143_0n[17], ifint_0n[17], itint_0n[17]);
  OR2 I701 (complete1143_0n[18], ifint_0n[18], itint_0n[18]);
  OR2 I702 (complete1143_0n[19], ifint_0n[19], itint_0n[19]);
  OR2 I703 (complete1143_0n[20], ifint_0n[20], itint_0n[20]);
  OR2 I704 (complete1143_0n[21], ifint_0n[21], itint_0n[21]);
  OR2 I705 (complete1143_0n[22], ifint_0n[22], itint_0n[22]);
  OR2 I706 (complete1143_0n[23], ifint_0n[23], itint_0n[23]);
  OR2 I707 (complete1143_0n[24], ifint_0n[24], itint_0n[24]);
  OR2 I708 (complete1143_0n[25], ifint_0n[25], itint_0n[25]);
  OR2 I709 (complete1143_0n[26], ifint_0n[26], itint_0n[26]);
  OR2 I710 (complete1143_0n[27], ifint_0n[27], itint_0n[27]);
  OR2 I711 (complete1143_0n[28], ifint_0n[28], itint_0n[28]);
  OR2 I712 (complete1143_0n[29], ifint_0n[29], itint_0n[29]);
  OR2 I713 (complete1143_0n[30], ifint_0n[30], itint_0n[30]);
  OR2 I714 (complete1143_0n[31], ifint_0n[31], itint_0n[31]);
  OR2 I715 (complete1143_0n[32], ifint_0n[32], itint_0n[32]);
  OR2 I716 (complete1143_0n[33], ifint_0n[33], itint_0n[33]);
  OR2 I717 (complete1143_0n[34], ifint_0n[34], itint_0n[34]);
  C3 I718 (matchi_2n, ifint_0n[33], ifint_0n[32], itint_0n[34]);
  assign sel_2n = matchi_2n;
  C3 I720 (matchi_1n, ifint_0n[34], ifint_0n[32], itint_0n[33]);
  assign sel_1n = matchi_1n;
  C3 I722 (matchi_0n, ifint_0n[34], ifint_0n[33], itint_0n[32]);
  assign sel_0n = matchi_0n;
endmodule

module AO22 (
  q,
  i0,
  i1,
  i2,
  i3
);
  output q;
  input i0;
  input i1;
  input i2;
  input i3;
  wire [1:0] int_0n;
  OR2 I0 (q, int_0n[0], int_0n[1]);
  AND2 I1 (int_0n[1], i2, i3);
  AND2 I2 (int_0n[0], i0, i1);
endmodule

module AC2 (
  q,
  i0,
  i1
);
  output q;
  input i0;
  input i1;
  AO22 I0 (q, i0, i1, i0, q);
endmodule

module GIVE_INIT (
  iout,
  initialise
);
  output iout;
  input initialise;
  assign iout = initialise;
endmodule

module BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rd_0r0d, rd_0r1d, rd_0a,
  initialise
);
  input wg_0r0d;
  input wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output rd_0r0d;
  output rd_0r1d;
  input rd_0a;
  input initialise;
  wire wf_0n;
  wire wt_0n;
  wire df_0n;
  wire dt_0n;
  wire rgrint_0n;
  wire wc_0n;
  wire wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire wgfint_0n;
  wire wgtint_0n;
  wire rgaint_0n;
  wire rdfint_0n;
  wire rdtint_0n;
  wire wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire gif_0n;
  wire git_0n;
  wire complete1162_0n;
  wire gt1161_0n;
  wire gf1160_0n;
  assign rgaint_0n = rd_0a;
  assign rd_0r0d = rdfint_0n;
  assign rd_0r1d = rdtint_0n;
  assign wg_0a = wgaint_0n;
  assign wgfint_0n = wg_0r0d;
  assign wgtint_0n = wg_0r1d;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I10 (nanyread_0n, rgrint_0n, rgaint_0n);
  AND2 I11 (rdtint_0n, rgrint_0n, dt_0n);
  AND2 I12 (rdfint_0n, rgrint_0n, df_0n);
  C2 I13 (wdrint_0n, wc_0n, wacks_0n);
  assign wen_0n = wc_0n;
  assign wt_0n = git_0n;
  assign wf_0n = gif_0n;
  AC2 I17 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I19 (git_0n, wgtint_0n, ig_0n);
  AND2 I20 (gif_0n, wgfint_0n, ig_0n);
  assign wc_0n = complete1162_0n;
  OR2 I22 (complete1162_0n, wgfint_0n, wgtint_0n);
  AO22 I23 (wacks_0n, gf1160_0n, df_0n, gt1161_0n, dt_0n);
  NOR2 I24 (dt_0n, df_0n, gf1160_0n);
  NOR3 I25 (df_0n, dt_0n, gt1161_0n, init_0n);
  AND2 I26 (gt1161_0n, wt_0n, wen_0n);
  AND2 I27 (gf1160_0n, wf_0n, wen_0n);
  GIVE_INIT I28 (init_0n, initialise);
endmodule

module BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m72m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  initialise
);
  input wg_0r0d;
  input wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output rd_0r0d;
  output rd_0r1d;
  input rd_0a;
  output rd_1r0d;
  output rd_1r1d;
  input rd_1a;
  input initialise;
  wire [1:0] internal_0n;
  wire wf_0n;
  wire wt_0n;
  wire df_0n;
  wire dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire wc_0n;
  wire wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire wgfint_0n;
  wire wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire rdfint_0n;
  wire rdfint_1n;
  wire rdtint_0n;
  wire rdtint_1n;
  wire wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire gif_0n;
  wire git_0n;
  wire complete1173_0n;
  wire gt1172_0n;
  wire gf1171_0n;
  assign rgaint_1n = rd_1a;
  assign rd_1r0d = rdfint_1n;
  assign rd_1r1d = rdtint_1n;
  assign rgaint_0n = rd_0a;
  assign rd_0r0d = rdfint_0n;
  assign rd_0r1d = rdtint_0n;
  assign wg_0a = wgaint_0n;
  assign wgfint_0n = wg_0r0d;
  assign wgtint_0n = wg_0r1d;
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I15 (internal_0n[0], rgrint_0n, rgrint_1n);
  NOR2 I16 (internal_0n[1], rgaint_0n, rgaint_1n);
  AND2 I17 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I18 (rdtint_1n, rgrint_1n, dt_0n);
  AND2 I19 (rdtint_0n, rgrint_0n, dt_0n);
  AND2 I20 (rdfint_1n, rgrint_1n, df_0n);
  AND2 I21 (rdfint_0n, rgrint_0n, df_0n);
  C2 I22 (wdrint_0n, wc_0n, wacks_0n);
  assign wen_0n = wc_0n;
  assign wt_0n = git_0n;
  assign wf_0n = gif_0n;
  AC2 I26 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I28 (git_0n, wgtint_0n, ig_0n);
  AND2 I29 (gif_0n, wgfint_0n, ig_0n);
  assign wc_0n = complete1173_0n;
  OR2 I31 (complete1173_0n, wgfint_0n, wgtint_0n);
  AO22 I32 (wacks_0n, gf1171_0n, df_0n, gt1172_0n, dt_0n);
  NOR2 I33 (dt_0n, df_0n, gf1171_0n);
  NOR3 I34 (df_0n, dt_0n, gt1172_0n, init_0n);
  AND2 I35 (gt1172_0n, wt_0n, wen_0n);
  AND2 I36 (gf1171_0n, wf_0n, wen_0n);
  GIVE_INIT I37 (init_0n, initialise);
endmodule

module BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m73m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rg_2r, rg_2a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  rd_2r0d, rd_2r1d, rd_2a,
  initialise
);
  input wg_0r0d;
  input wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output rd_0r0d;
  output rd_0r1d;
  input rd_0a;
  output rd_1r0d;
  output rd_1r1d;
  input rd_1a;
  output rd_2r0d;
  output rd_2r1d;
  input rd_2a;
  input initialise;
  wire [1:0] internal_0n;
  wire wf_0n;
  wire wt_0n;
  wire df_0n;
  wire dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire rgrint_2n;
  wire wc_0n;
  wire wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire wgfint_0n;
  wire wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire rgaint_2n;
  wire rdfint_0n;
  wire rdfint_1n;
  wire rdfint_2n;
  wire rdtint_0n;
  wire rdtint_1n;
  wire rdtint_2n;
  wire wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire gif_0n;
  wire git_0n;
  wire complete1188_0n;
  wire gt1187_0n;
  wire gf1186_0n;
  assign rgaint_2n = rd_2a;
  assign rd_2r0d = rdfint_2n;
  assign rd_2r1d = rdtint_2n;
  assign rgaint_1n = rd_1a;
  assign rd_1r0d = rdfint_1n;
  assign rd_1r1d = rdtint_1n;
  assign rgaint_0n = rd_0a;
  assign rd_0r0d = rdfint_0n;
  assign rd_0r1d = rdtint_0n;
  assign wg_0a = wgaint_0n;
  assign wgfint_0n = wg_0r0d;
  assign wgtint_0n = wg_0r1d;
  assign rg_2a = rgaint_2n;
  assign rgrint_2n = rg_2r;
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR3 I20 (internal_0n[0], rgrint_0n, rgrint_1n, rgrint_2n);
  NOR3 I21 (internal_0n[1], rgaint_0n, rgaint_1n, rgaint_2n);
  AND2 I22 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I23 (rdtint_2n, rgrint_2n, dt_0n);
  AND2 I24 (rdtint_1n, rgrint_1n, dt_0n);
  AND2 I25 (rdtint_0n, rgrint_0n, dt_0n);
  AND2 I26 (rdfint_2n, rgrint_2n, df_0n);
  AND2 I27 (rdfint_1n, rgrint_1n, df_0n);
  AND2 I28 (rdfint_0n, rgrint_0n, df_0n);
  C2 I29 (wdrint_0n, wc_0n, wacks_0n);
  assign wen_0n = wc_0n;
  assign wt_0n = git_0n;
  assign wf_0n = gif_0n;
  AC2 I33 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I35 (git_0n, wgtint_0n, ig_0n);
  AND2 I36 (gif_0n, wgfint_0n, ig_0n);
  assign wc_0n = complete1188_0n;
  OR2 I38 (complete1188_0n, wgfint_0n, wgtint_0n);
  AO22 I39 (wacks_0n, gf1186_0n, df_0n, gt1187_0n, dt_0n);
  NOR2 I40 (dt_0n, df_0n, gf1186_0n);
  NOR3 I41 (df_0n, dt_0n, gt1187_0n, init_0n);
  AND2 I42 (gt1187_0n, wt_0n, wen_0n);
  AND2 I43 (gf1186_0n, wf_0n, wen_0n);
  GIVE_INIT I44 (init_0n, initialise);
endmodule

module BrzV_1_l6__28_29_l43__28_28_280_201_29_29__m74m (
  wg_0r0d, wg_0r1d, wg_0a,
  wg_1r0d, wg_1r1d, wg_1a,
  wd_0r, wd_0a,
  wd_1r, wd_1a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  initialise
);
  input wg_0r0d;
  input wg_0r1d;
  output wg_0a;
  input wg_1r0d;
  input wg_1r1d;
  output wg_1a;
  output wd_0r;
  input wd_0a;
  output wd_1r;
  input wd_1a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output rd_0r0d;
  output rd_0r1d;
  input rd_0a;
  output rd_1r0d;
  output rd_1r1d;
  input rd_1a;
  input initialise;
  wire [1:0] internal_0n;
  wire wf_0n;
  wire wt_0n;
  wire df_0n;
  wire dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire wc_0n;
  wire wc_1n;
  wire wacks_0n;
  wire wdrint_0n;
  wire wdrint_1n;
  wire wgaint_0n;
  wire wgaint_1n;
  wire wgfint_0n;
  wire wgfint_1n;
  wire wgtint_0n;
  wire wgtint_1n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire rdfint_0n;
  wire rdfint_1n;
  wire rdtint_0n;
  wire rdtint_1n;
  wire wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire igc_1n;
  wire ig_0n;
  wire ig_1n;
  wire gif_0n;
  wire gif_1n;
  wire git_0n;
  wire git_1n;
  wire complete1208_0n;
  wire complete1207_0n;
  wire gt1206_0n;
  wire gf1205_0n;
  assign rgaint_1n = rd_1a;
  assign rd_1r0d = rdfint_1n;
  assign rd_1r1d = rdtint_1n;
  assign rgaint_0n = rd_0a;
  assign rd_0r0d = rdfint_0n;
  assign rd_0r1d = rdtint_0n;
  assign wg_1a = wgaint_1n;
  assign wgfint_1n = wg_1r0d;
  assign wgtint_1n = wg_1r1d;
  assign wg_0a = wgaint_0n;
  assign wgfint_0n = wg_0r0d;
  assign wgtint_0n = wg_0r1d;
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_1n = wd_1a;
  assign wd_1r = wdrint_1n;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I20 (internal_0n[0], rgrint_0n, rgrint_1n);
  NOR2 I21 (internal_0n[1], rgaint_0n, rgaint_1n);
  AND2 I22 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I23 (rdtint_1n, rgrint_1n, dt_0n);
  AND2 I24 (rdtint_0n, rgrint_0n, dt_0n);
  AND2 I25 (rdfint_1n, rgrint_1n, df_0n);
  AND2 I26 (rdfint_0n, rgrint_0n, df_0n);
  C2 I27 (wdrint_1n, wc_1n, wacks_0n);
  C2 I28 (wdrint_0n, wc_0n, wacks_0n);
  OR2 I29 (wen_0n, wc_1n, wc_0n);
  OR2 I30 (wt_0n, git_1n, git_0n);
  OR2 I31 (wf_0n, gif_1n, gif_0n);
  AC2 I32 (ig_0n, igc_0n, nanyread_0n);
  AC2 I33 (ig_1n, igc_1n, nanyread_0n);
  assign igc_0n = wc_0n;
  assign igc_1n = wc_1n;
  AND2 I36 (git_1n, wgtint_1n, ig_1n);
  AND2 I37 (git_0n, wgtint_0n, ig_0n);
  AND2 I38 (gif_1n, wgfint_1n, ig_1n);
  AND2 I39 (gif_0n, wgfint_0n, ig_0n);
  assign wc_1n = complete1208_0n;
  OR2 I41 (complete1208_0n, wgfint_1n, wgtint_1n);
  assign wc_0n = complete1207_0n;
  OR2 I43 (complete1207_0n, wgfint_0n, wgtint_0n);
  AO22 I44 (wacks_0n, gf1205_0n, df_0n, gt1206_0n, dt_0n);
  NOR2 I45 (dt_0n, df_0n, gf1205_0n);
  NOR3 I46 (df_0n, dt_0n, gt1206_0n, init_0n);
  AND2 I47 (gt1206_0n, wt_0n, wen_0n);
  AND2 I48 (gf1205_0n, wf_0n, wen_0n);
  GIVE_INIT I49 (init_0n, initialise);
endmodule

module BrzV_3_l6__28_29_l23__28_28_280_203_29_29__m75m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rg_2r, rg_2a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  rd_2r0d, rd_2r1d, rd_2a,
  initialise
);
  input [2:0] wg_0r0d;
  input [2:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [2:0] rd_0r0d;
  output [2:0] rd_0r1d;
  input rd_0a;
  output [2:0] rd_1r0d;
  output [2:0] rd_1r1d;
  input rd_1a;
  output [2:0] rd_2r0d;
  output [2:0] rd_2r1d;
  input rd_2a;
  input initialise;
  wire [3:0] internal_0n;
  wire [2:0] wf_0n;
  wire [2:0] wt_0n;
  wire [2:0] df_0n;
  wire [2:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire rgrint_2n;
  wire wc_0n;
  wire [2:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [2:0] wgfint_0n;
  wire [2:0] wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire rgaint_2n;
  wire [2:0] rdfint_0n;
  wire [2:0] rdfint_1n;
  wire [2:0] rdfint_2n;
  wire [2:0] rdtint_0n;
  wire [2:0] rdtint_1n;
  wire [2:0] rdtint_2n;
  wire [2:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [2:0] gif_0n;
  wire [2:0] git_0n;
  wire [2:0] complete1227_0n;
  wire [2:0] gt1226_0n;
  wire [2:0] gf1225_0n;
  assign rgaint_2n = rd_2a;
  assign rd_2r0d[0] = rdfint_2n[0];
  assign rd_2r0d[1] = rdfint_2n[1];
  assign rd_2r0d[2] = rdfint_2n[2];
  assign rd_2r1d[0] = rdtint_2n[0];
  assign rd_2r1d[1] = rdtint_2n[1];
  assign rd_2r1d[2] = rdtint_2n[2];
  assign rgaint_1n = rd_1a;
  assign rd_1r0d[0] = rdfint_1n[0];
  assign rd_1r0d[1] = rdfint_1n[1];
  assign rd_1r0d[2] = rdfint_1n[2];
  assign rd_1r1d[0] = rdtint_1n[0];
  assign rd_1r1d[1] = rdtint_1n[1];
  assign rd_1r1d[2] = rdtint_1n[2];
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign rg_2a = rgaint_2n;
  assign rgrint_2n = rg_2r;
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR3 I36 (internal_0n[0], rgrint_0n, rgrint_1n, rgrint_2n);
  NOR3 I37 (internal_0n[1], rgaint_0n, rgaint_1n, rgaint_2n);
  AND2 I38 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I39 (rdtint_2n[0], rgrint_2n, dt_0n[0]);
  AND2 I40 (rdtint_2n[1], rgrint_2n, dt_0n[1]);
  AND2 I41 (rdtint_2n[2], rgrint_2n, dt_0n[2]);
  AND2 I42 (rdtint_1n[0], rgrint_1n, dt_0n[0]);
  AND2 I43 (rdtint_1n[1], rgrint_1n, dt_0n[1]);
  AND2 I44 (rdtint_1n[2], rgrint_1n, dt_0n[2]);
  AND2 I45 (rdtint_0n[0], rgrint_0n, dt_0n[0]);
  AND2 I46 (rdtint_0n[1], rgrint_0n, dt_0n[1]);
  AND2 I47 (rdtint_0n[2], rgrint_0n, dt_0n[2]);
  AND2 I48 (rdfint_2n[0], rgrint_2n, df_0n[0]);
  AND2 I49 (rdfint_2n[1], rgrint_2n, df_0n[1]);
  AND2 I50 (rdfint_2n[2], rgrint_2n, df_0n[2]);
  AND2 I51 (rdfint_1n[0], rgrint_1n, df_0n[0]);
  AND2 I52 (rdfint_1n[1], rgrint_1n, df_0n[1]);
  AND2 I53 (rdfint_1n[2], rgrint_1n, df_0n[2]);
  AND2 I54 (rdfint_0n[0], rgrint_0n, df_0n[0]);
  AND2 I55 (rdfint_0n[1], rgrint_0n, df_0n[1]);
  AND2 I56 (rdfint_0n[2], rgrint_0n, df_0n[2]);
  C2 I57 (internal_0n[2], wc_0n, wacks_0n[2]);
  C2 I58 (internal_0n[3], wacks_0n[1], wacks_0n[0]);
  C2 I59 (wdrint_0n, internal_0n[2], internal_0n[3]);
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I69 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I71 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I72 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I73 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I74 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I75 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I76 (gif_0n[2], wgfint_0n[2], ig_0n);
  C3 I77 (wc_0n, complete1227_0n[0], complete1227_0n[1], complete1227_0n[2]);
  OR2 I78 (complete1227_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I79 (complete1227_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I80 (complete1227_0n[2], wgfint_0n[2], wgtint_0n[2]);
  AO22 I81 (wacks_0n[2], gf1225_0n[2], df_0n[2], gt1226_0n[2], dt_0n[2]);
  NOR2 I82 (dt_0n[2], df_0n[2], gf1225_0n[2]);
  NOR3 I83 (df_0n[2], dt_0n[2], gt1226_0n[2], init_0n);
  AND2 I84 (gt1226_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I85 (gf1225_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I86 (wacks_0n[1], gf1225_0n[1], df_0n[1], gt1226_0n[1], dt_0n[1]);
  NOR2 I87 (dt_0n[1], df_0n[1], gf1225_0n[1]);
  NOR3 I88 (df_0n[1], dt_0n[1], gt1226_0n[1], init_0n);
  AND2 I89 (gt1226_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I90 (gf1225_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I91 (wacks_0n[0], gf1225_0n[0], df_0n[0], gt1226_0n[0], dt_0n[0]);
  NOR2 I92 (dt_0n[0], df_0n[0], gf1225_0n[0]);
  NOR3 I93 (df_0n[0], dt_0n[0], gt1226_0n[0], init_0n);
  AND2 I94 (gt1226_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I95 (gf1225_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I96 (init_0n, initialise);
endmodule

module BrzV_3_l6__28_29_l23__28_28_280_203_29_29__m76m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rg_2r, rg_2a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  rd_2r0d, rd_2r1d, rd_2a,
  initialise
);
  input [2:0] wg_0r0d;
  input [2:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [2:0] rd_0r0d;
  output [2:0] rd_0r1d;
  input rd_0a;
  output rd_1r0d;
  output rd_1r1d;
  input rd_1a;
  output rd_2r0d;
  output rd_2r1d;
  input rd_2a;
  input initialise;
  wire [3:0] internal_0n;
  wire [2:0] wf_0n;
  wire [2:0] wt_0n;
  wire [2:0] df_0n;
  wire [2:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire rgrint_2n;
  wire wc_0n;
  wire [2:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [2:0] wgfint_0n;
  wire [2:0] wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire rgaint_2n;
  wire [2:0] rdfint_0n;
  wire rdfint_1n;
  wire rdfint_2n;
  wire [2:0] rdtint_0n;
  wire rdtint_1n;
  wire rdtint_2n;
  wire [2:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [2:0] gif_0n;
  wire [2:0] git_0n;
  wire [2:0] complete1246_0n;
  wire [2:0] gt1245_0n;
  wire [2:0] gf1244_0n;
  assign rgaint_2n = rd_2a;
  assign rd_2r0d = rdfint_2n;
  assign rd_2r1d = rdtint_2n;
  assign rgaint_1n = rd_1a;
  assign rd_1r0d = rdfint_1n;
  assign rd_1r1d = rdtint_1n;
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign rg_2a = rgaint_2n;
  assign rgrint_2n = rg_2r;
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR3 I28 (internal_0n[0], rgrint_0n, rgrint_1n, rgrint_2n);
  NOR3 I29 (internal_0n[1], rgaint_0n, rgaint_1n, rgaint_2n);
  AND2 I30 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I31 (rdtint_2n, rgrint_2n, dt_0n[0]);
  AND2 I32 (rdtint_1n, rgrint_1n, dt_0n[2]);
  AND2 I33 (rdtint_0n[0], rgrint_0n, dt_0n[0]);
  AND2 I34 (rdtint_0n[1], rgrint_0n, dt_0n[1]);
  AND2 I35 (rdtint_0n[2], rgrint_0n, dt_0n[2]);
  AND2 I36 (rdfint_2n, rgrint_2n, df_0n[0]);
  AND2 I37 (rdfint_1n, rgrint_1n, df_0n[2]);
  AND2 I38 (rdfint_0n[0], rgrint_0n, df_0n[0]);
  AND2 I39 (rdfint_0n[1], rgrint_0n, df_0n[1]);
  AND2 I40 (rdfint_0n[2], rgrint_0n, df_0n[2]);
  C2 I41 (internal_0n[2], wc_0n, wacks_0n[2]);
  C2 I42 (internal_0n[3], wacks_0n[1], wacks_0n[0]);
  C2 I43 (wdrint_0n, internal_0n[2], internal_0n[3]);
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I53 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I55 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I56 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I57 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I58 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I59 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I60 (gif_0n[2], wgfint_0n[2], ig_0n);
  C3 I61 (wc_0n, complete1246_0n[0], complete1246_0n[1], complete1246_0n[2]);
  OR2 I62 (complete1246_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I63 (complete1246_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I64 (complete1246_0n[2], wgfint_0n[2], wgtint_0n[2]);
  AO22 I65 (wacks_0n[2], gf1244_0n[2], df_0n[2], gt1245_0n[2], dt_0n[2]);
  NOR2 I66 (dt_0n[2], df_0n[2], gf1244_0n[2]);
  NOR3 I67 (df_0n[2], dt_0n[2], gt1245_0n[2], init_0n);
  AND2 I68 (gt1245_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I69 (gf1244_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I70 (wacks_0n[1], gf1244_0n[1], df_0n[1], gt1245_0n[1], dt_0n[1]);
  NOR2 I71 (dt_0n[1], df_0n[1], gf1244_0n[1]);
  NOR3 I72 (df_0n[1], dt_0n[1], gt1245_0n[1], init_0n);
  AND2 I73 (gt1245_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I74 (gf1244_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I75 (wacks_0n[0], gf1244_0n[0], df_0n[0], gt1245_0n[0], dt_0n[0]);
  NOR2 I76 (dt_0n[0], df_0n[0], gf1244_0n[0]);
  NOR3 I77 (df_0n[0], dt_0n[0], gt1245_0n[0], init_0n);
  AND2 I78 (gt1245_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I79 (gf1244_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I80 (init_0n, initialise);
endmodule

module BrzV_4_l6__28_29_l43__28_28_280_204_29_29__m77m (
  wg_0r0d, wg_0r1d, wg_0a,
  wg_1r0d, wg_1r1d, wg_1a,
  wd_0r, wd_0a,
  wd_1r, wd_1a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rg_2r, rg_2a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  rd_2r0d, rd_2r1d, rd_2a,
  initialise
);
  input [3:0] wg_0r0d;
  input [3:0] wg_0r1d;
  output wg_0a;
  input [3:0] wg_1r0d;
  input [3:0] wg_1r1d;
  output wg_1a;
  output wd_0r;
  input wd_0a;
  output wd_1r;
  input wd_1a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [3:0] rd_0r0d;
  output [3:0] rd_0r1d;
  input rd_0a;
  output [3:0] rd_1r0d;
  output [3:0] rd_1r1d;
  input rd_1a;
  output rd_2r0d;
  output rd_2r1d;
  input rd_2a;
  input initialise;
  wire [9:0] internal_0n;
  wire [3:0] wf_0n;
  wire [3:0] wt_0n;
  wire [3:0] df_0n;
  wire [3:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire rgrint_2n;
  wire wc_0n;
  wire wc_1n;
  wire [3:0] wacks_0n;
  wire wdrint_0n;
  wire wdrint_1n;
  wire wgaint_0n;
  wire wgaint_1n;
  wire [3:0] wgfint_0n;
  wire [3:0] wgfint_1n;
  wire [3:0] wgtint_0n;
  wire [3:0] wgtint_1n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire rgaint_2n;
  wire [3:0] rdfint_0n;
  wire [3:0] rdfint_1n;
  wire rdfint_2n;
  wire [3:0] rdtint_0n;
  wire [3:0] rdtint_1n;
  wire rdtint_2n;
  wire [3:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire igc_1n;
  wire ig_0n;
  wire ig_1n;
  wire [3:0] gif_0n;
  wire [3:0] gif_1n;
  wire [3:0] git_0n;
  wire [3:0] git_1n;
  wire [3:0] complete1266_0n;
  wire [3:0] complete1265_0n;
  wire [3:0] gt1264_0n;
  wire [3:0] gf1263_0n;
  assign rgaint_2n = rd_2a;
  assign rd_2r0d = rdfint_2n;
  assign rd_2r1d = rdtint_2n;
  assign rgaint_1n = rd_1a;
  assign rd_1r0d[0] = rdfint_1n[0];
  assign rd_1r0d[1] = rdfint_1n[1];
  assign rd_1r0d[2] = rdfint_1n[2];
  assign rd_1r0d[3] = rdfint_1n[3];
  assign rd_1r1d[0] = rdtint_1n[0];
  assign rd_1r1d[1] = rdtint_1n[1];
  assign rd_1r1d[2] = rdtint_1n[2];
  assign rd_1r1d[3] = rdtint_1n[3];
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign wg_1a = wgaint_1n;
  assign wgfint_1n[0] = wg_1r0d[0];
  assign wgfint_1n[1] = wg_1r0d[1];
  assign wgfint_1n[2] = wg_1r0d[2];
  assign wgfint_1n[3] = wg_1r0d[3];
  assign wgtint_1n[0] = wg_1r1d[0];
  assign wgtint_1n[1] = wg_1r1d[1];
  assign wgtint_1n[2] = wg_1r1d[2];
  assign wgtint_1n[3] = wg_1r1d[3];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign rg_2a = rgaint_2n;
  assign rgrint_2n = rg_2r;
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_1n = wd_1a;
  assign wd_1r = wdrint_1n;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR3 I49 (internal_0n[0], rgrint_0n, rgrint_1n, rgrint_2n);
  NOR3 I50 (internal_0n[1], rgaint_0n, rgaint_1n, rgaint_2n);
  AND2 I51 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I52 (rdtint_2n, rgrint_2n, dt_0n[3]);
  AND2 I53 (rdtint_1n[0], rgrint_1n, dt_0n[0]);
  AND2 I54 (rdtint_1n[1], rgrint_1n, dt_0n[1]);
  AND2 I55 (rdtint_1n[2], rgrint_1n, dt_0n[2]);
  AND2 I56 (rdtint_1n[3], rgrint_1n, dt_0n[3]);
  AND2 I57 (rdtint_0n[0], rgrint_0n, dt_0n[0]);
  AND2 I58 (rdtint_0n[1], rgrint_0n, dt_0n[1]);
  AND2 I59 (rdtint_0n[2], rgrint_0n, dt_0n[2]);
  AND2 I60 (rdtint_0n[3], rgrint_0n, dt_0n[3]);
  AND2 I61 (rdfint_2n, rgrint_2n, df_0n[3]);
  AND2 I62 (rdfint_1n[0], rgrint_1n, df_0n[0]);
  AND2 I63 (rdfint_1n[1], rgrint_1n, df_0n[1]);
  AND2 I64 (rdfint_1n[2], rgrint_1n, df_0n[2]);
  AND2 I65 (rdfint_1n[3], rgrint_1n, df_0n[3]);
  AND2 I66 (rdfint_0n[0], rgrint_0n, df_0n[0]);
  AND2 I67 (rdfint_0n[1], rgrint_0n, df_0n[1]);
  AND2 I68 (rdfint_0n[2], rgrint_0n, df_0n[2]);
  AND2 I69 (rdfint_0n[3], rgrint_0n, df_0n[3]);
  C3 I70 (internal_0n[2], wc_1n, wacks_0n[3], wacks_0n[2]);
  C2 I71 (internal_0n[3], wacks_0n[1], wacks_0n[0]);
  C2 I72 (wdrint_1n, internal_0n[2], internal_0n[3]);
  C3 I73 (internal_0n[4], wc_0n, wacks_0n[3], wacks_0n[2]);
  C2 I74 (internal_0n[5], wacks_0n[1], wacks_0n[0]);
  C2 I75 (wdrint_0n, internal_0n[4], internal_0n[5]);
  OR2 I76 (wen_0n[3], wc_1n, wc_0n);
  OR2 I77 (wen_0n[2], wc_1n, wc_0n);
  OR2 I78 (wen_0n[1], wc_1n, wc_0n);
  OR2 I79 (wen_0n[0], wc_1n, wc_0n);
  OR2 I80 (wt_0n[3], git_1n[3], git_0n[3]);
  OR2 I81 (wt_0n[2], git_1n[2], git_0n[2]);
  OR2 I82 (wt_0n[1], git_1n[1], git_0n[1]);
  OR2 I83 (wt_0n[0], git_1n[0], git_0n[0]);
  OR2 I84 (wf_0n[3], gif_1n[3], gif_0n[3]);
  OR2 I85 (wf_0n[2], gif_1n[2], gif_0n[2]);
  OR2 I86 (wf_0n[1], gif_1n[1], gif_0n[1]);
  OR2 I87 (wf_0n[0], gif_1n[0], gif_0n[0]);
  AC2 I88 (ig_0n, igc_0n, nanyread_0n);
  AC2 I89 (ig_1n, igc_1n, nanyread_0n);
  assign igc_0n = wc_0n;
  assign igc_1n = wc_1n;
  AND2 I92 (git_1n[0], wgtint_1n[0], ig_1n);
  AND2 I93 (git_1n[1], wgtint_1n[1], ig_1n);
  AND2 I94 (git_1n[2], wgtint_1n[2], ig_1n);
  AND2 I95 (git_1n[3], wgtint_1n[3], ig_1n);
  AND2 I96 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I97 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I98 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I99 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I100 (gif_1n[0], wgfint_1n[0], ig_1n);
  AND2 I101 (gif_1n[1], wgfint_1n[1], ig_1n);
  AND2 I102 (gif_1n[2], wgfint_1n[2], ig_1n);
  AND2 I103 (gif_1n[3], wgfint_1n[3], ig_1n);
  AND2 I104 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I105 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I106 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I107 (gif_0n[3], wgfint_0n[3], ig_0n);
  C2 I108 (internal_0n[6], complete1266_0n[0], complete1266_0n[1]);
  C2 I109 (internal_0n[7], complete1266_0n[2], complete1266_0n[3]);
  C2 I110 (wc_1n, internal_0n[6], internal_0n[7]);
  OR2 I111 (complete1266_0n[0], wgfint_1n[0], wgtint_1n[0]);
  OR2 I112 (complete1266_0n[1], wgfint_1n[1], wgtint_1n[1]);
  OR2 I113 (complete1266_0n[2], wgfint_1n[2], wgtint_1n[2]);
  OR2 I114 (complete1266_0n[3], wgfint_1n[3], wgtint_1n[3]);
  C2 I115 (internal_0n[8], complete1265_0n[0], complete1265_0n[1]);
  C2 I116 (internal_0n[9], complete1265_0n[2], complete1265_0n[3]);
  C2 I117 (wc_0n, internal_0n[8], internal_0n[9]);
  OR2 I118 (complete1265_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I119 (complete1265_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I120 (complete1265_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I121 (complete1265_0n[3], wgfint_0n[3], wgtint_0n[3]);
  AO22 I122 (wacks_0n[3], gf1263_0n[3], df_0n[3], gt1264_0n[3], dt_0n[3]);
  NOR2 I123 (dt_0n[3], df_0n[3], gf1263_0n[3]);
  NOR3 I124 (df_0n[3], dt_0n[3], gt1264_0n[3], init_0n);
  AND2 I125 (gt1264_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I126 (gf1263_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I127 (wacks_0n[2], gf1263_0n[2], df_0n[2], gt1264_0n[2], dt_0n[2]);
  NOR2 I128 (dt_0n[2], df_0n[2], gf1263_0n[2]);
  NOR3 I129 (df_0n[2], dt_0n[2], gt1264_0n[2], init_0n);
  AND2 I130 (gt1264_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I131 (gf1263_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I132 (wacks_0n[1], gf1263_0n[1], df_0n[1], gt1264_0n[1], dt_0n[1]);
  NOR2 I133 (dt_0n[1], df_0n[1], gf1263_0n[1]);
  NOR3 I134 (df_0n[1], dt_0n[1], gt1264_0n[1], init_0n);
  AND2 I135 (gt1264_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I136 (gf1263_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I137 (wacks_0n[0], gf1263_0n[0], df_0n[0], gt1264_0n[0], dt_0n[0]);
  NOR2 I138 (dt_0n[0], df_0n[0], gf1263_0n[0]);
  NOR3 I139 (df_0n[0], dt_0n[0], gt1264_0n[0], init_0n);
  AND2 I140 (gt1264_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I141 (gf1263_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I142 (init_0n, initialise);
endmodule

module BrzV_10_l6__28_29_l24__28_28_280_2010_29_2_m78m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rd_0r0d, rd_0r1d, rd_0a,
  initialise
);
  input [9:0] wg_0r0d;
  input [9:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [9:0] rd_0r0d;
  output [9:0] rd_0r1d;
  input rd_0a;
  input initialise;
  wire [11:0] internal_0n;
  wire [9:0] wf_0n;
  wire [9:0] wt_0n;
  wire [9:0] df_0n;
  wire [9:0] dt_0n;
  wire rgrint_0n;
  wire wc_0n;
  wire [9:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [9:0] wgfint_0n;
  wire [9:0] wgtint_0n;
  wire rgaint_0n;
  wire [9:0] rdfint_0n;
  wire [9:0] rdtint_0n;
  wire [9:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [9:0] gif_0n;
  wire [9:0] git_0n;
  wire [9:0] complete1289_0n;
  wire [9:0] gt1288_0n;
  wire [9:0] gf1287_0n;
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I46 (nanyread_0n, rgrint_0n, rgaint_0n);
  AND2 I47 (rdtint_0n[0], rgrint_0n, dt_0n[0]);
  AND2 I48 (rdtint_0n[1], rgrint_0n, dt_0n[1]);
  AND2 I49 (rdtint_0n[2], rgrint_0n, dt_0n[2]);
  AND2 I50 (rdtint_0n[3], rgrint_0n, dt_0n[3]);
  AND2 I51 (rdtint_0n[4], rgrint_0n, dt_0n[4]);
  AND2 I52 (rdtint_0n[5], rgrint_0n, dt_0n[5]);
  AND2 I53 (rdtint_0n[6], rgrint_0n, dt_0n[6]);
  AND2 I54 (rdtint_0n[7], rgrint_0n, dt_0n[7]);
  AND2 I55 (rdtint_0n[8], rgrint_0n, dt_0n[8]);
  AND2 I56 (rdtint_0n[9], rgrint_0n, dt_0n[9]);
  AND2 I57 (rdfint_0n[0], rgrint_0n, df_0n[0]);
  AND2 I58 (rdfint_0n[1], rgrint_0n, df_0n[1]);
  AND2 I59 (rdfint_0n[2], rgrint_0n, df_0n[2]);
  AND2 I60 (rdfint_0n[3], rgrint_0n, df_0n[3]);
  AND2 I61 (rdfint_0n[4], rgrint_0n, df_0n[4]);
  AND2 I62 (rdfint_0n[5], rgrint_0n, df_0n[5]);
  AND2 I63 (rdfint_0n[6], rgrint_0n, df_0n[6]);
  AND2 I64 (rdfint_0n[7], rgrint_0n, df_0n[7]);
  AND2 I65 (rdfint_0n[8], rgrint_0n, df_0n[8]);
  AND2 I66 (rdfint_0n[9], rgrint_0n, df_0n[9]);
  C3 I67 (internal_0n[0], wc_0n, wacks_0n[9], wacks_0n[8]);
  C3 I68 (internal_0n[1], wacks_0n[7], wacks_0n[6], wacks_0n[5]);
  C3 I69 (internal_0n[2], wacks_0n[4], wacks_0n[3], wacks_0n[2]);
  C2 I70 (internal_0n[3], wacks_0n[1], wacks_0n[0]);
  C2 I71 (internal_0n[4], internal_0n[0], internal_0n[1]);
  C2 I72 (internal_0n[5], internal_0n[2], internal_0n[3]);
  C2 I73 (wdrint_0n, internal_0n[4], internal_0n[5]);
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I104 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I106 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I107 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I108 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I109 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I110 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I111 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I112 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I113 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I114 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I115 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I116 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I117 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I118 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I119 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I120 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I121 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I122 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I123 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I124 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I125 (gif_0n[9], wgfint_0n[9], ig_0n);
  C3 I126 (internal_0n[6], complete1289_0n[0], complete1289_0n[1], complete1289_0n[2]);
  C3 I127 (internal_0n[7], complete1289_0n[3], complete1289_0n[4], complete1289_0n[5]);
  C2 I128 (internal_0n[8], complete1289_0n[6], complete1289_0n[7]);
  C2 I129 (internal_0n[9], complete1289_0n[8], complete1289_0n[9]);
  C2 I130 (internal_0n[10], internal_0n[6], internal_0n[7]);
  C2 I131 (internal_0n[11], internal_0n[8], internal_0n[9]);
  C2 I132 (wc_0n, internal_0n[10], internal_0n[11]);
  OR2 I133 (complete1289_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I134 (complete1289_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I135 (complete1289_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I136 (complete1289_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I137 (complete1289_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I138 (complete1289_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I139 (complete1289_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I140 (complete1289_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I141 (complete1289_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I142 (complete1289_0n[9], wgfint_0n[9], wgtint_0n[9]);
  AO22 I143 (wacks_0n[9], gf1287_0n[9], df_0n[9], gt1288_0n[9], dt_0n[9]);
  NOR2 I144 (dt_0n[9], df_0n[9], gf1287_0n[9]);
  NOR3 I145 (df_0n[9], dt_0n[9], gt1288_0n[9], init_0n);
  AND2 I146 (gt1288_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I147 (gf1287_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I148 (wacks_0n[8], gf1287_0n[8], df_0n[8], gt1288_0n[8], dt_0n[8]);
  NOR2 I149 (dt_0n[8], df_0n[8], gf1287_0n[8]);
  NOR3 I150 (df_0n[8], dt_0n[8], gt1288_0n[8], init_0n);
  AND2 I151 (gt1288_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I152 (gf1287_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I153 (wacks_0n[7], gf1287_0n[7], df_0n[7], gt1288_0n[7], dt_0n[7]);
  NOR2 I154 (dt_0n[7], df_0n[7], gf1287_0n[7]);
  NOR3 I155 (df_0n[7], dt_0n[7], gt1288_0n[7], init_0n);
  AND2 I156 (gt1288_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I157 (gf1287_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I158 (wacks_0n[6], gf1287_0n[6], df_0n[6], gt1288_0n[6], dt_0n[6]);
  NOR2 I159 (dt_0n[6], df_0n[6], gf1287_0n[6]);
  NOR3 I160 (df_0n[6], dt_0n[6], gt1288_0n[6], init_0n);
  AND2 I161 (gt1288_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I162 (gf1287_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I163 (wacks_0n[5], gf1287_0n[5], df_0n[5], gt1288_0n[5], dt_0n[5]);
  NOR2 I164 (dt_0n[5], df_0n[5], gf1287_0n[5]);
  NOR3 I165 (df_0n[5], dt_0n[5], gt1288_0n[5], init_0n);
  AND2 I166 (gt1288_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I167 (gf1287_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I168 (wacks_0n[4], gf1287_0n[4], df_0n[4], gt1288_0n[4], dt_0n[4]);
  NOR2 I169 (dt_0n[4], df_0n[4], gf1287_0n[4]);
  NOR3 I170 (df_0n[4], dt_0n[4], gt1288_0n[4], init_0n);
  AND2 I171 (gt1288_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I172 (gf1287_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I173 (wacks_0n[3], gf1287_0n[3], df_0n[3], gt1288_0n[3], dt_0n[3]);
  NOR2 I174 (dt_0n[3], df_0n[3], gf1287_0n[3]);
  NOR3 I175 (df_0n[3], dt_0n[3], gt1288_0n[3], init_0n);
  AND2 I176 (gt1288_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I177 (gf1287_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I178 (wacks_0n[2], gf1287_0n[2], df_0n[2], gt1288_0n[2], dt_0n[2]);
  NOR2 I179 (dt_0n[2], df_0n[2], gf1287_0n[2]);
  NOR3 I180 (df_0n[2], dt_0n[2], gt1288_0n[2], init_0n);
  AND2 I181 (gt1288_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I182 (gf1287_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I183 (wacks_0n[1], gf1287_0n[1], df_0n[1], gt1288_0n[1], dt_0n[1]);
  NOR2 I184 (dt_0n[1], df_0n[1], gf1287_0n[1]);
  NOR3 I185 (df_0n[1], dt_0n[1], gt1288_0n[1], init_0n);
  AND2 I186 (gt1288_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I187 (gf1287_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I188 (wacks_0n[0], gf1287_0n[0], df_0n[0], gt1288_0n[0], dt_0n[0]);
  NOR2 I189 (dt_0n[0], df_0n[0], gf1287_0n[0]);
  NOR3 I190 (df_0n[0], dt_0n[0], gt1288_0n[0], init_0n);
  AND2 I191 (gt1288_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I192 (gf1287_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I193 (init_0n, initialise);
endmodule

module BrzV_10_l6__28_29_l45__28_28_280_2010_29_2_m79m (
  wg_0r0d, wg_0r1d, wg_0a,
  wg_1r0d, wg_1r1d, wg_1a,
  wd_0r, wd_0a,
  wd_1r, wd_1a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  initialise
);
  input [9:0] wg_0r0d;
  input [9:0] wg_0r1d;
  output wg_0a;
  input [9:0] wg_1r0d;
  input [9:0] wg_1r1d;
  output wg_1a;
  output wd_0r;
  input wd_0a;
  output wd_1r;
  input wd_1a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [8:0] rd_0r0d;
  output [8:0] rd_0r1d;
  input rd_0a;
  output rd_1r0d;
  output rd_1r1d;
  input rd_1a;
  input initialise;
  wire [25:0] internal_0n;
  wire [9:0] wf_0n;
  wire [9:0] wt_0n;
  wire [9:0] df_0n;
  wire [9:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire wc_0n;
  wire wc_1n;
  wire [9:0] wacks_0n;
  wire wdrint_0n;
  wire wdrint_1n;
  wire wgaint_0n;
  wire wgaint_1n;
  wire [9:0] wgfint_0n;
  wire [9:0] wgfint_1n;
  wire [9:0] wgtint_0n;
  wire [9:0] wgtint_1n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire [8:0] rdfint_0n;
  wire rdfint_1n;
  wire [8:0] rdtint_0n;
  wire rdtint_1n;
  wire [9:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire igc_1n;
  wire ig_0n;
  wire ig_1n;
  wire [9:0] gif_0n;
  wire [9:0] gif_1n;
  wire [9:0] git_0n;
  wire [9:0] git_1n;
  wire [9:0] complete1301_0n;
  wire [9:0] complete1300_0n;
  wire [9:0] gt1299_0n;
  wire [9:0] gf1298_0n;
  assign rgaint_1n = rd_1a;
  assign rd_1r0d = rdfint_1n;
  assign rd_1r1d = rdtint_1n;
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign wg_1a = wgaint_1n;
  assign wgfint_1n[0] = wg_1r0d[0];
  assign wgfint_1n[1] = wg_1r0d[1];
  assign wgfint_1n[2] = wg_1r0d[2];
  assign wgfint_1n[3] = wg_1r0d[3];
  assign wgfint_1n[4] = wg_1r0d[4];
  assign wgfint_1n[5] = wg_1r0d[5];
  assign wgfint_1n[6] = wg_1r0d[6];
  assign wgfint_1n[7] = wg_1r0d[7];
  assign wgfint_1n[8] = wg_1r0d[8];
  assign wgfint_1n[9] = wg_1r0d[9];
  assign wgtint_1n[0] = wg_1r1d[0];
  assign wgtint_1n[1] = wg_1r1d[1];
  assign wgtint_1n[2] = wg_1r1d[2];
  assign wgtint_1n[3] = wg_1r1d[3];
  assign wgtint_1n[4] = wg_1r1d[4];
  assign wgtint_1n[5] = wg_1r1d[5];
  assign wgtint_1n[6] = wg_1r1d[6];
  assign wgtint_1n[7] = wg_1r1d[7];
  assign wgtint_1n[8] = wg_1r1d[8];
  assign wgtint_1n[9] = wg_1r1d[9];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_1n = wd_1a;
  assign wd_1r = wdrint_1n;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I72 (internal_0n[0], rgrint_0n, rgrint_1n);
  NOR2 I73 (internal_0n[1], rgaint_0n, rgaint_1n);
  AND2 I74 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I75 (rdtint_1n, rgrint_1n, dt_0n[0]);
  AND2 I76 (rdtint_0n[0], rgrint_0n, dt_0n[1]);
  AND2 I77 (rdtint_0n[1], rgrint_0n, dt_0n[2]);
  AND2 I78 (rdtint_0n[2], rgrint_0n, dt_0n[3]);
  AND2 I79 (rdtint_0n[3], rgrint_0n, dt_0n[4]);
  AND2 I80 (rdtint_0n[4], rgrint_0n, dt_0n[5]);
  AND2 I81 (rdtint_0n[5], rgrint_0n, dt_0n[6]);
  AND2 I82 (rdtint_0n[6], rgrint_0n, dt_0n[7]);
  AND2 I83 (rdtint_0n[7], rgrint_0n, dt_0n[8]);
  AND2 I84 (rdtint_0n[8], rgrint_0n, dt_0n[9]);
  AND2 I85 (rdfint_1n, rgrint_1n, df_0n[0]);
  AND2 I86 (rdfint_0n[0], rgrint_0n, df_0n[1]);
  AND2 I87 (rdfint_0n[1], rgrint_0n, df_0n[2]);
  AND2 I88 (rdfint_0n[2], rgrint_0n, df_0n[3]);
  AND2 I89 (rdfint_0n[3], rgrint_0n, df_0n[4]);
  AND2 I90 (rdfint_0n[4], rgrint_0n, df_0n[5]);
  AND2 I91 (rdfint_0n[5], rgrint_0n, df_0n[6]);
  AND2 I92 (rdfint_0n[6], rgrint_0n, df_0n[7]);
  AND2 I93 (rdfint_0n[7], rgrint_0n, df_0n[8]);
  AND2 I94 (rdfint_0n[8], rgrint_0n, df_0n[9]);
  C3 I95 (internal_0n[2], wc_1n, wacks_0n[9], wacks_0n[8]);
  C3 I96 (internal_0n[3], wacks_0n[7], wacks_0n[6], wacks_0n[5]);
  C3 I97 (internal_0n[4], wacks_0n[4], wacks_0n[3], wacks_0n[2]);
  C2 I98 (internal_0n[5], wacks_0n[1], wacks_0n[0]);
  C2 I99 (internal_0n[6], internal_0n[2], internal_0n[3]);
  C2 I100 (internal_0n[7], internal_0n[4], internal_0n[5]);
  C2 I101 (wdrint_1n, internal_0n[6], internal_0n[7]);
  C3 I102 (internal_0n[8], wc_0n, wacks_0n[9], wacks_0n[8]);
  C3 I103 (internal_0n[9], wacks_0n[7], wacks_0n[6], wacks_0n[5]);
  C3 I104 (internal_0n[10], wacks_0n[4], wacks_0n[3], wacks_0n[2]);
  C2 I105 (internal_0n[11], wacks_0n[1], wacks_0n[0]);
  C2 I106 (internal_0n[12], internal_0n[8], internal_0n[9]);
  C2 I107 (internal_0n[13], internal_0n[10], internal_0n[11]);
  C2 I108 (wdrint_0n, internal_0n[12], internal_0n[13]);
  OR2 I109 (wen_0n[9], wc_1n, wc_0n);
  OR2 I110 (wen_0n[8], wc_1n, wc_0n);
  OR2 I111 (wen_0n[7], wc_1n, wc_0n);
  OR2 I112 (wen_0n[6], wc_1n, wc_0n);
  OR2 I113 (wen_0n[5], wc_1n, wc_0n);
  OR2 I114 (wen_0n[4], wc_1n, wc_0n);
  OR2 I115 (wen_0n[3], wc_1n, wc_0n);
  OR2 I116 (wen_0n[2], wc_1n, wc_0n);
  OR2 I117 (wen_0n[1], wc_1n, wc_0n);
  OR2 I118 (wen_0n[0], wc_1n, wc_0n);
  OR2 I119 (wt_0n[9], git_1n[9], git_0n[9]);
  OR2 I120 (wt_0n[8], git_1n[8], git_0n[8]);
  OR2 I121 (wt_0n[7], git_1n[7], git_0n[7]);
  OR2 I122 (wt_0n[6], git_1n[6], git_0n[6]);
  OR2 I123 (wt_0n[5], git_1n[5], git_0n[5]);
  OR2 I124 (wt_0n[4], git_1n[4], git_0n[4]);
  OR2 I125 (wt_0n[3], git_1n[3], git_0n[3]);
  OR2 I126 (wt_0n[2], git_1n[2], git_0n[2]);
  OR2 I127 (wt_0n[1], git_1n[1], git_0n[1]);
  OR2 I128 (wt_0n[0], git_1n[0], git_0n[0]);
  OR2 I129 (wf_0n[9], gif_1n[9], gif_0n[9]);
  OR2 I130 (wf_0n[8], gif_1n[8], gif_0n[8]);
  OR2 I131 (wf_0n[7], gif_1n[7], gif_0n[7]);
  OR2 I132 (wf_0n[6], gif_1n[6], gif_0n[6]);
  OR2 I133 (wf_0n[5], gif_1n[5], gif_0n[5]);
  OR2 I134 (wf_0n[4], gif_1n[4], gif_0n[4]);
  OR2 I135 (wf_0n[3], gif_1n[3], gif_0n[3]);
  OR2 I136 (wf_0n[2], gif_1n[2], gif_0n[2]);
  OR2 I137 (wf_0n[1], gif_1n[1], gif_0n[1]);
  OR2 I138 (wf_0n[0], gif_1n[0], gif_0n[0]);
  AC2 I139 (ig_0n, igc_0n, nanyread_0n);
  AC2 I140 (ig_1n, igc_1n, nanyread_0n);
  assign igc_0n = wc_0n;
  assign igc_1n = wc_1n;
  AND2 I143 (git_1n[0], wgtint_1n[0], ig_1n);
  AND2 I144 (git_1n[1], wgtint_1n[1], ig_1n);
  AND2 I145 (git_1n[2], wgtint_1n[2], ig_1n);
  AND2 I146 (git_1n[3], wgtint_1n[3], ig_1n);
  AND2 I147 (git_1n[4], wgtint_1n[4], ig_1n);
  AND2 I148 (git_1n[5], wgtint_1n[5], ig_1n);
  AND2 I149 (git_1n[6], wgtint_1n[6], ig_1n);
  AND2 I150 (git_1n[7], wgtint_1n[7], ig_1n);
  AND2 I151 (git_1n[8], wgtint_1n[8], ig_1n);
  AND2 I152 (git_1n[9], wgtint_1n[9], ig_1n);
  AND2 I153 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I154 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I155 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I156 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I157 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I158 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I159 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I160 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I161 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I162 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I163 (gif_1n[0], wgfint_1n[0], ig_1n);
  AND2 I164 (gif_1n[1], wgfint_1n[1], ig_1n);
  AND2 I165 (gif_1n[2], wgfint_1n[2], ig_1n);
  AND2 I166 (gif_1n[3], wgfint_1n[3], ig_1n);
  AND2 I167 (gif_1n[4], wgfint_1n[4], ig_1n);
  AND2 I168 (gif_1n[5], wgfint_1n[5], ig_1n);
  AND2 I169 (gif_1n[6], wgfint_1n[6], ig_1n);
  AND2 I170 (gif_1n[7], wgfint_1n[7], ig_1n);
  AND2 I171 (gif_1n[8], wgfint_1n[8], ig_1n);
  AND2 I172 (gif_1n[9], wgfint_1n[9], ig_1n);
  AND2 I173 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I174 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I175 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I176 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I177 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I178 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I179 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I180 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I181 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I182 (gif_0n[9], wgfint_0n[9], ig_0n);
  C3 I183 (internal_0n[14], complete1301_0n[0], complete1301_0n[1], complete1301_0n[2]);
  C3 I184 (internal_0n[15], complete1301_0n[3], complete1301_0n[4], complete1301_0n[5]);
  C2 I185 (internal_0n[16], complete1301_0n[6], complete1301_0n[7]);
  C2 I186 (internal_0n[17], complete1301_0n[8], complete1301_0n[9]);
  C2 I187 (internal_0n[18], internal_0n[14], internal_0n[15]);
  C2 I188 (internal_0n[19], internal_0n[16], internal_0n[17]);
  C2 I189 (wc_1n, internal_0n[18], internal_0n[19]);
  OR2 I190 (complete1301_0n[0], wgfint_1n[0], wgtint_1n[0]);
  OR2 I191 (complete1301_0n[1], wgfint_1n[1], wgtint_1n[1]);
  OR2 I192 (complete1301_0n[2], wgfint_1n[2], wgtint_1n[2]);
  OR2 I193 (complete1301_0n[3], wgfint_1n[3], wgtint_1n[3]);
  OR2 I194 (complete1301_0n[4], wgfint_1n[4], wgtint_1n[4]);
  OR2 I195 (complete1301_0n[5], wgfint_1n[5], wgtint_1n[5]);
  OR2 I196 (complete1301_0n[6], wgfint_1n[6], wgtint_1n[6]);
  OR2 I197 (complete1301_0n[7], wgfint_1n[7], wgtint_1n[7]);
  OR2 I198 (complete1301_0n[8], wgfint_1n[8], wgtint_1n[8]);
  OR2 I199 (complete1301_0n[9], wgfint_1n[9], wgtint_1n[9]);
  C3 I200 (internal_0n[20], complete1300_0n[0], complete1300_0n[1], complete1300_0n[2]);
  C3 I201 (internal_0n[21], complete1300_0n[3], complete1300_0n[4], complete1300_0n[5]);
  C2 I202 (internal_0n[22], complete1300_0n[6], complete1300_0n[7]);
  C2 I203 (internal_0n[23], complete1300_0n[8], complete1300_0n[9]);
  C2 I204 (internal_0n[24], internal_0n[20], internal_0n[21]);
  C2 I205 (internal_0n[25], internal_0n[22], internal_0n[23]);
  C2 I206 (wc_0n, internal_0n[24], internal_0n[25]);
  OR2 I207 (complete1300_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I208 (complete1300_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I209 (complete1300_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I210 (complete1300_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I211 (complete1300_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I212 (complete1300_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I213 (complete1300_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I214 (complete1300_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I215 (complete1300_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I216 (complete1300_0n[9], wgfint_0n[9], wgtint_0n[9]);
  AO22 I217 (wacks_0n[9], gf1298_0n[9], df_0n[9], gt1299_0n[9], dt_0n[9]);
  NOR2 I218 (dt_0n[9], df_0n[9], gf1298_0n[9]);
  NOR3 I219 (df_0n[9], dt_0n[9], gt1299_0n[9], init_0n);
  AND2 I220 (gt1299_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I221 (gf1298_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I222 (wacks_0n[8], gf1298_0n[8], df_0n[8], gt1299_0n[8], dt_0n[8]);
  NOR2 I223 (dt_0n[8], df_0n[8], gf1298_0n[8]);
  NOR3 I224 (df_0n[8], dt_0n[8], gt1299_0n[8], init_0n);
  AND2 I225 (gt1299_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I226 (gf1298_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I227 (wacks_0n[7], gf1298_0n[7], df_0n[7], gt1299_0n[7], dt_0n[7]);
  NOR2 I228 (dt_0n[7], df_0n[7], gf1298_0n[7]);
  NOR3 I229 (df_0n[7], dt_0n[7], gt1299_0n[7], init_0n);
  AND2 I230 (gt1299_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I231 (gf1298_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I232 (wacks_0n[6], gf1298_0n[6], df_0n[6], gt1299_0n[6], dt_0n[6]);
  NOR2 I233 (dt_0n[6], df_0n[6], gf1298_0n[6]);
  NOR3 I234 (df_0n[6], dt_0n[6], gt1299_0n[6], init_0n);
  AND2 I235 (gt1299_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I236 (gf1298_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I237 (wacks_0n[5], gf1298_0n[5], df_0n[5], gt1299_0n[5], dt_0n[5]);
  NOR2 I238 (dt_0n[5], df_0n[5], gf1298_0n[5]);
  NOR3 I239 (df_0n[5], dt_0n[5], gt1299_0n[5], init_0n);
  AND2 I240 (gt1299_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I241 (gf1298_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I242 (wacks_0n[4], gf1298_0n[4], df_0n[4], gt1299_0n[4], dt_0n[4]);
  NOR2 I243 (dt_0n[4], df_0n[4], gf1298_0n[4]);
  NOR3 I244 (df_0n[4], dt_0n[4], gt1299_0n[4], init_0n);
  AND2 I245 (gt1299_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I246 (gf1298_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I247 (wacks_0n[3], gf1298_0n[3], df_0n[3], gt1299_0n[3], dt_0n[3]);
  NOR2 I248 (dt_0n[3], df_0n[3], gf1298_0n[3]);
  NOR3 I249 (df_0n[3], dt_0n[3], gt1299_0n[3], init_0n);
  AND2 I250 (gt1299_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I251 (gf1298_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I252 (wacks_0n[2], gf1298_0n[2], df_0n[2], gt1299_0n[2], dt_0n[2]);
  NOR2 I253 (dt_0n[2], df_0n[2], gf1298_0n[2]);
  NOR3 I254 (df_0n[2], dt_0n[2], gt1299_0n[2], init_0n);
  AND2 I255 (gt1299_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I256 (gf1298_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I257 (wacks_0n[1], gf1298_0n[1], df_0n[1], gt1299_0n[1], dt_0n[1]);
  NOR2 I258 (dt_0n[1], df_0n[1], gf1298_0n[1]);
  NOR3 I259 (df_0n[1], dt_0n[1], gt1299_0n[1], init_0n);
  AND2 I260 (gt1299_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I261 (gf1298_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I262 (wacks_0n[0], gf1298_0n[0], df_0n[0], gt1299_0n[0], dt_0n[0]);
  NOR2 I263 (dt_0n[0], df_0n[0], gf1298_0n[0]);
  NOR3 I264 (df_0n[0], dt_0n[0], gt1299_0n[0], init_0n);
  AND2 I265 (gt1299_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I266 (gf1298_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I267 (init_0n, initialise);
endmodule

module BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rd_0r0d, rd_0r1d, rd_0a,
  initialise
);
  input [31:0] wg_0r0d;
  input [31:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0d;
  output [31:0] rd_0r1d;
  input rd_0a;
  input initialise;
  wire [33:0] internal_0n;
  wire [31:0] wf_0n;
  wire [31:0] wt_0n;
  wire [31:0] df_0n;
  wire [31:0] dt_0n;
  wire rgrint_0n;
  wire wc_0n;
  wire [31:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [31:0] wgfint_0n;
  wire [31:0] wgtint_0n;
  wire rgaint_0n;
  wire [31:0] rdfint_0n;
  wire [31:0] rdtint_0n;
  wire [31:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [31:0] gif_0n;
  wire [31:0] git_0n;
  wire [31:0] complete1320_0n;
  wire [31:0] gt1319_0n;
  wire [31:0] gf1318_0n;
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r0d[10] = rdfint_0n[10];
  assign rd_0r0d[11] = rdfint_0n[11];
  assign rd_0r0d[12] = rdfint_0n[12];
  assign rd_0r0d[13] = rdfint_0n[13];
  assign rd_0r0d[14] = rdfint_0n[14];
  assign rd_0r0d[15] = rdfint_0n[15];
  assign rd_0r0d[16] = rdfint_0n[16];
  assign rd_0r0d[17] = rdfint_0n[17];
  assign rd_0r0d[18] = rdfint_0n[18];
  assign rd_0r0d[19] = rdfint_0n[19];
  assign rd_0r0d[20] = rdfint_0n[20];
  assign rd_0r0d[21] = rdfint_0n[21];
  assign rd_0r0d[22] = rdfint_0n[22];
  assign rd_0r0d[23] = rdfint_0n[23];
  assign rd_0r0d[24] = rdfint_0n[24];
  assign rd_0r0d[25] = rdfint_0n[25];
  assign rd_0r0d[26] = rdfint_0n[26];
  assign rd_0r0d[27] = rdfint_0n[27];
  assign rd_0r0d[28] = rdfint_0n[28];
  assign rd_0r0d[29] = rdfint_0n[29];
  assign rd_0r0d[30] = rdfint_0n[30];
  assign rd_0r0d[31] = rdfint_0n[31];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign rd_0r1d[10] = rdtint_0n[10];
  assign rd_0r1d[11] = rdtint_0n[11];
  assign rd_0r1d[12] = rdtint_0n[12];
  assign rd_0r1d[13] = rdtint_0n[13];
  assign rd_0r1d[14] = rdtint_0n[14];
  assign rd_0r1d[15] = rdtint_0n[15];
  assign rd_0r1d[16] = rdtint_0n[16];
  assign rd_0r1d[17] = rdtint_0n[17];
  assign rd_0r1d[18] = rdtint_0n[18];
  assign rd_0r1d[19] = rdtint_0n[19];
  assign rd_0r1d[20] = rdtint_0n[20];
  assign rd_0r1d[21] = rdtint_0n[21];
  assign rd_0r1d[22] = rdtint_0n[22];
  assign rd_0r1d[23] = rdtint_0n[23];
  assign rd_0r1d[24] = rdtint_0n[24];
  assign rd_0r1d[25] = rdtint_0n[25];
  assign rd_0r1d[26] = rdtint_0n[26];
  assign rd_0r1d[27] = rdtint_0n[27];
  assign rd_0r1d[28] = rdtint_0n[28];
  assign rd_0r1d[29] = rdtint_0n[29];
  assign rd_0r1d[30] = rdtint_0n[30];
  assign rd_0r1d[31] = rdtint_0n[31];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I134 (nanyread_0n, rgrint_0n, rgaint_0n);
  AND2 I135 (rdtint_0n[0], rgrint_0n, dt_0n[0]);
  AND2 I136 (rdtint_0n[1], rgrint_0n, dt_0n[1]);
  AND2 I137 (rdtint_0n[2], rgrint_0n, dt_0n[2]);
  AND2 I138 (rdtint_0n[3], rgrint_0n, dt_0n[3]);
  AND2 I139 (rdtint_0n[4], rgrint_0n, dt_0n[4]);
  AND2 I140 (rdtint_0n[5], rgrint_0n, dt_0n[5]);
  AND2 I141 (rdtint_0n[6], rgrint_0n, dt_0n[6]);
  AND2 I142 (rdtint_0n[7], rgrint_0n, dt_0n[7]);
  AND2 I143 (rdtint_0n[8], rgrint_0n, dt_0n[8]);
  AND2 I144 (rdtint_0n[9], rgrint_0n, dt_0n[9]);
  AND2 I145 (rdtint_0n[10], rgrint_0n, dt_0n[10]);
  AND2 I146 (rdtint_0n[11], rgrint_0n, dt_0n[11]);
  AND2 I147 (rdtint_0n[12], rgrint_0n, dt_0n[12]);
  AND2 I148 (rdtint_0n[13], rgrint_0n, dt_0n[13]);
  AND2 I149 (rdtint_0n[14], rgrint_0n, dt_0n[14]);
  AND2 I150 (rdtint_0n[15], rgrint_0n, dt_0n[15]);
  AND2 I151 (rdtint_0n[16], rgrint_0n, dt_0n[16]);
  AND2 I152 (rdtint_0n[17], rgrint_0n, dt_0n[17]);
  AND2 I153 (rdtint_0n[18], rgrint_0n, dt_0n[18]);
  AND2 I154 (rdtint_0n[19], rgrint_0n, dt_0n[19]);
  AND2 I155 (rdtint_0n[20], rgrint_0n, dt_0n[20]);
  AND2 I156 (rdtint_0n[21], rgrint_0n, dt_0n[21]);
  AND2 I157 (rdtint_0n[22], rgrint_0n, dt_0n[22]);
  AND2 I158 (rdtint_0n[23], rgrint_0n, dt_0n[23]);
  AND2 I159 (rdtint_0n[24], rgrint_0n, dt_0n[24]);
  AND2 I160 (rdtint_0n[25], rgrint_0n, dt_0n[25]);
  AND2 I161 (rdtint_0n[26], rgrint_0n, dt_0n[26]);
  AND2 I162 (rdtint_0n[27], rgrint_0n, dt_0n[27]);
  AND2 I163 (rdtint_0n[28], rgrint_0n, dt_0n[28]);
  AND2 I164 (rdtint_0n[29], rgrint_0n, dt_0n[29]);
  AND2 I165 (rdtint_0n[30], rgrint_0n, dt_0n[30]);
  AND2 I166 (rdtint_0n[31], rgrint_0n, dt_0n[31]);
  AND2 I167 (rdfint_0n[0], rgrint_0n, df_0n[0]);
  AND2 I168 (rdfint_0n[1], rgrint_0n, df_0n[1]);
  AND2 I169 (rdfint_0n[2], rgrint_0n, df_0n[2]);
  AND2 I170 (rdfint_0n[3], rgrint_0n, df_0n[3]);
  AND2 I171 (rdfint_0n[4], rgrint_0n, df_0n[4]);
  AND2 I172 (rdfint_0n[5], rgrint_0n, df_0n[5]);
  AND2 I173 (rdfint_0n[6], rgrint_0n, df_0n[6]);
  AND2 I174 (rdfint_0n[7], rgrint_0n, df_0n[7]);
  AND2 I175 (rdfint_0n[8], rgrint_0n, df_0n[8]);
  AND2 I176 (rdfint_0n[9], rgrint_0n, df_0n[9]);
  AND2 I177 (rdfint_0n[10], rgrint_0n, df_0n[10]);
  AND2 I178 (rdfint_0n[11], rgrint_0n, df_0n[11]);
  AND2 I179 (rdfint_0n[12], rgrint_0n, df_0n[12]);
  AND2 I180 (rdfint_0n[13], rgrint_0n, df_0n[13]);
  AND2 I181 (rdfint_0n[14], rgrint_0n, df_0n[14]);
  AND2 I182 (rdfint_0n[15], rgrint_0n, df_0n[15]);
  AND2 I183 (rdfint_0n[16], rgrint_0n, df_0n[16]);
  AND2 I184 (rdfint_0n[17], rgrint_0n, df_0n[17]);
  AND2 I185 (rdfint_0n[18], rgrint_0n, df_0n[18]);
  AND2 I186 (rdfint_0n[19], rgrint_0n, df_0n[19]);
  AND2 I187 (rdfint_0n[20], rgrint_0n, df_0n[20]);
  AND2 I188 (rdfint_0n[21], rgrint_0n, df_0n[21]);
  AND2 I189 (rdfint_0n[22], rgrint_0n, df_0n[22]);
  AND2 I190 (rdfint_0n[23], rgrint_0n, df_0n[23]);
  AND2 I191 (rdfint_0n[24], rgrint_0n, df_0n[24]);
  AND2 I192 (rdfint_0n[25], rgrint_0n, df_0n[25]);
  AND2 I193 (rdfint_0n[26], rgrint_0n, df_0n[26]);
  AND2 I194 (rdfint_0n[27], rgrint_0n, df_0n[27]);
  AND2 I195 (rdfint_0n[28], rgrint_0n, df_0n[28]);
  AND2 I196 (rdfint_0n[29], rgrint_0n, df_0n[29]);
  AND2 I197 (rdfint_0n[30], rgrint_0n, df_0n[30]);
  AND2 I198 (rdfint_0n[31], rgrint_0n, df_0n[31]);
  C3 I199 (internal_0n[0], wc_0n, wacks_0n[31], wacks_0n[30]);
  C3 I200 (internal_0n[1], wacks_0n[29], wacks_0n[28], wacks_0n[27]);
  C3 I201 (internal_0n[2], wacks_0n[26], wacks_0n[25], wacks_0n[24]);
  C3 I202 (internal_0n[3], wacks_0n[23], wacks_0n[22], wacks_0n[21]);
  C3 I203 (internal_0n[4], wacks_0n[20], wacks_0n[19], wacks_0n[18]);
  C3 I204 (internal_0n[5], wacks_0n[17], wacks_0n[16], wacks_0n[15]);
  C3 I205 (internal_0n[6], wacks_0n[14], wacks_0n[13], wacks_0n[12]);
  C3 I206 (internal_0n[7], wacks_0n[11], wacks_0n[10], wacks_0n[9]);
  C3 I207 (internal_0n[8], wacks_0n[8], wacks_0n[7], wacks_0n[6]);
  C3 I208 (internal_0n[9], wacks_0n[5], wacks_0n[4], wacks_0n[3]);
  C3 I209 (internal_0n[10], wacks_0n[2], wacks_0n[1], wacks_0n[0]);
  C3 I210 (internal_0n[11], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I211 (internal_0n[12], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I212 (internal_0n[13], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I213 (internal_0n[14], internal_0n[9], internal_0n[10]);
  C2 I214 (internal_0n[15], internal_0n[11], internal_0n[12]);
  C2 I215 (internal_0n[16], internal_0n[13], internal_0n[14]);
  C2 I216 (wdrint_0n, internal_0n[15], internal_0n[16]);
  assign wen_0n[31] = wc_0n;
  assign wen_0n[30] = wc_0n;
  assign wen_0n[29] = wc_0n;
  assign wen_0n[28] = wc_0n;
  assign wen_0n[27] = wc_0n;
  assign wen_0n[26] = wc_0n;
  assign wen_0n[25] = wc_0n;
  assign wen_0n[24] = wc_0n;
  assign wen_0n[23] = wc_0n;
  assign wen_0n[22] = wc_0n;
  assign wen_0n[21] = wc_0n;
  assign wen_0n[20] = wc_0n;
  assign wen_0n[19] = wc_0n;
  assign wen_0n[18] = wc_0n;
  assign wen_0n[17] = wc_0n;
  assign wen_0n[16] = wc_0n;
  assign wen_0n[15] = wc_0n;
  assign wen_0n[14] = wc_0n;
  assign wen_0n[13] = wc_0n;
  assign wen_0n[12] = wc_0n;
  assign wen_0n[11] = wc_0n;
  assign wen_0n[10] = wc_0n;
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[31] = git_0n[31];
  assign wt_0n[30] = git_0n[30];
  assign wt_0n[29] = git_0n[29];
  assign wt_0n[28] = git_0n[28];
  assign wt_0n[27] = git_0n[27];
  assign wt_0n[26] = git_0n[26];
  assign wt_0n[25] = git_0n[25];
  assign wt_0n[24] = git_0n[24];
  assign wt_0n[23] = git_0n[23];
  assign wt_0n[22] = git_0n[22];
  assign wt_0n[21] = git_0n[21];
  assign wt_0n[20] = git_0n[20];
  assign wt_0n[19] = git_0n[19];
  assign wt_0n[18] = git_0n[18];
  assign wt_0n[17] = git_0n[17];
  assign wt_0n[16] = git_0n[16];
  assign wt_0n[15] = git_0n[15];
  assign wt_0n[14] = git_0n[14];
  assign wt_0n[13] = git_0n[13];
  assign wt_0n[12] = git_0n[12];
  assign wt_0n[11] = git_0n[11];
  assign wt_0n[10] = git_0n[10];
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[31] = gif_0n[31];
  assign wf_0n[30] = gif_0n[30];
  assign wf_0n[29] = gif_0n[29];
  assign wf_0n[28] = gif_0n[28];
  assign wf_0n[27] = gif_0n[27];
  assign wf_0n[26] = gif_0n[26];
  assign wf_0n[25] = gif_0n[25];
  assign wf_0n[24] = gif_0n[24];
  assign wf_0n[23] = gif_0n[23];
  assign wf_0n[22] = gif_0n[22];
  assign wf_0n[21] = gif_0n[21];
  assign wf_0n[20] = gif_0n[20];
  assign wf_0n[19] = gif_0n[19];
  assign wf_0n[18] = gif_0n[18];
  assign wf_0n[17] = gif_0n[17];
  assign wf_0n[16] = gif_0n[16];
  assign wf_0n[15] = gif_0n[15];
  assign wf_0n[14] = gif_0n[14];
  assign wf_0n[13] = gif_0n[13];
  assign wf_0n[12] = gif_0n[12];
  assign wf_0n[11] = gif_0n[11];
  assign wf_0n[10] = gif_0n[10];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I313 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I315 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I316 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I317 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I318 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I319 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I320 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I321 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I322 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I323 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I324 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I325 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I326 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I327 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I328 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I329 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I330 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I331 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I332 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I333 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I334 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I335 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I336 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I337 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I338 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I339 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I340 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I341 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I342 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I343 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I344 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I345 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I346 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I347 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I348 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I349 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I350 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I351 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I352 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I353 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I354 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I355 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I356 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I357 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I358 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I359 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I360 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I361 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I362 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I363 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I364 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I365 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I366 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I367 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I368 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I369 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I370 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I371 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I372 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I373 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I374 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I375 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I376 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I377 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I378 (gif_0n[31], wgfint_0n[31], ig_0n);
  C3 I379 (internal_0n[17], complete1320_0n[0], complete1320_0n[1], complete1320_0n[2]);
  C3 I380 (internal_0n[18], complete1320_0n[3], complete1320_0n[4], complete1320_0n[5]);
  C3 I381 (internal_0n[19], complete1320_0n[6], complete1320_0n[7], complete1320_0n[8]);
  C3 I382 (internal_0n[20], complete1320_0n[9], complete1320_0n[10], complete1320_0n[11]);
  C3 I383 (internal_0n[21], complete1320_0n[12], complete1320_0n[13], complete1320_0n[14]);
  C3 I384 (internal_0n[22], complete1320_0n[15], complete1320_0n[16], complete1320_0n[17]);
  C3 I385 (internal_0n[23], complete1320_0n[18], complete1320_0n[19], complete1320_0n[20]);
  C3 I386 (internal_0n[24], complete1320_0n[21], complete1320_0n[22], complete1320_0n[23]);
  C3 I387 (internal_0n[25], complete1320_0n[24], complete1320_0n[25], complete1320_0n[26]);
  C3 I388 (internal_0n[26], complete1320_0n[27], complete1320_0n[28], complete1320_0n[29]);
  C2 I389 (internal_0n[27], complete1320_0n[30], complete1320_0n[31]);
  C3 I390 (internal_0n[28], internal_0n[17], internal_0n[18], internal_0n[19]);
  C3 I391 (internal_0n[29], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I392 (internal_0n[30], internal_0n[23], internal_0n[24], internal_0n[25]);
  C2 I393 (internal_0n[31], internal_0n[26], internal_0n[27]);
  C2 I394 (internal_0n[32], internal_0n[28], internal_0n[29]);
  C2 I395 (internal_0n[33], internal_0n[30], internal_0n[31]);
  C2 I396 (wc_0n, internal_0n[32], internal_0n[33]);
  OR2 I397 (complete1320_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I398 (complete1320_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I399 (complete1320_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I400 (complete1320_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I401 (complete1320_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I402 (complete1320_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I403 (complete1320_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I404 (complete1320_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I405 (complete1320_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I406 (complete1320_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I407 (complete1320_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I408 (complete1320_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I409 (complete1320_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I410 (complete1320_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I411 (complete1320_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I412 (complete1320_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I413 (complete1320_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I414 (complete1320_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I415 (complete1320_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I416 (complete1320_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I417 (complete1320_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I418 (complete1320_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I419 (complete1320_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I420 (complete1320_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I421 (complete1320_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I422 (complete1320_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I423 (complete1320_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I424 (complete1320_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I425 (complete1320_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I426 (complete1320_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I427 (complete1320_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I428 (complete1320_0n[31], wgfint_0n[31], wgtint_0n[31]);
  AO22 I429 (wacks_0n[31], gf1318_0n[31], df_0n[31], gt1319_0n[31], dt_0n[31]);
  NOR2 I430 (dt_0n[31], df_0n[31], gf1318_0n[31]);
  NOR3 I431 (df_0n[31], dt_0n[31], gt1319_0n[31], init_0n);
  AND2 I432 (gt1319_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I433 (gf1318_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I434 (wacks_0n[30], gf1318_0n[30], df_0n[30], gt1319_0n[30], dt_0n[30]);
  NOR2 I435 (dt_0n[30], df_0n[30], gf1318_0n[30]);
  NOR3 I436 (df_0n[30], dt_0n[30], gt1319_0n[30], init_0n);
  AND2 I437 (gt1319_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I438 (gf1318_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I439 (wacks_0n[29], gf1318_0n[29], df_0n[29], gt1319_0n[29], dt_0n[29]);
  NOR2 I440 (dt_0n[29], df_0n[29], gf1318_0n[29]);
  NOR3 I441 (df_0n[29], dt_0n[29], gt1319_0n[29], init_0n);
  AND2 I442 (gt1319_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I443 (gf1318_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I444 (wacks_0n[28], gf1318_0n[28], df_0n[28], gt1319_0n[28], dt_0n[28]);
  NOR2 I445 (dt_0n[28], df_0n[28], gf1318_0n[28]);
  NOR3 I446 (df_0n[28], dt_0n[28], gt1319_0n[28], init_0n);
  AND2 I447 (gt1319_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I448 (gf1318_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I449 (wacks_0n[27], gf1318_0n[27], df_0n[27], gt1319_0n[27], dt_0n[27]);
  NOR2 I450 (dt_0n[27], df_0n[27], gf1318_0n[27]);
  NOR3 I451 (df_0n[27], dt_0n[27], gt1319_0n[27], init_0n);
  AND2 I452 (gt1319_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I453 (gf1318_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I454 (wacks_0n[26], gf1318_0n[26], df_0n[26], gt1319_0n[26], dt_0n[26]);
  NOR2 I455 (dt_0n[26], df_0n[26], gf1318_0n[26]);
  NOR3 I456 (df_0n[26], dt_0n[26], gt1319_0n[26], init_0n);
  AND2 I457 (gt1319_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I458 (gf1318_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I459 (wacks_0n[25], gf1318_0n[25], df_0n[25], gt1319_0n[25], dt_0n[25]);
  NOR2 I460 (dt_0n[25], df_0n[25], gf1318_0n[25]);
  NOR3 I461 (df_0n[25], dt_0n[25], gt1319_0n[25], init_0n);
  AND2 I462 (gt1319_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I463 (gf1318_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I464 (wacks_0n[24], gf1318_0n[24], df_0n[24], gt1319_0n[24], dt_0n[24]);
  NOR2 I465 (dt_0n[24], df_0n[24], gf1318_0n[24]);
  NOR3 I466 (df_0n[24], dt_0n[24], gt1319_0n[24], init_0n);
  AND2 I467 (gt1319_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I468 (gf1318_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I469 (wacks_0n[23], gf1318_0n[23], df_0n[23], gt1319_0n[23], dt_0n[23]);
  NOR2 I470 (dt_0n[23], df_0n[23], gf1318_0n[23]);
  NOR3 I471 (df_0n[23], dt_0n[23], gt1319_0n[23], init_0n);
  AND2 I472 (gt1319_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I473 (gf1318_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I474 (wacks_0n[22], gf1318_0n[22], df_0n[22], gt1319_0n[22], dt_0n[22]);
  NOR2 I475 (dt_0n[22], df_0n[22], gf1318_0n[22]);
  NOR3 I476 (df_0n[22], dt_0n[22], gt1319_0n[22], init_0n);
  AND2 I477 (gt1319_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I478 (gf1318_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I479 (wacks_0n[21], gf1318_0n[21], df_0n[21], gt1319_0n[21], dt_0n[21]);
  NOR2 I480 (dt_0n[21], df_0n[21], gf1318_0n[21]);
  NOR3 I481 (df_0n[21], dt_0n[21], gt1319_0n[21], init_0n);
  AND2 I482 (gt1319_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I483 (gf1318_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I484 (wacks_0n[20], gf1318_0n[20], df_0n[20], gt1319_0n[20], dt_0n[20]);
  NOR2 I485 (dt_0n[20], df_0n[20], gf1318_0n[20]);
  NOR3 I486 (df_0n[20], dt_0n[20], gt1319_0n[20], init_0n);
  AND2 I487 (gt1319_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I488 (gf1318_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I489 (wacks_0n[19], gf1318_0n[19], df_0n[19], gt1319_0n[19], dt_0n[19]);
  NOR2 I490 (dt_0n[19], df_0n[19], gf1318_0n[19]);
  NOR3 I491 (df_0n[19], dt_0n[19], gt1319_0n[19], init_0n);
  AND2 I492 (gt1319_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I493 (gf1318_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I494 (wacks_0n[18], gf1318_0n[18], df_0n[18], gt1319_0n[18], dt_0n[18]);
  NOR2 I495 (dt_0n[18], df_0n[18], gf1318_0n[18]);
  NOR3 I496 (df_0n[18], dt_0n[18], gt1319_0n[18], init_0n);
  AND2 I497 (gt1319_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I498 (gf1318_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I499 (wacks_0n[17], gf1318_0n[17], df_0n[17], gt1319_0n[17], dt_0n[17]);
  NOR2 I500 (dt_0n[17], df_0n[17], gf1318_0n[17]);
  NOR3 I501 (df_0n[17], dt_0n[17], gt1319_0n[17], init_0n);
  AND2 I502 (gt1319_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I503 (gf1318_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I504 (wacks_0n[16], gf1318_0n[16], df_0n[16], gt1319_0n[16], dt_0n[16]);
  NOR2 I505 (dt_0n[16], df_0n[16], gf1318_0n[16]);
  NOR3 I506 (df_0n[16], dt_0n[16], gt1319_0n[16], init_0n);
  AND2 I507 (gt1319_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I508 (gf1318_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I509 (wacks_0n[15], gf1318_0n[15], df_0n[15], gt1319_0n[15], dt_0n[15]);
  NOR2 I510 (dt_0n[15], df_0n[15], gf1318_0n[15]);
  NOR3 I511 (df_0n[15], dt_0n[15], gt1319_0n[15], init_0n);
  AND2 I512 (gt1319_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I513 (gf1318_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I514 (wacks_0n[14], gf1318_0n[14], df_0n[14], gt1319_0n[14], dt_0n[14]);
  NOR2 I515 (dt_0n[14], df_0n[14], gf1318_0n[14]);
  NOR3 I516 (df_0n[14], dt_0n[14], gt1319_0n[14], init_0n);
  AND2 I517 (gt1319_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I518 (gf1318_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I519 (wacks_0n[13], gf1318_0n[13], df_0n[13], gt1319_0n[13], dt_0n[13]);
  NOR2 I520 (dt_0n[13], df_0n[13], gf1318_0n[13]);
  NOR3 I521 (df_0n[13], dt_0n[13], gt1319_0n[13], init_0n);
  AND2 I522 (gt1319_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I523 (gf1318_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I524 (wacks_0n[12], gf1318_0n[12], df_0n[12], gt1319_0n[12], dt_0n[12]);
  NOR2 I525 (dt_0n[12], df_0n[12], gf1318_0n[12]);
  NOR3 I526 (df_0n[12], dt_0n[12], gt1319_0n[12], init_0n);
  AND2 I527 (gt1319_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I528 (gf1318_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I529 (wacks_0n[11], gf1318_0n[11], df_0n[11], gt1319_0n[11], dt_0n[11]);
  NOR2 I530 (dt_0n[11], df_0n[11], gf1318_0n[11]);
  NOR3 I531 (df_0n[11], dt_0n[11], gt1319_0n[11], init_0n);
  AND2 I532 (gt1319_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I533 (gf1318_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I534 (wacks_0n[10], gf1318_0n[10], df_0n[10], gt1319_0n[10], dt_0n[10]);
  NOR2 I535 (dt_0n[10], df_0n[10], gf1318_0n[10]);
  NOR3 I536 (df_0n[10], dt_0n[10], gt1319_0n[10], init_0n);
  AND2 I537 (gt1319_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I538 (gf1318_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I539 (wacks_0n[9], gf1318_0n[9], df_0n[9], gt1319_0n[9], dt_0n[9]);
  NOR2 I540 (dt_0n[9], df_0n[9], gf1318_0n[9]);
  NOR3 I541 (df_0n[9], dt_0n[9], gt1319_0n[9], init_0n);
  AND2 I542 (gt1319_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I543 (gf1318_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I544 (wacks_0n[8], gf1318_0n[8], df_0n[8], gt1319_0n[8], dt_0n[8]);
  NOR2 I545 (dt_0n[8], df_0n[8], gf1318_0n[8]);
  NOR3 I546 (df_0n[8], dt_0n[8], gt1319_0n[8], init_0n);
  AND2 I547 (gt1319_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I548 (gf1318_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I549 (wacks_0n[7], gf1318_0n[7], df_0n[7], gt1319_0n[7], dt_0n[7]);
  NOR2 I550 (dt_0n[7], df_0n[7], gf1318_0n[7]);
  NOR3 I551 (df_0n[7], dt_0n[7], gt1319_0n[7], init_0n);
  AND2 I552 (gt1319_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I553 (gf1318_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I554 (wacks_0n[6], gf1318_0n[6], df_0n[6], gt1319_0n[6], dt_0n[6]);
  NOR2 I555 (dt_0n[6], df_0n[6], gf1318_0n[6]);
  NOR3 I556 (df_0n[6], dt_0n[6], gt1319_0n[6], init_0n);
  AND2 I557 (gt1319_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I558 (gf1318_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I559 (wacks_0n[5], gf1318_0n[5], df_0n[5], gt1319_0n[5], dt_0n[5]);
  NOR2 I560 (dt_0n[5], df_0n[5], gf1318_0n[5]);
  NOR3 I561 (df_0n[5], dt_0n[5], gt1319_0n[5], init_0n);
  AND2 I562 (gt1319_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I563 (gf1318_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I564 (wacks_0n[4], gf1318_0n[4], df_0n[4], gt1319_0n[4], dt_0n[4]);
  NOR2 I565 (dt_0n[4], df_0n[4], gf1318_0n[4]);
  NOR3 I566 (df_0n[4], dt_0n[4], gt1319_0n[4], init_0n);
  AND2 I567 (gt1319_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I568 (gf1318_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I569 (wacks_0n[3], gf1318_0n[3], df_0n[3], gt1319_0n[3], dt_0n[3]);
  NOR2 I570 (dt_0n[3], df_0n[3], gf1318_0n[3]);
  NOR3 I571 (df_0n[3], dt_0n[3], gt1319_0n[3], init_0n);
  AND2 I572 (gt1319_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I573 (gf1318_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I574 (wacks_0n[2], gf1318_0n[2], df_0n[2], gt1319_0n[2], dt_0n[2]);
  NOR2 I575 (dt_0n[2], df_0n[2], gf1318_0n[2]);
  NOR3 I576 (df_0n[2], dt_0n[2], gt1319_0n[2], init_0n);
  AND2 I577 (gt1319_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I578 (gf1318_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I579 (wacks_0n[1], gf1318_0n[1], df_0n[1], gt1319_0n[1], dt_0n[1]);
  NOR2 I580 (dt_0n[1], df_0n[1], gf1318_0n[1]);
  NOR3 I581 (df_0n[1], dt_0n[1], gt1319_0n[1], init_0n);
  AND2 I582 (gt1319_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I583 (gf1318_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I584 (wacks_0n[0], gf1318_0n[0], df_0n[0], gt1319_0n[0], dt_0n[0]);
  NOR2 I585 (dt_0n[0], df_0n[0], gf1318_0n[0]);
  NOR3 I586 (df_0n[0], dt_0n[0], gt1319_0n[0], init_0n);
  AND2 I587 (gt1319_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I588 (gf1318_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I589 (init_0n, initialise);
endmodule

module BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m81m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  initialise
);
  input [31:0] wg_0r0d;
  input [31:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [31:0] rd_0r0d;
  output [31:0] rd_0r1d;
  input rd_0a;
  output [31:0] rd_1r0d;
  output [31:0] rd_1r1d;
  input rd_1a;
  input initialise;
  wire [35:0] internal_0n;
  wire [31:0] wf_0n;
  wire [31:0] wt_0n;
  wire [31:0] df_0n;
  wire [31:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire wc_0n;
  wire [31:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [31:0] wgfint_0n;
  wire [31:0] wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire [31:0] rdfint_0n;
  wire [31:0] rdfint_1n;
  wire [31:0] rdtint_0n;
  wire [31:0] rdtint_1n;
  wire [31:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [31:0] gif_0n;
  wire [31:0] git_0n;
  wire [31:0] complete1331_0n;
  wire [31:0] gt1330_0n;
  wire [31:0] gf1329_0n;
  assign rgaint_1n = rd_1a;
  assign rd_1r0d[0] = rdfint_1n[0];
  assign rd_1r0d[1] = rdfint_1n[1];
  assign rd_1r0d[2] = rdfint_1n[2];
  assign rd_1r0d[3] = rdfint_1n[3];
  assign rd_1r0d[4] = rdfint_1n[4];
  assign rd_1r0d[5] = rdfint_1n[5];
  assign rd_1r0d[6] = rdfint_1n[6];
  assign rd_1r0d[7] = rdfint_1n[7];
  assign rd_1r0d[8] = rdfint_1n[8];
  assign rd_1r0d[9] = rdfint_1n[9];
  assign rd_1r0d[10] = rdfint_1n[10];
  assign rd_1r0d[11] = rdfint_1n[11];
  assign rd_1r0d[12] = rdfint_1n[12];
  assign rd_1r0d[13] = rdfint_1n[13];
  assign rd_1r0d[14] = rdfint_1n[14];
  assign rd_1r0d[15] = rdfint_1n[15];
  assign rd_1r0d[16] = rdfint_1n[16];
  assign rd_1r0d[17] = rdfint_1n[17];
  assign rd_1r0d[18] = rdfint_1n[18];
  assign rd_1r0d[19] = rdfint_1n[19];
  assign rd_1r0d[20] = rdfint_1n[20];
  assign rd_1r0d[21] = rdfint_1n[21];
  assign rd_1r0d[22] = rdfint_1n[22];
  assign rd_1r0d[23] = rdfint_1n[23];
  assign rd_1r0d[24] = rdfint_1n[24];
  assign rd_1r0d[25] = rdfint_1n[25];
  assign rd_1r0d[26] = rdfint_1n[26];
  assign rd_1r0d[27] = rdfint_1n[27];
  assign rd_1r0d[28] = rdfint_1n[28];
  assign rd_1r0d[29] = rdfint_1n[29];
  assign rd_1r0d[30] = rdfint_1n[30];
  assign rd_1r0d[31] = rdfint_1n[31];
  assign rd_1r1d[0] = rdtint_1n[0];
  assign rd_1r1d[1] = rdtint_1n[1];
  assign rd_1r1d[2] = rdtint_1n[2];
  assign rd_1r1d[3] = rdtint_1n[3];
  assign rd_1r1d[4] = rdtint_1n[4];
  assign rd_1r1d[5] = rdtint_1n[5];
  assign rd_1r1d[6] = rdtint_1n[6];
  assign rd_1r1d[7] = rdtint_1n[7];
  assign rd_1r1d[8] = rdtint_1n[8];
  assign rd_1r1d[9] = rdtint_1n[9];
  assign rd_1r1d[10] = rdtint_1n[10];
  assign rd_1r1d[11] = rdtint_1n[11];
  assign rd_1r1d[12] = rdtint_1n[12];
  assign rd_1r1d[13] = rdtint_1n[13];
  assign rd_1r1d[14] = rdtint_1n[14];
  assign rd_1r1d[15] = rdtint_1n[15];
  assign rd_1r1d[16] = rdtint_1n[16];
  assign rd_1r1d[17] = rdtint_1n[17];
  assign rd_1r1d[18] = rdtint_1n[18];
  assign rd_1r1d[19] = rdtint_1n[19];
  assign rd_1r1d[20] = rdtint_1n[20];
  assign rd_1r1d[21] = rdtint_1n[21];
  assign rd_1r1d[22] = rdtint_1n[22];
  assign rd_1r1d[23] = rdtint_1n[23];
  assign rd_1r1d[24] = rdtint_1n[24];
  assign rd_1r1d[25] = rdtint_1n[25];
  assign rd_1r1d[26] = rdtint_1n[26];
  assign rd_1r1d[27] = rdtint_1n[27];
  assign rd_1r1d[28] = rdtint_1n[28];
  assign rd_1r1d[29] = rdtint_1n[29];
  assign rd_1r1d[30] = rdtint_1n[30];
  assign rd_1r1d[31] = rdtint_1n[31];
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r0d[10] = rdfint_0n[10];
  assign rd_0r0d[11] = rdfint_0n[11];
  assign rd_0r0d[12] = rdfint_0n[12];
  assign rd_0r0d[13] = rdfint_0n[13];
  assign rd_0r0d[14] = rdfint_0n[14];
  assign rd_0r0d[15] = rdfint_0n[15];
  assign rd_0r0d[16] = rdfint_0n[16];
  assign rd_0r0d[17] = rdfint_0n[17];
  assign rd_0r0d[18] = rdfint_0n[18];
  assign rd_0r0d[19] = rdfint_0n[19];
  assign rd_0r0d[20] = rdfint_0n[20];
  assign rd_0r0d[21] = rdfint_0n[21];
  assign rd_0r0d[22] = rdfint_0n[22];
  assign rd_0r0d[23] = rdfint_0n[23];
  assign rd_0r0d[24] = rdfint_0n[24];
  assign rd_0r0d[25] = rdfint_0n[25];
  assign rd_0r0d[26] = rdfint_0n[26];
  assign rd_0r0d[27] = rdfint_0n[27];
  assign rd_0r0d[28] = rdfint_0n[28];
  assign rd_0r0d[29] = rdfint_0n[29];
  assign rd_0r0d[30] = rdfint_0n[30];
  assign rd_0r0d[31] = rdfint_0n[31];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign rd_0r1d[10] = rdtint_0n[10];
  assign rd_0r1d[11] = rdtint_0n[11];
  assign rd_0r1d[12] = rdtint_0n[12];
  assign rd_0r1d[13] = rdtint_0n[13];
  assign rd_0r1d[14] = rdtint_0n[14];
  assign rd_0r1d[15] = rdtint_0n[15];
  assign rd_0r1d[16] = rdtint_0n[16];
  assign rd_0r1d[17] = rdtint_0n[17];
  assign rd_0r1d[18] = rdtint_0n[18];
  assign rd_0r1d[19] = rdtint_0n[19];
  assign rd_0r1d[20] = rdtint_0n[20];
  assign rd_0r1d[21] = rdtint_0n[21];
  assign rd_0r1d[22] = rdtint_0n[22];
  assign rd_0r1d[23] = rdtint_0n[23];
  assign rd_0r1d[24] = rdtint_0n[24];
  assign rd_0r1d[25] = rdtint_0n[25];
  assign rd_0r1d[26] = rdtint_0n[26];
  assign rd_0r1d[27] = rdtint_0n[27];
  assign rd_0r1d[28] = rdtint_0n[28];
  assign rd_0r1d[29] = rdtint_0n[29];
  assign rd_0r1d[30] = rdtint_0n[30];
  assign rd_0r1d[31] = rdtint_0n[31];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I201 (internal_0n[0], rgrint_0n, rgrint_1n);
  NOR2 I202 (internal_0n[1], rgaint_0n, rgaint_1n);
  AND2 I203 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I204 (rdtint_1n[0], rgrint_1n, dt_0n[0]);
  AND2 I205 (rdtint_1n[1], rgrint_1n, dt_0n[1]);
  AND2 I206 (rdtint_1n[2], rgrint_1n, dt_0n[2]);
  AND2 I207 (rdtint_1n[3], rgrint_1n, dt_0n[3]);
  AND2 I208 (rdtint_1n[4], rgrint_1n, dt_0n[4]);
  AND2 I209 (rdtint_1n[5], rgrint_1n, dt_0n[5]);
  AND2 I210 (rdtint_1n[6], rgrint_1n, dt_0n[6]);
  AND2 I211 (rdtint_1n[7], rgrint_1n, dt_0n[7]);
  AND2 I212 (rdtint_1n[8], rgrint_1n, dt_0n[8]);
  AND2 I213 (rdtint_1n[9], rgrint_1n, dt_0n[9]);
  AND2 I214 (rdtint_1n[10], rgrint_1n, dt_0n[10]);
  AND2 I215 (rdtint_1n[11], rgrint_1n, dt_0n[11]);
  AND2 I216 (rdtint_1n[12], rgrint_1n, dt_0n[12]);
  AND2 I217 (rdtint_1n[13], rgrint_1n, dt_0n[13]);
  AND2 I218 (rdtint_1n[14], rgrint_1n, dt_0n[14]);
  AND2 I219 (rdtint_1n[15], rgrint_1n, dt_0n[15]);
  AND2 I220 (rdtint_1n[16], rgrint_1n, dt_0n[16]);
  AND2 I221 (rdtint_1n[17], rgrint_1n, dt_0n[17]);
  AND2 I222 (rdtint_1n[18], rgrint_1n, dt_0n[18]);
  AND2 I223 (rdtint_1n[19], rgrint_1n, dt_0n[19]);
  AND2 I224 (rdtint_1n[20], rgrint_1n, dt_0n[20]);
  AND2 I225 (rdtint_1n[21], rgrint_1n, dt_0n[21]);
  AND2 I226 (rdtint_1n[22], rgrint_1n, dt_0n[22]);
  AND2 I227 (rdtint_1n[23], rgrint_1n, dt_0n[23]);
  AND2 I228 (rdtint_1n[24], rgrint_1n, dt_0n[24]);
  AND2 I229 (rdtint_1n[25], rgrint_1n, dt_0n[25]);
  AND2 I230 (rdtint_1n[26], rgrint_1n, dt_0n[26]);
  AND2 I231 (rdtint_1n[27], rgrint_1n, dt_0n[27]);
  AND2 I232 (rdtint_1n[28], rgrint_1n, dt_0n[28]);
  AND2 I233 (rdtint_1n[29], rgrint_1n, dt_0n[29]);
  AND2 I234 (rdtint_1n[30], rgrint_1n, dt_0n[30]);
  AND2 I235 (rdtint_1n[31], rgrint_1n, dt_0n[31]);
  AND2 I236 (rdtint_0n[0], rgrint_0n, dt_0n[0]);
  AND2 I237 (rdtint_0n[1], rgrint_0n, dt_0n[1]);
  AND2 I238 (rdtint_0n[2], rgrint_0n, dt_0n[2]);
  AND2 I239 (rdtint_0n[3], rgrint_0n, dt_0n[3]);
  AND2 I240 (rdtint_0n[4], rgrint_0n, dt_0n[4]);
  AND2 I241 (rdtint_0n[5], rgrint_0n, dt_0n[5]);
  AND2 I242 (rdtint_0n[6], rgrint_0n, dt_0n[6]);
  AND2 I243 (rdtint_0n[7], rgrint_0n, dt_0n[7]);
  AND2 I244 (rdtint_0n[8], rgrint_0n, dt_0n[8]);
  AND2 I245 (rdtint_0n[9], rgrint_0n, dt_0n[9]);
  AND2 I246 (rdtint_0n[10], rgrint_0n, dt_0n[10]);
  AND2 I247 (rdtint_0n[11], rgrint_0n, dt_0n[11]);
  AND2 I248 (rdtint_0n[12], rgrint_0n, dt_0n[12]);
  AND2 I249 (rdtint_0n[13], rgrint_0n, dt_0n[13]);
  AND2 I250 (rdtint_0n[14], rgrint_0n, dt_0n[14]);
  AND2 I251 (rdtint_0n[15], rgrint_0n, dt_0n[15]);
  AND2 I252 (rdtint_0n[16], rgrint_0n, dt_0n[16]);
  AND2 I253 (rdtint_0n[17], rgrint_0n, dt_0n[17]);
  AND2 I254 (rdtint_0n[18], rgrint_0n, dt_0n[18]);
  AND2 I255 (rdtint_0n[19], rgrint_0n, dt_0n[19]);
  AND2 I256 (rdtint_0n[20], rgrint_0n, dt_0n[20]);
  AND2 I257 (rdtint_0n[21], rgrint_0n, dt_0n[21]);
  AND2 I258 (rdtint_0n[22], rgrint_0n, dt_0n[22]);
  AND2 I259 (rdtint_0n[23], rgrint_0n, dt_0n[23]);
  AND2 I260 (rdtint_0n[24], rgrint_0n, dt_0n[24]);
  AND2 I261 (rdtint_0n[25], rgrint_0n, dt_0n[25]);
  AND2 I262 (rdtint_0n[26], rgrint_0n, dt_0n[26]);
  AND2 I263 (rdtint_0n[27], rgrint_0n, dt_0n[27]);
  AND2 I264 (rdtint_0n[28], rgrint_0n, dt_0n[28]);
  AND2 I265 (rdtint_0n[29], rgrint_0n, dt_0n[29]);
  AND2 I266 (rdtint_0n[30], rgrint_0n, dt_0n[30]);
  AND2 I267 (rdtint_0n[31], rgrint_0n, dt_0n[31]);
  AND2 I268 (rdfint_1n[0], rgrint_1n, df_0n[0]);
  AND2 I269 (rdfint_1n[1], rgrint_1n, df_0n[1]);
  AND2 I270 (rdfint_1n[2], rgrint_1n, df_0n[2]);
  AND2 I271 (rdfint_1n[3], rgrint_1n, df_0n[3]);
  AND2 I272 (rdfint_1n[4], rgrint_1n, df_0n[4]);
  AND2 I273 (rdfint_1n[5], rgrint_1n, df_0n[5]);
  AND2 I274 (rdfint_1n[6], rgrint_1n, df_0n[6]);
  AND2 I275 (rdfint_1n[7], rgrint_1n, df_0n[7]);
  AND2 I276 (rdfint_1n[8], rgrint_1n, df_0n[8]);
  AND2 I277 (rdfint_1n[9], rgrint_1n, df_0n[9]);
  AND2 I278 (rdfint_1n[10], rgrint_1n, df_0n[10]);
  AND2 I279 (rdfint_1n[11], rgrint_1n, df_0n[11]);
  AND2 I280 (rdfint_1n[12], rgrint_1n, df_0n[12]);
  AND2 I281 (rdfint_1n[13], rgrint_1n, df_0n[13]);
  AND2 I282 (rdfint_1n[14], rgrint_1n, df_0n[14]);
  AND2 I283 (rdfint_1n[15], rgrint_1n, df_0n[15]);
  AND2 I284 (rdfint_1n[16], rgrint_1n, df_0n[16]);
  AND2 I285 (rdfint_1n[17], rgrint_1n, df_0n[17]);
  AND2 I286 (rdfint_1n[18], rgrint_1n, df_0n[18]);
  AND2 I287 (rdfint_1n[19], rgrint_1n, df_0n[19]);
  AND2 I288 (rdfint_1n[20], rgrint_1n, df_0n[20]);
  AND2 I289 (rdfint_1n[21], rgrint_1n, df_0n[21]);
  AND2 I290 (rdfint_1n[22], rgrint_1n, df_0n[22]);
  AND2 I291 (rdfint_1n[23], rgrint_1n, df_0n[23]);
  AND2 I292 (rdfint_1n[24], rgrint_1n, df_0n[24]);
  AND2 I293 (rdfint_1n[25], rgrint_1n, df_0n[25]);
  AND2 I294 (rdfint_1n[26], rgrint_1n, df_0n[26]);
  AND2 I295 (rdfint_1n[27], rgrint_1n, df_0n[27]);
  AND2 I296 (rdfint_1n[28], rgrint_1n, df_0n[28]);
  AND2 I297 (rdfint_1n[29], rgrint_1n, df_0n[29]);
  AND2 I298 (rdfint_1n[30], rgrint_1n, df_0n[30]);
  AND2 I299 (rdfint_1n[31], rgrint_1n, df_0n[31]);
  AND2 I300 (rdfint_0n[0], rgrint_0n, df_0n[0]);
  AND2 I301 (rdfint_0n[1], rgrint_0n, df_0n[1]);
  AND2 I302 (rdfint_0n[2], rgrint_0n, df_0n[2]);
  AND2 I303 (rdfint_0n[3], rgrint_0n, df_0n[3]);
  AND2 I304 (rdfint_0n[4], rgrint_0n, df_0n[4]);
  AND2 I305 (rdfint_0n[5], rgrint_0n, df_0n[5]);
  AND2 I306 (rdfint_0n[6], rgrint_0n, df_0n[6]);
  AND2 I307 (rdfint_0n[7], rgrint_0n, df_0n[7]);
  AND2 I308 (rdfint_0n[8], rgrint_0n, df_0n[8]);
  AND2 I309 (rdfint_0n[9], rgrint_0n, df_0n[9]);
  AND2 I310 (rdfint_0n[10], rgrint_0n, df_0n[10]);
  AND2 I311 (rdfint_0n[11], rgrint_0n, df_0n[11]);
  AND2 I312 (rdfint_0n[12], rgrint_0n, df_0n[12]);
  AND2 I313 (rdfint_0n[13], rgrint_0n, df_0n[13]);
  AND2 I314 (rdfint_0n[14], rgrint_0n, df_0n[14]);
  AND2 I315 (rdfint_0n[15], rgrint_0n, df_0n[15]);
  AND2 I316 (rdfint_0n[16], rgrint_0n, df_0n[16]);
  AND2 I317 (rdfint_0n[17], rgrint_0n, df_0n[17]);
  AND2 I318 (rdfint_0n[18], rgrint_0n, df_0n[18]);
  AND2 I319 (rdfint_0n[19], rgrint_0n, df_0n[19]);
  AND2 I320 (rdfint_0n[20], rgrint_0n, df_0n[20]);
  AND2 I321 (rdfint_0n[21], rgrint_0n, df_0n[21]);
  AND2 I322 (rdfint_0n[22], rgrint_0n, df_0n[22]);
  AND2 I323 (rdfint_0n[23], rgrint_0n, df_0n[23]);
  AND2 I324 (rdfint_0n[24], rgrint_0n, df_0n[24]);
  AND2 I325 (rdfint_0n[25], rgrint_0n, df_0n[25]);
  AND2 I326 (rdfint_0n[26], rgrint_0n, df_0n[26]);
  AND2 I327 (rdfint_0n[27], rgrint_0n, df_0n[27]);
  AND2 I328 (rdfint_0n[28], rgrint_0n, df_0n[28]);
  AND2 I329 (rdfint_0n[29], rgrint_0n, df_0n[29]);
  AND2 I330 (rdfint_0n[30], rgrint_0n, df_0n[30]);
  AND2 I331 (rdfint_0n[31], rgrint_0n, df_0n[31]);
  C3 I332 (internal_0n[2], wc_0n, wacks_0n[31], wacks_0n[30]);
  C3 I333 (internal_0n[3], wacks_0n[29], wacks_0n[28], wacks_0n[27]);
  C3 I334 (internal_0n[4], wacks_0n[26], wacks_0n[25], wacks_0n[24]);
  C3 I335 (internal_0n[5], wacks_0n[23], wacks_0n[22], wacks_0n[21]);
  C3 I336 (internal_0n[6], wacks_0n[20], wacks_0n[19], wacks_0n[18]);
  C3 I337 (internal_0n[7], wacks_0n[17], wacks_0n[16], wacks_0n[15]);
  C3 I338 (internal_0n[8], wacks_0n[14], wacks_0n[13], wacks_0n[12]);
  C3 I339 (internal_0n[9], wacks_0n[11], wacks_0n[10], wacks_0n[9]);
  C3 I340 (internal_0n[10], wacks_0n[8], wacks_0n[7], wacks_0n[6]);
  C3 I341 (internal_0n[11], wacks_0n[5], wacks_0n[4], wacks_0n[3]);
  C3 I342 (internal_0n[12], wacks_0n[2], wacks_0n[1], wacks_0n[0]);
  C3 I343 (internal_0n[13], internal_0n[2], internal_0n[3], internal_0n[4]);
  C3 I344 (internal_0n[14], internal_0n[5], internal_0n[6], internal_0n[7]);
  C3 I345 (internal_0n[15], internal_0n[8], internal_0n[9], internal_0n[10]);
  C2 I346 (internal_0n[16], internal_0n[11], internal_0n[12]);
  C2 I347 (internal_0n[17], internal_0n[13], internal_0n[14]);
  C2 I348 (internal_0n[18], internal_0n[15], internal_0n[16]);
  C2 I349 (wdrint_0n, internal_0n[17], internal_0n[18]);
  assign wen_0n[31] = wc_0n;
  assign wen_0n[30] = wc_0n;
  assign wen_0n[29] = wc_0n;
  assign wen_0n[28] = wc_0n;
  assign wen_0n[27] = wc_0n;
  assign wen_0n[26] = wc_0n;
  assign wen_0n[25] = wc_0n;
  assign wen_0n[24] = wc_0n;
  assign wen_0n[23] = wc_0n;
  assign wen_0n[22] = wc_0n;
  assign wen_0n[21] = wc_0n;
  assign wen_0n[20] = wc_0n;
  assign wen_0n[19] = wc_0n;
  assign wen_0n[18] = wc_0n;
  assign wen_0n[17] = wc_0n;
  assign wen_0n[16] = wc_0n;
  assign wen_0n[15] = wc_0n;
  assign wen_0n[14] = wc_0n;
  assign wen_0n[13] = wc_0n;
  assign wen_0n[12] = wc_0n;
  assign wen_0n[11] = wc_0n;
  assign wen_0n[10] = wc_0n;
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[31] = git_0n[31];
  assign wt_0n[30] = git_0n[30];
  assign wt_0n[29] = git_0n[29];
  assign wt_0n[28] = git_0n[28];
  assign wt_0n[27] = git_0n[27];
  assign wt_0n[26] = git_0n[26];
  assign wt_0n[25] = git_0n[25];
  assign wt_0n[24] = git_0n[24];
  assign wt_0n[23] = git_0n[23];
  assign wt_0n[22] = git_0n[22];
  assign wt_0n[21] = git_0n[21];
  assign wt_0n[20] = git_0n[20];
  assign wt_0n[19] = git_0n[19];
  assign wt_0n[18] = git_0n[18];
  assign wt_0n[17] = git_0n[17];
  assign wt_0n[16] = git_0n[16];
  assign wt_0n[15] = git_0n[15];
  assign wt_0n[14] = git_0n[14];
  assign wt_0n[13] = git_0n[13];
  assign wt_0n[12] = git_0n[12];
  assign wt_0n[11] = git_0n[11];
  assign wt_0n[10] = git_0n[10];
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[31] = gif_0n[31];
  assign wf_0n[30] = gif_0n[30];
  assign wf_0n[29] = gif_0n[29];
  assign wf_0n[28] = gif_0n[28];
  assign wf_0n[27] = gif_0n[27];
  assign wf_0n[26] = gif_0n[26];
  assign wf_0n[25] = gif_0n[25];
  assign wf_0n[24] = gif_0n[24];
  assign wf_0n[23] = gif_0n[23];
  assign wf_0n[22] = gif_0n[22];
  assign wf_0n[21] = gif_0n[21];
  assign wf_0n[20] = gif_0n[20];
  assign wf_0n[19] = gif_0n[19];
  assign wf_0n[18] = gif_0n[18];
  assign wf_0n[17] = gif_0n[17];
  assign wf_0n[16] = gif_0n[16];
  assign wf_0n[15] = gif_0n[15];
  assign wf_0n[14] = gif_0n[14];
  assign wf_0n[13] = gif_0n[13];
  assign wf_0n[12] = gif_0n[12];
  assign wf_0n[11] = gif_0n[11];
  assign wf_0n[10] = gif_0n[10];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I446 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I448 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I449 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I450 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I451 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I452 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I453 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I454 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I455 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I456 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I457 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I458 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I459 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I460 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I461 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I462 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I463 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I464 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I465 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I466 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I467 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I468 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I469 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I470 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I471 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I472 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I473 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I474 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I475 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I476 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I477 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I478 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I479 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I480 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I481 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I482 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I483 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I484 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I485 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I486 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I487 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I488 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I489 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I490 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I491 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I492 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I493 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I494 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I495 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I496 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I497 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I498 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I499 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I500 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I501 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I502 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I503 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I504 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I505 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I506 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I507 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I508 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I509 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I510 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I511 (gif_0n[31], wgfint_0n[31], ig_0n);
  C3 I512 (internal_0n[19], complete1331_0n[0], complete1331_0n[1], complete1331_0n[2]);
  C3 I513 (internal_0n[20], complete1331_0n[3], complete1331_0n[4], complete1331_0n[5]);
  C3 I514 (internal_0n[21], complete1331_0n[6], complete1331_0n[7], complete1331_0n[8]);
  C3 I515 (internal_0n[22], complete1331_0n[9], complete1331_0n[10], complete1331_0n[11]);
  C3 I516 (internal_0n[23], complete1331_0n[12], complete1331_0n[13], complete1331_0n[14]);
  C3 I517 (internal_0n[24], complete1331_0n[15], complete1331_0n[16], complete1331_0n[17]);
  C3 I518 (internal_0n[25], complete1331_0n[18], complete1331_0n[19], complete1331_0n[20]);
  C3 I519 (internal_0n[26], complete1331_0n[21], complete1331_0n[22], complete1331_0n[23]);
  C3 I520 (internal_0n[27], complete1331_0n[24], complete1331_0n[25], complete1331_0n[26]);
  C3 I521 (internal_0n[28], complete1331_0n[27], complete1331_0n[28], complete1331_0n[29]);
  C2 I522 (internal_0n[29], complete1331_0n[30], complete1331_0n[31]);
  C3 I523 (internal_0n[30], internal_0n[19], internal_0n[20], internal_0n[21]);
  C3 I524 (internal_0n[31], internal_0n[22], internal_0n[23], internal_0n[24]);
  C3 I525 (internal_0n[32], internal_0n[25], internal_0n[26], internal_0n[27]);
  C2 I526 (internal_0n[33], internal_0n[28], internal_0n[29]);
  C2 I527 (internal_0n[34], internal_0n[30], internal_0n[31]);
  C2 I528 (internal_0n[35], internal_0n[32], internal_0n[33]);
  C2 I529 (wc_0n, internal_0n[34], internal_0n[35]);
  OR2 I530 (complete1331_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I531 (complete1331_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I532 (complete1331_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I533 (complete1331_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I534 (complete1331_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I535 (complete1331_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I536 (complete1331_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I537 (complete1331_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I538 (complete1331_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I539 (complete1331_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I540 (complete1331_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I541 (complete1331_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I542 (complete1331_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I543 (complete1331_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I544 (complete1331_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I545 (complete1331_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I546 (complete1331_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I547 (complete1331_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I548 (complete1331_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I549 (complete1331_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I550 (complete1331_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I551 (complete1331_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I552 (complete1331_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I553 (complete1331_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I554 (complete1331_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I555 (complete1331_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I556 (complete1331_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I557 (complete1331_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I558 (complete1331_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I559 (complete1331_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I560 (complete1331_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I561 (complete1331_0n[31], wgfint_0n[31], wgtint_0n[31]);
  AO22 I562 (wacks_0n[31], gf1329_0n[31], df_0n[31], gt1330_0n[31], dt_0n[31]);
  NOR2 I563 (dt_0n[31], df_0n[31], gf1329_0n[31]);
  NOR3 I564 (df_0n[31], dt_0n[31], gt1330_0n[31], init_0n);
  AND2 I565 (gt1330_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I566 (gf1329_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I567 (wacks_0n[30], gf1329_0n[30], df_0n[30], gt1330_0n[30], dt_0n[30]);
  NOR2 I568 (dt_0n[30], df_0n[30], gf1329_0n[30]);
  NOR3 I569 (df_0n[30], dt_0n[30], gt1330_0n[30], init_0n);
  AND2 I570 (gt1330_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I571 (gf1329_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I572 (wacks_0n[29], gf1329_0n[29], df_0n[29], gt1330_0n[29], dt_0n[29]);
  NOR2 I573 (dt_0n[29], df_0n[29], gf1329_0n[29]);
  NOR3 I574 (df_0n[29], dt_0n[29], gt1330_0n[29], init_0n);
  AND2 I575 (gt1330_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I576 (gf1329_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I577 (wacks_0n[28], gf1329_0n[28], df_0n[28], gt1330_0n[28], dt_0n[28]);
  NOR2 I578 (dt_0n[28], df_0n[28], gf1329_0n[28]);
  NOR3 I579 (df_0n[28], dt_0n[28], gt1330_0n[28], init_0n);
  AND2 I580 (gt1330_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I581 (gf1329_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I582 (wacks_0n[27], gf1329_0n[27], df_0n[27], gt1330_0n[27], dt_0n[27]);
  NOR2 I583 (dt_0n[27], df_0n[27], gf1329_0n[27]);
  NOR3 I584 (df_0n[27], dt_0n[27], gt1330_0n[27], init_0n);
  AND2 I585 (gt1330_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I586 (gf1329_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I587 (wacks_0n[26], gf1329_0n[26], df_0n[26], gt1330_0n[26], dt_0n[26]);
  NOR2 I588 (dt_0n[26], df_0n[26], gf1329_0n[26]);
  NOR3 I589 (df_0n[26], dt_0n[26], gt1330_0n[26], init_0n);
  AND2 I590 (gt1330_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I591 (gf1329_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I592 (wacks_0n[25], gf1329_0n[25], df_0n[25], gt1330_0n[25], dt_0n[25]);
  NOR2 I593 (dt_0n[25], df_0n[25], gf1329_0n[25]);
  NOR3 I594 (df_0n[25], dt_0n[25], gt1330_0n[25], init_0n);
  AND2 I595 (gt1330_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I596 (gf1329_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I597 (wacks_0n[24], gf1329_0n[24], df_0n[24], gt1330_0n[24], dt_0n[24]);
  NOR2 I598 (dt_0n[24], df_0n[24], gf1329_0n[24]);
  NOR3 I599 (df_0n[24], dt_0n[24], gt1330_0n[24], init_0n);
  AND2 I600 (gt1330_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I601 (gf1329_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I602 (wacks_0n[23], gf1329_0n[23], df_0n[23], gt1330_0n[23], dt_0n[23]);
  NOR2 I603 (dt_0n[23], df_0n[23], gf1329_0n[23]);
  NOR3 I604 (df_0n[23], dt_0n[23], gt1330_0n[23], init_0n);
  AND2 I605 (gt1330_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I606 (gf1329_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I607 (wacks_0n[22], gf1329_0n[22], df_0n[22], gt1330_0n[22], dt_0n[22]);
  NOR2 I608 (dt_0n[22], df_0n[22], gf1329_0n[22]);
  NOR3 I609 (df_0n[22], dt_0n[22], gt1330_0n[22], init_0n);
  AND2 I610 (gt1330_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I611 (gf1329_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I612 (wacks_0n[21], gf1329_0n[21], df_0n[21], gt1330_0n[21], dt_0n[21]);
  NOR2 I613 (dt_0n[21], df_0n[21], gf1329_0n[21]);
  NOR3 I614 (df_0n[21], dt_0n[21], gt1330_0n[21], init_0n);
  AND2 I615 (gt1330_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I616 (gf1329_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I617 (wacks_0n[20], gf1329_0n[20], df_0n[20], gt1330_0n[20], dt_0n[20]);
  NOR2 I618 (dt_0n[20], df_0n[20], gf1329_0n[20]);
  NOR3 I619 (df_0n[20], dt_0n[20], gt1330_0n[20], init_0n);
  AND2 I620 (gt1330_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I621 (gf1329_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I622 (wacks_0n[19], gf1329_0n[19], df_0n[19], gt1330_0n[19], dt_0n[19]);
  NOR2 I623 (dt_0n[19], df_0n[19], gf1329_0n[19]);
  NOR3 I624 (df_0n[19], dt_0n[19], gt1330_0n[19], init_0n);
  AND2 I625 (gt1330_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I626 (gf1329_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I627 (wacks_0n[18], gf1329_0n[18], df_0n[18], gt1330_0n[18], dt_0n[18]);
  NOR2 I628 (dt_0n[18], df_0n[18], gf1329_0n[18]);
  NOR3 I629 (df_0n[18], dt_0n[18], gt1330_0n[18], init_0n);
  AND2 I630 (gt1330_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I631 (gf1329_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I632 (wacks_0n[17], gf1329_0n[17], df_0n[17], gt1330_0n[17], dt_0n[17]);
  NOR2 I633 (dt_0n[17], df_0n[17], gf1329_0n[17]);
  NOR3 I634 (df_0n[17], dt_0n[17], gt1330_0n[17], init_0n);
  AND2 I635 (gt1330_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I636 (gf1329_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I637 (wacks_0n[16], gf1329_0n[16], df_0n[16], gt1330_0n[16], dt_0n[16]);
  NOR2 I638 (dt_0n[16], df_0n[16], gf1329_0n[16]);
  NOR3 I639 (df_0n[16], dt_0n[16], gt1330_0n[16], init_0n);
  AND2 I640 (gt1330_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I641 (gf1329_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I642 (wacks_0n[15], gf1329_0n[15], df_0n[15], gt1330_0n[15], dt_0n[15]);
  NOR2 I643 (dt_0n[15], df_0n[15], gf1329_0n[15]);
  NOR3 I644 (df_0n[15], dt_0n[15], gt1330_0n[15], init_0n);
  AND2 I645 (gt1330_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I646 (gf1329_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I647 (wacks_0n[14], gf1329_0n[14], df_0n[14], gt1330_0n[14], dt_0n[14]);
  NOR2 I648 (dt_0n[14], df_0n[14], gf1329_0n[14]);
  NOR3 I649 (df_0n[14], dt_0n[14], gt1330_0n[14], init_0n);
  AND2 I650 (gt1330_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I651 (gf1329_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I652 (wacks_0n[13], gf1329_0n[13], df_0n[13], gt1330_0n[13], dt_0n[13]);
  NOR2 I653 (dt_0n[13], df_0n[13], gf1329_0n[13]);
  NOR3 I654 (df_0n[13], dt_0n[13], gt1330_0n[13], init_0n);
  AND2 I655 (gt1330_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I656 (gf1329_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I657 (wacks_0n[12], gf1329_0n[12], df_0n[12], gt1330_0n[12], dt_0n[12]);
  NOR2 I658 (dt_0n[12], df_0n[12], gf1329_0n[12]);
  NOR3 I659 (df_0n[12], dt_0n[12], gt1330_0n[12], init_0n);
  AND2 I660 (gt1330_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I661 (gf1329_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I662 (wacks_0n[11], gf1329_0n[11], df_0n[11], gt1330_0n[11], dt_0n[11]);
  NOR2 I663 (dt_0n[11], df_0n[11], gf1329_0n[11]);
  NOR3 I664 (df_0n[11], dt_0n[11], gt1330_0n[11], init_0n);
  AND2 I665 (gt1330_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I666 (gf1329_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I667 (wacks_0n[10], gf1329_0n[10], df_0n[10], gt1330_0n[10], dt_0n[10]);
  NOR2 I668 (dt_0n[10], df_0n[10], gf1329_0n[10]);
  NOR3 I669 (df_0n[10], dt_0n[10], gt1330_0n[10], init_0n);
  AND2 I670 (gt1330_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I671 (gf1329_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I672 (wacks_0n[9], gf1329_0n[9], df_0n[9], gt1330_0n[9], dt_0n[9]);
  NOR2 I673 (dt_0n[9], df_0n[9], gf1329_0n[9]);
  NOR3 I674 (df_0n[9], dt_0n[9], gt1330_0n[9], init_0n);
  AND2 I675 (gt1330_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I676 (gf1329_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I677 (wacks_0n[8], gf1329_0n[8], df_0n[8], gt1330_0n[8], dt_0n[8]);
  NOR2 I678 (dt_0n[8], df_0n[8], gf1329_0n[8]);
  NOR3 I679 (df_0n[8], dt_0n[8], gt1330_0n[8], init_0n);
  AND2 I680 (gt1330_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I681 (gf1329_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I682 (wacks_0n[7], gf1329_0n[7], df_0n[7], gt1330_0n[7], dt_0n[7]);
  NOR2 I683 (dt_0n[7], df_0n[7], gf1329_0n[7]);
  NOR3 I684 (df_0n[7], dt_0n[7], gt1330_0n[7], init_0n);
  AND2 I685 (gt1330_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I686 (gf1329_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I687 (wacks_0n[6], gf1329_0n[6], df_0n[6], gt1330_0n[6], dt_0n[6]);
  NOR2 I688 (dt_0n[6], df_0n[6], gf1329_0n[6]);
  NOR3 I689 (df_0n[6], dt_0n[6], gt1330_0n[6], init_0n);
  AND2 I690 (gt1330_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I691 (gf1329_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I692 (wacks_0n[5], gf1329_0n[5], df_0n[5], gt1330_0n[5], dt_0n[5]);
  NOR2 I693 (dt_0n[5], df_0n[5], gf1329_0n[5]);
  NOR3 I694 (df_0n[5], dt_0n[5], gt1330_0n[5], init_0n);
  AND2 I695 (gt1330_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I696 (gf1329_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I697 (wacks_0n[4], gf1329_0n[4], df_0n[4], gt1330_0n[4], dt_0n[4]);
  NOR2 I698 (dt_0n[4], df_0n[4], gf1329_0n[4]);
  NOR3 I699 (df_0n[4], dt_0n[4], gt1330_0n[4], init_0n);
  AND2 I700 (gt1330_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I701 (gf1329_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I702 (wacks_0n[3], gf1329_0n[3], df_0n[3], gt1330_0n[3], dt_0n[3]);
  NOR2 I703 (dt_0n[3], df_0n[3], gf1329_0n[3]);
  NOR3 I704 (df_0n[3], dt_0n[3], gt1330_0n[3], init_0n);
  AND2 I705 (gt1330_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I706 (gf1329_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I707 (wacks_0n[2], gf1329_0n[2], df_0n[2], gt1330_0n[2], dt_0n[2]);
  NOR2 I708 (dt_0n[2], df_0n[2], gf1329_0n[2]);
  NOR3 I709 (df_0n[2], dt_0n[2], gt1330_0n[2], init_0n);
  AND2 I710 (gt1330_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I711 (gf1329_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I712 (wacks_0n[1], gf1329_0n[1], df_0n[1], gt1330_0n[1], dt_0n[1]);
  NOR2 I713 (dt_0n[1], df_0n[1], gf1329_0n[1]);
  NOR3 I714 (df_0n[1], dt_0n[1], gt1330_0n[1], init_0n);
  AND2 I715 (gt1330_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I716 (gf1329_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I717 (wacks_0n[0], gf1329_0n[0], df_0n[0], gt1330_0n[0], dt_0n[0]);
  NOR2 I718 (dt_0n[0], df_0n[0], gf1329_0n[0]);
  NOR3 I719 (df_0n[0], dt_0n[0], gt1330_0n[0], init_0n);
  AND2 I720 (gt1330_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I721 (gf1329_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I722 (init_0n, initialise);
endmodule

module BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m82m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rg_2r, rg_2a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  rd_2r0d, rd_2r1d, rd_2a,
  initialise
);
  input [31:0] wg_0r0d;
  input [31:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0d;
  output [31:0] rd_0r1d;
  input rd_0a;
  output rd_1r0d;
  output rd_1r1d;
  input rd_1a;
  output [31:0] rd_2r0d;
  output [31:0] rd_2r1d;
  input rd_2a;
  input initialise;
  wire [35:0] internal_0n;
  wire [31:0] wf_0n;
  wire [31:0] wt_0n;
  wire [31:0] df_0n;
  wire [31:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire rgrint_2n;
  wire wc_0n;
  wire [31:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [31:0] wgfint_0n;
  wire [31:0] wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire rgaint_2n;
  wire [31:0] rdfint_0n;
  wire rdfint_1n;
  wire [31:0] rdfint_2n;
  wire [31:0] rdtint_0n;
  wire rdtint_1n;
  wire [31:0] rdtint_2n;
  wire [31:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [31:0] gif_0n;
  wire [31:0] git_0n;
  wire [31:0] complete1346_0n;
  wire [31:0] gt1345_0n;
  wire [31:0] gf1344_0n;
  assign rgaint_2n = rd_2a;
  assign rd_2r0d[0] = rdfint_2n[0];
  assign rd_2r0d[1] = rdfint_2n[1];
  assign rd_2r0d[2] = rdfint_2n[2];
  assign rd_2r0d[3] = rdfint_2n[3];
  assign rd_2r0d[4] = rdfint_2n[4];
  assign rd_2r0d[5] = rdfint_2n[5];
  assign rd_2r0d[6] = rdfint_2n[6];
  assign rd_2r0d[7] = rdfint_2n[7];
  assign rd_2r0d[8] = rdfint_2n[8];
  assign rd_2r0d[9] = rdfint_2n[9];
  assign rd_2r0d[10] = rdfint_2n[10];
  assign rd_2r0d[11] = rdfint_2n[11];
  assign rd_2r0d[12] = rdfint_2n[12];
  assign rd_2r0d[13] = rdfint_2n[13];
  assign rd_2r0d[14] = rdfint_2n[14];
  assign rd_2r0d[15] = rdfint_2n[15];
  assign rd_2r0d[16] = rdfint_2n[16];
  assign rd_2r0d[17] = rdfint_2n[17];
  assign rd_2r0d[18] = rdfint_2n[18];
  assign rd_2r0d[19] = rdfint_2n[19];
  assign rd_2r0d[20] = rdfint_2n[20];
  assign rd_2r0d[21] = rdfint_2n[21];
  assign rd_2r0d[22] = rdfint_2n[22];
  assign rd_2r0d[23] = rdfint_2n[23];
  assign rd_2r0d[24] = rdfint_2n[24];
  assign rd_2r0d[25] = rdfint_2n[25];
  assign rd_2r0d[26] = rdfint_2n[26];
  assign rd_2r0d[27] = rdfint_2n[27];
  assign rd_2r0d[28] = rdfint_2n[28];
  assign rd_2r0d[29] = rdfint_2n[29];
  assign rd_2r0d[30] = rdfint_2n[30];
  assign rd_2r0d[31] = rdfint_2n[31];
  assign rd_2r1d[0] = rdtint_2n[0];
  assign rd_2r1d[1] = rdtint_2n[1];
  assign rd_2r1d[2] = rdtint_2n[2];
  assign rd_2r1d[3] = rdtint_2n[3];
  assign rd_2r1d[4] = rdtint_2n[4];
  assign rd_2r1d[5] = rdtint_2n[5];
  assign rd_2r1d[6] = rdtint_2n[6];
  assign rd_2r1d[7] = rdtint_2n[7];
  assign rd_2r1d[8] = rdtint_2n[8];
  assign rd_2r1d[9] = rdtint_2n[9];
  assign rd_2r1d[10] = rdtint_2n[10];
  assign rd_2r1d[11] = rdtint_2n[11];
  assign rd_2r1d[12] = rdtint_2n[12];
  assign rd_2r1d[13] = rdtint_2n[13];
  assign rd_2r1d[14] = rdtint_2n[14];
  assign rd_2r1d[15] = rdtint_2n[15];
  assign rd_2r1d[16] = rdtint_2n[16];
  assign rd_2r1d[17] = rdtint_2n[17];
  assign rd_2r1d[18] = rdtint_2n[18];
  assign rd_2r1d[19] = rdtint_2n[19];
  assign rd_2r1d[20] = rdtint_2n[20];
  assign rd_2r1d[21] = rdtint_2n[21];
  assign rd_2r1d[22] = rdtint_2n[22];
  assign rd_2r1d[23] = rdtint_2n[23];
  assign rd_2r1d[24] = rdtint_2n[24];
  assign rd_2r1d[25] = rdtint_2n[25];
  assign rd_2r1d[26] = rdtint_2n[26];
  assign rd_2r1d[27] = rdtint_2n[27];
  assign rd_2r1d[28] = rdtint_2n[28];
  assign rd_2r1d[29] = rdtint_2n[29];
  assign rd_2r1d[30] = rdtint_2n[30];
  assign rd_2r1d[31] = rdtint_2n[31];
  assign rgaint_1n = rd_1a;
  assign rd_1r0d = rdfint_1n;
  assign rd_1r1d = rdtint_1n;
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r0d[10] = rdfint_0n[10];
  assign rd_0r0d[11] = rdfint_0n[11];
  assign rd_0r0d[12] = rdfint_0n[12];
  assign rd_0r0d[13] = rdfint_0n[13];
  assign rd_0r0d[14] = rdfint_0n[14];
  assign rd_0r0d[15] = rdfint_0n[15];
  assign rd_0r0d[16] = rdfint_0n[16];
  assign rd_0r0d[17] = rdfint_0n[17];
  assign rd_0r0d[18] = rdfint_0n[18];
  assign rd_0r0d[19] = rdfint_0n[19];
  assign rd_0r0d[20] = rdfint_0n[20];
  assign rd_0r0d[21] = rdfint_0n[21];
  assign rd_0r0d[22] = rdfint_0n[22];
  assign rd_0r0d[23] = rdfint_0n[23];
  assign rd_0r0d[24] = rdfint_0n[24];
  assign rd_0r0d[25] = rdfint_0n[25];
  assign rd_0r0d[26] = rdfint_0n[26];
  assign rd_0r0d[27] = rdfint_0n[27];
  assign rd_0r0d[28] = rdfint_0n[28];
  assign rd_0r0d[29] = rdfint_0n[29];
  assign rd_0r0d[30] = rdfint_0n[30];
  assign rd_0r0d[31] = rdfint_0n[31];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign rd_0r1d[10] = rdtint_0n[10];
  assign rd_0r1d[11] = rdtint_0n[11];
  assign rd_0r1d[12] = rdtint_0n[12];
  assign rd_0r1d[13] = rdtint_0n[13];
  assign rd_0r1d[14] = rdtint_0n[14];
  assign rd_0r1d[15] = rdtint_0n[15];
  assign rd_0r1d[16] = rdtint_0n[16];
  assign rd_0r1d[17] = rdtint_0n[17];
  assign rd_0r1d[18] = rdtint_0n[18];
  assign rd_0r1d[19] = rdtint_0n[19];
  assign rd_0r1d[20] = rdtint_0n[20];
  assign rd_0r1d[21] = rdtint_0n[21];
  assign rd_0r1d[22] = rdtint_0n[22];
  assign rd_0r1d[23] = rdtint_0n[23];
  assign rd_0r1d[24] = rdtint_0n[24];
  assign rd_0r1d[25] = rdtint_0n[25];
  assign rd_0r1d[26] = rdtint_0n[26];
  assign rd_0r1d[27] = rdtint_0n[27];
  assign rd_0r1d[28] = rdtint_0n[28];
  assign rd_0r1d[29] = rdtint_0n[29];
  assign rd_0r1d[30] = rdtint_0n[30];
  assign rd_0r1d[31] = rdtint_0n[31];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign rg_2a = rgaint_2n;
  assign rgrint_2n = rg_2r;
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR3 I206 (internal_0n[0], rgrint_0n, rgrint_1n, rgrint_2n);
  NOR3 I207 (internal_0n[1], rgaint_0n, rgaint_1n, rgaint_2n);
  AND2 I208 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I209 (rdtint_2n[0], rgrint_2n, dt_0n[0]);
  AND2 I210 (rdtint_2n[1], rgrint_2n, dt_0n[1]);
  AND2 I211 (rdtint_2n[2], rgrint_2n, dt_0n[2]);
  AND2 I212 (rdtint_2n[3], rgrint_2n, dt_0n[3]);
  AND2 I213 (rdtint_2n[4], rgrint_2n, dt_0n[4]);
  AND2 I214 (rdtint_2n[5], rgrint_2n, dt_0n[5]);
  AND2 I215 (rdtint_2n[6], rgrint_2n, dt_0n[6]);
  AND2 I216 (rdtint_2n[7], rgrint_2n, dt_0n[7]);
  AND2 I217 (rdtint_2n[8], rgrint_2n, dt_0n[8]);
  AND2 I218 (rdtint_2n[9], rgrint_2n, dt_0n[9]);
  AND2 I219 (rdtint_2n[10], rgrint_2n, dt_0n[10]);
  AND2 I220 (rdtint_2n[11], rgrint_2n, dt_0n[11]);
  AND2 I221 (rdtint_2n[12], rgrint_2n, dt_0n[12]);
  AND2 I222 (rdtint_2n[13], rgrint_2n, dt_0n[13]);
  AND2 I223 (rdtint_2n[14], rgrint_2n, dt_0n[14]);
  AND2 I224 (rdtint_2n[15], rgrint_2n, dt_0n[15]);
  AND2 I225 (rdtint_2n[16], rgrint_2n, dt_0n[16]);
  AND2 I226 (rdtint_2n[17], rgrint_2n, dt_0n[17]);
  AND2 I227 (rdtint_2n[18], rgrint_2n, dt_0n[18]);
  AND2 I228 (rdtint_2n[19], rgrint_2n, dt_0n[19]);
  AND2 I229 (rdtint_2n[20], rgrint_2n, dt_0n[20]);
  AND2 I230 (rdtint_2n[21], rgrint_2n, dt_0n[21]);
  AND2 I231 (rdtint_2n[22], rgrint_2n, dt_0n[22]);
  AND2 I232 (rdtint_2n[23], rgrint_2n, dt_0n[23]);
  AND2 I233 (rdtint_2n[24], rgrint_2n, dt_0n[24]);
  AND2 I234 (rdtint_2n[25], rgrint_2n, dt_0n[25]);
  AND2 I235 (rdtint_2n[26], rgrint_2n, dt_0n[26]);
  AND2 I236 (rdtint_2n[27], rgrint_2n, dt_0n[27]);
  AND2 I237 (rdtint_2n[28], rgrint_2n, dt_0n[28]);
  AND2 I238 (rdtint_2n[29], rgrint_2n, dt_0n[29]);
  AND2 I239 (rdtint_2n[30], rgrint_2n, dt_0n[30]);
  AND2 I240 (rdtint_2n[31], rgrint_2n, dt_0n[31]);
  AND2 I241 (rdtint_1n, rgrint_1n, dt_0n[31]);
  AND2 I242 (rdtint_0n[0], rgrint_0n, dt_0n[0]);
  AND2 I243 (rdtint_0n[1], rgrint_0n, dt_0n[1]);
  AND2 I244 (rdtint_0n[2], rgrint_0n, dt_0n[2]);
  AND2 I245 (rdtint_0n[3], rgrint_0n, dt_0n[3]);
  AND2 I246 (rdtint_0n[4], rgrint_0n, dt_0n[4]);
  AND2 I247 (rdtint_0n[5], rgrint_0n, dt_0n[5]);
  AND2 I248 (rdtint_0n[6], rgrint_0n, dt_0n[6]);
  AND2 I249 (rdtint_0n[7], rgrint_0n, dt_0n[7]);
  AND2 I250 (rdtint_0n[8], rgrint_0n, dt_0n[8]);
  AND2 I251 (rdtint_0n[9], rgrint_0n, dt_0n[9]);
  AND2 I252 (rdtint_0n[10], rgrint_0n, dt_0n[10]);
  AND2 I253 (rdtint_0n[11], rgrint_0n, dt_0n[11]);
  AND2 I254 (rdtint_0n[12], rgrint_0n, dt_0n[12]);
  AND2 I255 (rdtint_0n[13], rgrint_0n, dt_0n[13]);
  AND2 I256 (rdtint_0n[14], rgrint_0n, dt_0n[14]);
  AND2 I257 (rdtint_0n[15], rgrint_0n, dt_0n[15]);
  AND2 I258 (rdtint_0n[16], rgrint_0n, dt_0n[16]);
  AND2 I259 (rdtint_0n[17], rgrint_0n, dt_0n[17]);
  AND2 I260 (rdtint_0n[18], rgrint_0n, dt_0n[18]);
  AND2 I261 (rdtint_0n[19], rgrint_0n, dt_0n[19]);
  AND2 I262 (rdtint_0n[20], rgrint_0n, dt_0n[20]);
  AND2 I263 (rdtint_0n[21], rgrint_0n, dt_0n[21]);
  AND2 I264 (rdtint_0n[22], rgrint_0n, dt_0n[22]);
  AND2 I265 (rdtint_0n[23], rgrint_0n, dt_0n[23]);
  AND2 I266 (rdtint_0n[24], rgrint_0n, dt_0n[24]);
  AND2 I267 (rdtint_0n[25], rgrint_0n, dt_0n[25]);
  AND2 I268 (rdtint_0n[26], rgrint_0n, dt_0n[26]);
  AND2 I269 (rdtint_0n[27], rgrint_0n, dt_0n[27]);
  AND2 I270 (rdtint_0n[28], rgrint_0n, dt_0n[28]);
  AND2 I271 (rdtint_0n[29], rgrint_0n, dt_0n[29]);
  AND2 I272 (rdtint_0n[30], rgrint_0n, dt_0n[30]);
  AND2 I273 (rdtint_0n[31], rgrint_0n, dt_0n[31]);
  AND2 I274 (rdfint_2n[0], rgrint_2n, df_0n[0]);
  AND2 I275 (rdfint_2n[1], rgrint_2n, df_0n[1]);
  AND2 I276 (rdfint_2n[2], rgrint_2n, df_0n[2]);
  AND2 I277 (rdfint_2n[3], rgrint_2n, df_0n[3]);
  AND2 I278 (rdfint_2n[4], rgrint_2n, df_0n[4]);
  AND2 I279 (rdfint_2n[5], rgrint_2n, df_0n[5]);
  AND2 I280 (rdfint_2n[6], rgrint_2n, df_0n[6]);
  AND2 I281 (rdfint_2n[7], rgrint_2n, df_0n[7]);
  AND2 I282 (rdfint_2n[8], rgrint_2n, df_0n[8]);
  AND2 I283 (rdfint_2n[9], rgrint_2n, df_0n[9]);
  AND2 I284 (rdfint_2n[10], rgrint_2n, df_0n[10]);
  AND2 I285 (rdfint_2n[11], rgrint_2n, df_0n[11]);
  AND2 I286 (rdfint_2n[12], rgrint_2n, df_0n[12]);
  AND2 I287 (rdfint_2n[13], rgrint_2n, df_0n[13]);
  AND2 I288 (rdfint_2n[14], rgrint_2n, df_0n[14]);
  AND2 I289 (rdfint_2n[15], rgrint_2n, df_0n[15]);
  AND2 I290 (rdfint_2n[16], rgrint_2n, df_0n[16]);
  AND2 I291 (rdfint_2n[17], rgrint_2n, df_0n[17]);
  AND2 I292 (rdfint_2n[18], rgrint_2n, df_0n[18]);
  AND2 I293 (rdfint_2n[19], rgrint_2n, df_0n[19]);
  AND2 I294 (rdfint_2n[20], rgrint_2n, df_0n[20]);
  AND2 I295 (rdfint_2n[21], rgrint_2n, df_0n[21]);
  AND2 I296 (rdfint_2n[22], rgrint_2n, df_0n[22]);
  AND2 I297 (rdfint_2n[23], rgrint_2n, df_0n[23]);
  AND2 I298 (rdfint_2n[24], rgrint_2n, df_0n[24]);
  AND2 I299 (rdfint_2n[25], rgrint_2n, df_0n[25]);
  AND2 I300 (rdfint_2n[26], rgrint_2n, df_0n[26]);
  AND2 I301 (rdfint_2n[27], rgrint_2n, df_0n[27]);
  AND2 I302 (rdfint_2n[28], rgrint_2n, df_0n[28]);
  AND2 I303 (rdfint_2n[29], rgrint_2n, df_0n[29]);
  AND2 I304 (rdfint_2n[30], rgrint_2n, df_0n[30]);
  AND2 I305 (rdfint_2n[31], rgrint_2n, df_0n[31]);
  AND2 I306 (rdfint_1n, rgrint_1n, df_0n[31]);
  AND2 I307 (rdfint_0n[0], rgrint_0n, df_0n[0]);
  AND2 I308 (rdfint_0n[1], rgrint_0n, df_0n[1]);
  AND2 I309 (rdfint_0n[2], rgrint_0n, df_0n[2]);
  AND2 I310 (rdfint_0n[3], rgrint_0n, df_0n[3]);
  AND2 I311 (rdfint_0n[4], rgrint_0n, df_0n[4]);
  AND2 I312 (rdfint_0n[5], rgrint_0n, df_0n[5]);
  AND2 I313 (rdfint_0n[6], rgrint_0n, df_0n[6]);
  AND2 I314 (rdfint_0n[7], rgrint_0n, df_0n[7]);
  AND2 I315 (rdfint_0n[8], rgrint_0n, df_0n[8]);
  AND2 I316 (rdfint_0n[9], rgrint_0n, df_0n[9]);
  AND2 I317 (rdfint_0n[10], rgrint_0n, df_0n[10]);
  AND2 I318 (rdfint_0n[11], rgrint_0n, df_0n[11]);
  AND2 I319 (rdfint_0n[12], rgrint_0n, df_0n[12]);
  AND2 I320 (rdfint_0n[13], rgrint_0n, df_0n[13]);
  AND2 I321 (rdfint_0n[14], rgrint_0n, df_0n[14]);
  AND2 I322 (rdfint_0n[15], rgrint_0n, df_0n[15]);
  AND2 I323 (rdfint_0n[16], rgrint_0n, df_0n[16]);
  AND2 I324 (rdfint_0n[17], rgrint_0n, df_0n[17]);
  AND2 I325 (rdfint_0n[18], rgrint_0n, df_0n[18]);
  AND2 I326 (rdfint_0n[19], rgrint_0n, df_0n[19]);
  AND2 I327 (rdfint_0n[20], rgrint_0n, df_0n[20]);
  AND2 I328 (rdfint_0n[21], rgrint_0n, df_0n[21]);
  AND2 I329 (rdfint_0n[22], rgrint_0n, df_0n[22]);
  AND2 I330 (rdfint_0n[23], rgrint_0n, df_0n[23]);
  AND2 I331 (rdfint_0n[24], rgrint_0n, df_0n[24]);
  AND2 I332 (rdfint_0n[25], rgrint_0n, df_0n[25]);
  AND2 I333 (rdfint_0n[26], rgrint_0n, df_0n[26]);
  AND2 I334 (rdfint_0n[27], rgrint_0n, df_0n[27]);
  AND2 I335 (rdfint_0n[28], rgrint_0n, df_0n[28]);
  AND2 I336 (rdfint_0n[29], rgrint_0n, df_0n[29]);
  AND2 I337 (rdfint_0n[30], rgrint_0n, df_0n[30]);
  AND2 I338 (rdfint_0n[31], rgrint_0n, df_0n[31]);
  C3 I339 (internal_0n[2], wc_0n, wacks_0n[31], wacks_0n[30]);
  C3 I340 (internal_0n[3], wacks_0n[29], wacks_0n[28], wacks_0n[27]);
  C3 I341 (internal_0n[4], wacks_0n[26], wacks_0n[25], wacks_0n[24]);
  C3 I342 (internal_0n[5], wacks_0n[23], wacks_0n[22], wacks_0n[21]);
  C3 I343 (internal_0n[6], wacks_0n[20], wacks_0n[19], wacks_0n[18]);
  C3 I344 (internal_0n[7], wacks_0n[17], wacks_0n[16], wacks_0n[15]);
  C3 I345 (internal_0n[8], wacks_0n[14], wacks_0n[13], wacks_0n[12]);
  C3 I346 (internal_0n[9], wacks_0n[11], wacks_0n[10], wacks_0n[9]);
  C3 I347 (internal_0n[10], wacks_0n[8], wacks_0n[7], wacks_0n[6]);
  C3 I348 (internal_0n[11], wacks_0n[5], wacks_0n[4], wacks_0n[3]);
  C3 I349 (internal_0n[12], wacks_0n[2], wacks_0n[1], wacks_0n[0]);
  C3 I350 (internal_0n[13], internal_0n[2], internal_0n[3], internal_0n[4]);
  C3 I351 (internal_0n[14], internal_0n[5], internal_0n[6], internal_0n[7]);
  C3 I352 (internal_0n[15], internal_0n[8], internal_0n[9], internal_0n[10]);
  C2 I353 (internal_0n[16], internal_0n[11], internal_0n[12]);
  C2 I354 (internal_0n[17], internal_0n[13], internal_0n[14]);
  C2 I355 (internal_0n[18], internal_0n[15], internal_0n[16]);
  C2 I356 (wdrint_0n, internal_0n[17], internal_0n[18]);
  assign wen_0n[31] = wc_0n;
  assign wen_0n[30] = wc_0n;
  assign wen_0n[29] = wc_0n;
  assign wen_0n[28] = wc_0n;
  assign wen_0n[27] = wc_0n;
  assign wen_0n[26] = wc_0n;
  assign wen_0n[25] = wc_0n;
  assign wen_0n[24] = wc_0n;
  assign wen_0n[23] = wc_0n;
  assign wen_0n[22] = wc_0n;
  assign wen_0n[21] = wc_0n;
  assign wen_0n[20] = wc_0n;
  assign wen_0n[19] = wc_0n;
  assign wen_0n[18] = wc_0n;
  assign wen_0n[17] = wc_0n;
  assign wen_0n[16] = wc_0n;
  assign wen_0n[15] = wc_0n;
  assign wen_0n[14] = wc_0n;
  assign wen_0n[13] = wc_0n;
  assign wen_0n[12] = wc_0n;
  assign wen_0n[11] = wc_0n;
  assign wen_0n[10] = wc_0n;
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[31] = git_0n[31];
  assign wt_0n[30] = git_0n[30];
  assign wt_0n[29] = git_0n[29];
  assign wt_0n[28] = git_0n[28];
  assign wt_0n[27] = git_0n[27];
  assign wt_0n[26] = git_0n[26];
  assign wt_0n[25] = git_0n[25];
  assign wt_0n[24] = git_0n[24];
  assign wt_0n[23] = git_0n[23];
  assign wt_0n[22] = git_0n[22];
  assign wt_0n[21] = git_0n[21];
  assign wt_0n[20] = git_0n[20];
  assign wt_0n[19] = git_0n[19];
  assign wt_0n[18] = git_0n[18];
  assign wt_0n[17] = git_0n[17];
  assign wt_0n[16] = git_0n[16];
  assign wt_0n[15] = git_0n[15];
  assign wt_0n[14] = git_0n[14];
  assign wt_0n[13] = git_0n[13];
  assign wt_0n[12] = git_0n[12];
  assign wt_0n[11] = git_0n[11];
  assign wt_0n[10] = git_0n[10];
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[31] = gif_0n[31];
  assign wf_0n[30] = gif_0n[30];
  assign wf_0n[29] = gif_0n[29];
  assign wf_0n[28] = gif_0n[28];
  assign wf_0n[27] = gif_0n[27];
  assign wf_0n[26] = gif_0n[26];
  assign wf_0n[25] = gif_0n[25];
  assign wf_0n[24] = gif_0n[24];
  assign wf_0n[23] = gif_0n[23];
  assign wf_0n[22] = gif_0n[22];
  assign wf_0n[21] = gif_0n[21];
  assign wf_0n[20] = gif_0n[20];
  assign wf_0n[19] = gif_0n[19];
  assign wf_0n[18] = gif_0n[18];
  assign wf_0n[17] = gif_0n[17];
  assign wf_0n[16] = gif_0n[16];
  assign wf_0n[15] = gif_0n[15];
  assign wf_0n[14] = gif_0n[14];
  assign wf_0n[13] = gif_0n[13];
  assign wf_0n[12] = gif_0n[12];
  assign wf_0n[11] = gif_0n[11];
  assign wf_0n[10] = gif_0n[10];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I453 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I455 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I456 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I457 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I458 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I459 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I460 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I461 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I462 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I463 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I464 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I465 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I466 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I467 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I468 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I469 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I470 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I471 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I472 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I473 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I474 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I475 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I476 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I477 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I478 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I479 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I480 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I481 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I482 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I483 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I484 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I485 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I486 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I487 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I488 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I489 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I490 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I491 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I492 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I493 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I494 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I495 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I496 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I497 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I498 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I499 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I500 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I501 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I502 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I503 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I504 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I505 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I506 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I507 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I508 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I509 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I510 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I511 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I512 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I513 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I514 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I515 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I516 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I517 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I518 (gif_0n[31], wgfint_0n[31], ig_0n);
  C3 I519 (internal_0n[19], complete1346_0n[0], complete1346_0n[1], complete1346_0n[2]);
  C3 I520 (internal_0n[20], complete1346_0n[3], complete1346_0n[4], complete1346_0n[5]);
  C3 I521 (internal_0n[21], complete1346_0n[6], complete1346_0n[7], complete1346_0n[8]);
  C3 I522 (internal_0n[22], complete1346_0n[9], complete1346_0n[10], complete1346_0n[11]);
  C3 I523 (internal_0n[23], complete1346_0n[12], complete1346_0n[13], complete1346_0n[14]);
  C3 I524 (internal_0n[24], complete1346_0n[15], complete1346_0n[16], complete1346_0n[17]);
  C3 I525 (internal_0n[25], complete1346_0n[18], complete1346_0n[19], complete1346_0n[20]);
  C3 I526 (internal_0n[26], complete1346_0n[21], complete1346_0n[22], complete1346_0n[23]);
  C3 I527 (internal_0n[27], complete1346_0n[24], complete1346_0n[25], complete1346_0n[26]);
  C3 I528 (internal_0n[28], complete1346_0n[27], complete1346_0n[28], complete1346_0n[29]);
  C2 I529 (internal_0n[29], complete1346_0n[30], complete1346_0n[31]);
  C3 I530 (internal_0n[30], internal_0n[19], internal_0n[20], internal_0n[21]);
  C3 I531 (internal_0n[31], internal_0n[22], internal_0n[23], internal_0n[24]);
  C3 I532 (internal_0n[32], internal_0n[25], internal_0n[26], internal_0n[27]);
  C2 I533 (internal_0n[33], internal_0n[28], internal_0n[29]);
  C2 I534 (internal_0n[34], internal_0n[30], internal_0n[31]);
  C2 I535 (internal_0n[35], internal_0n[32], internal_0n[33]);
  C2 I536 (wc_0n, internal_0n[34], internal_0n[35]);
  OR2 I537 (complete1346_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I538 (complete1346_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I539 (complete1346_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I540 (complete1346_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I541 (complete1346_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I542 (complete1346_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I543 (complete1346_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I544 (complete1346_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I545 (complete1346_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I546 (complete1346_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I547 (complete1346_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I548 (complete1346_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I549 (complete1346_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I550 (complete1346_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I551 (complete1346_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I552 (complete1346_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I553 (complete1346_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I554 (complete1346_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I555 (complete1346_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I556 (complete1346_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I557 (complete1346_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I558 (complete1346_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I559 (complete1346_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I560 (complete1346_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I561 (complete1346_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I562 (complete1346_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I563 (complete1346_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I564 (complete1346_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I565 (complete1346_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I566 (complete1346_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I567 (complete1346_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I568 (complete1346_0n[31], wgfint_0n[31], wgtint_0n[31]);
  AO22 I569 (wacks_0n[31], gf1344_0n[31], df_0n[31], gt1345_0n[31], dt_0n[31]);
  NOR2 I570 (dt_0n[31], df_0n[31], gf1344_0n[31]);
  NOR3 I571 (df_0n[31], dt_0n[31], gt1345_0n[31], init_0n);
  AND2 I572 (gt1345_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I573 (gf1344_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I574 (wacks_0n[30], gf1344_0n[30], df_0n[30], gt1345_0n[30], dt_0n[30]);
  NOR2 I575 (dt_0n[30], df_0n[30], gf1344_0n[30]);
  NOR3 I576 (df_0n[30], dt_0n[30], gt1345_0n[30], init_0n);
  AND2 I577 (gt1345_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I578 (gf1344_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I579 (wacks_0n[29], gf1344_0n[29], df_0n[29], gt1345_0n[29], dt_0n[29]);
  NOR2 I580 (dt_0n[29], df_0n[29], gf1344_0n[29]);
  NOR3 I581 (df_0n[29], dt_0n[29], gt1345_0n[29], init_0n);
  AND2 I582 (gt1345_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I583 (gf1344_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I584 (wacks_0n[28], gf1344_0n[28], df_0n[28], gt1345_0n[28], dt_0n[28]);
  NOR2 I585 (dt_0n[28], df_0n[28], gf1344_0n[28]);
  NOR3 I586 (df_0n[28], dt_0n[28], gt1345_0n[28], init_0n);
  AND2 I587 (gt1345_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I588 (gf1344_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I589 (wacks_0n[27], gf1344_0n[27], df_0n[27], gt1345_0n[27], dt_0n[27]);
  NOR2 I590 (dt_0n[27], df_0n[27], gf1344_0n[27]);
  NOR3 I591 (df_0n[27], dt_0n[27], gt1345_0n[27], init_0n);
  AND2 I592 (gt1345_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I593 (gf1344_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I594 (wacks_0n[26], gf1344_0n[26], df_0n[26], gt1345_0n[26], dt_0n[26]);
  NOR2 I595 (dt_0n[26], df_0n[26], gf1344_0n[26]);
  NOR3 I596 (df_0n[26], dt_0n[26], gt1345_0n[26], init_0n);
  AND2 I597 (gt1345_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I598 (gf1344_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I599 (wacks_0n[25], gf1344_0n[25], df_0n[25], gt1345_0n[25], dt_0n[25]);
  NOR2 I600 (dt_0n[25], df_0n[25], gf1344_0n[25]);
  NOR3 I601 (df_0n[25], dt_0n[25], gt1345_0n[25], init_0n);
  AND2 I602 (gt1345_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I603 (gf1344_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I604 (wacks_0n[24], gf1344_0n[24], df_0n[24], gt1345_0n[24], dt_0n[24]);
  NOR2 I605 (dt_0n[24], df_0n[24], gf1344_0n[24]);
  NOR3 I606 (df_0n[24], dt_0n[24], gt1345_0n[24], init_0n);
  AND2 I607 (gt1345_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I608 (gf1344_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I609 (wacks_0n[23], gf1344_0n[23], df_0n[23], gt1345_0n[23], dt_0n[23]);
  NOR2 I610 (dt_0n[23], df_0n[23], gf1344_0n[23]);
  NOR3 I611 (df_0n[23], dt_0n[23], gt1345_0n[23], init_0n);
  AND2 I612 (gt1345_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I613 (gf1344_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I614 (wacks_0n[22], gf1344_0n[22], df_0n[22], gt1345_0n[22], dt_0n[22]);
  NOR2 I615 (dt_0n[22], df_0n[22], gf1344_0n[22]);
  NOR3 I616 (df_0n[22], dt_0n[22], gt1345_0n[22], init_0n);
  AND2 I617 (gt1345_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I618 (gf1344_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I619 (wacks_0n[21], gf1344_0n[21], df_0n[21], gt1345_0n[21], dt_0n[21]);
  NOR2 I620 (dt_0n[21], df_0n[21], gf1344_0n[21]);
  NOR3 I621 (df_0n[21], dt_0n[21], gt1345_0n[21], init_0n);
  AND2 I622 (gt1345_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I623 (gf1344_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I624 (wacks_0n[20], gf1344_0n[20], df_0n[20], gt1345_0n[20], dt_0n[20]);
  NOR2 I625 (dt_0n[20], df_0n[20], gf1344_0n[20]);
  NOR3 I626 (df_0n[20], dt_0n[20], gt1345_0n[20], init_0n);
  AND2 I627 (gt1345_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I628 (gf1344_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I629 (wacks_0n[19], gf1344_0n[19], df_0n[19], gt1345_0n[19], dt_0n[19]);
  NOR2 I630 (dt_0n[19], df_0n[19], gf1344_0n[19]);
  NOR3 I631 (df_0n[19], dt_0n[19], gt1345_0n[19], init_0n);
  AND2 I632 (gt1345_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I633 (gf1344_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I634 (wacks_0n[18], gf1344_0n[18], df_0n[18], gt1345_0n[18], dt_0n[18]);
  NOR2 I635 (dt_0n[18], df_0n[18], gf1344_0n[18]);
  NOR3 I636 (df_0n[18], dt_0n[18], gt1345_0n[18], init_0n);
  AND2 I637 (gt1345_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I638 (gf1344_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I639 (wacks_0n[17], gf1344_0n[17], df_0n[17], gt1345_0n[17], dt_0n[17]);
  NOR2 I640 (dt_0n[17], df_0n[17], gf1344_0n[17]);
  NOR3 I641 (df_0n[17], dt_0n[17], gt1345_0n[17], init_0n);
  AND2 I642 (gt1345_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I643 (gf1344_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I644 (wacks_0n[16], gf1344_0n[16], df_0n[16], gt1345_0n[16], dt_0n[16]);
  NOR2 I645 (dt_0n[16], df_0n[16], gf1344_0n[16]);
  NOR3 I646 (df_0n[16], dt_0n[16], gt1345_0n[16], init_0n);
  AND2 I647 (gt1345_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I648 (gf1344_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I649 (wacks_0n[15], gf1344_0n[15], df_0n[15], gt1345_0n[15], dt_0n[15]);
  NOR2 I650 (dt_0n[15], df_0n[15], gf1344_0n[15]);
  NOR3 I651 (df_0n[15], dt_0n[15], gt1345_0n[15], init_0n);
  AND2 I652 (gt1345_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I653 (gf1344_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I654 (wacks_0n[14], gf1344_0n[14], df_0n[14], gt1345_0n[14], dt_0n[14]);
  NOR2 I655 (dt_0n[14], df_0n[14], gf1344_0n[14]);
  NOR3 I656 (df_0n[14], dt_0n[14], gt1345_0n[14], init_0n);
  AND2 I657 (gt1345_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I658 (gf1344_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I659 (wacks_0n[13], gf1344_0n[13], df_0n[13], gt1345_0n[13], dt_0n[13]);
  NOR2 I660 (dt_0n[13], df_0n[13], gf1344_0n[13]);
  NOR3 I661 (df_0n[13], dt_0n[13], gt1345_0n[13], init_0n);
  AND2 I662 (gt1345_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I663 (gf1344_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I664 (wacks_0n[12], gf1344_0n[12], df_0n[12], gt1345_0n[12], dt_0n[12]);
  NOR2 I665 (dt_0n[12], df_0n[12], gf1344_0n[12]);
  NOR3 I666 (df_0n[12], dt_0n[12], gt1345_0n[12], init_0n);
  AND2 I667 (gt1345_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I668 (gf1344_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I669 (wacks_0n[11], gf1344_0n[11], df_0n[11], gt1345_0n[11], dt_0n[11]);
  NOR2 I670 (dt_0n[11], df_0n[11], gf1344_0n[11]);
  NOR3 I671 (df_0n[11], dt_0n[11], gt1345_0n[11], init_0n);
  AND2 I672 (gt1345_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I673 (gf1344_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I674 (wacks_0n[10], gf1344_0n[10], df_0n[10], gt1345_0n[10], dt_0n[10]);
  NOR2 I675 (dt_0n[10], df_0n[10], gf1344_0n[10]);
  NOR3 I676 (df_0n[10], dt_0n[10], gt1345_0n[10], init_0n);
  AND2 I677 (gt1345_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I678 (gf1344_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I679 (wacks_0n[9], gf1344_0n[9], df_0n[9], gt1345_0n[9], dt_0n[9]);
  NOR2 I680 (dt_0n[9], df_0n[9], gf1344_0n[9]);
  NOR3 I681 (df_0n[9], dt_0n[9], gt1345_0n[9], init_0n);
  AND2 I682 (gt1345_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I683 (gf1344_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I684 (wacks_0n[8], gf1344_0n[8], df_0n[8], gt1345_0n[8], dt_0n[8]);
  NOR2 I685 (dt_0n[8], df_0n[8], gf1344_0n[8]);
  NOR3 I686 (df_0n[8], dt_0n[8], gt1345_0n[8], init_0n);
  AND2 I687 (gt1345_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I688 (gf1344_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I689 (wacks_0n[7], gf1344_0n[7], df_0n[7], gt1345_0n[7], dt_0n[7]);
  NOR2 I690 (dt_0n[7], df_0n[7], gf1344_0n[7]);
  NOR3 I691 (df_0n[7], dt_0n[7], gt1345_0n[7], init_0n);
  AND2 I692 (gt1345_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I693 (gf1344_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I694 (wacks_0n[6], gf1344_0n[6], df_0n[6], gt1345_0n[6], dt_0n[6]);
  NOR2 I695 (dt_0n[6], df_0n[6], gf1344_0n[6]);
  NOR3 I696 (df_0n[6], dt_0n[6], gt1345_0n[6], init_0n);
  AND2 I697 (gt1345_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I698 (gf1344_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I699 (wacks_0n[5], gf1344_0n[5], df_0n[5], gt1345_0n[5], dt_0n[5]);
  NOR2 I700 (dt_0n[5], df_0n[5], gf1344_0n[5]);
  NOR3 I701 (df_0n[5], dt_0n[5], gt1345_0n[5], init_0n);
  AND2 I702 (gt1345_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I703 (gf1344_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I704 (wacks_0n[4], gf1344_0n[4], df_0n[4], gt1345_0n[4], dt_0n[4]);
  NOR2 I705 (dt_0n[4], df_0n[4], gf1344_0n[4]);
  NOR3 I706 (df_0n[4], dt_0n[4], gt1345_0n[4], init_0n);
  AND2 I707 (gt1345_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I708 (gf1344_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I709 (wacks_0n[3], gf1344_0n[3], df_0n[3], gt1345_0n[3], dt_0n[3]);
  NOR2 I710 (dt_0n[3], df_0n[3], gf1344_0n[3]);
  NOR3 I711 (df_0n[3], dt_0n[3], gt1345_0n[3], init_0n);
  AND2 I712 (gt1345_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I713 (gf1344_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I714 (wacks_0n[2], gf1344_0n[2], df_0n[2], gt1345_0n[2], dt_0n[2]);
  NOR2 I715 (dt_0n[2], df_0n[2], gf1344_0n[2]);
  NOR3 I716 (df_0n[2], dt_0n[2], gt1345_0n[2], init_0n);
  AND2 I717 (gt1345_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I718 (gf1344_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I719 (wacks_0n[1], gf1344_0n[1], df_0n[1], gt1345_0n[1], dt_0n[1]);
  NOR2 I720 (dt_0n[1], df_0n[1], gf1344_0n[1]);
  NOR3 I721 (df_0n[1], dt_0n[1], gt1345_0n[1], init_0n);
  AND2 I722 (gt1345_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I723 (gf1344_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I724 (wacks_0n[0], gf1344_0n[0], df_0n[0], gt1345_0n[0], dt_0n[0]);
  NOR2 I725 (dt_0n[0], df_0n[0], gf1344_0n[0]);
  NOR3 I726 (df_0n[0], dt_0n[0], gt1345_0n[0], init_0n);
  AND2 I727 (gt1345_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I728 (gf1344_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I729 (init_0n, initialise);
endmodule

module BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m83m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rg_2r, rg_2a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  rd_2r0d, rd_2r1d, rd_2a,
  initialise
);
  input [31:0] wg_0r0d;
  input [31:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output rd_0r0d;
  output rd_0r1d;
  input rd_0a;
  output [31:0] rd_1r0d;
  output [31:0] rd_1r1d;
  input rd_1a;
  output [31:0] rd_2r0d;
  output [31:0] rd_2r1d;
  input rd_2a;
  input initialise;
  wire [35:0] internal_0n;
  wire [31:0] wf_0n;
  wire [31:0] wt_0n;
  wire [31:0] df_0n;
  wire [31:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire rgrint_2n;
  wire wc_0n;
  wire [31:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [31:0] wgfint_0n;
  wire [31:0] wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire rgaint_2n;
  wire rdfint_0n;
  wire [31:0] rdfint_1n;
  wire [31:0] rdfint_2n;
  wire rdtint_0n;
  wire [31:0] rdtint_1n;
  wire [31:0] rdtint_2n;
  wire [31:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [31:0] gif_0n;
  wire [31:0] git_0n;
  wire [31:0] complete1365_0n;
  wire [31:0] gt1364_0n;
  wire [31:0] gf1363_0n;
  assign rgaint_2n = rd_2a;
  assign rd_2r0d[0] = rdfint_2n[0];
  assign rd_2r0d[1] = rdfint_2n[1];
  assign rd_2r0d[2] = rdfint_2n[2];
  assign rd_2r0d[3] = rdfint_2n[3];
  assign rd_2r0d[4] = rdfint_2n[4];
  assign rd_2r0d[5] = rdfint_2n[5];
  assign rd_2r0d[6] = rdfint_2n[6];
  assign rd_2r0d[7] = rdfint_2n[7];
  assign rd_2r0d[8] = rdfint_2n[8];
  assign rd_2r0d[9] = rdfint_2n[9];
  assign rd_2r0d[10] = rdfint_2n[10];
  assign rd_2r0d[11] = rdfint_2n[11];
  assign rd_2r0d[12] = rdfint_2n[12];
  assign rd_2r0d[13] = rdfint_2n[13];
  assign rd_2r0d[14] = rdfint_2n[14];
  assign rd_2r0d[15] = rdfint_2n[15];
  assign rd_2r0d[16] = rdfint_2n[16];
  assign rd_2r0d[17] = rdfint_2n[17];
  assign rd_2r0d[18] = rdfint_2n[18];
  assign rd_2r0d[19] = rdfint_2n[19];
  assign rd_2r0d[20] = rdfint_2n[20];
  assign rd_2r0d[21] = rdfint_2n[21];
  assign rd_2r0d[22] = rdfint_2n[22];
  assign rd_2r0d[23] = rdfint_2n[23];
  assign rd_2r0d[24] = rdfint_2n[24];
  assign rd_2r0d[25] = rdfint_2n[25];
  assign rd_2r0d[26] = rdfint_2n[26];
  assign rd_2r0d[27] = rdfint_2n[27];
  assign rd_2r0d[28] = rdfint_2n[28];
  assign rd_2r0d[29] = rdfint_2n[29];
  assign rd_2r0d[30] = rdfint_2n[30];
  assign rd_2r0d[31] = rdfint_2n[31];
  assign rd_2r1d[0] = rdtint_2n[0];
  assign rd_2r1d[1] = rdtint_2n[1];
  assign rd_2r1d[2] = rdtint_2n[2];
  assign rd_2r1d[3] = rdtint_2n[3];
  assign rd_2r1d[4] = rdtint_2n[4];
  assign rd_2r1d[5] = rdtint_2n[5];
  assign rd_2r1d[6] = rdtint_2n[6];
  assign rd_2r1d[7] = rdtint_2n[7];
  assign rd_2r1d[8] = rdtint_2n[8];
  assign rd_2r1d[9] = rdtint_2n[9];
  assign rd_2r1d[10] = rdtint_2n[10];
  assign rd_2r1d[11] = rdtint_2n[11];
  assign rd_2r1d[12] = rdtint_2n[12];
  assign rd_2r1d[13] = rdtint_2n[13];
  assign rd_2r1d[14] = rdtint_2n[14];
  assign rd_2r1d[15] = rdtint_2n[15];
  assign rd_2r1d[16] = rdtint_2n[16];
  assign rd_2r1d[17] = rdtint_2n[17];
  assign rd_2r1d[18] = rdtint_2n[18];
  assign rd_2r1d[19] = rdtint_2n[19];
  assign rd_2r1d[20] = rdtint_2n[20];
  assign rd_2r1d[21] = rdtint_2n[21];
  assign rd_2r1d[22] = rdtint_2n[22];
  assign rd_2r1d[23] = rdtint_2n[23];
  assign rd_2r1d[24] = rdtint_2n[24];
  assign rd_2r1d[25] = rdtint_2n[25];
  assign rd_2r1d[26] = rdtint_2n[26];
  assign rd_2r1d[27] = rdtint_2n[27];
  assign rd_2r1d[28] = rdtint_2n[28];
  assign rd_2r1d[29] = rdtint_2n[29];
  assign rd_2r1d[30] = rdtint_2n[30];
  assign rd_2r1d[31] = rdtint_2n[31];
  assign rgaint_1n = rd_1a;
  assign rd_1r0d[0] = rdfint_1n[0];
  assign rd_1r0d[1] = rdfint_1n[1];
  assign rd_1r0d[2] = rdfint_1n[2];
  assign rd_1r0d[3] = rdfint_1n[3];
  assign rd_1r0d[4] = rdfint_1n[4];
  assign rd_1r0d[5] = rdfint_1n[5];
  assign rd_1r0d[6] = rdfint_1n[6];
  assign rd_1r0d[7] = rdfint_1n[7];
  assign rd_1r0d[8] = rdfint_1n[8];
  assign rd_1r0d[9] = rdfint_1n[9];
  assign rd_1r0d[10] = rdfint_1n[10];
  assign rd_1r0d[11] = rdfint_1n[11];
  assign rd_1r0d[12] = rdfint_1n[12];
  assign rd_1r0d[13] = rdfint_1n[13];
  assign rd_1r0d[14] = rdfint_1n[14];
  assign rd_1r0d[15] = rdfint_1n[15];
  assign rd_1r0d[16] = rdfint_1n[16];
  assign rd_1r0d[17] = rdfint_1n[17];
  assign rd_1r0d[18] = rdfint_1n[18];
  assign rd_1r0d[19] = rdfint_1n[19];
  assign rd_1r0d[20] = rdfint_1n[20];
  assign rd_1r0d[21] = rdfint_1n[21];
  assign rd_1r0d[22] = rdfint_1n[22];
  assign rd_1r0d[23] = rdfint_1n[23];
  assign rd_1r0d[24] = rdfint_1n[24];
  assign rd_1r0d[25] = rdfint_1n[25];
  assign rd_1r0d[26] = rdfint_1n[26];
  assign rd_1r0d[27] = rdfint_1n[27];
  assign rd_1r0d[28] = rdfint_1n[28];
  assign rd_1r0d[29] = rdfint_1n[29];
  assign rd_1r0d[30] = rdfint_1n[30];
  assign rd_1r0d[31] = rdfint_1n[31];
  assign rd_1r1d[0] = rdtint_1n[0];
  assign rd_1r1d[1] = rdtint_1n[1];
  assign rd_1r1d[2] = rdtint_1n[2];
  assign rd_1r1d[3] = rdtint_1n[3];
  assign rd_1r1d[4] = rdtint_1n[4];
  assign rd_1r1d[5] = rdtint_1n[5];
  assign rd_1r1d[6] = rdtint_1n[6];
  assign rd_1r1d[7] = rdtint_1n[7];
  assign rd_1r1d[8] = rdtint_1n[8];
  assign rd_1r1d[9] = rdtint_1n[9];
  assign rd_1r1d[10] = rdtint_1n[10];
  assign rd_1r1d[11] = rdtint_1n[11];
  assign rd_1r1d[12] = rdtint_1n[12];
  assign rd_1r1d[13] = rdtint_1n[13];
  assign rd_1r1d[14] = rdtint_1n[14];
  assign rd_1r1d[15] = rdtint_1n[15];
  assign rd_1r1d[16] = rdtint_1n[16];
  assign rd_1r1d[17] = rdtint_1n[17];
  assign rd_1r1d[18] = rdtint_1n[18];
  assign rd_1r1d[19] = rdtint_1n[19];
  assign rd_1r1d[20] = rdtint_1n[20];
  assign rd_1r1d[21] = rdtint_1n[21];
  assign rd_1r1d[22] = rdtint_1n[22];
  assign rd_1r1d[23] = rdtint_1n[23];
  assign rd_1r1d[24] = rdtint_1n[24];
  assign rd_1r1d[25] = rdtint_1n[25];
  assign rd_1r1d[26] = rdtint_1n[26];
  assign rd_1r1d[27] = rdtint_1n[27];
  assign rd_1r1d[28] = rdtint_1n[28];
  assign rd_1r1d[29] = rdtint_1n[29];
  assign rd_1r1d[30] = rdtint_1n[30];
  assign rd_1r1d[31] = rdtint_1n[31];
  assign rgaint_0n = rd_0a;
  assign rd_0r0d = rdfint_0n;
  assign rd_0r1d = rdtint_0n;
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign rg_2a = rgaint_2n;
  assign rgrint_2n = rg_2r;
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR3 I206 (internal_0n[0], rgrint_0n, rgrint_1n, rgrint_2n);
  NOR3 I207 (internal_0n[1], rgaint_0n, rgaint_1n, rgaint_2n);
  AND2 I208 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I209 (rdtint_2n[0], rgrint_2n, dt_0n[0]);
  AND2 I210 (rdtint_2n[1], rgrint_2n, dt_0n[1]);
  AND2 I211 (rdtint_2n[2], rgrint_2n, dt_0n[2]);
  AND2 I212 (rdtint_2n[3], rgrint_2n, dt_0n[3]);
  AND2 I213 (rdtint_2n[4], rgrint_2n, dt_0n[4]);
  AND2 I214 (rdtint_2n[5], rgrint_2n, dt_0n[5]);
  AND2 I215 (rdtint_2n[6], rgrint_2n, dt_0n[6]);
  AND2 I216 (rdtint_2n[7], rgrint_2n, dt_0n[7]);
  AND2 I217 (rdtint_2n[8], rgrint_2n, dt_0n[8]);
  AND2 I218 (rdtint_2n[9], rgrint_2n, dt_0n[9]);
  AND2 I219 (rdtint_2n[10], rgrint_2n, dt_0n[10]);
  AND2 I220 (rdtint_2n[11], rgrint_2n, dt_0n[11]);
  AND2 I221 (rdtint_2n[12], rgrint_2n, dt_0n[12]);
  AND2 I222 (rdtint_2n[13], rgrint_2n, dt_0n[13]);
  AND2 I223 (rdtint_2n[14], rgrint_2n, dt_0n[14]);
  AND2 I224 (rdtint_2n[15], rgrint_2n, dt_0n[15]);
  AND2 I225 (rdtint_2n[16], rgrint_2n, dt_0n[16]);
  AND2 I226 (rdtint_2n[17], rgrint_2n, dt_0n[17]);
  AND2 I227 (rdtint_2n[18], rgrint_2n, dt_0n[18]);
  AND2 I228 (rdtint_2n[19], rgrint_2n, dt_0n[19]);
  AND2 I229 (rdtint_2n[20], rgrint_2n, dt_0n[20]);
  AND2 I230 (rdtint_2n[21], rgrint_2n, dt_0n[21]);
  AND2 I231 (rdtint_2n[22], rgrint_2n, dt_0n[22]);
  AND2 I232 (rdtint_2n[23], rgrint_2n, dt_0n[23]);
  AND2 I233 (rdtint_2n[24], rgrint_2n, dt_0n[24]);
  AND2 I234 (rdtint_2n[25], rgrint_2n, dt_0n[25]);
  AND2 I235 (rdtint_2n[26], rgrint_2n, dt_0n[26]);
  AND2 I236 (rdtint_2n[27], rgrint_2n, dt_0n[27]);
  AND2 I237 (rdtint_2n[28], rgrint_2n, dt_0n[28]);
  AND2 I238 (rdtint_2n[29], rgrint_2n, dt_0n[29]);
  AND2 I239 (rdtint_2n[30], rgrint_2n, dt_0n[30]);
  AND2 I240 (rdtint_2n[31], rgrint_2n, dt_0n[31]);
  AND2 I241 (rdtint_1n[0], rgrint_1n, dt_0n[0]);
  AND2 I242 (rdtint_1n[1], rgrint_1n, dt_0n[1]);
  AND2 I243 (rdtint_1n[2], rgrint_1n, dt_0n[2]);
  AND2 I244 (rdtint_1n[3], rgrint_1n, dt_0n[3]);
  AND2 I245 (rdtint_1n[4], rgrint_1n, dt_0n[4]);
  AND2 I246 (rdtint_1n[5], rgrint_1n, dt_0n[5]);
  AND2 I247 (rdtint_1n[6], rgrint_1n, dt_0n[6]);
  AND2 I248 (rdtint_1n[7], rgrint_1n, dt_0n[7]);
  AND2 I249 (rdtint_1n[8], rgrint_1n, dt_0n[8]);
  AND2 I250 (rdtint_1n[9], rgrint_1n, dt_0n[9]);
  AND2 I251 (rdtint_1n[10], rgrint_1n, dt_0n[10]);
  AND2 I252 (rdtint_1n[11], rgrint_1n, dt_0n[11]);
  AND2 I253 (rdtint_1n[12], rgrint_1n, dt_0n[12]);
  AND2 I254 (rdtint_1n[13], rgrint_1n, dt_0n[13]);
  AND2 I255 (rdtint_1n[14], rgrint_1n, dt_0n[14]);
  AND2 I256 (rdtint_1n[15], rgrint_1n, dt_0n[15]);
  AND2 I257 (rdtint_1n[16], rgrint_1n, dt_0n[16]);
  AND2 I258 (rdtint_1n[17], rgrint_1n, dt_0n[17]);
  AND2 I259 (rdtint_1n[18], rgrint_1n, dt_0n[18]);
  AND2 I260 (rdtint_1n[19], rgrint_1n, dt_0n[19]);
  AND2 I261 (rdtint_1n[20], rgrint_1n, dt_0n[20]);
  AND2 I262 (rdtint_1n[21], rgrint_1n, dt_0n[21]);
  AND2 I263 (rdtint_1n[22], rgrint_1n, dt_0n[22]);
  AND2 I264 (rdtint_1n[23], rgrint_1n, dt_0n[23]);
  AND2 I265 (rdtint_1n[24], rgrint_1n, dt_0n[24]);
  AND2 I266 (rdtint_1n[25], rgrint_1n, dt_0n[25]);
  AND2 I267 (rdtint_1n[26], rgrint_1n, dt_0n[26]);
  AND2 I268 (rdtint_1n[27], rgrint_1n, dt_0n[27]);
  AND2 I269 (rdtint_1n[28], rgrint_1n, dt_0n[28]);
  AND2 I270 (rdtint_1n[29], rgrint_1n, dt_0n[29]);
  AND2 I271 (rdtint_1n[30], rgrint_1n, dt_0n[30]);
  AND2 I272 (rdtint_1n[31], rgrint_1n, dt_0n[31]);
  AND2 I273 (rdtint_0n, rgrint_0n, dt_0n[31]);
  AND2 I274 (rdfint_2n[0], rgrint_2n, df_0n[0]);
  AND2 I275 (rdfint_2n[1], rgrint_2n, df_0n[1]);
  AND2 I276 (rdfint_2n[2], rgrint_2n, df_0n[2]);
  AND2 I277 (rdfint_2n[3], rgrint_2n, df_0n[3]);
  AND2 I278 (rdfint_2n[4], rgrint_2n, df_0n[4]);
  AND2 I279 (rdfint_2n[5], rgrint_2n, df_0n[5]);
  AND2 I280 (rdfint_2n[6], rgrint_2n, df_0n[6]);
  AND2 I281 (rdfint_2n[7], rgrint_2n, df_0n[7]);
  AND2 I282 (rdfint_2n[8], rgrint_2n, df_0n[8]);
  AND2 I283 (rdfint_2n[9], rgrint_2n, df_0n[9]);
  AND2 I284 (rdfint_2n[10], rgrint_2n, df_0n[10]);
  AND2 I285 (rdfint_2n[11], rgrint_2n, df_0n[11]);
  AND2 I286 (rdfint_2n[12], rgrint_2n, df_0n[12]);
  AND2 I287 (rdfint_2n[13], rgrint_2n, df_0n[13]);
  AND2 I288 (rdfint_2n[14], rgrint_2n, df_0n[14]);
  AND2 I289 (rdfint_2n[15], rgrint_2n, df_0n[15]);
  AND2 I290 (rdfint_2n[16], rgrint_2n, df_0n[16]);
  AND2 I291 (rdfint_2n[17], rgrint_2n, df_0n[17]);
  AND2 I292 (rdfint_2n[18], rgrint_2n, df_0n[18]);
  AND2 I293 (rdfint_2n[19], rgrint_2n, df_0n[19]);
  AND2 I294 (rdfint_2n[20], rgrint_2n, df_0n[20]);
  AND2 I295 (rdfint_2n[21], rgrint_2n, df_0n[21]);
  AND2 I296 (rdfint_2n[22], rgrint_2n, df_0n[22]);
  AND2 I297 (rdfint_2n[23], rgrint_2n, df_0n[23]);
  AND2 I298 (rdfint_2n[24], rgrint_2n, df_0n[24]);
  AND2 I299 (rdfint_2n[25], rgrint_2n, df_0n[25]);
  AND2 I300 (rdfint_2n[26], rgrint_2n, df_0n[26]);
  AND2 I301 (rdfint_2n[27], rgrint_2n, df_0n[27]);
  AND2 I302 (rdfint_2n[28], rgrint_2n, df_0n[28]);
  AND2 I303 (rdfint_2n[29], rgrint_2n, df_0n[29]);
  AND2 I304 (rdfint_2n[30], rgrint_2n, df_0n[30]);
  AND2 I305 (rdfint_2n[31], rgrint_2n, df_0n[31]);
  AND2 I306 (rdfint_1n[0], rgrint_1n, df_0n[0]);
  AND2 I307 (rdfint_1n[1], rgrint_1n, df_0n[1]);
  AND2 I308 (rdfint_1n[2], rgrint_1n, df_0n[2]);
  AND2 I309 (rdfint_1n[3], rgrint_1n, df_0n[3]);
  AND2 I310 (rdfint_1n[4], rgrint_1n, df_0n[4]);
  AND2 I311 (rdfint_1n[5], rgrint_1n, df_0n[5]);
  AND2 I312 (rdfint_1n[6], rgrint_1n, df_0n[6]);
  AND2 I313 (rdfint_1n[7], rgrint_1n, df_0n[7]);
  AND2 I314 (rdfint_1n[8], rgrint_1n, df_0n[8]);
  AND2 I315 (rdfint_1n[9], rgrint_1n, df_0n[9]);
  AND2 I316 (rdfint_1n[10], rgrint_1n, df_0n[10]);
  AND2 I317 (rdfint_1n[11], rgrint_1n, df_0n[11]);
  AND2 I318 (rdfint_1n[12], rgrint_1n, df_0n[12]);
  AND2 I319 (rdfint_1n[13], rgrint_1n, df_0n[13]);
  AND2 I320 (rdfint_1n[14], rgrint_1n, df_0n[14]);
  AND2 I321 (rdfint_1n[15], rgrint_1n, df_0n[15]);
  AND2 I322 (rdfint_1n[16], rgrint_1n, df_0n[16]);
  AND2 I323 (rdfint_1n[17], rgrint_1n, df_0n[17]);
  AND2 I324 (rdfint_1n[18], rgrint_1n, df_0n[18]);
  AND2 I325 (rdfint_1n[19], rgrint_1n, df_0n[19]);
  AND2 I326 (rdfint_1n[20], rgrint_1n, df_0n[20]);
  AND2 I327 (rdfint_1n[21], rgrint_1n, df_0n[21]);
  AND2 I328 (rdfint_1n[22], rgrint_1n, df_0n[22]);
  AND2 I329 (rdfint_1n[23], rgrint_1n, df_0n[23]);
  AND2 I330 (rdfint_1n[24], rgrint_1n, df_0n[24]);
  AND2 I331 (rdfint_1n[25], rgrint_1n, df_0n[25]);
  AND2 I332 (rdfint_1n[26], rgrint_1n, df_0n[26]);
  AND2 I333 (rdfint_1n[27], rgrint_1n, df_0n[27]);
  AND2 I334 (rdfint_1n[28], rgrint_1n, df_0n[28]);
  AND2 I335 (rdfint_1n[29], rgrint_1n, df_0n[29]);
  AND2 I336 (rdfint_1n[30], rgrint_1n, df_0n[30]);
  AND2 I337 (rdfint_1n[31], rgrint_1n, df_0n[31]);
  AND2 I338 (rdfint_0n, rgrint_0n, df_0n[31]);
  C3 I339 (internal_0n[2], wc_0n, wacks_0n[31], wacks_0n[30]);
  C3 I340 (internal_0n[3], wacks_0n[29], wacks_0n[28], wacks_0n[27]);
  C3 I341 (internal_0n[4], wacks_0n[26], wacks_0n[25], wacks_0n[24]);
  C3 I342 (internal_0n[5], wacks_0n[23], wacks_0n[22], wacks_0n[21]);
  C3 I343 (internal_0n[6], wacks_0n[20], wacks_0n[19], wacks_0n[18]);
  C3 I344 (internal_0n[7], wacks_0n[17], wacks_0n[16], wacks_0n[15]);
  C3 I345 (internal_0n[8], wacks_0n[14], wacks_0n[13], wacks_0n[12]);
  C3 I346 (internal_0n[9], wacks_0n[11], wacks_0n[10], wacks_0n[9]);
  C3 I347 (internal_0n[10], wacks_0n[8], wacks_0n[7], wacks_0n[6]);
  C3 I348 (internal_0n[11], wacks_0n[5], wacks_0n[4], wacks_0n[3]);
  C3 I349 (internal_0n[12], wacks_0n[2], wacks_0n[1], wacks_0n[0]);
  C3 I350 (internal_0n[13], internal_0n[2], internal_0n[3], internal_0n[4]);
  C3 I351 (internal_0n[14], internal_0n[5], internal_0n[6], internal_0n[7]);
  C3 I352 (internal_0n[15], internal_0n[8], internal_0n[9], internal_0n[10]);
  C2 I353 (internal_0n[16], internal_0n[11], internal_0n[12]);
  C2 I354 (internal_0n[17], internal_0n[13], internal_0n[14]);
  C2 I355 (internal_0n[18], internal_0n[15], internal_0n[16]);
  C2 I356 (wdrint_0n, internal_0n[17], internal_0n[18]);
  assign wen_0n[31] = wc_0n;
  assign wen_0n[30] = wc_0n;
  assign wen_0n[29] = wc_0n;
  assign wen_0n[28] = wc_0n;
  assign wen_0n[27] = wc_0n;
  assign wen_0n[26] = wc_0n;
  assign wen_0n[25] = wc_0n;
  assign wen_0n[24] = wc_0n;
  assign wen_0n[23] = wc_0n;
  assign wen_0n[22] = wc_0n;
  assign wen_0n[21] = wc_0n;
  assign wen_0n[20] = wc_0n;
  assign wen_0n[19] = wc_0n;
  assign wen_0n[18] = wc_0n;
  assign wen_0n[17] = wc_0n;
  assign wen_0n[16] = wc_0n;
  assign wen_0n[15] = wc_0n;
  assign wen_0n[14] = wc_0n;
  assign wen_0n[13] = wc_0n;
  assign wen_0n[12] = wc_0n;
  assign wen_0n[11] = wc_0n;
  assign wen_0n[10] = wc_0n;
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[31] = git_0n[31];
  assign wt_0n[30] = git_0n[30];
  assign wt_0n[29] = git_0n[29];
  assign wt_0n[28] = git_0n[28];
  assign wt_0n[27] = git_0n[27];
  assign wt_0n[26] = git_0n[26];
  assign wt_0n[25] = git_0n[25];
  assign wt_0n[24] = git_0n[24];
  assign wt_0n[23] = git_0n[23];
  assign wt_0n[22] = git_0n[22];
  assign wt_0n[21] = git_0n[21];
  assign wt_0n[20] = git_0n[20];
  assign wt_0n[19] = git_0n[19];
  assign wt_0n[18] = git_0n[18];
  assign wt_0n[17] = git_0n[17];
  assign wt_0n[16] = git_0n[16];
  assign wt_0n[15] = git_0n[15];
  assign wt_0n[14] = git_0n[14];
  assign wt_0n[13] = git_0n[13];
  assign wt_0n[12] = git_0n[12];
  assign wt_0n[11] = git_0n[11];
  assign wt_0n[10] = git_0n[10];
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[31] = gif_0n[31];
  assign wf_0n[30] = gif_0n[30];
  assign wf_0n[29] = gif_0n[29];
  assign wf_0n[28] = gif_0n[28];
  assign wf_0n[27] = gif_0n[27];
  assign wf_0n[26] = gif_0n[26];
  assign wf_0n[25] = gif_0n[25];
  assign wf_0n[24] = gif_0n[24];
  assign wf_0n[23] = gif_0n[23];
  assign wf_0n[22] = gif_0n[22];
  assign wf_0n[21] = gif_0n[21];
  assign wf_0n[20] = gif_0n[20];
  assign wf_0n[19] = gif_0n[19];
  assign wf_0n[18] = gif_0n[18];
  assign wf_0n[17] = gif_0n[17];
  assign wf_0n[16] = gif_0n[16];
  assign wf_0n[15] = gif_0n[15];
  assign wf_0n[14] = gif_0n[14];
  assign wf_0n[13] = gif_0n[13];
  assign wf_0n[12] = gif_0n[12];
  assign wf_0n[11] = gif_0n[11];
  assign wf_0n[10] = gif_0n[10];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I453 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I455 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I456 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I457 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I458 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I459 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I460 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I461 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I462 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I463 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I464 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I465 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I466 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I467 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I468 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I469 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I470 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I471 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I472 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I473 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I474 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I475 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I476 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I477 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I478 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I479 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I480 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I481 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I482 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I483 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I484 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I485 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I486 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I487 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I488 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I489 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I490 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I491 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I492 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I493 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I494 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I495 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I496 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I497 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I498 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I499 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I500 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I501 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I502 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I503 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I504 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I505 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I506 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I507 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I508 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I509 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I510 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I511 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I512 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I513 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I514 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I515 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I516 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I517 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I518 (gif_0n[31], wgfint_0n[31], ig_0n);
  C3 I519 (internal_0n[19], complete1365_0n[0], complete1365_0n[1], complete1365_0n[2]);
  C3 I520 (internal_0n[20], complete1365_0n[3], complete1365_0n[4], complete1365_0n[5]);
  C3 I521 (internal_0n[21], complete1365_0n[6], complete1365_0n[7], complete1365_0n[8]);
  C3 I522 (internal_0n[22], complete1365_0n[9], complete1365_0n[10], complete1365_0n[11]);
  C3 I523 (internal_0n[23], complete1365_0n[12], complete1365_0n[13], complete1365_0n[14]);
  C3 I524 (internal_0n[24], complete1365_0n[15], complete1365_0n[16], complete1365_0n[17]);
  C3 I525 (internal_0n[25], complete1365_0n[18], complete1365_0n[19], complete1365_0n[20]);
  C3 I526 (internal_0n[26], complete1365_0n[21], complete1365_0n[22], complete1365_0n[23]);
  C3 I527 (internal_0n[27], complete1365_0n[24], complete1365_0n[25], complete1365_0n[26]);
  C3 I528 (internal_0n[28], complete1365_0n[27], complete1365_0n[28], complete1365_0n[29]);
  C2 I529 (internal_0n[29], complete1365_0n[30], complete1365_0n[31]);
  C3 I530 (internal_0n[30], internal_0n[19], internal_0n[20], internal_0n[21]);
  C3 I531 (internal_0n[31], internal_0n[22], internal_0n[23], internal_0n[24]);
  C3 I532 (internal_0n[32], internal_0n[25], internal_0n[26], internal_0n[27]);
  C2 I533 (internal_0n[33], internal_0n[28], internal_0n[29]);
  C2 I534 (internal_0n[34], internal_0n[30], internal_0n[31]);
  C2 I535 (internal_0n[35], internal_0n[32], internal_0n[33]);
  C2 I536 (wc_0n, internal_0n[34], internal_0n[35]);
  OR2 I537 (complete1365_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I538 (complete1365_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I539 (complete1365_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I540 (complete1365_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I541 (complete1365_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I542 (complete1365_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I543 (complete1365_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I544 (complete1365_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I545 (complete1365_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I546 (complete1365_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I547 (complete1365_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I548 (complete1365_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I549 (complete1365_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I550 (complete1365_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I551 (complete1365_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I552 (complete1365_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I553 (complete1365_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I554 (complete1365_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I555 (complete1365_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I556 (complete1365_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I557 (complete1365_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I558 (complete1365_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I559 (complete1365_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I560 (complete1365_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I561 (complete1365_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I562 (complete1365_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I563 (complete1365_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I564 (complete1365_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I565 (complete1365_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I566 (complete1365_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I567 (complete1365_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I568 (complete1365_0n[31], wgfint_0n[31], wgtint_0n[31]);
  AO22 I569 (wacks_0n[31], gf1363_0n[31], df_0n[31], gt1364_0n[31], dt_0n[31]);
  NOR2 I570 (dt_0n[31], df_0n[31], gf1363_0n[31]);
  NOR3 I571 (df_0n[31], dt_0n[31], gt1364_0n[31], init_0n);
  AND2 I572 (gt1364_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I573 (gf1363_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I574 (wacks_0n[30], gf1363_0n[30], df_0n[30], gt1364_0n[30], dt_0n[30]);
  NOR2 I575 (dt_0n[30], df_0n[30], gf1363_0n[30]);
  NOR3 I576 (df_0n[30], dt_0n[30], gt1364_0n[30], init_0n);
  AND2 I577 (gt1364_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I578 (gf1363_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I579 (wacks_0n[29], gf1363_0n[29], df_0n[29], gt1364_0n[29], dt_0n[29]);
  NOR2 I580 (dt_0n[29], df_0n[29], gf1363_0n[29]);
  NOR3 I581 (df_0n[29], dt_0n[29], gt1364_0n[29], init_0n);
  AND2 I582 (gt1364_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I583 (gf1363_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I584 (wacks_0n[28], gf1363_0n[28], df_0n[28], gt1364_0n[28], dt_0n[28]);
  NOR2 I585 (dt_0n[28], df_0n[28], gf1363_0n[28]);
  NOR3 I586 (df_0n[28], dt_0n[28], gt1364_0n[28], init_0n);
  AND2 I587 (gt1364_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I588 (gf1363_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I589 (wacks_0n[27], gf1363_0n[27], df_0n[27], gt1364_0n[27], dt_0n[27]);
  NOR2 I590 (dt_0n[27], df_0n[27], gf1363_0n[27]);
  NOR3 I591 (df_0n[27], dt_0n[27], gt1364_0n[27], init_0n);
  AND2 I592 (gt1364_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I593 (gf1363_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I594 (wacks_0n[26], gf1363_0n[26], df_0n[26], gt1364_0n[26], dt_0n[26]);
  NOR2 I595 (dt_0n[26], df_0n[26], gf1363_0n[26]);
  NOR3 I596 (df_0n[26], dt_0n[26], gt1364_0n[26], init_0n);
  AND2 I597 (gt1364_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I598 (gf1363_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I599 (wacks_0n[25], gf1363_0n[25], df_0n[25], gt1364_0n[25], dt_0n[25]);
  NOR2 I600 (dt_0n[25], df_0n[25], gf1363_0n[25]);
  NOR3 I601 (df_0n[25], dt_0n[25], gt1364_0n[25], init_0n);
  AND2 I602 (gt1364_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I603 (gf1363_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I604 (wacks_0n[24], gf1363_0n[24], df_0n[24], gt1364_0n[24], dt_0n[24]);
  NOR2 I605 (dt_0n[24], df_0n[24], gf1363_0n[24]);
  NOR3 I606 (df_0n[24], dt_0n[24], gt1364_0n[24], init_0n);
  AND2 I607 (gt1364_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I608 (gf1363_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I609 (wacks_0n[23], gf1363_0n[23], df_0n[23], gt1364_0n[23], dt_0n[23]);
  NOR2 I610 (dt_0n[23], df_0n[23], gf1363_0n[23]);
  NOR3 I611 (df_0n[23], dt_0n[23], gt1364_0n[23], init_0n);
  AND2 I612 (gt1364_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I613 (gf1363_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I614 (wacks_0n[22], gf1363_0n[22], df_0n[22], gt1364_0n[22], dt_0n[22]);
  NOR2 I615 (dt_0n[22], df_0n[22], gf1363_0n[22]);
  NOR3 I616 (df_0n[22], dt_0n[22], gt1364_0n[22], init_0n);
  AND2 I617 (gt1364_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I618 (gf1363_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I619 (wacks_0n[21], gf1363_0n[21], df_0n[21], gt1364_0n[21], dt_0n[21]);
  NOR2 I620 (dt_0n[21], df_0n[21], gf1363_0n[21]);
  NOR3 I621 (df_0n[21], dt_0n[21], gt1364_0n[21], init_0n);
  AND2 I622 (gt1364_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I623 (gf1363_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I624 (wacks_0n[20], gf1363_0n[20], df_0n[20], gt1364_0n[20], dt_0n[20]);
  NOR2 I625 (dt_0n[20], df_0n[20], gf1363_0n[20]);
  NOR3 I626 (df_0n[20], dt_0n[20], gt1364_0n[20], init_0n);
  AND2 I627 (gt1364_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I628 (gf1363_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I629 (wacks_0n[19], gf1363_0n[19], df_0n[19], gt1364_0n[19], dt_0n[19]);
  NOR2 I630 (dt_0n[19], df_0n[19], gf1363_0n[19]);
  NOR3 I631 (df_0n[19], dt_0n[19], gt1364_0n[19], init_0n);
  AND2 I632 (gt1364_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I633 (gf1363_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I634 (wacks_0n[18], gf1363_0n[18], df_0n[18], gt1364_0n[18], dt_0n[18]);
  NOR2 I635 (dt_0n[18], df_0n[18], gf1363_0n[18]);
  NOR3 I636 (df_0n[18], dt_0n[18], gt1364_0n[18], init_0n);
  AND2 I637 (gt1364_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I638 (gf1363_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I639 (wacks_0n[17], gf1363_0n[17], df_0n[17], gt1364_0n[17], dt_0n[17]);
  NOR2 I640 (dt_0n[17], df_0n[17], gf1363_0n[17]);
  NOR3 I641 (df_0n[17], dt_0n[17], gt1364_0n[17], init_0n);
  AND2 I642 (gt1364_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I643 (gf1363_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I644 (wacks_0n[16], gf1363_0n[16], df_0n[16], gt1364_0n[16], dt_0n[16]);
  NOR2 I645 (dt_0n[16], df_0n[16], gf1363_0n[16]);
  NOR3 I646 (df_0n[16], dt_0n[16], gt1364_0n[16], init_0n);
  AND2 I647 (gt1364_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I648 (gf1363_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I649 (wacks_0n[15], gf1363_0n[15], df_0n[15], gt1364_0n[15], dt_0n[15]);
  NOR2 I650 (dt_0n[15], df_0n[15], gf1363_0n[15]);
  NOR3 I651 (df_0n[15], dt_0n[15], gt1364_0n[15], init_0n);
  AND2 I652 (gt1364_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I653 (gf1363_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I654 (wacks_0n[14], gf1363_0n[14], df_0n[14], gt1364_0n[14], dt_0n[14]);
  NOR2 I655 (dt_0n[14], df_0n[14], gf1363_0n[14]);
  NOR3 I656 (df_0n[14], dt_0n[14], gt1364_0n[14], init_0n);
  AND2 I657 (gt1364_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I658 (gf1363_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I659 (wacks_0n[13], gf1363_0n[13], df_0n[13], gt1364_0n[13], dt_0n[13]);
  NOR2 I660 (dt_0n[13], df_0n[13], gf1363_0n[13]);
  NOR3 I661 (df_0n[13], dt_0n[13], gt1364_0n[13], init_0n);
  AND2 I662 (gt1364_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I663 (gf1363_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I664 (wacks_0n[12], gf1363_0n[12], df_0n[12], gt1364_0n[12], dt_0n[12]);
  NOR2 I665 (dt_0n[12], df_0n[12], gf1363_0n[12]);
  NOR3 I666 (df_0n[12], dt_0n[12], gt1364_0n[12], init_0n);
  AND2 I667 (gt1364_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I668 (gf1363_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I669 (wacks_0n[11], gf1363_0n[11], df_0n[11], gt1364_0n[11], dt_0n[11]);
  NOR2 I670 (dt_0n[11], df_0n[11], gf1363_0n[11]);
  NOR3 I671 (df_0n[11], dt_0n[11], gt1364_0n[11], init_0n);
  AND2 I672 (gt1364_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I673 (gf1363_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I674 (wacks_0n[10], gf1363_0n[10], df_0n[10], gt1364_0n[10], dt_0n[10]);
  NOR2 I675 (dt_0n[10], df_0n[10], gf1363_0n[10]);
  NOR3 I676 (df_0n[10], dt_0n[10], gt1364_0n[10], init_0n);
  AND2 I677 (gt1364_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I678 (gf1363_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I679 (wacks_0n[9], gf1363_0n[9], df_0n[9], gt1364_0n[9], dt_0n[9]);
  NOR2 I680 (dt_0n[9], df_0n[9], gf1363_0n[9]);
  NOR3 I681 (df_0n[9], dt_0n[9], gt1364_0n[9], init_0n);
  AND2 I682 (gt1364_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I683 (gf1363_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I684 (wacks_0n[8], gf1363_0n[8], df_0n[8], gt1364_0n[8], dt_0n[8]);
  NOR2 I685 (dt_0n[8], df_0n[8], gf1363_0n[8]);
  NOR3 I686 (df_0n[8], dt_0n[8], gt1364_0n[8], init_0n);
  AND2 I687 (gt1364_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I688 (gf1363_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I689 (wacks_0n[7], gf1363_0n[7], df_0n[7], gt1364_0n[7], dt_0n[7]);
  NOR2 I690 (dt_0n[7], df_0n[7], gf1363_0n[7]);
  NOR3 I691 (df_0n[7], dt_0n[7], gt1364_0n[7], init_0n);
  AND2 I692 (gt1364_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I693 (gf1363_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I694 (wacks_0n[6], gf1363_0n[6], df_0n[6], gt1364_0n[6], dt_0n[6]);
  NOR2 I695 (dt_0n[6], df_0n[6], gf1363_0n[6]);
  NOR3 I696 (df_0n[6], dt_0n[6], gt1364_0n[6], init_0n);
  AND2 I697 (gt1364_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I698 (gf1363_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I699 (wacks_0n[5], gf1363_0n[5], df_0n[5], gt1364_0n[5], dt_0n[5]);
  NOR2 I700 (dt_0n[5], df_0n[5], gf1363_0n[5]);
  NOR3 I701 (df_0n[5], dt_0n[5], gt1364_0n[5], init_0n);
  AND2 I702 (gt1364_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I703 (gf1363_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I704 (wacks_0n[4], gf1363_0n[4], df_0n[4], gt1364_0n[4], dt_0n[4]);
  NOR2 I705 (dt_0n[4], df_0n[4], gf1363_0n[4]);
  NOR3 I706 (df_0n[4], dt_0n[4], gt1364_0n[4], init_0n);
  AND2 I707 (gt1364_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I708 (gf1363_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I709 (wacks_0n[3], gf1363_0n[3], df_0n[3], gt1364_0n[3], dt_0n[3]);
  NOR2 I710 (dt_0n[3], df_0n[3], gf1363_0n[3]);
  NOR3 I711 (df_0n[3], dt_0n[3], gt1364_0n[3], init_0n);
  AND2 I712 (gt1364_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I713 (gf1363_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I714 (wacks_0n[2], gf1363_0n[2], df_0n[2], gt1364_0n[2], dt_0n[2]);
  NOR2 I715 (dt_0n[2], df_0n[2], gf1363_0n[2]);
  NOR3 I716 (df_0n[2], dt_0n[2], gt1364_0n[2], init_0n);
  AND2 I717 (gt1364_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I718 (gf1363_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I719 (wacks_0n[1], gf1363_0n[1], df_0n[1], gt1364_0n[1], dt_0n[1]);
  NOR2 I720 (dt_0n[1], df_0n[1], gf1363_0n[1]);
  NOR3 I721 (df_0n[1], dt_0n[1], gt1364_0n[1], init_0n);
  AND2 I722 (gt1364_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I723 (gf1363_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I724 (wacks_0n[0], gf1363_0n[0], df_0n[0], gt1364_0n[0], dt_0n[0]);
  NOR2 I725 (dt_0n[0], df_0n[0], gf1363_0n[0]);
  NOR3 I726 (df_0n[0], dt_0n[0], gt1364_0n[0], init_0n);
  AND2 I727 (gt1364_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I728 (gf1363_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I729 (init_0n, initialise);
endmodule

module BrzV_33_l6__28_29_l24__28_28_280_2033_29_2_m84m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rd_0r0d, rd_0r1d, rd_0a,
  initialise
);
  input [32:0] wg_0r0d;
  input [32:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [32:0] rd_0r0d;
  output [32:0] rd_0r1d;
  input rd_0a;
  input initialise;
  wire [34:0] internal_0n;
  wire [32:0] wf_0n;
  wire [32:0] wt_0n;
  wire [32:0] df_0n;
  wire [32:0] dt_0n;
  wire rgrint_0n;
  wire wc_0n;
  wire [32:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [32:0] wgfint_0n;
  wire [32:0] wgtint_0n;
  wire rgaint_0n;
  wire [32:0] rdfint_0n;
  wire [32:0] rdtint_0n;
  wire [32:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [32:0] gif_0n;
  wire [32:0] git_0n;
  wire [32:0] complete1384_0n;
  wire [32:0] gt1383_0n;
  wire [32:0] gf1382_0n;
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r0d[10] = rdfint_0n[10];
  assign rd_0r0d[11] = rdfint_0n[11];
  assign rd_0r0d[12] = rdfint_0n[12];
  assign rd_0r0d[13] = rdfint_0n[13];
  assign rd_0r0d[14] = rdfint_0n[14];
  assign rd_0r0d[15] = rdfint_0n[15];
  assign rd_0r0d[16] = rdfint_0n[16];
  assign rd_0r0d[17] = rdfint_0n[17];
  assign rd_0r0d[18] = rdfint_0n[18];
  assign rd_0r0d[19] = rdfint_0n[19];
  assign rd_0r0d[20] = rdfint_0n[20];
  assign rd_0r0d[21] = rdfint_0n[21];
  assign rd_0r0d[22] = rdfint_0n[22];
  assign rd_0r0d[23] = rdfint_0n[23];
  assign rd_0r0d[24] = rdfint_0n[24];
  assign rd_0r0d[25] = rdfint_0n[25];
  assign rd_0r0d[26] = rdfint_0n[26];
  assign rd_0r0d[27] = rdfint_0n[27];
  assign rd_0r0d[28] = rdfint_0n[28];
  assign rd_0r0d[29] = rdfint_0n[29];
  assign rd_0r0d[30] = rdfint_0n[30];
  assign rd_0r0d[31] = rdfint_0n[31];
  assign rd_0r0d[32] = rdfint_0n[32];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign rd_0r1d[10] = rdtint_0n[10];
  assign rd_0r1d[11] = rdtint_0n[11];
  assign rd_0r1d[12] = rdtint_0n[12];
  assign rd_0r1d[13] = rdtint_0n[13];
  assign rd_0r1d[14] = rdtint_0n[14];
  assign rd_0r1d[15] = rdtint_0n[15];
  assign rd_0r1d[16] = rdtint_0n[16];
  assign rd_0r1d[17] = rdtint_0n[17];
  assign rd_0r1d[18] = rdtint_0n[18];
  assign rd_0r1d[19] = rdtint_0n[19];
  assign rd_0r1d[20] = rdtint_0n[20];
  assign rd_0r1d[21] = rdtint_0n[21];
  assign rd_0r1d[22] = rdtint_0n[22];
  assign rd_0r1d[23] = rdtint_0n[23];
  assign rd_0r1d[24] = rdtint_0n[24];
  assign rd_0r1d[25] = rdtint_0n[25];
  assign rd_0r1d[26] = rdtint_0n[26];
  assign rd_0r1d[27] = rdtint_0n[27];
  assign rd_0r1d[28] = rdtint_0n[28];
  assign rd_0r1d[29] = rdtint_0n[29];
  assign rd_0r1d[30] = rdtint_0n[30];
  assign rd_0r1d[31] = rdtint_0n[31];
  assign rd_0r1d[32] = rdtint_0n[32];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgfint_0n[32] = wg_0r0d[32];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign wgtint_0n[32] = wg_0r1d[32];
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I138 (nanyread_0n, rgrint_0n, rgaint_0n);
  AND2 I139 (rdtint_0n[0], rgrint_0n, dt_0n[0]);
  AND2 I140 (rdtint_0n[1], rgrint_0n, dt_0n[1]);
  AND2 I141 (rdtint_0n[2], rgrint_0n, dt_0n[2]);
  AND2 I142 (rdtint_0n[3], rgrint_0n, dt_0n[3]);
  AND2 I143 (rdtint_0n[4], rgrint_0n, dt_0n[4]);
  AND2 I144 (rdtint_0n[5], rgrint_0n, dt_0n[5]);
  AND2 I145 (rdtint_0n[6], rgrint_0n, dt_0n[6]);
  AND2 I146 (rdtint_0n[7], rgrint_0n, dt_0n[7]);
  AND2 I147 (rdtint_0n[8], rgrint_0n, dt_0n[8]);
  AND2 I148 (rdtint_0n[9], rgrint_0n, dt_0n[9]);
  AND2 I149 (rdtint_0n[10], rgrint_0n, dt_0n[10]);
  AND2 I150 (rdtint_0n[11], rgrint_0n, dt_0n[11]);
  AND2 I151 (rdtint_0n[12], rgrint_0n, dt_0n[12]);
  AND2 I152 (rdtint_0n[13], rgrint_0n, dt_0n[13]);
  AND2 I153 (rdtint_0n[14], rgrint_0n, dt_0n[14]);
  AND2 I154 (rdtint_0n[15], rgrint_0n, dt_0n[15]);
  AND2 I155 (rdtint_0n[16], rgrint_0n, dt_0n[16]);
  AND2 I156 (rdtint_0n[17], rgrint_0n, dt_0n[17]);
  AND2 I157 (rdtint_0n[18], rgrint_0n, dt_0n[18]);
  AND2 I158 (rdtint_0n[19], rgrint_0n, dt_0n[19]);
  AND2 I159 (rdtint_0n[20], rgrint_0n, dt_0n[20]);
  AND2 I160 (rdtint_0n[21], rgrint_0n, dt_0n[21]);
  AND2 I161 (rdtint_0n[22], rgrint_0n, dt_0n[22]);
  AND2 I162 (rdtint_0n[23], rgrint_0n, dt_0n[23]);
  AND2 I163 (rdtint_0n[24], rgrint_0n, dt_0n[24]);
  AND2 I164 (rdtint_0n[25], rgrint_0n, dt_0n[25]);
  AND2 I165 (rdtint_0n[26], rgrint_0n, dt_0n[26]);
  AND2 I166 (rdtint_0n[27], rgrint_0n, dt_0n[27]);
  AND2 I167 (rdtint_0n[28], rgrint_0n, dt_0n[28]);
  AND2 I168 (rdtint_0n[29], rgrint_0n, dt_0n[29]);
  AND2 I169 (rdtint_0n[30], rgrint_0n, dt_0n[30]);
  AND2 I170 (rdtint_0n[31], rgrint_0n, dt_0n[31]);
  AND2 I171 (rdtint_0n[32], rgrint_0n, dt_0n[32]);
  AND2 I172 (rdfint_0n[0], rgrint_0n, df_0n[0]);
  AND2 I173 (rdfint_0n[1], rgrint_0n, df_0n[1]);
  AND2 I174 (rdfint_0n[2], rgrint_0n, df_0n[2]);
  AND2 I175 (rdfint_0n[3], rgrint_0n, df_0n[3]);
  AND2 I176 (rdfint_0n[4], rgrint_0n, df_0n[4]);
  AND2 I177 (rdfint_0n[5], rgrint_0n, df_0n[5]);
  AND2 I178 (rdfint_0n[6], rgrint_0n, df_0n[6]);
  AND2 I179 (rdfint_0n[7], rgrint_0n, df_0n[7]);
  AND2 I180 (rdfint_0n[8], rgrint_0n, df_0n[8]);
  AND2 I181 (rdfint_0n[9], rgrint_0n, df_0n[9]);
  AND2 I182 (rdfint_0n[10], rgrint_0n, df_0n[10]);
  AND2 I183 (rdfint_0n[11], rgrint_0n, df_0n[11]);
  AND2 I184 (rdfint_0n[12], rgrint_0n, df_0n[12]);
  AND2 I185 (rdfint_0n[13], rgrint_0n, df_0n[13]);
  AND2 I186 (rdfint_0n[14], rgrint_0n, df_0n[14]);
  AND2 I187 (rdfint_0n[15], rgrint_0n, df_0n[15]);
  AND2 I188 (rdfint_0n[16], rgrint_0n, df_0n[16]);
  AND2 I189 (rdfint_0n[17], rgrint_0n, df_0n[17]);
  AND2 I190 (rdfint_0n[18], rgrint_0n, df_0n[18]);
  AND2 I191 (rdfint_0n[19], rgrint_0n, df_0n[19]);
  AND2 I192 (rdfint_0n[20], rgrint_0n, df_0n[20]);
  AND2 I193 (rdfint_0n[21], rgrint_0n, df_0n[21]);
  AND2 I194 (rdfint_0n[22], rgrint_0n, df_0n[22]);
  AND2 I195 (rdfint_0n[23], rgrint_0n, df_0n[23]);
  AND2 I196 (rdfint_0n[24], rgrint_0n, df_0n[24]);
  AND2 I197 (rdfint_0n[25], rgrint_0n, df_0n[25]);
  AND2 I198 (rdfint_0n[26], rgrint_0n, df_0n[26]);
  AND2 I199 (rdfint_0n[27], rgrint_0n, df_0n[27]);
  AND2 I200 (rdfint_0n[28], rgrint_0n, df_0n[28]);
  AND2 I201 (rdfint_0n[29], rgrint_0n, df_0n[29]);
  AND2 I202 (rdfint_0n[30], rgrint_0n, df_0n[30]);
  AND2 I203 (rdfint_0n[31], rgrint_0n, df_0n[31]);
  AND2 I204 (rdfint_0n[32], rgrint_0n, df_0n[32]);
  C3 I205 (internal_0n[0], wc_0n, wacks_0n[32], wacks_0n[31]);
  C3 I206 (internal_0n[1], wacks_0n[30], wacks_0n[29], wacks_0n[28]);
  C3 I207 (internal_0n[2], wacks_0n[27], wacks_0n[26], wacks_0n[25]);
  C3 I208 (internal_0n[3], wacks_0n[24], wacks_0n[23], wacks_0n[22]);
  C3 I209 (internal_0n[4], wacks_0n[21], wacks_0n[20], wacks_0n[19]);
  C3 I210 (internal_0n[5], wacks_0n[18], wacks_0n[17], wacks_0n[16]);
  C3 I211 (internal_0n[6], wacks_0n[15], wacks_0n[14], wacks_0n[13]);
  C3 I212 (internal_0n[7], wacks_0n[12], wacks_0n[11], wacks_0n[10]);
  C3 I213 (internal_0n[8], wacks_0n[9], wacks_0n[8], wacks_0n[7]);
  C3 I214 (internal_0n[9], wacks_0n[6], wacks_0n[5], wacks_0n[4]);
  C2 I215 (internal_0n[10], wacks_0n[3], wacks_0n[2]);
  C2 I216 (internal_0n[11], wacks_0n[1], wacks_0n[0]);
  C3 I217 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I218 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I219 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I220 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I221 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I222 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I223 (wdrint_0n, internal_0n[16], internal_0n[17]);
  assign wen_0n[32] = wc_0n;
  assign wen_0n[31] = wc_0n;
  assign wen_0n[30] = wc_0n;
  assign wen_0n[29] = wc_0n;
  assign wen_0n[28] = wc_0n;
  assign wen_0n[27] = wc_0n;
  assign wen_0n[26] = wc_0n;
  assign wen_0n[25] = wc_0n;
  assign wen_0n[24] = wc_0n;
  assign wen_0n[23] = wc_0n;
  assign wen_0n[22] = wc_0n;
  assign wen_0n[21] = wc_0n;
  assign wen_0n[20] = wc_0n;
  assign wen_0n[19] = wc_0n;
  assign wen_0n[18] = wc_0n;
  assign wen_0n[17] = wc_0n;
  assign wen_0n[16] = wc_0n;
  assign wen_0n[15] = wc_0n;
  assign wen_0n[14] = wc_0n;
  assign wen_0n[13] = wc_0n;
  assign wen_0n[12] = wc_0n;
  assign wen_0n[11] = wc_0n;
  assign wen_0n[10] = wc_0n;
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[32] = git_0n[32];
  assign wt_0n[31] = git_0n[31];
  assign wt_0n[30] = git_0n[30];
  assign wt_0n[29] = git_0n[29];
  assign wt_0n[28] = git_0n[28];
  assign wt_0n[27] = git_0n[27];
  assign wt_0n[26] = git_0n[26];
  assign wt_0n[25] = git_0n[25];
  assign wt_0n[24] = git_0n[24];
  assign wt_0n[23] = git_0n[23];
  assign wt_0n[22] = git_0n[22];
  assign wt_0n[21] = git_0n[21];
  assign wt_0n[20] = git_0n[20];
  assign wt_0n[19] = git_0n[19];
  assign wt_0n[18] = git_0n[18];
  assign wt_0n[17] = git_0n[17];
  assign wt_0n[16] = git_0n[16];
  assign wt_0n[15] = git_0n[15];
  assign wt_0n[14] = git_0n[14];
  assign wt_0n[13] = git_0n[13];
  assign wt_0n[12] = git_0n[12];
  assign wt_0n[11] = git_0n[11];
  assign wt_0n[10] = git_0n[10];
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[32] = gif_0n[32];
  assign wf_0n[31] = gif_0n[31];
  assign wf_0n[30] = gif_0n[30];
  assign wf_0n[29] = gif_0n[29];
  assign wf_0n[28] = gif_0n[28];
  assign wf_0n[27] = gif_0n[27];
  assign wf_0n[26] = gif_0n[26];
  assign wf_0n[25] = gif_0n[25];
  assign wf_0n[24] = gif_0n[24];
  assign wf_0n[23] = gif_0n[23];
  assign wf_0n[22] = gif_0n[22];
  assign wf_0n[21] = gif_0n[21];
  assign wf_0n[20] = gif_0n[20];
  assign wf_0n[19] = gif_0n[19];
  assign wf_0n[18] = gif_0n[18];
  assign wf_0n[17] = gif_0n[17];
  assign wf_0n[16] = gif_0n[16];
  assign wf_0n[15] = gif_0n[15];
  assign wf_0n[14] = gif_0n[14];
  assign wf_0n[13] = gif_0n[13];
  assign wf_0n[12] = gif_0n[12];
  assign wf_0n[11] = gif_0n[11];
  assign wf_0n[10] = gif_0n[10];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I323 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I325 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I326 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I327 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I328 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I329 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I330 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I331 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I332 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I333 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I334 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I335 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I336 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I337 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I338 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I339 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I340 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I341 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I342 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I343 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I344 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I345 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I346 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I347 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I348 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I349 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I350 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I351 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I352 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I353 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I354 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I355 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I356 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I357 (git_0n[32], wgtint_0n[32], ig_0n);
  AND2 I358 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I359 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I360 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I361 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I362 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I363 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I364 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I365 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I366 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I367 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I368 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I369 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I370 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I371 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I372 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I373 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I374 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I375 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I376 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I377 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I378 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I379 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I380 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I381 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I382 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I383 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I384 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I385 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I386 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I387 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I388 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I389 (gif_0n[31], wgfint_0n[31], ig_0n);
  AND2 I390 (gif_0n[32], wgfint_0n[32], ig_0n);
  C3 I391 (internal_0n[18], complete1384_0n[0], complete1384_0n[1], complete1384_0n[2]);
  C3 I392 (internal_0n[19], complete1384_0n[3], complete1384_0n[4], complete1384_0n[5]);
  C3 I393 (internal_0n[20], complete1384_0n[6], complete1384_0n[7], complete1384_0n[8]);
  C3 I394 (internal_0n[21], complete1384_0n[9], complete1384_0n[10], complete1384_0n[11]);
  C3 I395 (internal_0n[22], complete1384_0n[12], complete1384_0n[13], complete1384_0n[14]);
  C3 I396 (internal_0n[23], complete1384_0n[15], complete1384_0n[16], complete1384_0n[17]);
  C3 I397 (internal_0n[24], complete1384_0n[18], complete1384_0n[19], complete1384_0n[20]);
  C3 I398 (internal_0n[25], complete1384_0n[21], complete1384_0n[22], complete1384_0n[23]);
  C3 I399 (internal_0n[26], complete1384_0n[24], complete1384_0n[25], complete1384_0n[26]);
  C3 I400 (internal_0n[27], complete1384_0n[27], complete1384_0n[28], complete1384_0n[29]);
  C3 I401 (internal_0n[28], complete1384_0n[30], complete1384_0n[31], complete1384_0n[32]);
  C3 I402 (internal_0n[29], internal_0n[18], internal_0n[19], internal_0n[20]);
  C3 I403 (internal_0n[30], internal_0n[21], internal_0n[22], internal_0n[23]);
  C3 I404 (internal_0n[31], internal_0n[24], internal_0n[25], internal_0n[26]);
  C2 I405 (internal_0n[32], internal_0n[27], internal_0n[28]);
  C2 I406 (internal_0n[33], internal_0n[29], internal_0n[30]);
  C2 I407 (internal_0n[34], internal_0n[31], internal_0n[32]);
  C2 I408 (wc_0n, internal_0n[33], internal_0n[34]);
  OR2 I409 (complete1384_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I410 (complete1384_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I411 (complete1384_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I412 (complete1384_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I413 (complete1384_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I414 (complete1384_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I415 (complete1384_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I416 (complete1384_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I417 (complete1384_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I418 (complete1384_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I419 (complete1384_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I420 (complete1384_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I421 (complete1384_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I422 (complete1384_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I423 (complete1384_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I424 (complete1384_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I425 (complete1384_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I426 (complete1384_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I427 (complete1384_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I428 (complete1384_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I429 (complete1384_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I430 (complete1384_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I431 (complete1384_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I432 (complete1384_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I433 (complete1384_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I434 (complete1384_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I435 (complete1384_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I436 (complete1384_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I437 (complete1384_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I438 (complete1384_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I439 (complete1384_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I440 (complete1384_0n[31], wgfint_0n[31], wgtint_0n[31]);
  OR2 I441 (complete1384_0n[32], wgfint_0n[32], wgtint_0n[32]);
  AO22 I442 (wacks_0n[32], gf1382_0n[32], df_0n[32], gt1383_0n[32], dt_0n[32]);
  NOR2 I443 (dt_0n[32], df_0n[32], gf1382_0n[32]);
  NOR3 I444 (df_0n[32], dt_0n[32], gt1383_0n[32], init_0n);
  AND2 I445 (gt1383_0n[32], wt_0n[32], wen_0n[32]);
  AND2 I446 (gf1382_0n[32], wf_0n[32], wen_0n[32]);
  AO22 I447 (wacks_0n[31], gf1382_0n[31], df_0n[31], gt1383_0n[31], dt_0n[31]);
  NOR2 I448 (dt_0n[31], df_0n[31], gf1382_0n[31]);
  NOR3 I449 (df_0n[31], dt_0n[31], gt1383_0n[31], init_0n);
  AND2 I450 (gt1383_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I451 (gf1382_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I452 (wacks_0n[30], gf1382_0n[30], df_0n[30], gt1383_0n[30], dt_0n[30]);
  NOR2 I453 (dt_0n[30], df_0n[30], gf1382_0n[30]);
  NOR3 I454 (df_0n[30], dt_0n[30], gt1383_0n[30], init_0n);
  AND2 I455 (gt1383_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I456 (gf1382_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I457 (wacks_0n[29], gf1382_0n[29], df_0n[29], gt1383_0n[29], dt_0n[29]);
  NOR2 I458 (dt_0n[29], df_0n[29], gf1382_0n[29]);
  NOR3 I459 (df_0n[29], dt_0n[29], gt1383_0n[29], init_0n);
  AND2 I460 (gt1383_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I461 (gf1382_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I462 (wacks_0n[28], gf1382_0n[28], df_0n[28], gt1383_0n[28], dt_0n[28]);
  NOR2 I463 (dt_0n[28], df_0n[28], gf1382_0n[28]);
  NOR3 I464 (df_0n[28], dt_0n[28], gt1383_0n[28], init_0n);
  AND2 I465 (gt1383_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I466 (gf1382_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I467 (wacks_0n[27], gf1382_0n[27], df_0n[27], gt1383_0n[27], dt_0n[27]);
  NOR2 I468 (dt_0n[27], df_0n[27], gf1382_0n[27]);
  NOR3 I469 (df_0n[27], dt_0n[27], gt1383_0n[27], init_0n);
  AND2 I470 (gt1383_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I471 (gf1382_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I472 (wacks_0n[26], gf1382_0n[26], df_0n[26], gt1383_0n[26], dt_0n[26]);
  NOR2 I473 (dt_0n[26], df_0n[26], gf1382_0n[26]);
  NOR3 I474 (df_0n[26], dt_0n[26], gt1383_0n[26], init_0n);
  AND2 I475 (gt1383_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I476 (gf1382_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I477 (wacks_0n[25], gf1382_0n[25], df_0n[25], gt1383_0n[25], dt_0n[25]);
  NOR2 I478 (dt_0n[25], df_0n[25], gf1382_0n[25]);
  NOR3 I479 (df_0n[25], dt_0n[25], gt1383_0n[25], init_0n);
  AND2 I480 (gt1383_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I481 (gf1382_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I482 (wacks_0n[24], gf1382_0n[24], df_0n[24], gt1383_0n[24], dt_0n[24]);
  NOR2 I483 (dt_0n[24], df_0n[24], gf1382_0n[24]);
  NOR3 I484 (df_0n[24], dt_0n[24], gt1383_0n[24], init_0n);
  AND2 I485 (gt1383_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I486 (gf1382_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I487 (wacks_0n[23], gf1382_0n[23], df_0n[23], gt1383_0n[23], dt_0n[23]);
  NOR2 I488 (dt_0n[23], df_0n[23], gf1382_0n[23]);
  NOR3 I489 (df_0n[23], dt_0n[23], gt1383_0n[23], init_0n);
  AND2 I490 (gt1383_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I491 (gf1382_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I492 (wacks_0n[22], gf1382_0n[22], df_0n[22], gt1383_0n[22], dt_0n[22]);
  NOR2 I493 (dt_0n[22], df_0n[22], gf1382_0n[22]);
  NOR3 I494 (df_0n[22], dt_0n[22], gt1383_0n[22], init_0n);
  AND2 I495 (gt1383_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I496 (gf1382_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I497 (wacks_0n[21], gf1382_0n[21], df_0n[21], gt1383_0n[21], dt_0n[21]);
  NOR2 I498 (dt_0n[21], df_0n[21], gf1382_0n[21]);
  NOR3 I499 (df_0n[21], dt_0n[21], gt1383_0n[21], init_0n);
  AND2 I500 (gt1383_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I501 (gf1382_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I502 (wacks_0n[20], gf1382_0n[20], df_0n[20], gt1383_0n[20], dt_0n[20]);
  NOR2 I503 (dt_0n[20], df_0n[20], gf1382_0n[20]);
  NOR3 I504 (df_0n[20], dt_0n[20], gt1383_0n[20], init_0n);
  AND2 I505 (gt1383_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I506 (gf1382_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I507 (wacks_0n[19], gf1382_0n[19], df_0n[19], gt1383_0n[19], dt_0n[19]);
  NOR2 I508 (dt_0n[19], df_0n[19], gf1382_0n[19]);
  NOR3 I509 (df_0n[19], dt_0n[19], gt1383_0n[19], init_0n);
  AND2 I510 (gt1383_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I511 (gf1382_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I512 (wacks_0n[18], gf1382_0n[18], df_0n[18], gt1383_0n[18], dt_0n[18]);
  NOR2 I513 (dt_0n[18], df_0n[18], gf1382_0n[18]);
  NOR3 I514 (df_0n[18], dt_0n[18], gt1383_0n[18], init_0n);
  AND2 I515 (gt1383_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I516 (gf1382_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I517 (wacks_0n[17], gf1382_0n[17], df_0n[17], gt1383_0n[17], dt_0n[17]);
  NOR2 I518 (dt_0n[17], df_0n[17], gf1382_0n[17]);
  NOR3 I519 (df_0n[17], dt_0n[17], gt1383_0n[17], init_0n);
  AND2 I520 (gt1383_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I521 (gf1382_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I522 (wacks_0n[16], gf1382_0n[16], df_0n[16], gt1383_0n[16], dt_0n[16]);
  NOR2 I523 (dt_0n[16], df_0n[16], gf1382_0n[16]);
  NOR3 I524 (df_0n[16], dt_0n[16], gt1383_0n[16], init_0n);
  AND2 I525 (gt1383_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I526 (gf1382_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I527 (wacks_0n[15], gf1382_0n[15], df_0n[15], gt1383_0n[15], dt_0n[15]);
  NOR2 I528 (dt_0n[15], df_0n[15], gf1382_0n[15]);
  NOR3 I529 (df_0n[15], dt_0n[15], gt1383_0n[15], init_0n);
  AND2 I530 (gt1383_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I531 (gf1382_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I532 (wacks_0n[14], gf1382_0n[14], df_0n[14], gt1383_0n[14], dt_0n[14]);
  NOR2 I533 (dt_0n[14], df_0n[14], gf1382_0n[14]);
  NOR3 I534 (df_0n[14], dt_0n[14], gt1383_0n[14], init_0n);
  AND2 I535 (gt1383_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I536 (gf1382_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I537 (wacks_0n[13], gf1382_0n[13], df_0n[13], gt1383_0n[13], dt_0n[13]);
  NOR2 I538 (dt_0n[13], df_0n[13], gf1382_0n[13]);
  NOR3 I539 (df_0n[13], dt_0n[13], gt1383_0n[13], init_0n);
  AND2 I540 (gt1383_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I541 (gf1382_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I542 (wacks_0n[12], gf1382_0n[12], df_0n[12], gt1383_0n[12], dt_0n[12]);
  NOR2 I543 (dt_0n[12], df_0n[12], gf1382_0n[12]);
  NOR3 I544 (df_0n[12], dt_0n[12], gt1383_0n[12], init_0n);
  AND2 I545 (gt1383_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I546 (gf1382_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I547 (wacks_0n[11], gf1382_0n[11], df_0n[11], gt1383_0n[11], dt_0n[11]);
  NOR2 I548 (dt_0n[11], df_0n[11], gf1382_0n[11]);
  NOR3 I549 (df_0n[11], dt_0n[11], gt1383_0n[11], init_0n);
  AND2 I550 (gt1383_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I551 (gf1382_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I552 (wacks_0n[10], gf1382_0n[10], df_0n[10], gt1383_0n[10], dt_0n[10]);
  NOR2 I553 (dt_0n[10], df_0n[10], gf1382_0n[10]);
  NOR3 I554 (df_0n[10], dt_0n[10], gt1383_0n[10], init_0n);
  AND2 I555 (gt1383_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I556 (gf1382_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I557 (wacks_0n[9], gf1382_0n[9], df_0n[9], gt1383_0n[9], dt_0n[9]);
  NOR2 I558 (dt_0n[9], df_0n[9], gf1382_0n[9]);
  NOR3 I559 (df_0n[9], dt_0n[9], gt1383_0n[9], init_0n);
  AND2 I560 (gt1383_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I561 (gf1382_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I562 (wacks_0n[8], gf1382_0n[8], df_0n[8], gt1383_0n[8], dt_0n[8]);
  NOR2 I563 (dt_0n[8], df_0n[8], gf1382_0n[8]);
  NOR3 I564 (df_0n[8], dt_0n[8], gt1383_0n[8], init_0n);
  AND2 I565 (gt1383_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I566 (gf1382_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I567 (wacks_0n[7], gf1382_0n[7], df_0n[7], gt1383_0n[7], dt_0n[7]);
  NOR2 I568 (dt_0n[7], df_0n[7], gf1382_0n[7]);
  NOR3 I569 (df_0n[7], dt_0n[7], gt1383_0n[7], init_0n);
  AND2 I570 (gt1383_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I571 (gf1382_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I572 (wacks_0n[6], gf1382_0n[6], df_0n[6], gt1383_0n[6], dt_0n[6]);
  NOR2 I573 (dt_0n[6], df_0n[6], gf1382_0n[6]);
  NOR3 I574 (df_0n[6], dt_0n[6], gt1383_0n[6], init_0n);
  AND2 I575 (gt1383_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I576 (gf1382_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I577 (wacks_0n[5], gf1382_0n[5], df_0n[5], gt1383_0n[5], dt_0n[5]);
  NOR2 I578 (dt_0n[5], df_0n[5], gf1382_0n[5]);
  NOR3 I579 (df_0n[5], dt_0n[5], gt1383_0n[5], init_0n);
  AND2 I580 (gt1383_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I581 (gf1382_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I582 (wacks_0n[4], gf1382_0n[4], df_0n[4], gt1383_0n[4], dt_0n[4]);
  NOR2 I583 (dt_0n[4], df_0n[4], gf1382_0n[4]);
  NOR3 I584 (df_0n[4], dt_0n[4], gt1383_0n[4], init_0n);
  AND2 I585 (gt1383_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I586 (gf1382_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I587 (wacks_0n[3], gf1382_0n[3], df_0n[3], gt1383_0n[3], dt_0n[3]);
  NOR2 I588 (dt_0n[3], df_0n[3], gf1382_0n[3]);
  NOR3 I589 (df_0n[3], dt_0n[3], gt1383_0n[3], init_0n);
  AND2 I590 (gt1383_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I591 (gf1382_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I592 (wacks_0n[2], gf1382_0n[2], df_0n[2], gt1383_0n[2], dt_0n[2]);
  NOR2 I593 (dt_0n[2], df_0n[2], gf1382_0n[2]);
  NOR3 I594 (df_0n[2], dt_0n[2], gt1383_0n[2], init_0n);
  AND2 I595 (gt1383_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I596 (gf1382_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I597 (wacks_0n[1], gf1382_0n[1], df_0n[1], gt1383_0n[1], dt_0n[1]);
  NOR2 I598 (dt_0n[1], df_0n[1], gf1382_0n[1]);
  NOR3 I599 (df_0n[1], dt_0n[1], gt1383_0n[1], init_0n);
  AND2 I600 (gt1383_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I601 (gf1382_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I602 (wacks_0n[0], gf1382_0n[0], df_0n[0], gt1383_0n[0], dt_0n[0]);
  NOR2 I603 (dt_0n[0], df_0n[0], gf1382_0n[0]);
  NOR3 I604 (df_0n[0], dt_0n[0], gt1383_0n[0], init_0n);
  AND2 I605 (gt1383_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I606 (gf1382_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I607 (init_0n, initialise);
endmodule

module BrzV_34_l6__28_29_l24__28_28_280_2034_29_2_m85m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  initialise
);
  input [33:0] wg_0r0d;
  input [33:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [31:0] rd_0r0d;
  output [31:0] rd_0r1d;
  input rd_0a;
  output rd_1r0d;
  output rd_1r1d;
  input rd_1a;
  input initialise;
  wire [37:0] internal_0n;
  wire [33:0] wf_0n;
  wire [33:0] wt_0n;
  wire [33:0] df_0n;
  wire [33:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire wc_0n;
  wire [33:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [33:0] wgfint_0n;
  wire [33:0] wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire [31:0] rdfint_0n;
  wire rdfint_1n;
  wire [31:0] rdtint_0n;
  wire rdtint_1n;
  wire [33:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [33:0] gif_0n;
  wire [33:0] git_0n;
  wire [33:0] complete1395_0n;
  wire [33:0] gt1394_0n;
  wire [33:0] gf1393_0n;
  assign rgaint_1n = rd_1a;
  assign rd_1r0d = rdfint_1n;
  assign rd_1r1d = rdtint_1n;
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r0d[10] = rdfint_0n[10];
  assign rd_0r0d[11] = rdfint_0n[11];
  assign rd_0r0d[12] = rdfint_0n[12];
  assign rd_0r0d[13] = rdfint_0n[13];
  assign rd_0r0d[14] = rdfint_0n[14];
  assign rd_0r0d[15] = rdfint_0n[15];
  assign rd_0r0d[16] = rdfint_0n[16];
  assign rd_0r0d[17] = rdfint_0n[17];
  assign rd_0r0d[18] = rdfint_0n[18];
  assign rd_0r0d[19] = rdfint_0n[19];
  assign rd_0r0d[20] = rdfint_0n[20];
  assign rd_0r0d[21] = rdfint_0n[21];
  assign rd_0r0d[22] = rdfint_0n[22];
  assign rd_0r0d[23] = rdfint_0n[23];
  assign rd_0r0d[24] = rdfint_0n[24];
  assign rd_0r0d[25] = rdfint_0n[25];
  assign rd_0r0d[26] = rdfint_0n[26];
  assign rd_0r0d[27] = rdfint_0n[27];
  assign rd_0r0d[28] = rdfint_0n[28];
  assign rd_0r0d[29] = rdfint_0n[29];
  assign rd_0r0d[30] = rdfint_0n[30];
  assign rd_0r0d[31] = rdfint_0n[31];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign rd_0r1d[10] = rdtint_0n[10];
  assign rd_0r1d[11] = rdtint_0n[11];
  assign rd_0r1d[12] = rdtint_0n[12];
  assign rd_0r1d[13] = rdtint_0n[13];
  assign rd_0r1d[14] = rdtint_0n[14];
  assign rd_0r1d[15] = rdtint_0n[15];
  assign rd_0r1d[16] = rdtint_0n[16];
  assign rd_0r1d[17] = rdtint_0n[17];
  assign rd_0r1d[18] = rdtint_0n[18];
  assign rd_0r1d[19] = rdtint_0n[19];
  assign rd_0r1d[20] = rdtint_0n[20];
  assign rd_0r1d[21] = rdtint_0n[21];
  assign rd_0r1d[22] = rdtint_0n[22];
  assign rd_0r1d[23] = rdtint_0n[23];
  assign rd_0r1d[24] = rdtint_0n[24];
  assign rd_0r1d[25] = rdtint_0n[25];
  assign rd_0r1d[26] = rdtint_0n[26];
  assign rd_0r1d[27] = rdtint_0n[27];
  assign rd_0r1d[28] = rdtint_0n[28];
  assign rd_0r1d[29] = rdtint_0n[29];
  assign rd_0r1d[30] = rdtint_0n[30];
  assign rd_0r1d[31] = rdtint_0n[31];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgfint_0n[32] = wg_0r0d[32];
  assign wgfint_0n[33] = wg_0r0d[33];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign wgtint_0n[32] = wg_0r1d[32];
  assign wgtint_0n[33] = wg_0r1d[33];
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I143 (internal_0n[0], rgrint_0n, rgrint_1n);
  NOR2 I144 (internal_0n[1], rgaint_0n, rgaint_1n);
  AND2 I145 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I146 (rdtint_1n, rgrint_1n, dt_0n[33]);
  AND2 I147 (rdtint_0n[0], rgrint_0n, dt_0n[1]);
  AND2 I148 (rdtint_0n[1], rgrint_0n, dt_0n[2]);
  AND2 I149 (rdtint_0n[2], rgrint_0n, dt_0n[3]);
  AND2 I150 (rdtint_0n[3], rgrint_0n, dt_0n[4]);
  AND2 I151 (rdtint_0n[4], rgrint_0n, dt_0n[5]);
  AND2 I152 (rdtint_0n[5], rgrint_0n, dt_0n[6]);
  AND2 I153 (rdtint_0n[6], rgrint_0n, dt_0n[7]);
  AND2 I154 (rdtint_0n[7], rgrint_0n, dt_0n[8]);
  AND2 I155 (rdtint_0n[8], rgrint_0n, dt_0n[9]);
  AND2 I156 (rdtint_0n[9], rgrint_0n, dt_0n[10]);
  AND2 I157 (rdtint_0n[10], rgrint_0n, dt_0n[11]);
  AND2 I158 (rdtint_0n[11], rgrint_0n, dt_0n[12]);
  AND2 I159 (rdtint_0n[12], rgrint_0n, dt_0n[13]);
  AND2 I160 (rdtint_0n[13], rgrint_0n, dt_0n[14]);
  AND2 I161 (rdtint_0n[14], rgrint_0n, dt_0n[15]);
  AND2 I162 (rdtint_0n[15], rgrint_0n, dt_0n[16]);
  AND2 I163 (rdtint_0n[16], rgrint_0n, dt_0n[17]);
  AND2 I164 (rdtint_0n[17], rgrint_0n, dt_0n[18]);
  AND2 I165 (rdtint_0n[18], rgrint_0n, dt_0n[19]);
  AND2 I166 (rdtint_0n[19], rgrint_0n, dt_0n[20]);
  AND2 I167 (rdtint_0n[20], rgrint_0n, dt_0n[21]);
  AND2 I168 (rdtint_0n[21], rgrint_0n, dt_0n[22]);
  AND2 I169 (rdtint_0n[22], rgrint_0n, dt_0n[23]);
  AND2 I170 (rdtint_0n[23], rgrint_0n, dt_0n[24]);
  AND2 I171 (rdtint_0n[24], rgrint_0n, dt_0n[25]);
  AND2 I172 (rdtint_0n[25], rgrint_0n, dt_0n[26]);
  AND2 I173 (rdtint_0n[26], rgrint_0n, dt_0n[27]);
  AND2 I174 (rdtint_0n[27], rgrint_0n, dt_0n[28]);
  AND2 I175 (rdtint_0n[28], rgrint_0n, dt_0n[29]);
  AND2 I176 (rdtint_0n[29], rgrint_0n, dt_0n[30]);
  AND2 I177 (rdtint_0n[30], rgrint_0n, dt_0n[31]);
  AND2 I178 (rdtint_0n[31], rgrint_0n, dt_0n[32]);
  AND2 I179 (rdfint_1n, rgrint_1n, df_0n[33]);
  AND2 I180 (rdfint_0n[0], rgrint_0n, df_0n[1]);
  AND2 I181 (rdfint_0n[1], rgrint_0n, df_0n[2]);
  AND2 I182 (rdfint_0n[2], rgrint_0n, df_0n[3]);
  AND2 I183 (rdfint_0n[3], rgrint_0n, df_0n[4]);
  AND2 I184 (rdfint_0n[4], rgrint_0n, df_0n[5]);
  AND2 I185 (rdfint_0n[5], rgrint_0n, df_0n[6]);
  AND2 I186 (rdfint_0n[6], rgrint_0n, df_0n[7]);
  AND2 I187 (rdfint_0n[7], rgrint_0n, df_0n[8]);
  AND2 I188 (rdfint_0n[8], rgrint_0n, df_0n[9]);
  AND2 I189 (rdfint_0n[9], rgrint_0n, df_0n[10]);
  AND2 I190 (rdfint_0n[10], rgrint_0n, df_0n[11]);
  AND2 I191 (rdfint_0n[11], rgrint_0n, df_0n[12]);
  AND2 I192 (rdfint_0n[12], rgrint_0n, df_0n[13]);
  AND2 I193 (rdfint_0n[13], rgrint_0n, df_0n[14]);
  AND2 I194 (rdfint_0n[14], rgrint_0n, df_0n[15]);
  AND2 I195 (rdfint_0n[15], rgrint_0n, df_0n[16]);
  AND2 I196 (rdfint_0n[16], rgrint_0n, df_0n[17]);
  AND2 I197 (rdfint_0n[17], rgrint_0n, df_0n[18]);
  AND2 I198 (rdfint_0n[18], rgrint_0n, df_0n[19]);
  AND2 I199 (rdfint_0n[19], rgrint_0n, df_0n[20]);
  AND2 I200 (rdfint_0n[20], rgrint_0n, df_0n[21]);
  AND2 I201 (rdfint_0n[21], rgrint_0n, df_0n[22]);
  AND2 I202 (rdfint_0n[22], rgrint_0n, df_0n[23]);
  AND2 I203 (rdfint_0n[23], rgrint_0n, df_0n[24]);
  AND2 I204 (rdfint_0n[24], rgrint_0n, df_0n[25]);
  AND2 I205 (rdfint_0n[25], rgrint_0n, df_0n[26]);
  AND2 I206 (rdfint_0n[26], rgrint_0n, df_0n[27]);
  AND2 I207 (rdfint_0n[27], rgrint_0n, df_0n[28]);
  AND2 I208 (rdfint_0n[28], rgrint_0n, df_0n[29]);
  AND2 I209 (rdfint_0n[29], rgrint_0n, df_0n[30]);
  AND2 I210 (rdfint_0n[30], rgrint_0n, df_0n[31]);
  AND2 I211 (rdfint_0n[31], rgrint_0n, df_0n[32]);
  C3 I212 (internal_0n[2], wc_0n, wacks_0n[33], wacks_0n[32]);
  C3 I213 (internal_0n[3], wacks_0n[31], wacks_0n[30], wacks_0n[29]);
  C3 I214 (internal_0n[4], wacks_0n[28], wacks_0n[27], wacks_0n[26]);
  C3 I215 (internal_0n[5], wacks_0n[25], wacks_0n[24], wacks_0n[23]);
  C3 I216 (internal_0n[6], wacks_0n[22], wacks_0n[21], wacks_0n[20]);
  C3 I217 (internal_0n[7], wacks_0n[19], wacks_0n[18], wacks_0n[17]);
  C3 I218 (internal_0n[8], wacks_0n[16], wacks_0n[15], wacks_0n[14]);
  C3 I219 (internal_0n[9], wacks_0n[13], wacks_0n[12], wacks_0n[11]);
  C3 I220 (internal_0n[10], wacks_0n[10], wacks_0n[9], wacks_0n[8]);
  C3 I221 (internal_0n[11], wacks_0n[7], wacks_0n[6], wacks_0n[5]);
  C3 I222 (internal_0n[12], wacks_0n[4], wacks_0n[3], wacks_0n[2]);
  C2 I223 (internal_0n[13], wacks_0n[1], wacks_0n[0]);
  C3 I224 (internal_0n[14], internal_0n[2], internal_0n[3], internal_0n[4]);
  C3 I225 (internal_0n[15], internal_0n[5], internal_0n[6], internal_0n[7]);
  C3 I226 (internal_0n[16], internal_0n[8], internal_0n[9], internal_0n[10]);
  C3 I227 (internal_0n[17], internal_0n[11], internal_0n[12], internal_0n[13]);
  C2 I228 (internal_0n[18], internal_0n[14], internal_0n[15]);
  C2 I229 (internal_0n[19], internal_0n[16], internal_0n[17]);
  C2 I230 (wdrint_0n, internal_0n[18], internal_0n[19]);
  assign wen_0n[33] = wc_0n;
  assign wen_0n[32] = wc_0n;
  assign wen_0n[31] = wc_0n;
  assign wen_0n[30] = wc_0n;
  assign wen_0n[29] = wc_0n;
  assign wen_0n[28] = wc_0n;
  assign wen_0n[27] = wc_0n;
  assign wen_0n[26] = wc_0n;
  assign wen_0n[25] = wc_0n;
  assign wen_0n[24] = wc_0n;
  assign wen_0n[23] = wc_0n;
  assign wen_0n[22] = wc_0n;
  assign wen_0n[21] = wc_0n;
  assign wen_0n[20] = wc_0n;
  assign wen_0n[19] = wc_0n;
  assign wen_0n[18] = wc_0n;
  assign wen_0n[17] = wc_0n;
  assign wen_0n[16] = wc_0n;
  assign wen_0n[15] = wc_0n;
  assign wen_0n[14] = wc_0n;
  assign wen_0n[13] = wc_0n;
  assign wen_0n[12] = wc_0n;
  assign wen_0n[11] = wc_0n;
  assign wen_0n[10] = wc_0n;
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[33] = git_0n[33];
  assign wt_0n[32] = git_0n[32];
  assign wt_0n[31] = git_0n[31];
  assign wt_0n[30] = git_0n[30];
  assign wt_0n[29] = git_0n[29];
  assign wt_0n[28] = git_0n[28];
  assign wt_0n[27] = git_0n[27];
  assign wt_0n[26] = git_0n[26];
  assign wt_0n[25] = git_0n[25];
  assign wt_0n[24] = git_0n[24];
  assign wt_0n[23] = git_0n[23];
  assign wt_0n[22] = git_0n[22];
  assign wt_0n[21] = git_0n[21];
  assign wt_0n[20] = git_0n[20];
  assign wt_0n[19] = git_0n[19];
  assign wt_0n[18] = git_0n[18];
  assign wt_0n[17] = git_0n[17];
  assign wt_0n[16] = git_0n[16];
  assign wt_0n[15] = git_0n[15];
  assign wt_0n[14] = git_0n[14];
  assign wt_0n[13] = git_0n[13];
  assign wt_0n[12] = git_0n[12];
  assign wt_0n[11] = git_0n[11];
  assign wt_0n[10] = git_0n[10];
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[33] = gif_0n[33];
  assign wf_0n[32] = gif_0n[32];
  assign wf_0n[31] = gif_0n[31];
  assign wf_0n[30] = gif_0n[30];
  assign wf_0n[29] = gif_0n[29];
  assign wf_0n[28] = gif_0n[28];
  assign wf_0n[27] = gif_0n[27];
  assign wf_0n[26] = gif_0n[26];
  assign wf_0n[25] = gif_0n[25];
  assign wf_0n[24] = gif_0n[24];
  assign wf_0n[23] = gif_0n[23];
  assign wf_0n[22] = gif_0n[22];
  assign wf_0n[21] = gif_0n[21];
  assign wf_0n[20] = gif_0n[20];
  assign wf_0n[19] = gif_0n[19];
  assign wf_0n[18] = gif_0n[18];
  assign wf_0n[17] = gif_0n[17];
  assign wf_0n[16] = gif_0n[16];
  assign wf_0n[15] = gif_0n[15];
  assign wf_0n[14] = gif_0n[14];
  assign wf_0n[13] = gif_0n[13];
  assign wf_0n[12] = gif_0n[12];
  assign wf_0n[11] = gif_0n[11];
  assign wf_0n[10] = gif_0n[10];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I333 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I335 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I336 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I337 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I338 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I339 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I340 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I341 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I342 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I343 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I344 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I345 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I346 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I347 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I348 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I349 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I350 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I351 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I352 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I353 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I354 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I355 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I356 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I357 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I358 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I359 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I360 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I361 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I362 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I363 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I364 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I365 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I366 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I367 (git_0n[32], wgtint_0n[32], ig_0n);
  AND2 I368 (git_0n[33], wgtint_0n[33], ig_0n);
  AND2 I369 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I370 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I371 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I372 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I373 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I374 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I375 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I376 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I377 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I378 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I379 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I380 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I381 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I382 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I383 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I384 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I385 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I386 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I387 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I388 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I389 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I390 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I391 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I392 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I393 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I394 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I395 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I396 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I397 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I398 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I399 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I400 (gif_0n[31], wgfint_0n[31], ig_0n);
  AND2 I401 (gif_0n[32], wgfint_0n[32], ig_0n);
  AND2 I402 (gif_0n[33], wgfint_0n[33], ig_0n);
  C3 I403 (internal_0n[20], complete1395_0n[0], complete1395_0n[1], complete1395_0n[2]);
  C3 I404 (internal_0n[21], complete1395_0n[3], complete1395_0n[4], complete1395_0n[5]);
  C3 I405 (internal_0n[22], complete1395_0n[6], complete1395_0n[7], complete1395_0n[8]);
  C3 I406 (internal_0n[23], complete1395_0n[9], complete1395_0n[10], complete1395_0n[11]);
  C3 I407 (internal_0n[24], complete1395_0n[12], complete1395_0n[13], complete1395_0n[14]);
  C3 I408 (internal_0n[25], complete1395_0n[15], complete1395_0n[16], complete1395_0n[17]);
  C3 I409 (internal_0n[26], complete1395_0n[18], complete1395_0n[19], complete1395_0n[20]);
  C3 I410 (internal_0n[27], complete1395_0n[21], complete1395_0n[22], complete1395_0n[23]);
  C3 I411 (internal_0n[28], complete1395_0n[24], complete1395_0n[25], complete1395_0n[26]);
  C3 I412 (internal_0n[29], complete1395_0n[27], complete1395_0n[28], complete1395_0n[29]);
  C2 I413 (internal_0n[30], complete1395_0n[30], complete1395_0n[31]);
  C2 I414 (internal_0n[31], complete1395_0n[32], complete1395_0n[33]);
  C3 I415 (internal_0n[32], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I416 (internal_0n[33], internal_0n[23], internal_0n[24], internal_0n[25]);
  C3 I417 (internal_0n[34], internal_0n[26], internal_0n[27], internal_0n[28]);
  C3 I418 (internal_0n[35], internal_0n[29], internal_0n[30], internal_0n[31]);
  C2 I419 (internal_0n[36], internal_0n[32], internal_0n[33]);
  C2 I420 (internal_0n[37], internal_0n[34], internal_0n[35]);
  C2 I421 (wc_0n, internal_0n[36], internal_0n[37]);
  OR2 I422 (complete1395_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I423 (complete1395_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I424 (complete1395_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I425 (complete1395_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I426 (complete1395_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I427 (complete1395_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I428 (complete1395_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I429 (complete1395_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I430 (complete1395_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I431 (complete1395_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I432 (complete1395_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I433 (complete1395_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I434 (complete1395_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I435 (complete1395_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I436 (complete1395_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I437 (complete1395_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I438 (complete1395_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I439 (complete1395_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I440 (complete1395_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I441 (complete1395_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I442 (complete1395_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I443 (complete1395_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I444 (complete1395_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I445 (complete1395_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I446 (complete1395_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I447 (complete1395_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I448 (complete1395_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I449 (complete1395_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I450 (complete1395_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I451 (complete1395_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I452 (complete1395_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I453 (complete1395_0n[31], wgfint_0n[31], wgtint_0n[31]);
  OR2 I454 (complete1395_0n[32], wgfint_0n[32], wgtint_0n[32]);
  OR2 I455 (complete1395_0n[33], wgfint_0n[33], wgtint_0n[33]);
  AO22 I456 (wacks_0n[33], gf1393_0n[33], df_0n[33], gt1394_0n[33], dt_0n[33]);
  NOR2 I457 (dt_0n[33], df_0n[33], gf1393_0n[33]);
  NOR3 I458 (df_0n[33], dt_0n[33], gt1394_0n[33], init_0n);
  AND2 I459 (gt1394_0n[33], wt_0n[33], wen_0n[33]);
  AND2 I460 (gf1393_0n[33], wf_0n[33], wen_0n[33]);
  AO22 I461 (wacks_0n[32], gf1393_0n[32], df_0n[32], gt1394_0n[32], dt_0n[32]);
  NOR2 I462 (dt_0n[32], df_0n[32], gf1393_0n[32]);
  NOR3 I463 (df_0n[32], dt_0n[32], gt1394_0n[32], init_0n);
  AND2 I464 (gt1394_0n[32], wt_0n[32], wen_0n[32]);
  AND2 I465 (gf1393_0n[32], wf_0n[32], wen_0n[32]);
  AO22 I466 (wacks_0n[31], gf1393_0n[31], df_0n[31], gt1394_0n[31], dt_0n[31]);
  NOR2 I467 (dt_0n[31], df_0n[31], gf1393_0n[31]);
  NOR3 I468 (df_0n[31], dt_0n[31], gt1394_0n[31], init_0n);
  AND2 I469 (gt1394_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I470 (gf1393_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I471 (wacks_0n[30], gf1393_0n[30], df_0n[30], gt1394_0n[30], dt_0n[30]);
  NOR2 I472 (dt_0n[30], df_0n[30], gf1393_0n[30]);
  NOR3 I473 (df_0n[30], dt_0n[30], gt1394_0n[30], init_0n);
  AND2 I474 (gt1394_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I475 (gf1393_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I476 (wacks_0n[29], gf1393_0n[29], df_0n[29], gt1394_0n[29], dt_0n[29]);
  NOR2 I477 (dt_0n[29], df_0n[29], gf1393_0n[29]);
  NOR3 I478 (df_0n[29], dt_0n[29], gt1394_0n[29], init_0n);
  AND2 I479 (gt1394_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I480 (gf1393_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I481 (wacks_0n[28], gf1393_0n[28], df_0n[28], gt1394_0n[28], dt_0n[28]);
  NOR2 I482 (dt_0n[28], df_0n[28], gf1393_0n[28]);
  NOR3 I483 (df_0n[28], dt_0n[28], gt1394_0n[28], init_0n);
  AND2 I484 (gt1394_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I485 (gf1393_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I486 (wacks_0n[27], gf1393_0n[27], df_0n[27], gt1394_0n[27], dt_0n[27]);
  NOR2 I487 (dt_0n[27], df_0n[27], gf1393_0n[27]);
  NOR3 I488 (df_0n[27], dt_0n[27], gt1394_0n[27], init_0n);
  AND2 I489 (gt1394_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I490 (gf1393_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I491 (wacks_0n[26], gf1393_0n[26], df_0n[26], gt1394_0n[26], dt_0n[26]);
  NOR2 I492 (dt_0n[26], df_0n[26], gf1393_0n[26]);
  NOR3 I493 (df_0n[26], dt_0n[26], gt1394_0n[26], init_0n);
  AND2 I494 (gt1394_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I495 (gf1393_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I496 (wacks_0n[25], gf1393_0n[25], df_0n[25], gt1394_0n[25], dt_0n[25]);
  NOR2 I497 (dt_0n[25], df_0n[25], gf1393_0n[25]);
  NOR3 I498 (df_0n[25], dt_0n[25], gt1394_0n[25], init_0n);
  AND2 I499 (gt1394_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I500 (gf1393_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I501 (wacks_0n[24], gf1393_0n[24], df_0n[24], gt1394_0n[24], dt_0n[24]);
  NOR2 I502 (dt_0n[24], df_0n[24], gf1393_0n[24]);
  NOR3 I503 (df_0n[24], dt_0n[24], gt1394_0n[24], init_0n);
  AND2 I504 (gt1394_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I505 (gf1393_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I506 (wacks_0n[23], gf1393_0n[23], df_0n[23], gt1394_0n[23], dt_0n[23]);
  NOR2 I507 (dt_0n[23], df_0n[23], gf1393_0n[23]);
  NOR3 I508 (df_0n[23], dt_0n[23], gt1394_0n[23], init_0n);
  AND2 I509 (gt1394_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I510 (gf1393_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I511 (wacks_0n[22], gf1393_0n[22], df_0n[22], gt1394_0n[22], dt_0n[22]);
  NOR2 I512 (dt_0n[22], df_0n[22], gf1393_0n[22]);
  NOR3 I513 (df_0n[22], dt_0n[22], gt1394_0n[22], init_0n);
  AND2 I514 (gt1394_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I515 (gf1393_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I516 (wacks_0n[21], gf1393_0n[21], df_0n[21], gt1394_0n[21], dt_0n[21]);
  NOR2 I517 (dt_0n[21], df_0n[21], gf1393_0n[21]);
  NOR3 I518 (df_0n[21], dt_0n[21], gt1394_0n[21], init_0n);
  AND2 I519 (gt1394_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I520 (gf1393_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I521 (wacks_0n[20], gf1393_0n[20], df_0n[20], gt1394_0n[20], dt_0n[20]);
  NOR2 I522 (dt_0n[20], df_0n[20], gf1393_0n[20]);
  NOR3 I523 (df_0n[20], dt_0n[20], gt1394_0n[20], init_0n);
  AND2 I524 (gt1394_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I525 (gf1393_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I526 (wacks_0n[19], gf1393_0n[19], df_0n[19], gt1394_0n[19], dt_0n[19]);
  NOR2 I527 (dt_0n[19], df_0n[19], gf1393_0n[19]);
  NOR3 I528 (df_0n[19], dt_0n[19], gt1394_0n[19], init_0n);
  AND2 I529 (gt1394_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I530 (gf1393_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I531 (wacks_0n[18], gf1393_0n[18], df_0n[18], gt1394_0n[18], dt_0n[18]);
  NOR2 I532 (dt_0n[18], df_0n[18], gf1393_0n[18]);
  NOR3 I533 (df_0n[18], dt_0n[18], gt1394_0n[18], init_0n);
  AND2 I534 (gt1394_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I535 (gf1393_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I536 (wacks_0n[17], gf1393_0n[17], df_0n[17], gt1394_0n[17], dt_0n[17]);
  NOR2 I537 (dt_0n[17], df_0n[17], gf1393_0n[17]);
  NOR3 I538 (df_0n[17], dt_0n[17], gt1394_0n[17], init_0n);
  AND2 I539 (gt1394_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I540 (gf1393_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I541 (wacks_0n[16], gf1393_0n[16], df_0n[16], gt1394_0n[16], dt_0n[16]);
  NOR2 I542 (dt_0n[16], df_0n[16], gf1393_0n[16]);
  NOR3 I543 (df_0n[16], dt_0n[16], gt1394_0n[16], init_0n);
  AND2 I544 (gt1394_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I545 (gf1393_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I546 (wacks_0n[15], gf1393_0n[15], df_0n[15], gt1394_0n[15], dt_0n[15]);
  NOR2 I547 (dt_0n[15], df_0n[15], gf1393_0n[15]);
  NOR3 I548 (df_0n[15], dt_0n[15], gt1394_0n[15], init_0n);
  AND2 I549 (gt1394_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I550 (gf1393_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I551 (wacks_0n[14], gf1393_0n[14], df_0n[14], gt1394_0n[14], dt_0n[14]);
  NOR2 I552 (dt_0n[14], df_0n[14], gf1393_0n[14]);
  NOR3 I553 (df_0n[14], dt_0n[14], gt1394_0n[14], init_0n);
  AND2 I554 (gt1394_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I555 (gf1393_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I556 (wacks_0n[13], gf1393_0n[13], df_0n[13], gt1394_0n[13], dt_0n[13]);
  NOR2 I557 (dt_0n[13], df_0n[13], gf1393_0n[13]);
  NOR3 I558 (df_0n[13], dt_0n[13], gt1394_0n[13], init_0n);
  AND2 I559 (gt1394_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I560 (gf1393_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I561 (wacks_0n[12], gf1393_0n[12], df_0n[12], gt1394_0n[12], dt_0n[12]);
  NOR2 I562 (dt_0n[12], df_0n[12], gf1393_0n[12]);
  NOR3 I563 (df_0n[12], dt_0n[12], gt1394_0n[12], init_0n);
  AND2 I564 (gt1394_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I565 (gf1393_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I566 (wacks_0n[11], gf1393_0n[11], df_0n[11], gt1394_0n[11], dt_0n[11]);
  NOR2 I567 (dt_0n[11], df_0n[11], gf1393_0n[11]);
  NOR3 I568 (df_0n[11], dt_0n[11], gt1394_0n[11], init_0n);
  AND2 I569 (gt1394_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I570 (gf1393_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I571 (wacks_0n[10], gf1393_0n[10], df_0n[10], gt1394_0n[10], dt_0n[10]);
  NOR2 I572 (dt_0n[10], df_0n[10], gf1393_0n[10]);
  NOR3 I573 (df_0n[10], dt_0n[10], gt1394_0n[10], init_0n);
  AND2 I574 (gt1394_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I575 (gf1393_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I576 (wacks_0n[9], gf1393_0n[9], df_0n[9], gt1394_0n[9], dt_0n[9]);
  NOR2 I577 (dt_0n[9], df_0n[9], gf1393_0n[9]);
  NOR3 I578 (df_0n[9], dt_0n[9], gt1394_0n[9], init_0n);
  AND2 I579 (gt1394_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I580 (gf1393_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I581 (wacks_0n[8], gf1393_0n[8], df_0n[8], gt1394_0n[8], dt_0n[8]);
  NOR2 I582 (dt_0n[8], df_0n[8], gf1393_0n[8]);
  NOR3 I583 (df_0n[8], dt_0n[8], gt1394_0n[8], init_0n);
  AND2 I584 (gt1394_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I585 (gf1393_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I586 (wacks_0n[7], gf1393_0n[7], df_0n[7], gt1394_0n[7], dt_0n[7]);
  NOR2 I587 (dt_0n[7], df_0n[7], gf1393_0n[7]);
  NOR3 I588 (df_0n[7], dt_0n[7], gt1394_0n[7], init_0n);
  AND2 I589 (gt1394_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I590 (gf1393_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I591 (wacks_0n[6], gf1393_0n[6], df_0n[6], gt1394_0n[6], dt_0n[6]);
  NOR2 I592 (dt_0n[6], df_0n[6], gf1393_0n[6]);
  NOR3 I593 (df_0n[6], dt_0n[6], gt1394_0n[6], init_0n);
  AND2 I594 (gt1394_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I595 (gf1393_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I596 (wacks_0n[5], gf1393_0n[5], df_0n[5], gt1394_0n[5], dt_0n[5]);
  NOR2 I597 (dt_0n[5], df_0n[5], gf1393_0n[5]);
  NOR3 I598 (df_0n[5], dt_0n[5], gt1394_0n[5], init_0n);
  AND2 I599 (gt1394_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I600 (gf1393_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I601 (wacks_0n[4], gf1393_0n[4], df_0n[4], gt1394_0n[4], dt_0n[4]);
  NOR2 I602 (dt_0n[4], df_0n[4], gf1393_0n[4]);
  NOR3 I603 (df_0n[4], dt_0n[4], gt1394_0n[4], init_0n);
  AND2 I604 (gt1394_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I605 (gf1393_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I606 (wacks_0n[3], gf1393_0n[3], df_0n[3], gt1394_0n[3], dt_0n[3]);
  NOR2 I607 (dt_0n[3], df_0n[3], gf1393_0n[3]);
  NOR3 I608 (df_0n[3], dt_0n[3], gt1394_0n[3], init_0n);
  AND2 I609 (gt1394_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I610 (gf1393_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I611 (wacks_0n[2], gf1393_0n[2], df_0n[2], gt1394_0n[2], dt_0n[2]);
  NOR2 I612 (dt_0n[2], df_0n[2], gf1393_0n[2]);
  NOR3 I613 (df_0n[2], dt_0n[2], gt1394_0n[2], init_0n);
  AND2 I614 (gt1394_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I615 (gf1393_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I616 (wacks_0n[1], gf1393_0n[1], df_0n[1], gt1394_0n[1], dt_0n[1]);
  NOR2 I617 (dt_0n[1], df_0n[1], gf1393_0n[1]);
  NOR3 I618 (df_0n[1], dt_0n[1], gt1394_0n[1], init_0n);
  AND2 I619 (gt1394_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I620 (gf1393_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I621 (wacks_0n[0], gf1393_0n[0], df_0n[0], gt1394_0n[0], dt_0n[0]);
  NOR2 I622 (dt_0n[0], df_0n[0], gf1393_0n[0]);
  NOR3 I623 (df_0n[0], dt_0n[0], gt1394_0n[0], init_0n);
  AND2 I624 (gt1394_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I625 (gf1393_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I626 (init_0n, initialise);
endmodule

module BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m86m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  initialise
);
  input [34:0] wg_0r0d;
  input [34:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [30:0] rd_0r0d;
  output [30:0] rd_0r1d;
  input rd_0a;
  output [34:0] rd_1r0d;
  output [34:0] rd_1r1d;
  input rd_1a;
  input initialise;
  wire [37:0] internal_0n;
  wire [34:0] wf_0n;
  wire [34:0] wt_0n;
  wire [34:0] df_0n;
  wire [34:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire wc_0n;
  wire [34:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [34:0] wgfint_0n;
  wire [34:0] wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire [30:0] rdfint_0n;
  wire [34:0] rdfint_1n;
  wire [30:0] rdtint_0n;
  wire [34:0] rdtint_1n;
  wire [34:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [34:0] gif_0n;
  wire [34:0] git_0n;
  wire [34:0] complete1410_0n;
  wire [34:0] gt1409_0n;
  wire [34:0] gf1408_0n;
  assign rgaint_1n = rd_1a;
  assign rd_1r0d[0] = rdfint_1n[0];
  assign rd_1r0d[1] = rdfint_1n[1];
  assign rd_1r0d[2] = rdfint_1n[2];
  assign rd_1r0d[3] = rdfint_1n[3];
  assign rd_1r0d[4] = rdfint_1n[4];
  assign rd_1r0d[5] = rdfint_1n[5];
  assign rd_1r0d[6] = rdfint_1n[6];
  assign rd_1r0d[7] = rdfint_1n[7];
  assign rd_1r0d[8] = rdfint_1n[8];
  assign rd_1r0d[9] = rdfint_1n[9];
  assign rd_1r0d[10] = rdfint_1n[10];
  assign rd_1r0d[11] = rdfint_1n[11];
  assign rd_1r0d[12] = rdfint_1n[12];
  assign rd_1r0d[13] = rdfint_1n[13];
  assign rd_1r0d[14] = rdfint_1n[14];
  assign rd_1r0d[15] = rdfint_1n[15];
  assign rd_1r0d[16] = rdfint_1n[16];
  assign rd_1r0d[17] = rdfint_1n[17];
  assign rd_1r0d[18] = rdfint_1n[18];
  assign rd_1r0d[19] = rdfint_1n[19];
  assign rd_1r0d[20] = rdfint_1n[20];
  assign rd_1r0d[21] = rdfint_1n[21];
  assign rd_1r0d[22] = rdfint_1n[22];
  assign rd_1r0d[23] = rdfint_1n[23];
  assign rd_1r0d[24] = rdfint_1n[24];
  assign rd_1r0d[25] = rdfint_1n[25];
  assign rd_1r0d[26] = rdfint_1n[26];
  assign rd_1r0d[27] = rdfint_1n[27];
  assign rd_1r0d[28] = rdfint_1n[28];
  assign rd_1r0d[29] = rdfint_1n[29];
  assign rd_1r0d[30] = rdfint_1n[30];
  assign rd_1r0d[31] = rdfint_1n[31];
  assign rd_1r0d[32] = rdfint_1n[32];
  assign rd_1r0d[33] = rdfint_1n[33];
  assign rd_1r0d[34] = rdfint_1n[34];
  assign rd_1r1d[0] = rdtint_1n[0];
  assign rd_1r1d[1] = rdtint_1n[1];
  assign rd_1r1d[2] = rdtint_1n[2];
  assign rd_1r1d[3] = rdtint_1n[3];
  assign rd_1r1d[4] = rdtint_1n[4];
  assign rd_1r1d[5] = rdtint_1n[5];
  assign rd_1r1d[6] = rdtint_1n[6];
  assign rd_1r1d[7] = rdtint_1n[7];
  assign rd_1r1d[8] = rdtint_1n[8];
  assign rd_1r1d[9] = rdtint_1n[9];
  assign rd_1r1d[10] = rdtint_1n[10];
  assign rd_1r1d[11] = rdtint_1n[11];
  assign rd_1r1d[12] = rdtint_1n[12];
  assign rd_1r1d[13] = rdtint_1n[13];
  assign rd_1r1d[14] = rdtint_1n[14];
  assign rd_1r1d[15] = rdtint_1n[15];
  assign rd_1r1d[16] = rdtint_1n[16];
  assign rd_1r1d[17] = rdtint_1n[17];
  assign rd_1r1d[18] = rdtint_1n[18];
  assign rd_1r1d[19] = rdtint_1n[19];
  assign rd_1r1d[20] = rdtint_1n[20];
  assign rd_1r1d[21] = rdtint_1n[21];
  assign rd_1r1d[22] = rdtint_1n[22];
  assign rd_1r1d[23] = rdtint_1n[23];
  assign rd_1r1d[24] = rdtint_1n[24];
  assign rd_1r1d[25] = rdtint_1n[25];
  assign rd_1r1d[26] = rdtint_1n[26];
  assign rd_1r1d[27] = rdtint_1n[27];
  assign rd_1r1d[28] = rdtint_1n[28];
  assign rd_1r1d[29] = rdtint_1n[29];
  assign rd_1r1d[30] = rdtint_1n[30];
  assign rd_1r1d[31] = rdtint_1n[31];
  assign rd_1r1d[32] = rdtint_1n[32];
  assign rd_1r1d[33] = rdtint_1n[33];
  assign rd_1r1d[34] = rdtint_1n[34];
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r0d[10] = rdfint_0n[10];
  assign rd_0r0d[11] = rdfint_0n[11];
  assign rd_0r0d[12] = rdfint_0n[12];
  assign rd_0r0d[13] = rdfint_0n[13];
  assign rd_0r0d[14] = rdfint_0n[14];
  assign rd_0r0d[15] = rdfint_0n[15];
  assign rd_0r0d[16] = rdfint_0n[16];
  assign rd_0r0d[17] = rdfint_0n[17];
  assign rd_0r0d[18] = rdfint_0n[18];
  assign rd_0r0d[19] = rdfint_0n[19];
  assign rd_0r0d[20] = rdfint_0n[20];
  assign rd_0r0d[21] = rdfint_0n[21];
  assign rd_0r0d[22] = rdfint_0n[22];
  assign rd_0r0d[23] = rdfint_0n[23];
  assign rd_0r0d[24] = rdfint_0n[24];
  assign rd_0r0d[25] = rdfint_0n[25];
  assign rd_0r0d[26] = rdfint_0n[26];
  assign rd_0r0d[27] = rdfint_0n[27];
  assign rd_0r0d[28] = rdfint_0n[28];
  assign rd_0r0d[29] = rdfint_0n[29];
  assign rd_0r0d[30] = rdfint_0n[30];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign rd_0r1d[10] = rdtint_0n[10];
  assign rd_0r1d[11] = rdtint_0n[11];
  assign rd_0r1d[12] = rdtint_0n[12];
  assign rd_0r1d[13] = rdtint_0n[13];
  assign rd_0r1d[14] = rdtint_0n[14];
  assign rd_0r1d[15] = rdtint_0n[15];
  assign rd_0r1d[16] = rdtint_0n[16];
  assign rd_0r1d[17] = rdtint_0n[17];
  assign rd_0r1d[18] = rdtint_0n[18];
  assign rd_0r1d[19] = rdtint_0n[19];
  assign rd_0r1d[20] = rdtint_0n[20];
  assign rd_0r1d[21] = rdtint_0n[21];
  assign rd_0r1d[22] = rdtint_0n[22];
  assign rd_0r1d[23] = rdtint_0n[23];
  assign rd_0r1d[24] = rdtint_0n[24];
  assign rd_0r1d[25] = rdtint_0n[25];
  assign rd_0r1d[26] = rdtint_0n[26];
  assign rd_0r1d[27] = rdtint_0n[27];
  assign rd_0r1d[28] = rdtint_0n[28];
  assign rd_0r1d[29] = rdtint_0n[29];
  assign rd_0r1d[30] = rdtint_0n[30];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgfint_0n[32] = wg_0r0d[32];
  assign wgfint_0n[33] = wg_0r0d[33];
  assign wgfint_0n[34] = wg_0r0d[34];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign wgtint_0n[32] = wg_0r1d[32];
  assign wgtint_0n[33] = wg_0r1d[33];
  assign wgtint_0n[34] = wg_0r1d[34];
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I211 (internal_0n[0], rgrint_0n, rgrint_1n);
  NOR2 I212 (internal_0n[1], rgaint_0n, rgaint_1n);
  AND2 I213 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I214 (rdtint_1n[0], rgrint_1n, dt_0n[0]);
  AND2 I215 (rdtint_1n[1], rgrint_1n, dt_0n[1]);
  AND2 I216 (rdtint_1n[2], rgrint_1n, dt_0n[2]);
  AND2 I217 (rdtint_1n[3], rgrint_1n, dt_0n[3]);
  AND2 I218 (rdtint_1n[4], rgrint_1n, dt_0n[4]);
  AND2 I219 (rdtint_1n[5], rgrint_1n, dt_0n[5]);
  AND2 I220 (rdtint_1n[6], rgrint_1n, dt_0n[6]);
  AND2 I221 (rdtint_1n[7], rgrint_1n, dt_0n[7]);
  AND2 I222 (rdtint_1n[8], rgrint_1n, dt_0n[8]);
  AND2 I223 (rdtint_1n[9], rgrint_1n, dt_0n[9]);
  AND2 I224 (rdtint_1n[10], rgrint_1n, dt_0n[10]);
  AND2 I225 (rdtint_1n[11], rgrint_1n, dt_0n[11]);
  AND2 I226 (rdtint_1n[12], rgrint_1n, dt_0n[12]);
  AND2 I227 (rdtint_1n[13], rgrint_1n, dt_0n[13]);
  AND2 I228 (rdtint_1n[14], rgrint_1n, dt_0n[14]);
  AND2 I229 (rdtint_1n[15], rgrint_1n, dt_0n[15]);
  AND2 I230 (rdtint_1n[16], rgrint_1n, dt_0n[16]);
  AND2 I231 (rdtint_1n[17], rgrint_1n, dt_0n[17]);
  AND2 I232 (rdtint_1n[18], rgrint_1n, dt_0n[18]);
  AND2 I233 (rdtint_1n[19], rgrint_1n, dt_0n[19]);
  AND2 I234 (rdtint_1n[20], rgrint_1n, dt_0n[20]);
  AND2 I235 (rdtint_1n[21], rgrint_1n, dt_0n[21]);
  AND2 I236 (rdtint_1n[22], rgrint_1n, dt_0n[22]);
  AND2 I237 (rdtint_1n[23], rgrint_1n, dt_0n[23]);
  AND2 I238 (rdtint_1n[24], rgrint_1n, dt_0n[24]);
  AND2 I239 (rdtint_1n[25], rgrint_1n, dt_0n[25]);
  AND2 I240 (rdtint_1n[26], rgrint_1n, dt_0n[26]);
  AND2 I241 (rdtint_1n[27], rgrint_1n, dt_0n[27]);
  AND2 I242 (rdtint_1n[28], rgrint_1n, dt_0n[28]);
  AND2 I243 (rdtint_1n[29], rgrint_1n, dt_0n[29]);
  AND2 I244 (rdtint_1n[30], rgrint_1n, dt_0n[30]);
  AND2 I245 (rdtint_1n[31], rgrint_1n, dt_0n[31]);
  AND2 I246 (rdtint_1n[32], rgrint_1n, dt_0n[32]);
  AND2 I247 (rdtint_1n[33], rgrint_1n, dt_0n[33]);
  AND2 I248 (rdtint_1n[34], rgrint_1n, dt_0n[34]);
  AND2 I249 (rdtint_0n[0], rgrint_0n, dt_0n[0]);
  AND2 I250 (rdtint_0n[1], rgrint_0n, dt_0n[1]);
  AND2 I251 (rdtint_0n[2], rgrint_0n, dt_0n[2]);
  AND2 I252 (rdtint_0n[3], rgrint_0n, dt_0n[3]);
  AND2 I253 (rdtint_0n[4], rgrint_0n, dt_0n[4]);
  AND2 I254 (rdtint_0n[5], rgrint_0n, dt_0n[5]);
  AND2 I255 (rdtint_0n[6], rgrint_0n, dt_0n[6]);
  AND2 I256 (rdtint_0n[7], rgrint_0n, dt_0n[7]);
  AND2 I257 (rdtint_0n[8], rgrint_0n, dt_0n[8]);
  AND2 I258 (rdtint_0n[9], rgrint_0n, dt_0n[9]);
  AND2 I259 (rdtint_0n[10], rgrint_0n, dt_0n[10]);
  AND2 I260 (rdtint_0n[11], rgrint_0n, dt_0n[11]);
  AND2 I261 (rdtint_0n[12], rgrint_0n, dt_0n[12]);
  AND2 I262 (rdtint_0n[13], rgrint_0n, dt_0n[13]);
  AND2 I263 (rdtint_0n[14], rgrint_0n, dt_0n[14]);
  AND2 I264 (rdtint_0n[15], rgrint_0n, dt_0n[15]);
  AND2 I265 (rdtint_0n[16], rgrint_0n, dt_0n[16]);
  AND2 I266 (rdtint_0n[17], rgrint_0n, dt_0n[17]);
  AND2 I267 (rdtint_0n[18], rgrint_0n, dt_0n[18]);
  AND2 I268 (rdtint_0n[19], rgrint_0n, dt_0n[19]);
  AND2 I269 (rdtint_0n[20], rgrint_0n, dt_0n[20]);
  AND2 I270 (rdtint_0n[21], rgrint_0n, dt_0n[21]);
  AND2 I271 (rdtint_0n[22], rgrint_0n, dt_0n[22]);
  AND2 I272 (rdtint_0n[23], rgrint_0n, dt_0n[23]);
  AND2 I273 (rdtint_0n[24], rgrint_0n, dt_0n[24]);
  AND2 I274 (rdtint_0n[25], rgrint_0n, dt_0n[25]);
  AND2 I275 (rdtint_0n[26], rgrint_0n, dt_0n[26]);
  AND2 I276 (rdtint_0n[27], rgrint_0n, dt_0n[27]);
  AND2 I277 (rdtint_0n[28], rgrint_0n, dt_0n[28]);
  AND2 I278 (rdtint_0n[29], rgrint_0n, dt_0n[29]);
  AND2 I279 (rdtint_0n[30], rgrint_0n, dt_0n[30]);
  AND2 I280 (rdfint_1n[0], rgrint_1n, df_0n[0]);
  AND2 I281 (rdfint_1n[1], rgrint_1n, df_0n[1]);
  AND2 I282 (rdfint_1n[2], rgrint_1n, df_0n[2]);
  AND2 I283 (rdfint_1n[3], rgrint_1n, df_0n[3]);
  AND2 I284 (rdfint_1n[4], rgrint_1n, df_0n[4]);
  AND2 I285 (rdfint_1n[5], rgrint_1n, df_0n[5]);
  AND2 I286 (rdfint_1n[6], rgrint_1n, df_0n[6]);
  AND2 I287 (rdfint_1n[7], rgrint_1n, df_0n[7]);
  AND2 I288 (rdfint_1n[8], rgrint_1n, df_0n[8]);
  AND2 I289 (rdfint_1n[9], rgrint_1n, df_0n[9]);
  AND2 I290 (rdfint_1n[10], rgrint_1n, df_0n[10]);
  AND2 I291 (rdfint_1n[11], rgrint_1n, df_0n[11]);
  AND2 I292 (rdfint_1n[12], rgrint_1n, df_0n[12]);
  AND2 I293 (rdfint_1n[13], rgrint_1n, df_0n[13]);
  AND2 I294 (rdfint_1n[14], rgrint_1n, df_0n[14]);
  AND2 I295 (rdfint_1n[15], rgrint_1n, df_0n[15]);
  AND2 I296 (rdfint_1n[16], rgrint_1n, df_0n[16]);
  AND2 I297 (rdfint_1n[17], rgrint_1n, df_0n[17]);
  AND2 I298 (rdfint_1n[18], rgrint_1n, df_0n[18]);
  AND2 I299 (rdfint_1n[19], rgrint_1n, df_0n[19]);
  AND2 I300 (rdfint_1n[20], rgrint_1n, df_0n[20]);
  AND2 I301 (rdfint_1n[21], rgrint_1n, df_0n[21]);
  AND2 I302 (rdfint_1n[22], rgrint_1n, df_0n[22]);
  AND2 I303 (rdfint_1n[23], rgrint_1n, df_0n[23]);
  AND2 I304 (rdfint_1n[24], rgrint_1n, df_0n[24]);
  AND2 I305 (rdfint_1n[25], rgrint_1n, df_0n[25]);
  AND2 I306 (rdfint_1n[26], rgrint_1n, df_0n[26]);
  AND2 I307 (rdfint_1n[27], rgrint_1n, df_0n[27]);
  AND2 I308 (rdfint_1n[28], rgrint_1n, df_0n[28]);
  AND2 I309 (rdfint_1n[29], rgrint_1n, df_0n[29]);
  AND2 I310 (rdfint_1n[30], rgrint_1n, df_0n[30]);
  AND2 I311 (rdfint_1n[31], rgrint_1n, df_0n[31]);
  AND2 I312 (rdfint_1n[32], rgrint_1n, df_0n[32]);
  AND2 I313 (rdfint_1n[33], rgrint_1n, df_0n[33]);
  AND2 I314 (rdfint_1n[34], rgrint_1n, df_0n[34]);
  AND2 I315 (rdfint_0n[0], rgrint_0n, df_0n[0]);
  AND2 I316 (rdfint_0n[1], rgrint_0n, df_0n[1]);
  AND2 I317 (rdfint_0n[2], rgrint_0n, df_0n[2]);
  AND2 I318 (rdfint_0n[3], rgrint_0n, df_0n[3]);
  AND2 I319 (rdfint_0n[4], rgrint_0n, df_0n[4]);
  AND2 I320 (rdfint_0n[5], rgrint_0n, df_0n[5]);
  AND2 I321 (rdfint_0n[6], rgrint_0n, df_0n[6]);
  AND2 I322 (rdfint_0n[7], rgrint_0n, df_0n[7]);
  AND2 I323 (rdfint_0n[8], rgrint_0n, df_0n[8]);
  AND2 I324 (rdfint_0n[9], rgrint_0n, df_0n[9]);
  AND2 I325 (rdfint_0n[10], rgrint_0n, df_0n[10]);
  AND2 I326 (rdfint_0n[11], rgrint_0n, df_0n[11]);
  AND2 I327 (rdfint_0n[12], rgrint_0n, df_0n[12]);
  AND2 I328 (rdfint_0n[13], rgrint_0n, df_0n[13]);
  AND2 I329 (rdfint_0n[14], rgrint_0n, df_0n[14]);
  AND2 I330 (rdfint_0n[15], rgrint_0n, df_0n[15]);
  AND2 I331 (rdfint_0n[16], rgrint_0n, df_0n[16]);
  AND2 I332 (rdfint_0n[17], rgrint_0n, df_0n[17]);
  AND2 I333 (rdfint_0n[18], rgrint_0n, df_0n[18]);
  AND2 I334 (rdfint_0n[19], rgrint_0n, df_0n[19]);
  AND2 I335 (rdfint_0n[20], rgrint_0n, df_0n[20]);
  AND2 I336 (rdfint_0n[21], rgrint_0n, df_0n[21]);
  AND2 I337 (rdfint_0n[22], rgrint_0n, df_0n[22]);
  AND2 I338 (rdfint_0n[23], rgrint_0n, df_0n[23]);
  AND2 I339 (rdfint_0n[24], rgrint_0n, df_0n[24]);
  AND2 I340 (rdfint_0n[25], rgrint_0n, df_0n[25]);
  AND2 I341 (rdfint_0n[26], rgrint_0n, df_0n[26]);
  AND2 I342 (rdfint_0n[27], rgrint_0n, df_0n[27]);
  AND2 I343 (rdfint_0n[28], rgrint_0n, df_0n[28]);
  AND2 I344 (rdfint_0n[29], rgrint_0n, df_0n[29]);
  AND2 I345 (rdfint_0n[30], rgrint_0n, df_0n[30]);
  C3 I346 (internal_0n[2], wc_0n, wacks_0n[34], wacks_0n[33]);
  C3 I347 (internal_0n[3], wacks_0n[32], wacks_0n[31], wacks_0n[30]);
  C3 I348 (internal_0n[4], wacks_0n[29], wacks_0n[28], wacks_0n[27]);
  C3 I349 (internal_0n[5], wacks_0n[26], wacks_0n[25], wacks_0n[24]);
  C3 I350 (internal_0n[6], wacks_0n[23], wacks_0n[22], wacks_0n[21]);
  C3 I351 (internal_0n[7], wacks_0n[20], wacks_0n[19], wacks_0n[18]);
  C3 I352 (internal_0n[8], wacks_0n[17], wacks_0n[16], wacks_0n[15]);
  C3 I353 (internal_0n[9], wacks_0n[14], wacks_0n[13], wacks_0n[12]);
  C3 I354 (internal_0n[10], wacks_0n[11], wacks_0n[10], wacks_0n[9]);
  C3 I355 (internal_0n[11], wacks_0n[8], wacks_0n[7], wacks_0n[6]);
  C3 I356 (internal_0n[12], wacks_0n[5], wacks_0n[4], wacks_0n[3]);
  C3 I357 (internal_0n[13], wacks_0n[2], wacks_0n[1], wacks_0n[0]);
  C3 I358 (internal_0n[14], internal_0n[2], internal_0n[3], internal_0n[4]);
  C3 I359 (internal_0n[15], internal_0n[5], internal_0n[6], internal_0n[7]);
  C3 I360 (internal_0n[16], internal_0n[8], internal_0n[9], internal_0n[10]);
  C3 I361 (internal_0n[17], internal_0n[11], internal_0n[12], internal_0n[13]);
  C2 I362 (internal_0n[18], internal_0n[14], internal_0n[15]);
  C2 I363 (internal_0n[19], internal_0n[16], internal_0n[17]);
  C2 I364 (wdrint_0n, internal_0n[18], internal_0n[19]);
  assign wen_0n[34] = wc_0n;
  assign wen_0n[33] = wc_0n;
  assign wen_0n[32] = wc_0n;
  assign wen_0n[31] = wc_0n;
  assign wen_0n[30] = wc_0n;
  assign wen_0n[29] = wc_0n;
  assign wen_0n[28] = wc_0n;
  assign wen_0n[27] = wc_0n;
  assign wen_0n[26] = wc_0n;
  assign wen_0n[25] = wc_0n;
  assign wen_0n[24] = wc_0n;
  assign wen_0n[23] = wc_0n;
  assign wen_0n[22] = wc_0n;
  assign wen_0n[21] = wc_0n;
  assign wen_0n[20] = wc_0n;
  assign wen_0n[19] = wc_0n;
  assign wen_0n[18] = wc_0n;
  assign wen_0n[17] = wc_0n;
  assign wen_0n[16] = wc_0n;
  assign wen_0n[15] = wc_0n;
  assign wen_0n[14] = wc_0n;
  assign wen_0n[13] = wc_0n;
  assign wen_0n[12] = wc_0n;
  assign wen_0n[11] = wc_0n;
  assign wen_0n[10] = wc_0n;
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[34] = git_0n[34];
  assign wt_0n[33] = git_0n[33];
  assign wt_0n[32] = git_0n[32];
  assign wt_0n[31] = git_0n[31];
  assign wt_0n[30] = git_0n[30];
  assign wt_0n[29] = git_0n[29];
  assign wt_0n[28] = git_0n[28];
  assign wt_0n[27] = git_0n[27];
  assign wt_0n[26] = git_0n[26];
  assign wt_0n[25] = git_0n[25];
  assign wt_0n[24] = git_0n[24];
  assign wt_0n[23] = git_0n[23];
  assign wt_0n[22] = git_0n[22];
  assign wt_0n[21] = git_0n[21];
  assign wt_0n[20] = git_0n[20];
  assign wt_0n[19] = git_0n[19];
  assign wt_0n[18] = git_0n[18];
  assign wt_0n[17] = git_0n[17];
  assign wt_0n[16] = git_0n[16];
  assign wt_0n[15] = git_0n[15];
  assign wt_0n[14] = git_0n[14];
  assign wt_0n[13] = git_0n[13];
  assign wt_0n[12] = git_0n[12];
  assign wt_0n[11] = git_0n[11];
  assign wt_0n[10] = git_0n[10];
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[34] = gif_0n[34];
  assign wf_0n[33] = gif_0n[33];
  assign wf_0n[32] = gif_0n[32];
  assign wf_0n[31] = gif_0n[31];
  assign wf_0n[30] = gif_0n[30];
  assign wf_0n[29] = gif_0n[29];
  assign wf_0n[28] = gif_0n[28];
  assign wf_0n[27] = gif_0n[27];
  assign wf_0n[26] = gif_0n[26];
  assign wf_0n[25] = gif_0n[25];
  assign wf_0n[24] = gif_0n[24];
  assign wf_0n[23] = gif_0n[23];
  assign wf_0n[22] = gif_0n[22];
  assign wf_0n[21] = gif_0n[21];
  assign wf_0n[20] = gif_0n[20];
  assign wf_0n[19] = gif_0n[19];
  assign wf_0n[18] = gif_0n[18];
  assign wf_0n[17] = gif_0n[17];
  assign wf_0n[16] = gif_0n[16];
  assign wf_0n[15] = gif_0n[15];
  assign wf_0n[14] = gif_0n[14];
  assign wf_0n[13] = gif_0n[13];
  assign wf_0n[12] = gif_0n[12];
  assign wf_0n[11] = gif_0n[11];
  assign wf_0n[10] = gif_0n[10];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I470 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I472 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I473 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I474 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I475 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I476 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I477 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I478 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I479 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I480 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I481 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I482 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I483 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I484 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I485 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I486 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I487 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I488 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I489 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I490 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I491 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I492 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I493 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I494 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I495 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I496 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I497 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I498 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I499 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I500 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I501 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I502 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I503 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I504 (git_0n[32], wgtint_0n[32], ig_0n);
  AND2 I505 (git_0n[33], wgtint_0n[33], ig_0n);
  AND2 I506 (git_0n[34], wgtint_0n[34], ig_0n);
  AND2 I507 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I508 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I509 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I510 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I511 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I512 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I513 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I514 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I515 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I516 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I517 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I518 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I519 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I520 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I521 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I522 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I523 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I524 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I525 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I526 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I527 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I528 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I529 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I530 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I531 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I532 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I533 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I534 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I535 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I536 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I537 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I538 (gif_0n[31], wgfint_0n[31], ig_0n);
  AND2 I539 (gif_0n[32], wgfint_0n[32], ig_0n);
  AND2 I540 (gif_0n[33], wgfint_0n[33], ig_0n);
  AND2 I541 (gif_0n[34], wgfint_0n[34], ig_0n);
  C3 I542 (internal_0n[20], complete1410_0n[0], complete1410_0n[1], complete1410_0n[2]);
  C3 I543 (internal_0n[21], complete1410_0n[3], complete1410_0n[4], complete1410_0n[5]);
  C3 I544 (internal_0n[22], complete1410_0n[6], complete1410_0n[7], complete1410_0n[8]);
  C3 I545 (internal_0n[23], complete1410_0n[9], complete1410_0n[10], complete1410_0n[11]);
  C3 I546 (internal_0n[24], complete1410_0n[12], complete1410_0n[13], complete1410_0n[14]);
  C3 I547 (internal_0n[25], complete1410_0n[15], complete1410_0n[16], complete1410_0n[17]);
  C3 I548 (internal_0n[26], complete1410_0n[18], complete1410_0n[19], complete1410_0n[20]);
  C3 I549 (internal_0n[27], complete1410_0n[21], complete1410_0n[22], complete1410_0n[23]);
  C3 I550 (internal_0n[28], complete1410_0n[24], complete1410_0n[25], complete1410_0n[26]);
  C3 I551 (internal_0n[29], complete1410_0n[27], complete1410_0n[28], complete1410_0n[29]);
  C3 I552 (internal_0n[30], complete1410_0n[30], complete1410_0n[31], complete1410_0n[32]);
  C2 I553 (internal_0n[31], complete1410_0n[33], complete1410_0n[34]);
  C3 I554 (internal_0n[32], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I555 (internal_0n[33], internal_0n[23], internal_0n[24], internal_0n[25]);
  C3 I556 (internal_0n[34], internal_0n[26], internal_0n[27], internal_0n[28]);
  C3 I557 (internal_0n[35], internal_0n[29], internal_0n[30], internal_0n[31]);
  C2 I558 (internal_0n[36], internal_0n[32], internal_0n[33]);
  C2 I559 (internal_0n[37], internal_0n[34], internal_0n[35]);
  C2 I560 (wc_0n, internal_0n[36], internal_0n[37]);
  OR2 I561 (complete1410_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I562 (complete1410_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I563 (complete1410_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I564 (complete1410_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I565 (complete1410_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I566 (complete1410_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I567 (complete1410_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I568 (complete1410_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I569 (complete1410_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I570 (complete1410_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I571 (complete1410_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I572 (complete1410_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I573 (complete1410_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I574 (complete1410_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I575 (complete1410_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I576 (complete1410_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I577 (complete1410_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I578 (complete1410_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I579 (complete1410_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I580 (complete1410_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I581 (complete1410_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I582 (complete1410_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I583 (complete1410_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I584 (complete1410_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I585 (complete1410_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I586 (complete1410_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I587 (complete1410_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I588 (complete1410_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I589 (complete1410_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I590 (complete1410_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I591 (complete1410_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I592 (complete1410_0n[31], wgfint_0n[31], wgtint_0n[31]);
  OR2 I593 (complete1410_0n[32], wgfint_0n[32], wgtint_0n[32]);
  OR2 I594 (complete1410_0n[33], wgfint_0n[33], wgtint_0n[33]);
  OR2 I595 (complete1410_0n[34], wgfint_0n[34], wgtint_0n[34]);
  AO22 I596 (wacks_0n[34], gf1408_0n[34], df_0n[34], gt1409_0n[34], dt_0n[34]);
  NOR2 I597 (dt_0n[34], df_0n[34], gf1408_0n[34]);
  NOR3 I598 (df_0n[34], dt_0n[34], gt1409_0n[34], init_0n);
  AND2 I599 (gt1409_0n[34], wt_0n[34], wen_0n[34]);
  AND2 I600 (gf1408_0n[34], wf_0n[34], wen_0n[34]);
  AO22 I601 (wacks_0n[33], gf1408_0n[33], df_0n[33], gt1409_0n[33], dt_0n[33]);
  NOR2 I602 (dt_0n[33], df_0n[33], gf1408_0n[33]);
  NOR3 I603 (df_0n[33], dt_0n[33], gt1409_0n[33], init_0n);
  AND2 I604 (gt1409_0n[33], wt_0n[33], wen_0n[33]);
  AND2 I605 (gf1408_0n[33], wf_0n[33], wen_0n[33]);
  AO22 I606 (wacks_0n[32], gf1408_0n[32], df_0n[32], gt1409_0n[32], dt_0n[32]);
  NOR2 I607 (dt_0n[32], df_0n[32], gf1408_0n[32]);
  NOR3 I608 (df_0n[32], dt_0n[32], gt1409_0n[32], init_0n);
  AND2 I609 (gt1409_0n[32], wt_0n[32], wen_0n[32]);
  AND2 I610 (gf1408_0n[32], wf_0n[32], wen_0n[32]);
  AO22 I611 (wacks_0n[31], gf1408_0n[31], df_0n[31], gt1409_0n[31], dt_0n[31]);
  NOR2 I612 (dt_0n[31], df_0n[31], gf1408_0n[31]);
  NOR3 I613 (df_0n[31], dt_0n[31], gt1409_0n[31], init_0n);
  AND2 I614 (gt1409_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I615 (gf1408_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I616 (wacks_0n[30], gf1408_0n[30], df_0n[30], gt1409_0n[30], dt_0n[30]);
  NOR2 I617 (dt_0n[30], df_0n[30], gf1408_0n[30]);
  NOR3 I618 (df_0n[30], dt_0n[30], gt1409_0n[30], init_0n);
  AND2 I619 (gt1409_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I620 (gf1408_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I621 (wacks_0n[29], gf1408_0n[29], df_0n[29], gt1409_0n[29], dt_0n[29]);
  NOR2 I622 (dt_0n[29], df_0n[29], gf1408_0n[29]);
  NOR3 I623 (df_0n[29], dt_0n[29], gt1409_0n[29], init_0n);
  AND2 I624 (gt1409_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I625 (gf1408_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I626 (wacks_0n[28], gf1408_0n[28], df_0n[28], gt1409_0n[28], dt_0n[28]);
  NOR2 I627 (dt_0n[28], df_0n[28], gf1408_0n[28]);
  NOR3 I628 (df_0n[28], dt_0n[28], gt1409_0n[28], init_0n);
  AND2 I629 (gt1409_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I630 (gf1408_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I631 (wacks_0n[27], gf1408_0n[27], df_0n[27], gt1409_0n[27], dt_0n[27]);
  NOR2 I632 (dt_0n[27], df_0n[27], gf1408_0n[27]);
  NOR3 I633 (df_0n[27], dt_0n[27], gt1409_0n[27], init_0n);
  AND2 I634 (gt1409_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I635 (gf1408_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I636 (wacks_0n[26], gf1408_0n[26], df_0n[26], gt1409_0n[26], dt_0n[26]);
  NOR2 I637 (dt_0n[26], df_0n[26], gf1408_0n[26]);
  NOR3 I638 (df_0n[26], dt_0n[26], gt1409_0n[26], init_0n);
  AND2 I639 (gt1409_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I640 (gf1408_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I641 (wacks_0n[25], gf1408_0n[25], df_0n[25], gt1409_0n[25], dt_0n[25]);
  NOR2 I642 (dt_0n[25], df_0n[25], gf1408_0n[25]);
  NOR3 I643 (df_0n[25], dt_0n[25], gt1409_0n[25], init_0n);
  AND2 I644 (gt1409_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I645 (gf1408_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I646 (wacks_0n[24], gf1408_0n[24], df_0n[24], gt1409_0n[24], dt_0n[24]);
  NOR2 I647 (dt_0n[24], df_0n[24], gf1408_0n[24]);
  NOR3 I648 (df_0n[24], dt_0n[24], gt1409_0n[24], init_0n);
  AND2 I649 (gt1409_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I650 (gf1408_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I651 (wacks_0n[23], gf1408_0n[23], df_0n[23], gt1409_0n[23], dt_0n[23]);
  NOR2 I652 (dt_0n[23], df_0n[23], gf1408_0n[23]);
  NOR3 I653 (df_0n[23], dt_0n[23], gt1409_0n[23], init_0n);
  AND2 I654 (gt1409_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I655 (gf1408_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I656 (wacks_0n[22], gf1408_0n[22], df_0n[22], gt1409_0n[22], dt_0n[22]);
  NOR2 I657 (dt_0n[22], df_0n[22], gf1408_0n[22]);
  NOR3 I658 (df_0n[22], dt_0n[22], gt1409_0n[22], init_0n);
  AND2 I659 (gt1409_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I660 (gf1408_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I661 (wacks_0n[21], gf1408_0n[21], df_0n[21], gt1409_0n[21], dt_0n[21]);
  NOR2 I662 (dt_0n[21], df_0n[21], gf1408_0n[21]);
  NOR3 I663 (df_0n[21], dt_0n[21], gt1409_0n[21], init_0n);
  AND2 I664 (gt1409_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I665 (gf1408_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I666 (wacks_0n[20], gf1408_0n[20], df_0n[20], gt1409_0n[20], dt_0n[20]);
  NOR2 I667 (dt_0n[20], df_0n[20], gf1408_0n[20]);
  NOR3 I668 (df_0n[20], dt_0n[20], gt1409_0n[20], init_0n);
  AND2 I669 (gt1409_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I670 (gf1408_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I671 (wacks_0n[19], gf1408_0n[19], df_0n[19], gt1409_0n[19], dt_0n[19]);
  NOR2 I672 (dt_0n[19], df_0n[19], gf1408_0n[19]);
  NOR3 I673 (df_0n[19], dt_0n[19], gt1409_0n[19], init_0n);
  AND2 I674 (gt1409_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I675 (gf1408_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I676 (wacks_0n[18], gf1408_0n[18], df_0n[18], gt1409_0n[18], dt_0n[18]);
  NOR2 I677 (dt_0n[18], df_0n[18], gf1408_0n[18]);
  NOR3 I678 (df_0n[18], dt_0n[18], gt1409_0n[18], init_0n);
  AND2 I679 (gt1409_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I680 (gf1408_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I681 (wacks_0n[17], gf1408_0n[17], df_0n[17], gt1409_0n[17], dt_0n[17]);
  NOR2 I682 (dt_0n[17], df_0n[17], gf1408_0n[17]);
  NOR3 I683 (df_0n[17], dt_0n[17], gt1409_0n[17], init_0n);
  AND2 I684 (gt1409_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I685 (gf1408_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I686 (wacks_0n[16], gf1408_0n[16], df_0n[16], gt1409_0n[16], dt_0n[16]);
  NOR2 I687 (dt_0n[16], df_0n[16], gf1408_0n[16]);
  NOR3 I688 (df_0n[16], dt_0n[16], gt1409_0n[16], init_0n);
  AND2 I689 (gt1409_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I690 (gf1408_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I691 (wacks_0n[15], gf1408_0n[15], df_0n[15], gt1409_0n[15], dt_0n[15]);
  NOR2 I692 (dt_0n[15], df_0n[15], gf1408_0n[15]);
  NOR3 I693 (df_0n[15], dt_0n[15], gt1409_0n[15], init_0n);
  AND2 I694 (gt1409_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I695 (gf1408_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I696 (wacks_0n[14], gf1408_0n[14], df_0n[14], gt1409_0n[14], dt_0n[14]);
  NOR2 I697 (dt_0n[14], df_0n[14], gf1408_0n[14]);
  NOR3 I698 (df_0n[14], dt_0n[14], gt1409_0n[14], init_0n);
  AND2 I699 (gt1409_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I700 (gf1408_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I701 (wacks_0n[13], gf1408_0n[13], df_0n[13], gt1409_0n[13], dt_0n[13]);
  NOR2 I702 (dt_0n[13], df_0n[13], gf1408_0n[13]);
  NOR3 I703 (df_0n[13], dt_0n[13], gt1409_0n[13], init_0n);
  AND2 I704 (gt1409_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I705 (gf1408_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I706 (wacks_0n[12], gf1408_0n[12], df_0n[12], gt1409_0n[12], dt_0n[12]);
  NOR2 I707 (dt_0n[12], df_0n[12], gf1408_0n[12]);
  NOR3 I708 (df_0n[12], dt_0n[12], gt1409_0n[12], init_0n);
  AND2 I709 (gt1409_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I710 (gf1408_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I711 (wacks_0n[11], gf1408_0n[11], df_0n[11], gt1409_0n[11], dt_0n[11]);
  NOR2 I712 (dt_0n[11], df_0n[11], gf1408_0n[11]);
  NOR3 I713 (df_0n[11], dt_0n[11], gt1409_0n[11], init_0n);
  AND2 I714 (gt1409_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I715 (gf1408_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I716 (wacks_0n[10], gf1408_0n[10], df_0n[10], gt1409_0n[10], dt_0n[10]);
  NOR2 I717 (dt_0n[10], df_0n[10], gf1408_0n[10]);
  NOR3 I718 (df_0n[10], dt_0n[10], gt1409_0n[10], init_0n);
  AND2 I719 (gt1409_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I720 (gf1408_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I721 (wacks_0n[9], gf1408_0n[9], df_0n[9], gt1409_0n[9], dt_0n[9]);
  NOR2 I722 (dt_0n[9], df_0n[9], gf1408_0n[9]);
  NOR3 I723 (df_0n[9], dt_0n[9], gt1409_0n[9], init_0n);
  AND2 I724 (gt1409_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I725 (gf1408_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I726 (wacks_0n[8], gf1408_0n[8], df_0n[8], gt1409_0n[8], dt_0n[8]);
  NOR2 I727 (dt_0n[8], df_0n[8], gf1408_0n[8]);
  NOR3 I728 (df_0n[8], dt_0n[8], gt1409_0n[8], init_0n);
  AND2 I729 (gt1409_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I730 (gf1408_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I731 (wacks_0n[7], gf1408_0n[7], df_0n[7], gt1409_0n[7], dt_0n[7]);
  NOR2 I732 (dt_0n[7], df_0n[7], gf1408_0n[7]);
  NOR3 I733 (df_0n[7], dt_0n[7], gt1409_0n[7], init_0n);
  AND2 I734 (gt1409_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I735 (gf1408_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I736 (wacks_0n[6], gf1408_0n[6], df_0n[6], gt1409_0n[6], dt_0n[6]);
  NOR2 I737 (dt_0n[6], df_0n[6], gf1408_0n[6]);
  NOR3 I738 (df_0n[6], dt_0n[6], gt1409_0n[6], init_0n);
  AND2 I739 (gt1409_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I740 (gf1408_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I741 (wacks_0n[5], gf1408_0n[5], df_0n[5], gt1409_0n[5], dt_0n[5]);
  NOR2 I742 (dt_0n[5], df_0n[5], gf1408_0n[5]);
  NOR3 I743 (df_0n[5], dt_0n[5], gt1409_0n[5], init_0n);
  AND2 I744 (gt1409_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I745 (gf1408_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I746 (wacks_0n[4], gf1408_0n[4], df_0n[4], gt1409_0n[4], dt_0n[4]);
  NOR2 I747 (dt_0n[4], df_0n[4], gf1408_0n[4]);
  NOR3 I748 (df_0n[4], dt_0n[4], gt1409_0n[4], init_0n);
  AND2 I749 (gt1409_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I750 (gf1408_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I751 (wacks_0n[3], gf1408_0n[3], df_0n[3], gt1409_0n[3], dt_0n[3]);
  NOR2 I752 (dt_0n[3], df_0n[3], gf1408_0n[3]);
  NOR3 I753 (df_0n[3], dt_0n[3], gt1409_0n[3], init_0n);
  AND2 I754 (gt1409_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I755 (gf1408_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I756 (wacks_0n[2], gf1408_0n[2], df_0n[2], gt1409_0n[2], dt_0n[2]);
  NOR2 I757 (dt_0n[2], df_0n[2], gf1408_0n[2]);
  NOR3 I758 (df_0n[2], dt_0n[2], gt1409_0n[2], init_0n);
  AND2 I759 (gt1409_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I760 (gf1408_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I761 (wacks_0n[1], gf1408_0n[1], df_0n[1], gt1409_0n[1], dt_0n[1]);
  NOR2 I762 (dt_0n[1], df_0n[1], gf1408_0n[1]);
  NOR3 I763 (df_0n[1], dt_0n[1], gt1409_0n[1], init_0n);
  AND2 I764 (gt1409_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I765 (gf1408_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I766 (wacks_0n[0], gf1408_0n[0], df_0n[0], gt1409_0n[0], dt_0n[0]);
  NOR2 I767 (dt_0n[0], df_0n[0], gf1408_0n[0]);
  NOR3 I768 (df_0n[0], dt_0n[0], gt1409_0n[0], init_0n);
  AND2 I769 (gt1409_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I770 (gf1408_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I771 (init_0n, initialise);
endmodule

module BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rd_0r0d, rd_0r1d, rd_0a,
  initialise
);
  input [34:0] wg_0r0d;
  input [34:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [34:0] rd_0r0d;
  output [34:0] rd_0r1d;
  input rd_0a;
  input initialise;
  wire [35:0] internal_0n;
  wire [34:0] wf_0n;
  wire [34:0] wt_0n;
  wire [34:0] df_0n;
  wire [34:0] dt_0n;
  wire rgrint_0n;
  wire wc_0n;
  wire [34:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [34:0] wgfint_0n;
  wire [34:0] wgtint_0n;
  wire rgaint_0n;
  wire [34:0] rdfint_0n;
  wire [34:0] rdtint_0n;
  wire [34:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [34:0] gif_0n;
  wire [34:0] git_0n;
  wire [34:0] complete1425_0n;
  wire [34:0] gt1424_0n;
  wire [34:0] gf1423_0n;
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r0d[10] = rdfint_0n[10];
  assign rd_0r0d[11] = rdfint_0n[11];
  assign rd_0r0d[12] = rdfint_0n[12];
  assign rd_0r0d[13] = rdfint_0n[13];
  assign rd_0r0d[14] = rdfint_0n[14];
  assign rd_0r0d[15] = rdfint_0n[15];
  assign rd_0r0d[16] = rdfint_0n[16];
  assign rd_0r0d[17] = rdfint_0n[17];
  assign rd_0r0d[18] = rdfint_0n[18];
  assign rd_0r0d[19] = rdfint_0n[19];
  assign rd_0r0d[20] = rdfint_0n[20];
  assign rd_0r0d[21] = rdfint_0n[21];
  assign rd_0r0d[22] = rdfint_0n[22];
  assign rd_0r0d[23] = rdfint_0n[23];
  assign rd_0r0d[24] = rdfint_0n[24];
  assign rd_0r0d[25] = rdfint_0n[25];
  assign rd_0r0d[26] = rdfint_0n[26];
  assign rd_0r0d[27] = rdfint_0n[27];
  assign rd_0r0d[28] = rdfint_0n[28];
  assign rd_0r0d[29] = rdfint_0n[29];
  assign rd_0r0d[30] = rdfint_0n[30];
  assign rd_0r0d[31] = rdfint_0n[31];
  assign rd_0r0d[32] = rdfint_0n[32];
  assign rd_0r0d[33] = rdfint_0n[33];
  assign rd_0r0d[34] = rdfint_0n[34];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign rd_0r1d[10] = rdtint_0n[10];
  assign rd_0r1d[11] = rdtint_0n[11];
  assign rd_0r1d[12] = rdtint_0n[12];
  assign rd_0r1d[13] = rdtint_0n[13];
  assign rd_0r1d[14] = rdtint_0n[14];
  assign rd_0r1d[15] = rdtint_0n[15];
  assign rd_0r1d[16] = rdtint_0n[16];
  assign rd_0r1d[17] = rdtint_0n[17];
  assign rd_0r1d[18] = rdtint_0n[18];
  assign rd_0r1d[19] = rdtint_0n[19];
  assign rd_0r1d[20] = rdtint_0n[20];
  assign rd_0r1d[21] = rdtint_0n[21];
  assign rd_0r1d[22] = rdtint_0n[22];
  assign rd_0r1d[23] = rdtint_0n[23];
  assign rd_0r1d[24] = rdtint_0n[24];
  assign rd_0r1d[25] = rdtint_0n[25];
  assign rd_0r1d[26] = rdtint_0n[26];
  assign rd_0r1d[27] = rdtint_0n[27];
  assign rd_0r1d[28] = rdtint_0n[28];
  assign rd_0r1d[29] = rdtint_0n[29];
  assign rd_0r1d[30] = rdtint_0n[30];
  assign rd_0r1d[31] = rdtint_0n[31];
  assign rd_0r1d[32] = rdtint_0n[32];
  assign rd_0r1d[33] = rdtint_0n[33];
  assign rd_0r1d[34] = rdtint_0n[34];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgfint_0n[32] = wg_0r0d[32];
  assign wgfint_0n[33] = wg_0r0d[33];
  assign wgfint_0n[34] = wg_0r0d[34];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign wgtint_0n[32] = wg_0r1d[32];
  assign wgtint_0n[33] = wg_0r1d[33];
  assign wgtint_0n[34] = wg_0r1d[34];
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I146 (nanyread_0n, rgrint_0n, rgaint_0n);
  AND2 I147 (rdtint_0n[0], rgrint_0n, dt_0n[0]);
  AND2 I148 (rdtint_0n[1], rgrint_0n, dt_0n[1]);
  AND2 I149 (rdtint_0n[2], rgrint_0n, dt_0n[2]);
  AND2 I150 (rdtint_0n[3], rgrint_0n, dt_0n[3]);
  AND2 I151 (rdtint_0n[4], rgrint_0n, dt_0n[4]);
  AND2 I152 (rdtint_0n[5], rgrint_0n, dt_0n[5]);
  AND2 I153 (rdtint_0n[6], rgrint_0n, dt_0n[6]);
  AND2 I154 (rdtint_0n[7], rgrint_0n, dt_0n[7]);
  AND2 I155 (rdtint_0n[8], rgrint_0n, dt_0n[8]);
  AND2 I156 (rdtint_0n[9], rgrint_0n, dt_0n[9]);
  AND2 I157 (rdtint_0n[10], rgrint_0n, dt_0n[10]);
  AND2 I158 (rdtint_0n[11], rgrint_0n, dt_0n[11]);
  AND2 I159 (rdtint_0n[12], rgrint_0n, dt_0n[12]);
  AND2 I160 (rdtint_0n[13], rgrint_0n, dt_0n[13]);
  AND2 I161 (rdtint_0n[14], rgrint_0n, dt_0n[14]);
  AND2 I162 (rdtint_0n[15], rgrint_0n, dt_0n[15]);
  AND2 I163 (rdtint_0n[16], rgrint_0n, dt_0n[16]);
  AND2 I164 (rdtint_0n[17], rgrint_0n, dt_0n[17]);
  AND2 I165 (rdtint_0n[18], rgrint_0n, dt_0n[18]);
  AND2 I166 (rdtint_0n[19], rgrint_0n, dt_0n[19]);
  AND2 I167 (rdtint_0n[20], rgrint_0n, dt_0n[20]);
  AND2 I168 (rdtint_0n[21], rgrint_0n, dt_0n[21]);
  AND2 I169 (rdtint_0n[22], rgrint_0n, dt_0n[22]);
  AND2 I170 (rdtint_0n[23], rgrint_0n, dt_0n[23]);
  AND2 I171 (rdtint_0n[24], rgrint_0n, dt_0n[24]);
  AND2 I172 (rdtint_0n[25], rgrint_0n, dt_0n[25]);
  AND2 I173 (rdtint_0n[26], rgrint_0n, dt_0n[26]);
  AND2 I174 (rdtint_0n[27], rgrint_0n, dt_0n[27]);
  AND2 I175 (rdtint_0n[28], rgrint_0n, dt_0n[28]);
  AND2 I176 (rdtint_0n[29], rgrint_0n, dt_0n[29]);
  AND2 I177 (rdtint_0n[30], rgrint_0n, dt_0n[30]);
  AND2 I178 (rdtint_0n[31], rgrint_0n, dt_0n[31]);
  AND2 I179 (rdtint_0n[32], rgrint_0n, dt_0n[32]);
  AND2 I180 (rdtint_0n[33], rgrint_0n, dt_0n[33]);
  AND2 I181 (rdtint_0n[34], rgrint_0n, dt_0n[34]);
  AND2 I182 (rdfint_0n[0], rgrint_0n, df_0n[0]);
  AND2 I183 (rdfint_0n[1], rgrint_0n, df_0n[1]);
  AND2 I184 (rdfint_0n[2], rgrint_0n, df_0n[2]);
  AND2 I185 (rdfint_0n[3], rgrint_0n, df_0n[3]);
  AND2 I186 (rdfint_0n[4], rgrint_0n, df_0n[4]);
  AND2 I187 (rdfint_0n[5], rgrint_0n, df_0n[5]);
  AND2 I188 (rdfint_0n[6], rgrint_0n, df_0n[6]);
  AND2 I189 (rdfint_0n[7], rgrint_0n, df_0n[7]);
  AND2 I190 (rdfint_0n[8], rgrint_0n, df_0n[8]);
  AND2 I191 (rdfint_0n[9], rgrint_0n, df_0n[9]);
  AND2 I192 (rdfint_0n[10], rgrint_0n, df_0n[10]);
  AND2 I193 (rdfint_0n[11], rgrint_0n, df_0n[11]);
  AND2 I194 (rdfint_0n[12], rgrint_0n, df_0n[12]);
  AND2 I195 (rdfint_0n[13], rgrint_0n, df_0n[13]);
  AND2 I196 (rdfint_0n[14], rgrint_0n, df_0n[14]);
  AND2 I197 (rdfint_0n[15], rgrint_0n, df_0n[15]);
  AND2 I198 (rdfint_0n[16], rgrint_0n, df_0n[16]);
  AND2 I199 (rdfint_0n[17], rgrint_0n, df_0n[17]);
  AND2 I200 (rdfint_0n[18], rgrint_0n, df_0n[18]);
  AND2 I201 (rdfint_0n[19], rgrint_0n, df_0n[19]);
  AND2 I202 (rdfint_0n[20], rgrint_0n, df_0n[20]);
  AND2 I203 (rdfint_0n[21], rgrint_0n, df_0n[21]);
  AND2 I204 (rdfint_0n[22], rgrint_0n, df_0n[22]);
  AND2 I205 (rdfint_0n[23], rgrint_0n, df_0n[23]);
  AND2 I206 (rdfint_0n[24], rgrint_0n, df_0n[24]);
  AND2 I207 (rdfint_0n[25], rgrint_0n, df_0n[25]);
  AND2 I208 (rdfint_0n[26], rgrint_0n, df_0n[26]);
  AND2 I209 (rdfint_0n[27], rgrint_0n, df_0n[27]);
  AND2 I210 (rdfint_0n[28], rgrint_0n, df_0n[28]);
  AND2 I211 (rdfint_0n[29], rgrint_0n, df_0n[29]);
  AND2 I212 (rdfint_0n[30], rgrint_0n, df_0n[30]);
  AND2 I213 (rdfint_0n[31], rgrint_0n, df_0n[31]);
  AND2 I214 (rdfint_0n[32], rgrint_0n, df_0n[32]);
  AND2 I215 (rdfint_0n[33], rgrint_0n, df_0n[33]);
  AND2 I216 (rdfint_0n[34], rgrint_0n, df_0n[34]);
  C3 I217 (internal_0n[0], wc_0n, wacks_0n[34], wacks_0n[33]);
  C3 I218 (internal_0n[1], wacks_0n[32], wacks_0n[31], wacks_0n[30]);
  C3 I219 (internal_0n[2], wacks_0n[29], wacks_0n[28], wacks_0n[27]);
  C3 I220 (internal_0n[3], wacks_0n[26], wacks_0n[25], wacks_0n[24]);
  C3 I221 (internal_0n[4], wacks_0n[23], wacks_0n[22], wacks_0n[21]);
  C3 I222 (internal_0n[5], wacks_0n[20], wacks_0n[19], wacks_0n[18]);
  C3 I223 (internal_0n[6], wacks_0n[17], wacks_0n[16], wacks_0n[15]);
  C3 I224 (internal_0n[7], wacks_0n[14], wacks_0n[13], wacks_0n[12]);
  C3 I225 (internal_0n[8], wacks_0n[11], wacks_0n[10], wacks_0n[9]);
  C3 I226 (internal_0n[9], wacks_0n[8], wacks_0n[7], wacks_0n[6]);
  C3 I227 (internal_0n[10], wacks_0n[5], wacks_0n[4], wacks_0n[3]);
  C3 I228 (internal_0n[11], wacks_0n[2], wacks_0n[1], wacks_0n[0]);
  C3 I229 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I230 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I231 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I232 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I233 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I234 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I235 (wdrint_0n, internal_0n[16], internal_0n[17]);
  assign wen_0n[34] = wc_0n;
  assign wen_0n[33] = wc_0n;
  assign wen_0n[32] = wc_0n;
  assign wen_0n[31] = wc_0n;
  assign wen_0n[30] = wc_0n;
  assign wen_0n[29] = wc_0n;
  assign wen_0n[28] = wc_0n;
  assign wen_0n[27] = wc_0n;
  assign wen_0n[26] = wc_0n;
  assign wen_0n[25] = wc_0n;
  assign wen_0n[24] = wc_0n;
  assign wen_0n[23] = wc_0n;
  assign wen_0n[22] = wc_0n;
  assign wen_0n[21] = wc_0n;
  assign wen_0n[20] = wc_0n;
  assign wen_0n[19] = wc_0n;
  assign wen_0n[18] = wc_0n;
  assign wen_0n[17] = wc_0n;
  assign wen_0n[16] = wc_0n;
  assign wen_0n[15] = wc_0n;
  assign wen_0n[14] = wc_0n;
  assign wen_0n[13] = wc_0n;
  assign wen_0n[12] = wc_0n;
  assign wen_0n[11] = wc_0n;
  assign wen_0n[10] = wc_0n;
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[34] = git_0n[34];
  assign wt_0n[33] = git_0n[33];
  assign wt_0n[32] = git_0n[32];
  assign wt_0n[31] = git_0n[31];
  assign wt_0n[30] = git_0n[30];
  assign wt_0n[29] = git_0n[29];
  assign wt_0n[28] = git_0n[28];
  assign wt_0n[27] = git_0n[27];
  assign wt_0n[26] = git_0n[26];
  assign wt_0n[25] = git_0n[25];
  assign wt_0n[24] = git_0n[24];
  assign wt_0n[23] = git_0n[23];
  assign wt_0n[22] = git_0n[22];
  assign wt_0n[21] = git_0n[21];
  assign wt_0n[20] = git_0n[20];
  assign wt_0n[19] = git_0n[19];
  assign wt_0n[18] = git_0n[18];
  assign wt_0n[17] = git_0n[17];
  assign wt_0n[16] = git_0n[16];
  assign wt_0n[15] = git_0n[15];
  assign wt_0n[14] = git_0n[14];
  assign wt_0n[13] = git_0n[13];
  assign wt_0n[12] = git_0n[12];
  assign wt_0n[11] = git_0n[11];
  assign wt_0n[10] = git_0n[10];
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[34] = gif_0n[34];
  assign wf_0n[33] = gif_0n[33];
  assign wf_0n[32] = gif_0n[32];
  assign wf_0n[31] = gif_0n[31];
  assign wf_0n[30] = gif_0n[30];
  assign wf_0n[29] = gif_0n[29];
  assign wf_0n[28] = gif_0n[28];
  assign wf_0n[27] = gif_0n[27];
  assign wf_0n[26] = gif_0n[26];
  assign wf_0n[25] = gif_0n[25];
  assign wf_0n[24] = gif_0n[24];
  assign wf_0n[23] = gif_0n[23];
  assign wf_0n[22] = gif_0n[22];
  assign wf_0n[21] = gif_0n[21];
  assign wf_0n[20] = gif_0n[20];
  assign wf_0n[19] = gif_0n[19];
  assign wf_0n[18] = gif_0n[18];
  assign wf_0n[17] = gif_0n[17];
  assign wf_0n[16] = gif_0n[16];
  assign wf_0n[15] = gif_0n[15];
  assign wf_0n[14] = gif_0n[14];
  assign wf_0n[13] = gif_0n[13];
  assign wf_0n[12] = gif_0n[12];
  assign wf_0n[11] = gif_0n[11];
  assign wf_0n[10] = gif_0n[10];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I341 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I343 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I344 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I345 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I346 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I347 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I348 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I349 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I350 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I351 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I352 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I353 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I354 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I355 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I356 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I357 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I358 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I359 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I360 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I361 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I362 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I363 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I364 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I365 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I366 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I367 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I368 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I369 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I370 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I371 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I372 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I373 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I374 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I375 (git_0n[32], wgtint_0n[32], ig_0n);
  AND2 I376 (git_0n[33], wgtint_0n[33], ig_0n);
  AND2 I377 (git_0n[34], wgtint_0n[34], ig_0n);
  AND2 I378 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I379 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I380 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I381 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I382 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I383 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I384 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I385 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I386 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I387 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I388 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I389 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I390 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I391 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I392 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I393 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I394 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I395 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I396 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I397 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I398 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I399 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I400 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I401 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I402 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I403 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I404 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I405 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I406 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I407 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I408 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I409 (gif_0n[31], wgfint_0n[31], ig_0n);
  AND2 I410 (gif_0n[32], wgfint_0n[32], ig_0n);
  AND2 I411 (gif_0n[33], wgfint_0n[33], ig_0n);
  AND2 I412 (gif_0n[34], wgfint_0n[34], ig_0n);
  C3 I413 (internal_0n[18], complete1425_0n[0], complete1425_0n[1], complete1425_0n[2]);
  C3 I414 (internal_0n[19], complete1425_0n[3], complete1425_0n[4], complete1425_0n[5]);
  C3 I415 (internal_0n[20], complete1425_0n[6], complete1425_0n[7], complete1425_0n[8]);
  C3 I416 (internal_0n[21], complete1425_0n[9], complete1425_0n[10], complete1425_0n[11]);
  C3 I417 (internal_0n[22], complete1425_0n[12], complete1425_0n[13], complete1425_0n[14]);
  C3 I418 (internal_0n[23], complete1425_0n[15], complete1425_0n[16], complete1425_0n[17]);
  C3 I419 (internal_0n[24], complete1425_0n[18], complete1425_0n[19], complete1425_0n[20]);
  C3 I420 (internal_0n[25], complete1425_0n[21], complete1425_0n[22], complete1425_0n[23]);
  C3 I421 (internal_0n[26], complete1425_0n[24], complete1425_0n[25], complete1425_0n[26]);
  C3 I422 (internal_0n[27], complete1425_0n[27], complete1425_0n[28], complete1425_0n[29]);
  C3 I423 (internal_0n[28], complete1425_0n[30], complete1425_0n[31], complete1425_0n[32]);
  C2 I424 (internal_0n[29], complete1425_0n[33], complete1425_0n[34]);
  C3 I425 (internal_0n[30], internal_0n[18], internal_0n[19], internal_0n[20]);
  C3 I426 (internal_0n[31], internal_0n[21], internal_0n[22], internal_0n[23]);
  C3 I427 (internal_0n[32], internal_0n[24], internal_0n[25], internal_0n[26]);
  C3 I428 (internal_0n[33], internal_0n[27], internal_0n[28], internal_0n[29]);
  C2 I429 (internal_0n[34], internal_0n[30], internal_0n[31]);
  C2 I430 (internal_0n[35], internal_0n[32], internal_0n[33]);
  C2 I431 (wc_0n, internal_0n[34], internal_0n[35]);
  OR2 I432 (complete1425_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I433 (complete1425_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I434 (complete1425_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I435 (complete1425_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I436 (complete1425_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I437 (complete1425_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I438 (complete1425_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I439 (complete1425_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I440 (complete1425_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I441 (complete1425_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I442 (complete1425_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I443 (complete1425_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I444 (complete1425_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I445 (complete1425_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I446 (complete1425_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I447 (complete1425_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I448 (complete1425_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I449 (complete1425_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I450 (complete1425_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I451 (complete1425_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I452 (complete1425_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I453 (complete1425_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I454 (complete1425_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I455 (complete1425_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I456 (complete1425_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I457 (complete1425_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I458 (complete1425_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I459 (complete1425_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I460 (complete1425_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I461 (complete1425_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I462 (complete1425_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I463 (complete1425_0n[31], wgfint_0n[31], wgtint_0n[31]);
  OR2 I464 (complete1425_0n[32], wgfint_0n[32], wgtint_0n[32]);
  OR2 I465 (complete1425_0n[33], wgfint_0n[33], wgtint_0n[33]);
  OR2 I466 (complete1425_0n[34], wgfint_0n[34], wgtint_0n[34]);
  AO22 I467 (wacks_0n[34], gf1423_0n[34], df_0n[34], gt1424_0n[34], dt_0n[34]);
  NOR2 I468 (dt_0n[34], df_0n[34], gf1423_0n[34]);
  NOR3 I469 (df_0n[34], dt_0n[34], gt1424_0n[34], init_0n);
  AND2 I470 (gt1424_0n[34], wt_0n[34], wen_0n[34]);
  AND2 I471 (gf1423_0n[34], wf_0n[34], wen_0n[34]);
  AO22 I472 (wacks_0n[33], gf1423_0n[33], df_0n[33], gt1424_0n[33], dt_0n[33]);
  NOR2 I473 (dt_0n[33], df_0n[33], gf1423_0n[33]);
  NOR3 I474 (df_0n[33], dt_0n[33], gt1424_0n[33], init_0n);
  AND2 I475 (gt1424_0n[33], wt_0n[33], wen_0n[33]);
  AND2 I476 (gf1423_0n[33], wf_0n[33], wen_0n[33]);
  AO22 I477 (wacks_0n[32], gf1423_0n[32], df_0n[32], gt1424_0n[32], dt_0n[32]);
  NOR2 I478 (dt_0n[32], df_0n[32], gf1423_0n[32]);
  NOR3 I479 (df_0n[32], dt_0n[32], gt1424_0n[32], init_0n);
  AND2 I480 (gt1424_0n[32], wt_0n[32], wen_0n[32]);
  AND2 I481 (gf1423_0n[32], wf_0n[32], wen_0n[32]);
  AO22 I482 (wacks_0n[31], gf1423_0n[31], df_0n[31], gt1424_0n[31], dt_0n[31]);
  NOR2 I483 (dt_0n[31], df_0n[31], gf1423_0n[31]);
  NOR3 I484 (df_0n[31], dt_0n[31], gt1424_0n[31], init_0n);
  AND2 I485 (gt1424_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I486 (gf1423_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I487 (wacks_0n[30], gf1423_0n[30], df_0n[30], gt1424_0n[30], dt_0n[30]);
  NOR2 I488 (dt_0n[30], df_0n[30], gf1423_0n[30]);
  NOR3 I489 (df_0n[30], dt_0n[30], gt1424_0n[30], init_0n);
  AND2 I490 (gt1424_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I491 (gf1423_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I492 (wacks_0n[29], gf1423_0n[29], df_0n[29], gt1424_0n[29], dt_0n[29]);
  NOR2 I493 (dt_0n[29], df_0n[29], gf1423_0n[29]);
  NOR3 I494 (df_0n[29], dt_0n[29], gt1424_0n[29], init_0n);
  AND2 I495 (gt1424_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I496 (gf1423_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I497 (wacks_0n[28], gf1423_0n[28], df_0n[28], gt1424_0n[28], dt_0n[28]);
  NOR2 I498 (dt_0n[28], df_0n[28], gf1423_0n[28]);
  NOR3 I499 (df_0n[28], dt_0n[28], gt1424_0n[28], init_0n);
  AND2 I500 (gt1424_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I501 (gf1423_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I502 (wacks_0n[27], gf1423_0n[27], df_0n[27], gt1424_0n[27], dt_0n[27]);
  NOR2 I503 (dt_0n[27], df_0n[27], gf1423_0n[27]);
  NOR3 I504 (df_0n[27], dt_0n[27], gt1424_0n[27], init_0n);
  AND2 I505 (gt1424_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I506 (gf1423_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I507 (wacks_0n[26], gf1423_0n[26], df_0n[26], gt1424_0n[26], dt_0n[26]);
  NOR2 I508 (dt_0n[26], df_0n[26], gf1423_0n[26]);
  NOR3 I509 (df_0n[26], dt_0n[26], gt1424_0n[26], init_0n);
  AND2 I510 (gt1424_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I511 (gf1423_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I512 (wacks_0n[25], gf1423_0n[25], df_0n[25], gt1424_0n[25], dt_0n[25]);
  NOR2 I513 (dt_0n[25], df_0n[25], gf1423_0n[25]);
  NOR3 I514 (df_0n[25], dt_0n[25], gt1424_0n[25], init_0n);
  AND2 I515 (gt1424_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I516 (gf1423_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I517 (wacks_0n[24], gf1423_0n[24], df_0n[24], gt1424_0n[24], dt_0n[24]);
  NOR2 I518 (dt_0n[24], df_0n[24], gf1423_0n[24]);
  NOR3 I519 (df_0n[24], dt_0n[24], gt1424_0n[24], init_0n);
  AND2 I520 (gt1424_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I521 (gf1423_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I522 (wacks_0n[23], gf1423_0n[23], df_0n[23], gt1424_0n[23], dt_0n[23]);
  NOR2 I523 (dt_0n[23], df_0n[23], gf1423_0n[23]);
  NOR3 I524 (df_0n[23], dt_0n[23], gt1424_0n[23], init_0n);
  AND2 I525 (gt1424_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I526 (gf1423_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I527 (wacks_0n[22], gf1423_0n[22], df_0n[22], gt1424_0n[22], dt_0n[22]);
  NOR2 I528 (dt_0n[22], df_0n[22], gf1423_0n[22]);
  NOR3 I529 (df_0n[22], dt_0n[22], gt1424_0n[22], init_0n);
  AND2 I530 (gt1424_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I531 (gf1423_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I532 (wacks_0n[21], gf1423_0n[21], df_0n[21], gt1424_0n[21], dt_0n[21]);
  NOR2 I533 (dt_0n[21], df_0n[21], gf1423_0n[21]);
  NOR3 I534 (df_0n[21], dt_0n[21], gt1424_0n[21], init_0n);
  AND2 I535 (gt1424_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I536 (gf1423_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I537 (wacks_0n[20], gf1423_0n[20], df_0n[20], gt1424_0n[20], dt_0n[20]);
  NOR2 I538 (dt_0n[20], df_0n[20], gf1423_0n[20]);
  NOR3 I539 (df_0n[20], dt_0n[20], gt1424_0n[20], init_0n);
  AND2 I540 (gt1424_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I541 (gf1423_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I542 (wacks_0n[19], gf1423_0n[19], df_0n[19], gt1424_0n[19], dt_0n[19]);
  NOR2 I543 (dt_0n[19], df_0n[19], gf1423_0n[19]);
  NOR3 I544 (df_0n[19], dt_0n[19], gt1424_0n[19], init_0n);
  AND2 I545 (gt1424_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I546 (gf1423_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I547 (wacks_0n[18], gf1423_0n[18], df_0n[18], gt1424_0n[18], dt_0n[18]);
  NOR2 I548 (dt_0n[18], df_0n[18], gf1423_0n[18]);
  NOR3 I549 (df_0n[18], dt_0n[18], gt1424_0n[18], init_0n);
  AND2 I550 (gt1424_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I551 (gf1423_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I552 (wacks_0n[17], gf1423_0n[17], df_0n[17], gt1424_0n[17], dt_0n[17]);
  NOR2 I553 (dt_0n[17], df_0n[17], gf1423_0n[17]);
  NOR3 I554 (df_0n[17], dt_0n[17], gt1424_0n[17], init_0n);
  AND2 I555 (gt1424_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I556 (gf1423_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I557 (wacks_0n[16], gf1423_0n[16], df_0n[16], gt1424_0n[16], dt_0n[16]);
  NOR2 I558 (dt_0n[16], df_0n[16], gf1423_0n[16]);
  NOR3 I559 (df_0n[16], dt_0n[16], gt1424_0n[16], init_0n);
  AND2 I560 (gt1424_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I561 (gf1423_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I562 (wacks_0n[15], gf1423_0n[15], df_0n[15], gt1424_0n[15], dt_0n[15]);
  NOR2 I563 (dt_0n[15], df_0n[15], gf1423_0n[15]);
  NOR3 I564 (df_0n[15], dt_0n[15], gt1424_0n[15], init_0n);
  AND2 I565 (gt1424_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I566 (gf1423_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I567 (wacks_0n[14], gf1423_0n[14], df_0n[14], gt1424_0n[14], dt_0n[14]);
  NOR2 I568 (dt_0n[14], df_0n[14], gf1423_0n[14]);
  NOR3 I569 (df_0n[14], dt_0n[14], gt1424_0n[14], init_0n);
  AND2 I570 (gt1424_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I571 (gf1423_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I572 (wacks_0n[13], gf1423_0n[13], df_0n[13], gt1424_0n[13], dt_0n[13]);
  NOR2 I573 (dt_0n[13], df_0n[13], gf1423_0n[13]);
  NOR3 I574 (df_0n[13], dt_0n[13], gt1424_0n[13], init_0n);
  AND2 I575 (gt1424_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I576 (gf1423_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I577 (wacks_0n[12], gf1423_0n[12], df_0n[12], gt1424_0n[12], dt_0n[12]);
  NOR2 I578 (dt_0n[12], df_0n[12], gf1423_0n[12]);
  NOR3 I579 (df_0n[12], dt_0n[12], gt1424_0n[12], init_0n);
  AND2 I580 (gt1424_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I581 (gf1423_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I582 (wacks_0n[11], gf1423_0n[11], df_0n[11], gt1424_0n[11], dt_0n[11]);
  NOR2 I583 (dt_0n[11], df_0n[11], gf1423_0n[11]);
  NOR3 I584 (df_0n[11], dt_0n[11], gt1424_0n[11], init_0n);
  AND2 I585 (gt1424_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I586 (gf1423_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I587 (wacks_0n[10], gf1423_0n[10], df_0n[10], gt1424_0n[10], dt_0n[10]);
  NOR2 I588 (dt_0n[10], df_0n[10], gf1423_0n[10]);
  NOR3 I589 (df_0n[10], dt_0n[10], gt1424_0n[10], init_0n);
  AND2 I590 (gt1424_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I591 (gf1423_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I592 (wacks_0n[9], gf1423_0n[9], df_0n[9], gt1424_0n[9], dt_0n[9]);
  NOR2 I593 (dt_0n[9], df_0n[9], gf1423_0n[9]);
  NOR3 I594 (df_0n[9], dt_0n[9], gt1424_0n[9], init_0n);
  AND2 I595 (gt1424_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I596 (gf1423_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I597 (wacks_0n[8], gf1423_0n[8], df_0n[8], gt1424_0n[8], dt_0n[8]);
  NOR2 I598 (dt_0n[8], df_0n[8], gf1423_0n[8]);
  NOR3 I599 (df_0n[8], dt_0n[8], gt1424_0n[8], init_0n);
  AND2 I600 (gt1424_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I601 (gf1423_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I602 (wacks_0n[7], gf1423_0n[7], df_0n[7], gt1424_0n[7], dt_0n[7]);
  NOR2 I603 (dt_0n[7], df_0n[7], gf1423_0n[7]);
  NOR3 I604 (df_0n[7], dt_0n[7], gt1424_0n[7], init_0n);
  AND2 I605 (gt1424_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I606 (gf1423_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I607 (wacks_0n[6], gf1423_0n[6], df_0n[6], gt1424_0n[6], dt_0n[6]);
  NOR2 I608 (dt_0n[6], df_0n[6], gf1423_0n[6]);
  NOR3 I609 (df_0n[6], dt_0n[6], gt1424_0n[6], init_0n);
  AND2 I610 (gt1424_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I611 (gf1423_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I612 (wacks_0n[5], gf1423_0n[5], df_0n[5], gt1424_0n[5], dt_0n[5]);
  NOR2 I613 (dt_0n[5], df_0n[5], gf1423_0n[5]);
  NOR3 I614 (df_0n[5], dt_0n[5], gt1424_0n[5], init_0n);
  AND2 I615 (gt1424_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I616 (gf1423_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I617 (wacks_0n[4], gf1423_0n[4], df_0n[4], gt1424_0n[4], dt_0n[4]);
  NOR2 I618 (dt_0n[4], df_0n[4], gf1423_0n[4]);
  NOR3 I619 (df_0n[4], dt_0n[4], gt1424_0n[4], init_0n);
  AND2 I620 (gt1424_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I621 (gf1423_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I622 (wacks_0n[3], gf1423_0n[3], df_0n[3], gt1424_0n[3], dt_0n[3]);
  NOR2 I623 (dt_0n[3], df_0n[3], gf1423_0n[3]);
  NOR3 I624 (df_0n[3], dt_0n[3], gt1424_0n[3], init_0n);
  AND2 I625 (gt1424_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I626 (gf1423_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I627 (wacks_0n[2], gf1423_0n[2], df_0n[2], gt1424_0n[2], dt_0n[2]);
  NOR2 I628 (dt_0n[2], df_0n[2], gf1423_0n[2]);
  NOR3 I629 (df_0n[2], dt_0n[2], gt1424_0n[2], init_0n);
  AND2 I630 (gt1424_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I631 (gf1423_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I632 (wacks_0n[1], gf1423_0n[1], df_0n[1], gt1424_0n[1], dt_0n[1]);
  NOR2 I633 (dt_0n[1], df_0n[1], gf1423_0n[1]);
  NOR3 I634 (df_0n[1], dt_0n[1], gt1424_0n[1], init_0n);
  AND2 I635 (gt1424_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I636 (gf1423_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I637 (wacks_0n[0], gf1423_0n[0], df_0n[0], gt1424_0n[0], dt_0n[0]);
  NOR2 I638 (dt_0n[0], df_0n[0], gf1423_0n[0]);
  NOR3 I639 (df_0n[0], dt_0n[0], gt1424_0n[0], init_0n);
  AND2 I640 (gt1424_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I641 (gf1423_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I642 (init_0n, initialise);
endmodule

module BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m88m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  initialise
);
  input [34:0] wg_0r0d;
  input [34:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [34:0] rd_0r0d;
  output [34:0] rd_0r1d;
  input rd_0a;
  output [1:0] rd_1r0d;
  output [1:0] rd_1r1d;
  input rd_1a;
  input initialise;
  wire [37:0] internal_0n;
  wire [34:0] wf_0n;
  wire [34:0] wt_0n;
  wire [34:0] df_0n;
  wire [34:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire wc_0n;
  wire [34:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [34:0] wgfint_0n;
  wire [34:0] wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire [34:0] rdfint_0n;
  wire [1:0] rdfint_1n;
  wire [34:0] rdtint_0n;
  wire [1:0] rdtint_1n;
  wire [34:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [34:0] gif_0n;
  wire [34:0] git_0n;
  wire [34:0] complete1436_0n;
  wire [34:0] gt1435_0n;
  wire [34:0] gf1434_0n;
  assign rgaint_1n = rd_1a;
  assign rd_1r0d[0] = rdfint_1n[0];
  assign rd_1r0d[1] = rdfint_1n[1];
  assign rd_1r1d[0] = rdtint_1n[0];
  assign rd_1r1d[1] = rdtint_1n[1];
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r0d[10] = rdfint_0n[10];
  assign rd_0r0d[11] = rdfint_0n[11];
  assign rd_0r0d[12] = rdfint_0n[12];
  assign rd_0r0d[13] = rdfint_0n[13];
  assign rd_0r0d[14] = rdfint_0n[14];
  assign rd_0r0d[15] = rdfint_0n[15];
  assign rd_0r0d[16] = rdfint_0n[16];
  assign rd_0r0d[17] = rdfint_0n[17];
  assign rd_0r0d[18] = rdfint_0n[18];
  assign rd_0r0d[19] = rdfint_0n[19];
  assign rd_0r0d[20] = rdfint_0n[20];
  assign rd_0r0d[21] = rdfint_0n[21];
  assign rd_0r0d[22] = rdfint_0n[22];
  assign rd_0r0d[23] = rdfint_0n[23];
  assign rd_0r0d[24] = rdfint_0n[24];
  assign rd_0r0d[25] = rdfint_0n[25];
  assign rd_0r0d[26] = rdfint_0n[26];
  assign rd_0r0d[27] = rdfint_0n[27];
  assign rd_0r0d[28] = rdfint_0n[28];
  assign rd_0r0d[29] = rdfint_0n[29];
  assign rd_0r0d[30] = rdfint_0n[30];
  assign rd_0r0d[31] = rdfint_0n[31];
  assign rd_0r0d[32] = rdfint_0n[32];
  assign rd_0r0d[33] = rdfint_0n[33];
  assign rd_0r0d[34] = rdfint_0n[34];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign rd_0r1d[10] = rdtint_0n[10];
  assign rd_0r1d[11] = rdtint_0n[11];
  assign rd_0r1d[12] = rdtint_0n[12];
  assign rd_0r1d[13] = rdtint_0n[13];
  assign rd_0r1d[14] = rdtint_0n[14];
  assign rd_0r1d[15] = rdtint_0n[15];
  assign rd_0r1d[16] = rdtint_0n[16];
  assign rd_0r1d[17] = rdtint_0n[17];
  assign rd_0r1d[18] = rdtint_0n[18];
  assign rd_0r1d[19] = rdtint_0n[19];
  assign rd_0r1d[20] = rdtint_0n[20];
  assign rd_0r1d[21] = rdtint_0n[21];
  assign rd_0r1d[22] = rdtint_0n[22];
  assign rd_0r1d[23] = rdtint_0n[23];
  assign rd_0r1d[24] = rdtint_0n[24];
  assign rd_0r1d[25] = rdtint_0n[25];
  assign rd_0r1d[26] = rdtint_0n[26];
  assign rd_0r1d[27] = rdtint_0n[27];
  assign rd_0r1d[28] = rdtint_0n[28];
  assign rd_0r1d[29] = rdtint_0n[29];
  assign rd_0r1d[30] = rdtint_0n[30];
  assign rd_0r1d[31] = rdtint_0n[31];
  assign rd_0r1d[32] = rdtint_0n[32];
  assign rd_0r1d[33] = rdtint_0n[33];
  assign rd_0r1d[34] = rdtint_0n[34];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgfint_0n[32] = wg_0r0d[32];
  assign wgfint_0n[33] = wg_0r0d[33];
  assign wgfint_0n[34] = wg_0r0d[34];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign wgtint_0n[32] = wg_0r1d[32];
  assign wgtint_0n[33] = wg_0r1d[33];
  assign wgtint_0n[34] = wg_0r1d[34];
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I153 (internal_0n[0], rgrint_0n, rgrint_1n);
  NOR2 I154 (internal_0n[1], rgaint_0n, rgaint_1n);
  AND2 I155 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I156 (rdtint_1n[0], rgrint_1n, dt_0n[0]);
  AND2 I157 (rdtint_1n[1], rgrint_1n, dt_0n[1]);
  AND2 I158 (rdtint_0n[0], rgrint_0n, dt_0n[0]);
  AND2 I159 (rdtint_0n[1], rgrint_0n, dt_0n[1]);
  AND2 I160 (rdtint_0n[2], rgrint_0n, dt_0n[2]);
  AND2 I161 (rdtint_0n[3], rgrint_0n, dt_0n[3]);
  AND2 I162 (rdtint_0n[4], rgrint_0n, dt_0n[4]);
  AND2 I163 (rdtint_0n[5], rgrint_0n, dt_0n[5]);
  AND2 I164 (rdtint_0n[6], rgrint_0n, dt_0n[6]);
  AND2 I165 (rdtint_0n[7], rgrint_0n, dt_0n[7]);
  AND2 I166 (rdtint_0n[8], rgrint_0n, dt_0n[8]);
  AND2 I167 (rdtint_0n[9], rgrint_0n, dt_0n[9]);
  AND2 I168 (rdtint_0n[10], rgrint_0n, dt_0n[10]);
  AND2 I169 (rdtint_0n[11], rgrint_0n, dt_0n[11]);
  AND2 I170 (rdtint_0n[12], rgrint_0n, dt_0n[12]);
  AND2 I171 (rdtint_0n[13], rgrint_0n, dt_0n[13]);
  AND2 I172 (rdtint_0n[14], rgrint_0n, dt_0n[14]);
  AND2 I173 (rdtint_0n[15], rgrint_0n, dt_0n[15]);
  AND2 I174 (rdtint_0n[16], rgrint_0n, dt_0n[16]);
  AND2 I175 (rdtint_0n[17], rgrint_0n, dt_0n[17]);
  AND2 I176 (rdtint_0n[18], rgrint_0n, dt_0n[18]);
  AND2 I177 (rdtint_0n[19], rgrint_0n, dt_0n[19]);
  AND2 I178 (rdtint_0n[20], rgrint_0n, dt_0n[20]);
  AND2 I179 (rdtint_0n[21], rgrint_0n, dt_0n[21]);
  AND2 I180 (rdtint_0n[22], rgrint_0n, dt_0n[22]);
  AND2 I181 (rdtint_0n[23], rgrint_0n, dt_0n[23]);
  AND2 I182 (rdtint_0n[24], rgrint_0n, dt_0n[24]);
  AND2 I183 (rdtint_0n[25], rgrint_0n, dt_0n[25]);
  AND2 I184 (rdtint_0n[26], rgrint_0n, dt_0n[26]);
  AND2 I185 (rdtint_0n[27], rgrint_0n, dt_0n[27]);
  AND2 I186 (rdtint_0n[28], rgrint_0n, dt_0n[28]);
  AND2 I187 (rdtint_0n[29], rgrint_0n, dt_0n[29]);
  AND2 I188 (rdtint_0n[30], rgrint_0n, dt_0n[30]);
  AND2 I189 (rdtint_0n[31], rgrint_0n, dt_0n[31]);
  AND2 I190 (rdtint_0n[32], rgrint_0n, dt_0n[32]);
  AND2 I191 (rdtint_0n[33], rgrint_0n, dt_0n[33]);
  AND2 I192 (rdtint_0n[34], rgrint_0n, dt_0n[34]);
  AND2 I193 (rdfint_1n[0], rgrint_1n, df_0n[0]);
  AND2 I194 (rdfint_1n[1], rgrint_1n, df_0n[1]);
  AND2 I195 (rdfint_0n[0], rgrint_0n, df_0n[0]);
  AND2 I196 (rdfint_0n[1], rgrint_0n, df_0n[1]);
  AND2 I197 (rdfint_0n[2], rgrint_0n, df_0n[2]);
  AND2 I198 (rdfint_0n[3], rgrint_0n, df_0n[3]);
  AND2 I199 (rdfint_0n[4], rgrint_0n, df_0n[4]);
  AND2 I200 (rdfint_0n[5], rgrint_0n, df_0n[5]);
  AND2 I201 (rdfint_0n[6], rgrint_0n, df_0n[6]);
  AND2 I202 (rdfint_0n[7], rgrint_0n, df_0n[7]);
  AND2 I203 (rdfint_0n[8], rgrint_0n, df_0n[8]);
  AND2 I204 (rdfint_0n[9], rgrint_0n, df_0n[9]);
  AND2 I205 (rdfint_0n[10], rgrint_0n, df_0n[10]);
  AND2 I206 (rdfint_0n[11], rgrint_0n, df_0n[11]);
  AND2 I207 (rdfint_0n[12], rgrint_0n, df_0n[12]);
  AND2 I208 (rdfint_0n[13], rgrint_0n, df_0n[13]);
  AND2 I209 (rdfint_0n[14], rgrint_0n, df_0n[14]);
  AND2 I210 (rdfint_0n[15], rgrint_0n, df_0n[15]);
  AND2 I211 (rdfint_0n[16], rgrint_0n, df_0n[16]);
  AND2 I212 (rdfint_0n[17], rgrint_0n, df_0n[17]);
  AND2 I213 (rdfint_0n[18], rgrint_0n, df_0n[18]);
  AND2 I214 (rdfint_0n[19], rgrint_0n, df_0n[19]);
  AND2 I215 (rdfint_0n[20], rgrint_0n, df_0n[20]);
  AND2 I216 (rdfint_0n[21], rgrint_0n, df_0n[21]);
  AND2 I217 (rdfint_0n[22], rgrint_0n, df_0n[22]);
  AND2 I218 (rdfint_0n[23], rgrint_0n, df_0n[23]);
  AND2 I219 (rdfint_0n[24], rgrint_0n, df_0n[24]);
  AND2 I220 (rdfint_0n[25], rgrint_0n, df_0n[25]);
  AND2 I221 (rdfint_0n[26], rgrint_0n, df_0n[26]);
  AND2 I222 (rdfint_0n[27], rgrint_0n, df_0n[27]);
  AND2 I223 (rdfint_0n[28], rgrint_0n, df_0n[28]);
  AND2 I224 (rdfint_0n[29], rgrint_0n, df_0n[29]);
  AND2 I225 (rdfint_0n[30], rgrint_0n, df_0n[30]);
  AND2 I226 (rdfint_0n[31], rgrint_0n, df_0n[31]);
  AND2 I227 (rdfint_0n[32], rgrint_0n, df_0n[32]);
  AND2 I228 (rdfint_0n[33], rgrint_0n, df_0n[33]);
  AND2 I229 (rdfint_0n[34], rgrint_0n, df_0n[34]);
  C3 I230 (internal_0n[2], wc_0n, wacks_0n[34], wacks_0n[33]);
  C3 I231 (internal_0n[3], wacks_0n[32], wacks_0n[31], wacks_0n[30]);
  C3 I232 (internal_0n[4], wacks_0n[29], wacks_0n[28], wacks_0n[27]);
  C3 I233 (internal_0n[5], wacks_0n[26], wacks_0n[25], wacks_0n[24]);
  C3 I234 (internal_0n[6], wacks_0n[23], wacks_0n[22], wacks_0n[21]);
  C3 I235 (internal_0n[7], wacks_0n[20], wacks_0n[19], wacks_0n[18]);
  C3 I236 (internal_0n[8], wacks_0n[17], wacks_0n[16], wacks_0n[15]);
  C3 I237 (internal_0n[9], wacks_0n[14], wacks_0n[13], wacks_0n[12]);
  C3 I238 (internal_0n[10], wacks_0n[11], wacks_0n[10], wacks_0n[9]);
  C3 I239 (internal_0n[11], wacks_0n[8], wacks_0n[7], wacks_0n[6]);
  C3 I240 (internal_0n[12], wacks_0n[5], wacks_0n[4], wacks_0n[3]);
  C3 I241 (internal_0n[13], wacks_0n[2], wacks_0n[1], wacks_0n[0]);
  C3 I242 (internal_0n[14], internal_0n[2], internal_0n[3], internal_0n[4]);
  C3 I243 (internal_0n[15], internal_0n[5], internal_0n[6], internal_0n[7]);
  C3 I244 (internal_0n[16], internal_0n[8], internal_0n[9], internal_0n[10]);
  C3 I245 (internal_0n[17], internal_0n[11], internal_0n[12], internal_0n[13]);
  C2 I246 (internal_0n[18], internal_0n[14], internal_0n[15]);
  C2 I247 (internal_0n[19], internal_0n[16], internal_0n[17]);
  C2 I248 (wdrint_0n, internal_0n[18], internal_0n[19]);
  assign wen_0n[34] = wc_0n;
  assign wen_0n[33] = wc_0n;
  assign wen_0n[32] = wc_0n;
  assign wen_0n[31] = wc_0n;
  assign wen_0n[30] = wc_0n;
  assign wen_0n[29] = wc_0n;
  assign wen_0n[28] = wc_0n;
  assign wen_0n[27] = wc_0n;
  assign wen_0n[26] = wc_0n;
  assign wen_0n[25] = wc_0n;
  assign wen_0n[24] = wc_0n;
  assign wen_0n[23] = wc_0n;
  assign wen_0n[22] = wc_0n;
  assign wen_0n[21] = wc_0n;
  assign wen_0n[20] = wc_0n;
  assign wen_0n[19] = wc_0n;
  assign wen_0n[18] = wc_0n;
  assign wen_0n[17] = wc_0n;
  assign wen_0n[16] = wc_0n;
  assign wen_0n[15] = wc_0n;
  assign wen_0n[14] = wc_0n;
  assign wen_0n[13] = wc_0n;
  assign wen_0n[12] = wc_0n;
  assign wen_0n[11] = wc_0n;
  assign wen_0n[10] = wc_0n;
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[34] = git_0n[34];
  assign wt_0n[33] = git_0n[33];
  assign wt_0n[32] = git_0n[32];
  assign wt_0n[31] = git_0n[31];
  assign wt_0n[30] = git_0n[30];
  assign wt_0n[29] = git_0n[29];
  assign wt_0n[28] = git_0n[28];
  assign wt_0n[27] = git_0n[27];
  assign wt_0n[26] = git_0n[26];
  assign wt_0n[25] = git_0n[25];
  assign wt_0n[24] = git_0n[24];
  assign wt_0n[23] = git_0n[23];
  assign wt_0n[22] = git_0n[22];
  assign wt_0n[21] = git_0n[21];
  assign wt_0n[20] = git_0n[20];
  assign wt_0n[19] = git_0n[19];
  assign wt_0n[18] = git_0n[18];
  assign wt_0n[17] = git_0n[17];
  assign wt_0n[16] = git_0n[16];
  assign wt_0n[15] = git_0n[15];
  assign wt_0n[14] = git_0n[14];
  assign wt_0n[13] = git_0n[13];
  assign wt_0n[12] = git_0n[12];
  assign wt_0n[11] = git_0n[11];
  assign wt_0n[10] = git_0n[10];
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[34] = gif_0n[34];
  assign wf_0n[33] = gif_0n[33];
  assign wf_0n[32] = gif_0n[32];
  assign wf_0n[31] = gif_0n[31];
  assign wf_0n[30] = gif_0n[30];
  assign wf_0n[29] = gif_0n[29];
  assign wf_0n[28] = gif_0n[28];
  assign wf_0n[27] = gif_0n[27];
  assign wf_0n[26] = gif_0n[26];
  assign wf_0n[25] = gif_0n[25];
  assign wf_0n[24] = gif_0n[24];
  assign wf_0n[23] = gif_0n[23];
  assign wf_0n[22] = gif_0n[22];
  assign wf_0n[21] = gif_0n[21];
  assign wf_0n[20] = gif_0n[20];
  assign wf_0n[19] = gif_0n[19];
  assign wf_0n[18] = gif_0n[18];
  assign wf_0n[17] = gif_0n[17];
  assign wf_0n[16] = gif_0n[16];
  assign wf_0n[15] = gif_0n[15];
  assign wf_0n[14] = gif_0n[14];
  assign wf_0n[13] = gif_0n[13];
  assign wf_0n[12] = gif_0n[12];
  assign wf_0n[11] = gif_0n[11];
  assign wf_0n[10] = gif_0n[10];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I354 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I356 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I357 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I358 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I359 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I360 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I361 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I362 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I363 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I364 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I365 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I366 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I367 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I368 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I369 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I370 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I371 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I372 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I373 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I374 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I375 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I376 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I377 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I378 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I379 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I380 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I381 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I382 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I383 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I384 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I385 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I386 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I387 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I388 (git_0n[32], wgtint_0n[32], ig_0n);
  AND2 I389 (git_0n[33], wgtint_0n[33], ig_0n);
  AND2 I390 (git_0n[34], wgtint_0n[34], ig_0n);
  AND2 I391 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I392 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I393 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I394 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I395 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I396 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I397 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I398 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I399 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I400 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I401 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I402 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I403 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I404 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I405 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I406 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I407 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I408 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I409 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I410 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I411 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I412 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I413 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I414 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I415 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I416 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I417 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I418 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I419 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I420 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I421 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I422 (gif_0n[31], wgfint_0n[31], ig_0n);
  AND2 I423 (gif_0n[32], wgfint_0n[32], ig_0n);
  AND2 I424 (gif_0n[33], wgfint_0n[33], ig_0n);
  AND2 I425 (gif_0n[34], wgfint_0n[34], ig_0n);
  C3 I426 (internal_0n[20], complete1436_0n[0], complete1436_0n[1], complete1436_0n[2]);
  C3 I427 (internal_0n[21], complete1436_0n[3], complete1436_0n[4], complete1436_0n[5]);
  C3 I428 (internal_0n[22], complete1436_0n[6], complete1436_0n[7], complete1436_0n[8]);
  C3 I429 (internal_0n[23], complete1436_0n[9], complete1436_0n[10], complete1436_0n[11]);
  C3 I430 (internal_0n[24], complete1436_0n[12], complete1436_0n[13], complete1436_0n[14]);
  C3 I431 (internal_0n[25], complete1436_0n[15], complete1436_0n[16], complete1436_0n[17]);
  C3 I432 (internal_0n[26], complete1436_0n[18], complete1436_0n[19], complete1436_0n[20]);
  C3 I433 (internal_0n[27], complete1436_0n[21], complete1436_0n[22], complete1436_0n[23]);
  C3 I434 (internal_0n[28], complete1436_0n[24], complete1436_0n[25], complete1436_0n[26]);
  C3 I435 (internal_0n[29], complete1436_0n[27], complete1436_0n[28], complete1436_0n[29]);
  C3 I436 (internal_0n[30], complete1436_0n[30], complete1436_0n[31], complete1436_0n[32]);
  C2 I437 (internal_0n[31], complete1436_0n[33], complete1436_0n[34]);
  C3 I438 (internal_0n[32], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I439 (internal_0n[33], internal_0n[23], internal_0n[24], internal_0n[25]);
  C3 I440 (internal_0n[34], internal_0n[26], internal_0n[27], internal_0n[28]);
  C3 I441 (internal_0n[35], internal_0n[29], internal_0n[30], internal_0n[31]);
  C2 I442 (internal_0n[36], internal_0n[32], internal_0n[33]);
  C2 I443 (internal_0n[37], internal_0n[34], internal_0n[35]);
  C2 I444 (wc_0n, internal_0n[36], internal_0n[37]);
  OR2 I445 (complete1436_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I446 (complete1436_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I447 (complete1436_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I448 (complete1436_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I449 (complete1436_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I450 (complete1436_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I451 (complete1436_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I452 (complete1436_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I453 (complete1436_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I454 (complete1436_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I455 (complete1436_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I456 (complete1436_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I457 (complete1436_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I458 (complete1436_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I459 (complete1436_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I460 (complete1436_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I461 (complete1436_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I462 (complete1436_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I463 (complete1436_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I464 (complete1436_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I465 (complete1436_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I466 (complete1436_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I467 (complete1436_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I468 (complete1436_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I469 (complete1436_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I470 (complete1436_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I471 (complete1436_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I472 (complete1436_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I473 (complete1436_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I474 (complete1436_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I475 (complete1436_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I476 (complete1436_0n[31], wgfint_0n[31], wgtint_0n[31]);
  OR2 I477 (complete1436_0n[32], wgfint_0n[32], wgtint_0n[32]);
  OR2 I478 (complete1436_0n[33], wgfint_0n[33], wgtint_0n[33]);
  OR2 I479 (complete1436_0n[34], wgfint_0n[34], wgtint_0n[34]);
  AO22 I480 (wacks_0n[34], gf1434_0n[34], df_0n[34], gt1435_0n[34], dt_0n[34]);
  NOR2 I481 (dt_0n[34], df_0n[34], gf1434_0n[34]);
  NOR3 I482 (df_0n[34], dt_0n[34], gt1435_0n[34], init_0n);
  AND2 I483 (gt1435_0n[34], wt_0n[34], wen_0n[34]);
  AND2 I484 (gf1434_0n[34], wf_0n[34], wen_0n[34]);
  AO22 I485 (wacks_0n[33], gf1434_0n[33], df_0n[33], gt1435_0n[33], dt_0n[33]);
  NOR2 I486 (dt_0n[33], df_0n[33], gf1434_0n[33]);
  NOR3 I487 (df_0n[33], dt_0n[33], gt1435_0n[33], init_0n);
  AND2 I488 (gt1435_0n[33], wt_0n[33], wen_0n[33]);
  AND2 I489 (gf1434_0n[33], wf_0n[33], wen_0n[33]);
  AO22 I490 (wacks_0n[32], gf1434_0n[32], df_0n[32], gt1435_0n[32], dt_0n[32]);
  NOR2 I491 (dt_0n[32], df_0n[32], gf1434_0n[32]);
  NOR3 I492 (df_0n[32], dt_0n[32], gt1435_0n[32], init_0n);
  AND2 I493 (gt1435_0n[32], wt_0n[32], wen_0n[32]);
  AND2 I494 (gf1434_0n[32], wf_0n[32], wen_0n[32]);
  AO22 I495 (wacks_0n[31], gf1434_0n[31], df_0n[31], gt1435_0n[31], dt_0n[31]);
  NOR2 I496 (dt_0n[31], df_0n[31], gf1434_0n[31]);
  NOR3 I497 (df_0n[31], dt_0n[31], gt1435_0n[31], init_0n);
  AND2 I498 (gt1435_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I499 (gf1434_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I500 (wacks_0n[30], gf1434_0n[30], df_0n[30], gt1435_0n[30], dt_0n[30]);
  NOR2 I501 (dt_0n[30], df_0n[30], gf1434_0n[30]);
  NOR3 I502 (df_0n[30], dt_0n[30], gt1435_0n[30], init_0n);
  AND2 I503 (gt1435_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I504 (gf1434_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I505 (wacks_0n[29], gf1434_0n[29], df_0n[29], gt1435_0n[29], dt_0n[29]);
  NOR2 I506 (dt_0n[29], df_0n[29], gf1434_0n[29]);
  NOR3 I507 (df_0n[29], dt_0n[29], gt1435_0n[29], init_0n);
  AND2 I508 (gt1435_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I509 (gf1434_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I510 (wacks_0n[28], gf1434_0n[28], df_0n[28], gt1435_0n[28], dt_0n[28]);
  NOR2 I511 (dt_0n[28], df_0n[28], gf1434_0n[28]);
  NOR3 I512 (df_0n[28], dt_0n[28], gt1435_0n[28], init_0n);
  AND2 I513 (gt1435_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I514 (gf1434_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I515 (wacks_0n[27], gf1434_0n[27], df_0n[27], gt1435_0n[27], dt_0n[27]);
  NOR2 I516 (dt_0n[27], df_0n[27], gf1434_0n[27]);
  NOR3 I517 (df_0n[27], dt_0n[27], gt1435_0n[27], init_0n);
  AND2 I518 (gt1435_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I519 (gf1434_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I520 (wacks_0n[26], gf1434_0n[26], df_0n[26], gt1435_0n[26], dt_0n[26]);
  NOR2 I521 (dt_0n[26], df_0n[26], gf1434_0n[26]);
  NOR3 I522 (df_0n[26], dt_0n[26], gt1435_0n[26], init_0n);
  AND2 I523 (gt1435_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I524 (gf1434_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I525 (wacks_0n[25], gf1434_0n[25], df_0n[25], gt1435_0n[25], dt_0n[25]);
  NOR2 I526 (dt_0n[25], df_0n[25], gf1434_0n[25]);
  NOR3 I527 (df_0n[25], dt_0n[25], gt1435_0n[25], init_0n);
  AND2 I528 (gt1435_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I529 (gf1434_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I530 (wacks_0n[24], gf1434_0n[24], df_0n[24], gt1435_0n[24], dt_0n[24]);
  NOR2 I531 (dt_0n[24], df_0n[24], gf1434_0n[24]);
  NOR3 I532 (df_0n[24], dt_0n[24], gt1435_0n[24], init_0n);
  AND2 I533 (gt1435_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I534 (gf1434_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I535 (wacks_0n[23], gf1434_0n[23], df_0n[23], gt1435_0n[23], dt_0n[23]);
  NOR2 I536 (dt_0n[23], df_0n[23], gf1434_0n[23]);
  NOR3 I537 (df_0n[23], dt_0n[23], gt1435_0n[23], init_0n);
  AND2 I538 (gt1435_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I539 (gf1434_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I540 (wacks_0n[22], gf1434_0n[22], df_0n[22], gt1435_0n[22], dt_0n[22]);
  NOR2 I541 (dt_0n[22], df_0n[22], gf1434_0n[22]);
  NOR3 I542 (df_0n[22], dt_0n[22], gt1435_0n[22], init_0n);
  AND2 I543 (gt1435_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I544 (gf1434_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I545 (wacks_0n[21], gf1434_0n[21], df_0n[21], gt1435_0n[21], dt_0n[21]);
  NOR2 I546 (dt_0n[21], df_0n[21], gf1434_0n[21]);
  NOR3 I547 (df_0n[21], dt_0n[21], gt1435_0n[21], init_0n);
  AND2 I548 (gt1435_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I549 (gf1434_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I550 (wacks_0n[20], gf1434_0n[20], df_0n[20], gt1435_0n[20], dt_0n[20]);
  NOR2 I551 (dt_0n[20], df_0n[20], gf1434_0n[20]);
  NOR3 I552 (df_0n[20], dt_0n[20], gt1435_0n[20], init_0n);
  AND2 I553 (gt1435_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I554 (gf1434_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I555 (wacks_0n[19], gf1434_0n[19], df_0n[19], gt1435_0n[19], dt_0n[19]);
  NOR2 I556 (dt_0n[19], df_0n[19], gf1434_0n[19]);
  NOR3 I557 (df_0n[19], dt_0n[19], gt1435_0n[19], init_0n);
  AND2 I558 (gt1435_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I559 (gf1434_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I560 (wacks_0n[18], gf1434_0n[18], df_0n[18], gt1435_0n[18], dt_0n[18]);
  NOR2 I561 (dt_0n[18], df_0n[18], gf1434_0n[18]);
  NOR3 I562 (df_0n[18], dt_0n[18], gt1435_0n[18], init_0n);
  AND2 I563 (gt1435_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I564 (gf1434_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I565 (wacks_0n[17], gf1434_0n[17], df_0n[17], gt1435_0n[17], dt_0n[17]);
  NOR2 I566 (dt_0n[17], df_0n[17], gf1434_0n[17]);
  NOR3 I567 (df_0n[17], dt_0n[17], gt1435_0n[17], init_0n);
  AND2 I568 (gt1435_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I569 (gf1434_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I570 (wacks_0n[16], gf1434_0n[16], df_0n[16], gt1435_0n[16], dt_0n[16]);
  NOR2 I571 (dt_0n[16], df_0n[16], gf1434_0n[16]);
  NOR3 I572 (df_0n[16], dt_0n[16], gt1435_0n[16], init_0n);
  AND2 I573 (gt1435_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I574 (gf1434_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I575 (wacks_0n[15], gf1434_0n[15], df_0n[15], gt1435_0n[15], dt_0n[15]);
  NOR2 I576 (dt_0n[15], df_0n[15], gf1434_0n[15]);
  NOR3 I577 (df_0n[15], dt_0n[15], gt1435_0n[15], init_0n);
  AND2 I578 (gt1435_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I579 (gf1434_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I580 (wacks_0n[14], gf1434_0n[14], df_0n[14], gt1435_0n[14], dt_0n[14]);
  NOR2 I581 (dt_0n[14], df_0n[14], gf1434_0n[14]);
  NOR3 I582 (df_0n[14], dt_0n[14], gt1435_0n[14], init_0n);
  AND2 I583 (gt1435_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I584 (gf1434_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I585 (wacks_0n[13], gf1434_0n[13], df_0n[13], gt1435_0n[13], dt_0n[13]);
  NOR2 I586 (dt_0n[13], df_0n[13], gf1434_0n[13]);
  NOR3 I587 (df_0n[13], dt_0n[13], gt1435_0n[13], init_0n);
  AND2 I588 (gt1435_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I589 (gf1434_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I590 (wacks_0n[12], gf1434_0n[12], df_0n[12], gt1435_0n[12], dt_0n[12]);
  NOR2 I591 (dt_0n[12], df_0n[12], gf1434_0n[12]);
  NOR3 I592 (df_0n[12], dt_0n[12], gt1435_0n[12], init_0n);
  AND2 I593 (gt1435_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I594 (gf1434_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I595 (wacks_0n[11], gf1434_0n[11], df_0n[11], gt1435_0n[11], dt_0n[11]);
  NOR2 I596 (dt_0n[11], df_0n[11], gf1434_0n[11]);
  NOR3 I597 (df_0n[11], dt_0n[11], gt1435_0n[11], init_0n);
  AND2 I598 (gt1435_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I599 (gf1434_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I600 (wacks_0n[10], gf1434_0n[10], df_0n[10], gt1435_0n[10], dt_0n[10]);
  NOR2 I601 (dt_0n[10], df_0n[10], gf1434_0n[10]);
  NOR3 I602 (df_0n[10], dt_0n[10], gt1435_0n[10], init_0n);
  AND2 I603 (gt1435_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I604 (gf1434_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I605 (wacks_0n[9], gf1434_0n[9], df_0n[9], gt1435_0n[9], dt_0n[9]);
  NOR2 I606 (dt_0n[9], df_0n[9], gf1434_0n[9]);
  NOR3 I607 (df_0n[9], dt_0n[9], gt1435_0n[9], init_0n);
  AND2 I608 (gt1435_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I609 (gf1434_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I610 (wacks_0n[8], gf1434_0n[8], df_0n[8], gt1435_0n[8], dt_0n[8]);
  NOR2 I611 (dt_0n[8], df_0n[8], gf1434_0n[8]);
  NOR3 I612 (df_0n[8], dt_0n[8], gt1435_0n[8], init_0n);
  AND2 I613 (gt1435_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I614 (gf1434_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I615 (wacks_0n[7], gf1434_0n[7], df_0n[7], gt1435_0n[7], dt_0n[7]);
  NOR2 I616 (dt_0n[7], df_0n[7], gf1434_0n[7]);
  NOR3 I617 (df_0n[7], dt_0n[7], gt1435_0n[7], init_0n);
  AND2 I618 (gt1435_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I619 (gf1434_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I620 (wacks_0n[6], gf1434_0n[6], df_0n[6], gt1435_0n[6], dt_0n[6]);
  NOR2 I621 (dt_0n[6], df_0n[6], gf1434_0n[6]);
  NOR3 I622 (df_0n[6], dt_0n[6], gt1435_0n[6], init_0n);
  AND2 I623 (gt1435_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I624 (gf1434_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I625 (wacks_0n[5], gf1434_0n[5], df_0n[5], gt1435_0n[5], dt_0n[5]);
  NOR2 I626 (dt_0n[5], df_0n[5], gf1434_0n[5]);
  NOR3 I627 (df_0n[5], dt_0n[5], gt1435_0n[5], init_0n);
  AND2 I628 (gt1435_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I629 (gf1434_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I630 (wacks_0n[4], gf1434_0n[4], df_0n[4], gt1435_0n[4], dt_0n[4]);
  NOR2 I631 (dt_0n[4], df_0n[4], gf1434_0n[4]);
  NOR3 I632 (df_0n[4], dt_0n[4], gt1435_0n[4], init_0n);
  AND2 I633 (gt1435_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I634 (gf1434_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I635 (wacks_0n[3], gf1434_0n[3], df_0n[3], gt1435_0n[3], dt_0n[3]);
  NOR2 I636 (dt_0n[3], df_0n[3], gf1434_0n[3]);
  NOR3 I637 (df_0n[3], dt_0n[3], gt1435_0n[3], init_0n);
  AND2 I638 (gt1435_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I639 (gf1434_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I640 (wacks_0n[2], gf1434_0n[2], df_0n[2], gt1435_0n[2], dt_0n[2]);
  NOR2 I641 (dt_0n[2], df_0n[2], gf1434_0n[2]);
  NOR3 I642 (df_0n[2], dt_0n[2], gt1435_0n[2], init_0n);
  AND2 I643 (gt1435_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I644 (gf1434_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I645 (wacks_0n[1], gf1434_0n[1], df_0n[1], gt1435_0n[1], dt_0n[1]);
  NOR2 I646 (dt_0n[1], df_0n[1], gf1434_0n[1]);
  NOR3 I647 (df_0n[1], dt_0n[1], gt1435_0n[1], init_0n);
  AND2 I648 (gt1435_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I649 (gf1434_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I650 (wacks_0n[0], gf1434_0n[0], df_0n[0], gt1435_0n[0], dt_0n[0]);
  NOR2 I651 (dt_0n[0], df_0n[0], gf1434_0n[0]);
  NOR3 I652 (df_0n[0], dt_0n[0], gt1435_0n[0], init_0n);
  AND2 I653 (gt1435_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I654 (gf1434_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I655 (init_0n, initialise);
endmodule

module BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m89m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rg_2r, rg_2a,
  rg_3r, rg_3a,
  rg_4r, rg_4a,
  rg_5r, rg_5a,
  rg_6r, rg_6a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  rd_2r0d, rd_2r1d, rd_2a,
  rd_3r0d, rd_3r1d, rd_3a,
  rd_4r0d, rd_4r1d, rd_4a,
  rd_5r0d, rd_5r1d, rd_5a,
  rd_6r0d, rd_6r1d, rd_6a,
  initialise
);
  input [34:0] wg_0r0d;
  input [34:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  input rg_5r;
  output rg_5a;
  input rg_6r;
  output rg_6a;
  output [34:0] rd_0r0d;
  output [34:0] rd_0r1d;
  input rd_0a;
  output [33:0] rd_1r0d;
  output [33:0] rd_1r1d;
  input rd_1a;
  output [32:0] rd_2r0d;
  output [32:0] rd_2r1d;
  input rd_2a;
  output [31:0] rd_3r0d;
  output [31:0] rd_3r1d;
  input rd_3a;
  output [31:0] rd_4r0d;
  output [31:0] rd_4r1d;
  input rd_4a;
  output rd_5r0d;
  output rd_5r1d;
  input rd_5a;
  output rd_6r0d;
  output rd_6r1d;
  input rd_6a;
  input initialise;
  wire [42:0] internal_0n;
  wire [34:0] wf_0n;
  wire [34:0] wt_0n;
  wire [34:0] df_0n;
  wire [34:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire rgrint_2n;
  wire rgrint_3n;
  wire rgrint_4n;
  wire rgrint_5n;
  wire rgrint_6n;
  wire wc_0n;
  wire [34:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [34:0] wgfint_0n;
  wire [34:0] wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire rgaint_2n;
  wire rgaint_3n;
  wire rgaint_4n;
  wire rgaint_5n;
  wire rgaint_6n;
  wire [34:0] rdfint_0n;
  wire [33:0] rdfint_1n;
  wire [32:0] rdfint_2n;
  wire [31:0] rdfint_3n;
  wire [31:0] rdfint_4n;
  wire rdfint_5n;
  wire rdfint_6n;
  wire [34:0] rdtint_0n;
  wire [33:0] rdtint_1n;
  wire [32:0] rdtint_2n;
  wire [31:0] rdtint_3n;
  wire [31:0] rdtint_4n;
  wire rdtint_5n;
  wire rdtint_6n;
  wire [34:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [34:0] gif_0n;
  wire [34:0] git_0n;
  wire [34:0] complete1451_0n;
  wire [34:0] gt1450_0n;
  wire [34:0] gf1449_0n;
  assign rgaint_6n = rd_6a;
  assign rd_6r0d = rdfint_6n;
  assign rd_6r1d = rdtint_6n;
  assign rgaint_5n = rd_5a;
  assign rd_5r0d = rdfint_5n;
  assign rd_5r1d = rdtint_5n;
  assign rgaint_4n = rd_4a;
  assign rd_4r0d[0] = rdfint_4n[0];
  assign rd_4r0d[1] = rdfint_4n[1];
  assign rd_4r0d[2] = rdfint_4n[2];
  assign rd_4r0d[3] = rdfint_4n[3];
  assign rd_4r0d[4] = rdfint_4n[4];
  assign rd_4r0d[5] = rdfint_4n[5];
  assign rd_4r0d[6] = rdfint_4n[6];
  assign rd_4r0d[7] = rdfint_4n[7];
  assign rd_4r0d[8] = rdfint_4n[8];
  assign rd_4r0d[9] = rdfint_4n[9];
  assign rd_4r0d[10] = rdfint_4n[10];
  assign rd_4r0d[11] = rdfint_4n[11];
  assign rd_4r0d[12] = rdfint_4n[12];
  assign rd_4r0d[13] = rdfint_4n[13];
  assign rd_4r0d[14] = rdfint_4n[14];
  assign rd_4r0d[15] = rdfint_4n[15];
  assign rd_4r0d[16] = rdfint_4n[16];
  assign rd_4r0d[17] = rdfint_4n[17];
  assign rd_4r0d[18] = rdfint_4n[18];
  assign rd_4r0d[19] = rdfint_4n[19];
  assign rd_4r0d[20] = rdfint_4n[20];
  assign rd_4r0d[21] = rdfint_4n[21];
  assign rd_4r0d[22] = rdfint_4n[22];
  assign rd_4r0d[23] = rdfint_4n[23];
  assign rd_4r0d[24] = rdfint_4n[24];
  assign rd_4r0d[25] = rdfint_4n[25];
  assign rd_4r0d[26] = rdfint_4n[26];
  assign rd_4r0d[27] = rdfint_4n[27];
  assign rd_4r0d[28] = rdfint_4n[28];
  assign rd_4r0d[29] = rdfint_4n[29];
  assign rd_4r0d[30] = rdfint_4n[30];
  assign rd_4r0d[31] = rdfint_4n[31];
  assign rd_4r1d[0] = rdtint_4n[0];
  assign rd_4r1d[1] = rdtint_4n[1];
  assign rd_4r1d[2] = rdtint_4n[2];
  assign rd_4r1d[3] = rdtint_4n[3];
  assign rd_4r1d[4] = rdtint_4n[4];
  assign rd_4r1d[5] = rdtint_4n[5];
  assign rd_4r1d[6] = rdtint_4n[6];
  assign rd_4r1d[7] = rdtint_4n[7];
  assign rd_4r1d[8] = rdtint_4n[8];
  assign rd_4r1d[9] = rdtint_4n[9];
  assign rd_4r1d[10] = rdtint_4n[10];
  assign rd_4r1d[11] = rdtint_4n[11];
  assign rd_4r1d[12] = rdtint_4n[12];
  assign rd_4r1d[13] = rdtint_4n[13];
  assign rd_4r1d[14] = rdtint_4n[14];
  assign rd_4r1d[15] = rdtint_4n[15];
  assign rd_4r1d[16] = rdtint_4n[16];
  assign rd_4r1d[17] = rdtint_4n[17];
  assign rd_4r1d[18] = rdtint_4n[18];
  assign rd_4r1d[19] = rdtint_4n[19];
  assign rd_4r1d[20] = rdtint_4n[20];
  assign rd_4r1d[21] = rdtint_4n[21];
  assign rd_4r1d[22] = rdtint_4n[22];
  assign rd_4r1d[23] = rdtint_4n[23];
  assign rd_4r1d[24] = rdtint_4n[24];
  assign rd_4r1d[25] = rdtint_4n[25];
  assign rd_4r1d[26] = rdtint_4n[26];
  assign rd_4r1d[27] = rdtint_4n[27];
  assign rd_4r1d[28] = rdtint_4n[28];
  assign rd_4r1d[29] = rdtint_4n[29];
  assign rd_4r1d[30] = rdtint_4n[30];
  assign rd_4r1d[31] = rdtint_4n[31];
  assign rgaint_3n = rd_3a;
  assign rd_3r0d[0] = rdfint_3n[0];
  assign rd_3r0d[1] = rdfint_3n[1];
  assign rd_3r0d[2] = rdfint_3n[2];
  assign rd_3r0d[3] = rdfint_3n[3];
  assign rd_3r0d[4] = rdfint_3n[4];
  assign rd_3r0d[5] = rdfint_3n[5];
  assign rd_3r0d[6] = rdfint_3n[6];
  assign rd_3r0d[7] = rdfint_3n[7];
  assign rd_3r0d[8] = rdfint_3n[8];
  assign rd_3r0d[9] = rdfint_3n[9];
  assign rd_3r0d[10] = rdfint_3n[10];
  assign rd_3r0d[11] = rdfint_3n[11];
  assign rd_3r0d[12] = rdfint_3n[12];
  assign rd_3r0d[13] = rdfint_3n[13];
  assign rd_3r0d[14] = rdfint_3n[14];
  assign rd_3r0d[15] = rdfint_3n[15];
  assign rd_3r0d[16] = rdfint_3n[16];
  assign rd_3r0d[17] = rdfint_3n[17];
  assign rd_3r0d[18] = rdfint_3n[18];
  assign rd_3r0d[19] = rdfint_3n[19];
  assign rd_3r0d[20] = rdfint_3n[20];
  assign rd_3r0d[21] = rdfint_3n[21];
  assign rd_3r0d[22] = rdfint_3n[22];
  assign rd_3r0d[23] = rdfint_3n[23];
  assign rd_3r0d[24] = rdfint_3n[24];
  assign rd_3r0d[25] = rdfint_3n[25];
  assign rd_3r0d[26] = rdfint_3n[26];
  assign rd_3r0d[27] = rdfint_3n[27];
  assign rd_3r0d[28] = rdfint_3n[28];
  assign rd_3r0d[29] = rdfint_3n[29];
  assign rd_3r0d[30] = rdfint_3n[30];
  assign rd_3r0d[31] = rdfint_3n[31];
  assign rd_3r1d[0] = rdtint_3n[0];
  assign rd_3r1d[1] = rdtint_3n[1];
  assign rd_3r1d[2] = rdtint_3n[2];
  assign rd_3r1d[3] = rdtint_3n[3];
  assign rd_3r1d[4] = rdtint_3n[4];
  assign rd_3r1d[5] = rdtint_3n[5];
  assign rd_3r1d[6] = rdtint_3n[6];
  assign rd_3r1d[7] = rdtint_3n[7];
  assign rd_3r1d[8] = rdtint_3n[8];
  assign rd_3r1d[9] = rdtint_3n[9];
  assign rd_3r1d[10] = rdtint_3n[10];
  assign rd_3r1d[11] = rdtint_3n[11];
  assign rd_3r1d[12] = rdtint_3n[12];
  assign rd_3r1d[13] = rdtint_3n[13];
  assign rd_3r1d[14] = rdtint_3n[14];
  assign rd_3r1d[15] = rdtint_3n[15];
  assign rd_3r1d[16] = rdtint_3n[16];
  assign rd_3r1d[17] = rdtint_3n[17];
  assign rd_3r1d[18] = rdtint_3n[18];
  assign rd_3r1d[19] = rdtint_3n[19];
  assign rd_3r1d[20] = rdtint_3n[20];
  assign rd_3r1d[21] = rdtint_3n[21];
  assign rd_3r1d[22] = rdtint_3n[22];
  assign rd_3r1d[23] = rdtint_3n[23];
  assign rd_3r1d[24] = rdtint_3n[24];
  assign rd_3r1d[25] = rdtint_3n[25];
  assign rd_3r1d[26] = rdtint_3n[26];
  assign rd_3r1d[27] = rdtint_3n[27];
  assign rd_3r1d[28] = rdtint_3n[28];
  assign rd_3r1d[29] = rdtint_3n[29];
  assign rd_3r1d[30] = rdtint_3n[30];
  assign rd_3r1d[31] = rdtint_3n[31];
  assign rgaint_2n = rd_2a;
  assign rd_2r0d[0] = rdfint_2n[0];
  assign rd_2r0d[1] = rdfint_2n[1];
  assign rd_2r0d[2] = rdfint_2n[2];
  assign rd_2r0d[3] = rdfint_2n[3];
  assign rd_2r0d[4] = rdfint_2n[4];
  assign rd_2r0d[5] = rdfint_2n[5];
  assign rd_2r0d[6] = rdfint_2n[6];
  assign rd_2r0d[7] = rdfint_2n[7];
  assign rd_2r0d[8] = rdfint_2n[8];
  assign rd_2r0d[9] = rdfint_2n[9];
  assign rd_2r0d[10] = rdfint_2n[10];
  assign rd_2r0d[11] = rdfint_2n[11];
  assign rd_2r0d[12] = rdfint_2n[12];
  assign rd_2r0d[13] = rdfint_2n[13];
  assign rd_2r0d[14] = rdfint_2n[14];
  assign rd_2r0d[15] = rdfint_2n[15];
  assign rd_2r0d[16] = rdfint_2n[16];
  assign rd_2r0d[17] = rdfint_2n[17];
  assign rd_2r0d[18] = rdfint_2n[18];
  assign rd_2r0d[19] = rdfint_2n[19];
  assign rd_2r0d[20] = rdfint_2n[20];
  assign rd_2r0d[21] = rdfint_2n[21];
  assign rd_2r0d[22] = rdfint_2n[22];
  assign rd_2r0d[23] = rdfint_2n[23];
  assign rd_2r0d[24] = rdfint_2n[24];
  assign rd_2r0d[25] = rdfint_2n[25];
  assign rd_2r0d[26] = rdfint_2n[26];
  assign rd_2r0d[27] = rdfint_2n[27];
  assign rd_2r0d[28] = rdfint_2n[28];
  assign rd_2r0d[29] = rdfint_2n[29];
  assign rd_2r0d[30] = rdfint_2n[30];
  assign rd_2r0d[31] = rdfint_2n[31];
  assign rd_2r0d[32] = rdfint_2n[32];
  assign rd_2r1d[0] = rdtint_2n[0];
  assign rd_2r1d[1] = rdtint_2n[1];
  assign rd_2r1d[2] = rdtint_2n[2];
  assign rd_2r1d[3] = rdtint_2n[3];
  assign rd_2r1d[4] = rdtint_2n[4];
  assign rd_2r1d[5] = rdtint_2n[5];
  assign rd_2r1d[6] = rdtint_2n[6];
  assign rd_2r1d[7] = rdtint_2n[7];
  assign rd_2r1d[8] = rdtint_2n[8];
  assign rd_2r1d[9] = rdtint_2n[9];
  assign rd_2r1d[10] = rdtint_2n[10];
  assign rd_2r1d[11] = rdtint_2n[11];
  assign rd_2r1d[12] = rdtint_2n[12];
  assign rd_2r1d[13] = rdtint_2n[13];
  assign rd_2r1d[14] = rdtint_2n[14];
  assign rd_2r1d[15] = rdtint_2n[15];
  assign rd_2r1d[16] = rdtint_2n[16];
  assign rd_2r1d[17] = rdtint_2n[17];
  assign rd_2r1d[18] = rdtint_2n[18];
  assign rd_2r1d[19] = rdtint_2n[19];
  assign rd_2r1d[20] = rdtint_2n[20];
  assign rd_2r1d[21] = rdtint_2n[21];
  assign rd_2r1d[22] = rdtint_2n[22];
  assign rd_2r1d[23] = rdtint_2n[23];
  assign rd_2r1d[24] = rdtint_2n[24];
  assign rd_2r1d[25] = rdtint_2n[25];
  assign rd_2r1d[26] = rdtint_2n[26];
  assign rd_2r1d[27] = rdtint_2n[27];
  assign rd_2r1d[28] = rdtint_2n[28];
  assign rd_2r1d[29] = rdtint_2n[29];
  assign rd_2r1d[30] = rdtint_2n[30];
  assign rd_2r1d[31] = rdtint_2n[31];
  assign rd_2r1d[32] = rdtint_2n[32];
  assign rgaint_1n = rd_1a;
  assign rd_1r0d[0] = rdfint_1n[0];
  assign rd_1r0d[1] = rdfint_1n[1];
  assign rd_1r0d[2] = rdfint_1n[2];
  assign rd_1r0d[3] = rdfint_1n[3];
  assign rd_1r0d[4] = rdfint_1n[4];
  assign rd_1r0d[5] = rdfint_1n[5];
  assign rd_1r0d[6] = rdfint_1n[6];
  assign rd_1r0d[7] = rdfint_1n[7];
  assign rd_1r0d[8] = rdfint_1n[8];
  assign rd_1r0d[9] = rdfint_1n[9];
  assign rd_1r0d[10] = rdfint_1n[10];
  assign rd_1r0d[11] = rdfint_1n[11];
  assign rd_1r0d[12] = rdfint_1n[12];
  assign rd_1r0d[13] = rdfint_1n[13];
  assign rd_1r0d[14] = rdfint_1n[14];
  assign rd_1r0d[15] = rdfint_1n[15];
  assign rd_1r0d[16] = rdfint_1n[16];
  assign rd_1r0d[17] = rdfint_1n[17];
  assign rd_1r0d[18] = rdfint_1n[18];
  assign rd_1r0d[19] = rdfint_1n[19];
  assign rd_1r0d[20] = rdfint_1n[20];
  assign rd_1r0d[21] = rdfint_1n[21];
  assign rd_1r0d[22] = rdfint_1n[22];
  assign rd_1r0d[23] = rdfint_1n[23];
  assign rd_1r0d[24] = rdfint_1n[24];
  assign rd_1r0d[25] = rdfint_1n[25];
  assign rd_1r0d[26] = rdfint_1n[26];
  assign rd_1r0d[27] = rdfint_1n[27];
  assign rd_1r0d[28] = rdfint_1n[28];
  assign rd_1r0d[29] = rdfint_1n[29];
  assign rd_1r0d[30] = rdfint_1n[30];
  assign rd_1r0d[31] = rdfint_1n[31];
  assign rd_1r0d[32] = rdfint_1n[32];
  assign rd_1r0d[33] = rdfint_1n[33];
  assign rd_1r1d[0] = rdtint_1n[0];
  assign rd_1r1d[1] = rdtint_1n[1];
  assign rd_1r1d[2] = rdtint_1n[2];
  assign rd_1r1d[3] = rdtint_1n[3];
  assign rd_1r1d[4] = rdtint_1n[4];
  assign rd_1r1d[5] = rdtint_1n[5];
  assign rd_1r1d[6] = rdtint_1n[6];
  assign rd_1r1d[7] = rdtint_1n[7];
  assign rd_1r1d[8] = rdtint_1n[8];
  assign rd_1r1d[9] = rdtint_1n[9];
  assign rd_1r1d[10] = rdtint_1n[10];
  assign rd_1r1d[11] = rdtint_1n[11];
  assign rd_1r1d[12] = rdtint_1n[12];
  assign rd_1r1d[13] = rdtint_1n[13];
  assign rd_1r1d[14] = rdtint_1n[14];
  assign rd_1r1d[15] = rdtint_1n[15];
  assign rd_1r1d[16] = rdtint_1n[16];
  assign rd_1r1d[17] = rdtint_1n[17];
  assign rd_1r1d[18] = rdtint_1n[18];
  assign rd_1r1d[19] = rdtint_1n[19];
  assign rd_1r1d[20] = rdtint_1n[20];
  assign rd_1r1d[21] = rdtint_1n[21];
  assign rd_1r1d[22] = rdtint_1n[22];
  assign rd_1r1d[23] = rdtint_1n[23];
  assign rd_1r1d[24] = rdtint_1n[24];
  assign rd_1r1d[25] = rdtint_1n[25];
  assign rd_1r1d[26] = rdtint_1n[26];
  assign rd_1r1d[27] = rdtint_1n[27];
  assign rd_1r1d[28] = rdtint_1n[28];
  assign rd_1r1d[29] = rdtint_1n[29];
  assign rd_1r1d[30] = rdtint_1n[30];
  assign rd_1r1d[31] = rdtint_1n[31];
  assign rd_1r1d[32] = rdtint_1n[32];
  assign rd_1r1d[33] = rdtint_1n[33];
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r0d[10] = rdfint_0n[10];
  assign rd_0r0d[11] = rdfint_0n[11];
  assign rd_0r0d[12] = rdfint_0n[12];
  assign rd_0r0d[13] = rdfint_0n[13];
  assign rd_0r0d[14] = rdfint_0n[14];
  assign rd_0r0d[15] = rdfint_0n[15];
  assign rd_0r0d[16] = rdfint_0n[16];
  assign rd_0r0d[17] = rdfint_0n[17];
  assign rd_0r0d[18] = rdfint_0n[18];
  assign rd_0r0d[19] = rdfint_0n[19];
  assign rd_0r0d[20] = rdfint_0n[20];
  assign rd_0r0d[21] = rdfint_0n[21];
  assign rd_0r0d[22] = rdfint_0n[22];
  assign rd_0r0d[23] = rdfint_0n[23];
  assign rd_0r0d[24] = rdfint_0n[24];
  assign rd_0r0d[25] = rdfint_0n[25];
  assign rd_0r0d[26] = rdfint_0n[26];
  assign rd_0r0d[27] = rdfint_0n[27];
  assign rd_0r0d[28] = rdfint_0n[28];
  assign rd_0r0d[29] = rdfint_0n[29];
  assign rd_0r0d[30] = rdfint_0n[30];
  assign rd_0r0d[31] = rdfint_0n[31];
  assign rd_0r0d[32] = rdfint_0n[32];
  assign rd_0r0d[33] = rdfint_0n[33];
  assign rd_0r0d[34] = rdfint_0n[34];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign rd_0r1d[10] = rdtint_0n[10];
  assign rd_0r1d[11] = rdtint_0n[11];
  assign rd_0r1d[12] = rdtint_0n[12];
  assign rd_0r1d[13] = rdtint_0n[13];
  assign rd_0r1d[14] = rdtint_0n[14];
  assign rd_0r1d[15] = rdtint_0n[15];
  assign rd_0r1d[16] = rdtint_0n[16];
  assign rd_0r1d[17] = rdtint_0n[17];
  assign rd_0r1d[18] = rdtint_0n[18];
  assign rd_0r1d[19] = rdtint_0n[19];
  assign rd_0r1d[20] = rdtint_0n[20];
  assign rd_0r1d[21] = rdtint_0n[21];
  assign rd_0r1d[22] = rdtint_0n[22];
  assign rd_0r1d[23] = rdtint_0n[23];
  assign rd_0r1d[24] = rdtint_0n[24];
  assign rd_0r1d[25] = rdtint_0n[25];
  assign rd_0r1d[26] = rdtint_0n[26];
  assign rd_0r1d[27] = rdtint_0n[27];
  assign rd_0r1d[28] = rdtint_0n[28];
  assign rd_0r1d[29] = rdtint_0n[29];
  assign rd_0r1d[30] = rdtint_0n[30];
  assign rd_0r1d[31] = rdtint_0n[31];
  assign rd_0r1d[32] = rdtint_0n[32];
  assign rd_0r1d[33] = rdtint_0n[33];
  assign rd_0r1d[34] = rdtint_0n[34];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgfint_0n[32] = wg_0r0d[32];
  assign wgfint_0n[33] = wg_0r0d[33];
  assign wgfint_0n[34] = wg_0r0d[34];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign wgtint_0n[32] = wg_0r1d[32];
  assign wgtint_0n[33] = wg_0r1d[33];
  assign wgtint_0n[34] = wg_0r1d[34];
  assign rg_6a = rgaint_6n;
  assign rgrint_6n = rg_6r;
  assign rg_5a = rgaint_5n;
  assign rgrint_5n = rg_5r;
  assign rg_4a = rgaint_4n;
  assign rgrint_4n = rg_4r;
  assign rg_3a = rgaint_3n;
  assign rgrint_3n = rg_3r;
  assign rg_2a = rgaint_2n;
  assign rgrint_2n = rg_2r;
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR3 I430 (internal_0n[0], rgrint_0n, rgrint_1n, rgrint_2n);
  NOR3 I431 (internal_0n[1], rgrint_3n, rgrint_4n, rgrint_5n);
  NOR3 I432 (internal_0n[2], rgrint_6n, rgaint_0n, rgaint_1n);
  NOR3 I433 (internal_0n[3], rgaint_2n, rgaint_3n, rgaint_4n);
  NOR2 I434 (internal_0n[4], rgaint_5n, rgaint_6n);
  NAND3 I435 (internal_0n[5], internal_0n[0], internal_0n[1], internal_0n[2]);
  NAND2 I436 (internal_0n[6], internal_0n[3], internal_0n[4]);
  NOR2 I437 (nanyread_0n, internal_0n[5], internal_0n[6]);
  AND2 I438 (rdtint_6n, rgrint_6n, dt_0n[32]);
  AND2 I439 (rdtint_5n, rgrint_5n, dt_0n[0]);
  AND2 I440 (rdtint_4n[0], rgrint_4n, dt_0n[0]);
  AND2 I441 (rdtint_4n[1], rgrint_4n, dt_0n[1]);
  AND2 I442 (rdtint_4n[2], rgrint_4n, dt_0n[2]);
  AND2 I443 (rdtint_4n[3], rgrint_4n, dt_0n[3]);
  AND2 I444 (rdtint_4n[4], rgrint_4n, dt_0n[4]);
  AND2 I445 (rdtint_4n[5], rgrint_4n, dt_0n[5]);
  AND2 I446 (rdtint_4n[6], rgrint_4n, dt_0n[6]);
  AND2 I447 (rdtint_4n[7], rgrint_4n, dt_0n[7]);
  AND2 I448 (rdtint_4n[8], rgrint_4n, dt_0n[8]);
  AND2 I449 (rdtint_4n[9], rgrint_4n, dt_0n[9]);
  AND2 I450 (rdtint_4n[10], rgrint_4n, dt_0n[10]);
  AND2 I451 (rdtint_4n[11], rgrint_4n, dt_0n[11]);
  AND2 I452 (rdtint_4n[12], rgrint_4n, dt_0n[12]);
  AND2 I453 (rdtint_4n[13], rgrint_4n, dt_0n[13]);
  AND2 I454 (rdtint_4n[14], rgrint_4n, dt_0n[14]);
  AND2 I455 (rdtint_4n[15], rgrint_4n, dt_0n[15]);
  AND2 I456 (rdtint_4n[16], rgrint_4n, dt_0n[16]);
  AND2 I457 (rdtint_4n[17], rgrint_4n, dt_0n[17]);
  AND2 I458 (rdtint_4n[18], rgrint_4n, dt_0n[18]);
  AND2 I459 (rdtint_4n[19], rgrint_4n, dt_0n[19]);
  AND2 I460 (rdtint_4n[20], rgrint_4n, dt_0n[20]);
  AND2 I461 (rdtint_4n[21], rgrint_4n, dt_0n[21]);
  AND2 I462 (rdtint_4n[22], rgrint_4n, dt_0n[22]);
  AND2 I463 (rdtint_4n[23], rgrint_4n, dt_0n[23]);
  AND2 I464 (rdtint_4n[24], rgrint_4n, dt_0n[24]);
  AND2 I465 (rdtint_4n[25], rgrint_4n, dt_0n[25]);
  AND2 I466 (rdtint_4n[26], rgrint_4n, dt_0n[26]);
  AND2 I467 (rdtint_4n[27], rgrint_4n, dt_0n[27]);
  AND2 I468 (rdtint_4n[28], rgrint_4n, dt_0n[28]);
  AND2 I469 (rdtint_4n[29], rgrint_4n, dt_0n[29]);
  AND2 I470 (rdtint_4n[30], rgrint_4n, dt_0n[30]);
  AND2 I471 (rdtint_4n[31], rgrint_4n, dt_0n[31]);
  AND2 I472 (rdtint_3n[0], rgrint_3n, dt_0n[1]);
  AND2 I473 (rdtint_3n[1], rgrint_3n, dt_0n[2]);
  AND2 I474 (rdtint_3n[2], rgrint_3n, dt_0n[3]);
  AND2 I475 (rdtint_3n[3], rgrint_3n, dt_0n[4]);
  AND2 I476 (rdtint_3n[4], rgrint_3n, dt_0n[5]);
  AND2 I477 (rdtint_3n[5], rgrint_3n, dt_0n[6]);
  AND2 I478 (rdtint_3n[6], rgrint_3n, dt_0n[7]);
  AND2 I479 (rdtint_3n[7], rgrint_3n, dt_0n[8]);
  AND2 I480 (rdtint_3n[8], rgrint_3n, dt_0n[9]);
  AND2 I481 (rdtint_3n[9], rgrint_3n, dt_0n[10]);
  AND2 I482 (rdtint_3n[10], rgrint_3n, dt_0n[11]);
  AND2 I483 (rdtint_3n[11], rgrint_3n, dt_0n[12]);
  AND2 I484 (rdtint_3n[12], rgrint_3n, dt_0n[13]);
  AND2 I485 (rdtint_3n[13], rgrint_3n, dt_0n[14]);
  AND2 I486 (rdtint_3n[14], rgrint_3n, dt_0n[15]);
  AND2 I487 (rdtint_3n[15], rgrint_3n, dt_0n[16]);
  AND2 I488 (rdtint_3n[16], rgrint_3n, dt_0n[17]);
  AND2 I489 (rdtint_3n[17], rgrint_3n, dt_0n[18]);
  AND2 I490 (rdtint_3n[18], rgrint_3n, dt_0n[19]);
  AND2 I491 (rdtint_3n[19], rgrint_3n, dt_0n[20]);
  AND2 I492 (rdtint_3n[20], rgrint_3n, dt_0n[21]);
  AND2 I493 (rdtint_3n[21], rgrint_3n, dt_0n[22]);
  AND2 I494 (rdtint_3n[22], rgrint_3n, dt_0n[23]);
  AND2 I495 (rdtint_3n[23], rgrint_3n, dt_0n[24]);
  AND2 I496 (rdtint_3n[24], rgrint_3n, dt_0n[25]);
  AND2 I497 (rdtint_3n[25], rgrint_3n, dt_0n[26]);
  AND2 I498 (rdtint_3n[26], rgrint_3n, dt_0n[27]);
  AND2 I499 (rdtint_3n[27], rgrint_3n, dt_0n[28]);
  AND2 I500 (rdtint_3n[28], rgrint_3n, dt_0n[29]);
  AND2 I501 (rdtint_3n[29], rgrint_3n, dt_0n[30]);
  AND2 I502 (rdtint_3n[30], rgrint_3n, dt_0n[31]);
  AND2 I503 (rdtint_3n[31], rgrint_3n, dt_0n[32]);
  AND2 I504 (rdtint_2n[0], rgrint_2n, dt_0n[0]);
  AND2 I505 (rdtint_2n[1], rgrint_2n, dt_0n[1]);
  AND2 I506 (rdtint_2n[2], rgrint_2n, dt_0n[2]);
  AND2 I507 (rdtint_2n[3], rgrint_2n, dt_0n[3]);
  AND2 I508 (rdtint_2n[4], rgrint_2n, dt_0n[4]);
  AND2 I509 (rdtint_2n[5], rgrint_2n, dt_0n[5]);
  AND2 I510 (rdtint_2n[6], rgrint_2n, dt_0n[6]);
  AND2 I511 (rdtint_2n[7], rgrint_2n, dt_0n[7]);
  AND2 I512 (rdtint_2n[8], rgrint_2n, dt_0n[8]);
  AND2 I513 (rdtint_2n[9], rgrint_2n, dt_0n[9]);
  AND2 I514 (rdtint_2n[10], rgrint_2n, dt_0n[10]);
  AND2 I515 (rdtint_2n[11], rgrint_2n, dt_0n[11]);
  AND2 I516 (rdtint_2n[12], rgrint_2n, dt_0n[12]);
  AND2 I517 (rdtint_2n[13], rgrint_2n, dt_0n[13]);
  AND2 I518 (rdtint_2n[14], rgrint_2n, dt_0n[14]);
  AND2 I519 (rdtint_2n[15], rgrint_2n, dt_0n[15]);
  AND2 I520 (rdtint_2n[16], rgrint_2n, dt_0n[16]);
  AND2 I521 (rdtint_2n[17], rgrint_2n, dt_0n[17]);
  AND2 I522 (rdtint_2n[18], rgrint_2n, dt_0n[18]);
  AND2 I523 (rdtint_2n[19], rgrint_2n, dt_0n[19]);
  AND2 I524 (rdtint_2n[20], rgrint_2n, dt_0n[20]);
  AND2 I525 (rdtint_2n[21], rgrint_2n, dt_0n[21]);
  AND2 I526 (rdtint_2n[22], rgrint_2n, dt_0n[22]);
  AND2 I527 (rdtint_2n[23], rgrint_2n, dt_0n[23]);
  AND2 I528 (rdtint_2n[24], rgrint_2n, dt_0n[24]);
  AND2 I529 (rdtint_2n[25], rgrint_2n, dt_0n[25]);
  AND2 I530 (rdtint_2n[26], rgrint_2n, dt_0n[26]);
  AND2 I531 (rdtint_2n[27], rgrint_2n, dt_0n[27]);
  AND2 I532 (rdtint_2n[28], rgrint_2n, dt_0n[28]);
  AND2 I533 (rdtint_2n[29], rgrint_2n, dt_0n[29]);
  AND2 I534 (rdtint_2n[30], rgrint_2n, dt_0n[30]);
  AND2 I535 (rdtint_2n[31], rgrint_2n, dt_0n[31]);
  AND2 I536 (rdtint_2n[32], rgrint_2n, dt_0n[32]);
  AND2 I537 (rdtint_1n[0], rgrint_1n, dt_0n[0]);
  AND2 I538 (rdtint_1n[1], rgrint_1n, dt_0n[1]);
  AND2 I539 (rdtint_1n[2], rgrint_1n, dt_0n[2]);
  AND2 I540 (rdtint_1n[3], rgrint_1n, dt_0n[3]);
  AND2 I541 (rdtint_1n[4], rgrint_1n, dt_0n[4]);
  AND2 I542 (rdtint_1n[5], rgrint_1n, dt_0n[5]);
  AND2 I543 (rdtint_1n[6], rgrint_1n, dt_0n[6]);
  AND2 I544 (rdtint_1n[7], rgrint_1n, dt_0n[7]);
  AND2 I545 (rdtint_1n[8], rgrint_1n, dt_0n[8]);
  AND2 I546 (rdtint_1n[9], rgrint_1n, dt_0n[9]);
  AND2 I547 (rdtint_1n[10], rgrint_1n, dt_0n[10]);
  AND2 I548 (rdtint_1n[11], rgrint_1n, dt_0n[11]);
  AND2 I549 (rdtint_1n[12], rgrint_1n, dt_0n[12]);
  AND2 I550 (rdtint_1n[13], rgrint_1n, dt_0n[13]);
  AND2 I551 (rdtint_1n[14], rgrint_1n, dt_0n[14]);
  AND2 I552 (rdtint_1n[15], rgrint_1n, dt_0n[15]);
  AND2 I553 (rdtint_1n[16], rgrint_1n, dt_0n[16]);
  AND2 I554 (rdtint_1n[17], rgrint_1n, dt_0n[17]);
  AND2 I555 (rdtint_1n[18], rgrint_1n, dt_0n[18]);
  AND2 I556 (rdtint_1n[19], rgrint_1n, dt_0n[19]);
  AND2 I557 (rdtint_1n[20], rgrint_1n, dt_0n[20]);
  AND2 I558 (rdtint_1n[21], rgrint_1n, dt_0n[21]);
  AND2 I559 (rdtint_1n[22], rgrint_1n, dt_0n[22]);
  AND2 I560 (rdtint_1n[23], rgrint_1n, dt_0n[23]);
  AND2 I561 (rdtint_1n[24], rgrint_1n, dt_0n[24]);
  AND2 I562 (rdtint_1n[25], rgrint_1n, dt_0n[25]);
  AND2 I563 (rdtint_1n[26], rgrint_1n, dt_0n[26]);
  AND2 I564 (rdtint_1n[27], rgrint_1n, dt_0n[27]);
  AND2 I565 (rdtint_1n[28], rgrint_1n, dt_0n[28]);
  AND2 I566 (rdtint_1n[29], rgrint_1n, dt_0n[29]);
  AND2 I567 (rdtint_1n[30], rgrint_1n, dt_0n[30]);
  AND2 I568 (rdtint_1n[31], rgrint_1n, dt_0n[31]);
  AND2 I569 (rdtint_1n[32], rgrint_1n, dt_0n[32]);
  AND2 I570 (rdtint_1n[33], rgrint_1n, dt_0n[33]);
  AND2 I571 (rdtint_0n[0], rgrint_0n, dt_0n[0]);
  AND2 I572 (rdtint_0n[1], rgrint_0n, dt_0n[1]);
  AND2 I573 (rdtint_0n[2], rgrint_0n, dt_0n[2]);
  AND2 I574 (rdtint_0n[3], rgrint_0n, dt_0n[3]);
  AND2 I575 (rdtint_0n[4], rgrint_0n, dt_0n[4]);
  AND2 I576 (rdtint_0n[5], rgrint_0n, dt_0n[5]);
  AND2 I577 (rdtint_0n[6], rgrint_0n, dt_0n[6]);
  AND2 I578 (rdtint_0n[7], rgrint_0n, dt_0n[7]);
  AND2 I579 (rdtint_0n[8], rgrint_0n, dt_0n[8]);
  AND2 I580 (rdtint_0n[9], rgrint_0n, dt_0n[9]);
  AND2 I581 (rdtint_0n[10], rgrint_0n, dt_0n[10]);
  AND2 I582 (rdtint_0n[11], rgrint_0n, dt_0n[11]);
  AND2 I583 (rdtint_0n[12], rgrint_0n, dt_0n[12]);
  AND2 I584 (rdtint_0n[13], rgrint_0n, dt_0n[13]);
  AND2 I585 (rdtint_0n[14], rgrint_0n, dt_0n[14]);
  AND2 I586 (rdtint_0n[15], rgrint_0n, dt_0n[15]);
  AND2 I587 (rdtint_0n[16], rgrint_0n, dt_0n[16]);
  AND2 I588 (rdtint_0n[17], rgrint_0n, dt_0n[17]);
  AND2 I589 (rdtint_0n[18], rgrint_0n, dt_0n[18]);
  AND2 I590 (rdtint_0n[19], rgrint_0n, dt_0n[19]);
  AND2 I591 (rdtint_0n[20], rgrint_0n, dt_0n[20]);
  AND2 I592 (rdtint_0n[21], rgrint_0n, dt_0n[21]);
  AND2 I593 (rdtint_0n[22], rgrint_0n, dt_0n[22]);
  AND2 I594 (rdtint_0n[23], rgrint_0n, dt_0n[23]);
  AND2 I595 (rdtint_0n[24], rgrint_0n, dt_0n[24]);
  AND2 I596 (rdtint_0n[25], rgrint_0n, dt_0n[25]);
  AND2 I597 (rdtint_0n[26], rgrint_0n, dt_0n[26]);
  AND2 I598 (rdtint_0n[27], rgrint_0n, dt_0n[27]);
  AND2 I599 (rdtint_0n[28], rgrint_0n, dt_0n[28]);
  AND2 I600 (rdtint_0n[29], rgrint_0n, dt_0n[29]);
  AND2 I601 (rdtint_0n[30], rgrint_0n, dt_0n[30]);
  AND2 I602 (rdtint_0n[31], rgrint_0n, dt_0n[31]);
  AND2 I603 (rdtint_0n[32], rgrint_0n, dt_0n[32]);
  AND2 I604 (rdtint_0n[33], rgrint_0n, dt_0n[33]);
  AND2 I605 (rdtint_0n[34], rgrint_0n, dt_0n[34]);
  AND2 I606 (rdfint_6n, rgrint_6n, df_0n[32]);
  AND2 I607 (rdfint_5n, rgrint_5n, df_0n[0]);
  AND2 I608 (rdfint_4n[0], rgrint_4n, df_0n[0]);
  AND2 I609 (rdfint_4n[1], rgrint_4n, df_0n[1]);
  AND2 I610 (rdfint_4n[2], rgrint_4n, df_0n[2]);
  AND2 I611 (rdfint_4n[3], rgrint_4n, df_0n[3]);
  AND2 I612 (rdfint_4n[4], rgrint_4n, df_0n[4]);
  AND2 I613 (rdfint_4n[5], rgrint_4n, df_0n[5]);
  AND2 I614 (rdfint_4n[6], rgrint_4n, df_0n[6]);
  AND2 I615 (rdfint_4n[7], rgrint_4n, df_0n[7]);
  AND2 I616 (rdfint_4n[8], rgrint_4n, df_0n[8]);
  AND2 I617 (rdfint_4n[9], rgrint_4n, df_0n[9]);
  AND2 I618 (rdfint_4n[10], rgrint_4n, df_0n[10]);
  AND2 I619 (rdfint_4n[11], rgrint_4n, df_0n[11]);
  AND2 I620 (rdfint_4n[12], rgrint_4n, df_0n[12]);
  AND2 I621 (rdfint_4n[13], rgrint_4n, df_0n[13]);
  AND2 I622 (rdfint_4n[14], rgrint_4n, df_0n[14]);
  AND2 I623 (rdfint_4n[15], rgrint_4n, df_0n[15]);
  AND2 I624 (rdfint_4n[16], rgrint_4n, df_0n[16]);
  AND2 I625 (rdfint_4n[17], rgrint_4n, df_0n[17]);
  AND2 I626 (rdfint_4n[18], rgrint_4n, df_0n[18]);
  AND2 I627 (rdfint_4n[19], rgrint_4n, df_0n[19]);
  AND2 I628 (rdfint_4n[20], rgrint_4n, df_0n[20]);
  AND2 I629 (rdfint_4n[21], rgrint_4n, df_0n[21]);
  AND2 I630 (rdfint_4n[22], rgrint_4n, df_0n[22]);
  AND2 I631 (rdfint_4n[23], rgrint_4n, df_0n[23]);
  AND2 I632 (rdfint_4n[24], rgrint_4n, df_0n[24]);
  AND2 I633 (rdfint_4n[25], rgrint_4n, df_0n[25]);
  AND2 I634 (rdfint_4n[26], rgrint_4n, df_0n[26]);
  AND2 I635 (rdfint_4n[27], rgrint_4n, df_0n[27]);
  AND2 I636 (rdfint_4n[28], rgrint_4n, df_0n[28]);
  AND2 I637 (rdfint_4n[29], rgrint_4n, df_0n[29]);
  AND2 I638 (rdfint_4n[30], rgrint_4n, df_0n[30]);
  AND2 I639 (rdfint_4n[31], rgrint_4n, df_0n[31]);
  AND2 I640 (rdfint_3n[0], rgrint_3n, df_0n[1]);
  AND2 I641 (rdfint_3n[1], rgrint_3n, df_0n[2]);
  AND2 I642 (rdfint_3n[2], rgrint_3n, df_0n[3]);
  AND2 I643 (rdfint_3n[3], rgrint_3n, df_0n[4]);
  AND2 I644 (rdfint_3n[4], rgrint_3n, df_0n[5]);
  AND2 I645 (rdfint_3n[5], rgrint_3n, df_0n[6]);
  AND2 I646 (rdfint_3n[6], rgrint_3n, df_0n[7]);
  AND2 I647 (rdfint_3n[7], rgrint_3n, df_0n[8]);
  AND2 I648 (rdfint_3n[8], rgrint_3n, df_0n[9]);
  AND2 I649 (rdfint_3n[9], rgrint_3n, df_0n[10]);
  AND2 I650 (rdfint_3n[10], rgrint_3n, df_0n[11]);
  AND2 I651 (rdfint_3n[11], rgrint_3n, df_0n[12]);
  AND2 I652 (rdfint_3n[12], rgrint_3n, df_0n[13]);
  AND2 I653 (rdfint_3n[13], rgrint_3n, df_0n[14]);
  AND2 I654 (rdfint_3n[14], rgrint_3n, df_0n[15]);
  AND2 I655 (rdfint_3n[15], rgrint_3n, df_0n[16]);
  AND2 I656 (rdfint_3n[16], rgrint_3n, df_0n[17]);
  AND2 I657 (rdfint_3n[17], rgrint_3n, df_0n[18]);
  AND2 I658 (rdfint_3n[18], rgrint_3n, df_0n[19]);
  AND2 I659 (rdfint_3n[19], rgrint_3n, df_0n[20]);
  AND2 I660 (rdfint_3n[20], rgrint_3n, df_0n[21]);
  AND2 I661 (rdfint_3n[21], rgrint_3n, df_0n[22]);
  AND2 I662 (rdfint_3n[22], rgrint_3n, df_0n[23]);
  AND2 I663 (rdfint_3n[23], rgrint_3n, df_0n[24]);
  AND2 I664 (rdfint_3n[24], rgrint_3n, df_0n[25]);
  AND2 I665 (rdfint_3n[25], rgrint_3n, df_0n[26]);
  AND2 I666 (rdfint_3n[26], rgrint_3n, df_0n[27]);
  AND2 I667 (rdfint_3n[27], rgrint_3n, df_0n[28]);
  AND2 I668 (rdfint_3n[28], rgrint_3n, df_0n[29]);
  AND2 I669 (rdfint_3n[29], rgrint_3n, df_0n[30]);
  AND2 I670 (rdfint_3n[30], rgrint_3n, df_0n[31]);
  AND2 I671 (rdfint_3n[31], rgrint_3n, df_0n[32]);
  AND2 I672 (rdfint_2n[0], rgrint_2n, df_0n[0]);
  AND2 I673 (rdfint_2n[1], rgrint_2n, df_0n[1]);
  AND2 I674 (rdfint_2n[2], rgrint_2n, df_0n[2]);
  AND2 I675 (rdfint_2n[3], rgrint_2n, df_0n[3]);
  AND2 I676 (rdfint_2n[4], rgrint_2n, df_0n[4]);
  AND2 I677 (rdfint_2n[5], rgrint_2n, df_0n[5]);
  AND2 I678 (rdfint_2n[6], rgrint_2n, df_0n[6]);
  AND2 I679 (rdfint_2n[7], rgrint_2n, df_0n[7]);
  AND2 I680 (rdfint_2n[8], rgrint_2n, df_0n[8]);
  AND2 I681 (rdfint_2n[9], rgrint_2n, df_0n[9]);
  AND2 I682 (rdfint_2n[10], rgrint_2n, df_0n[10]);
  AND2 I683 (rdfint_2n[11], rgrint_2n, df_0n[11]);
  AND2 I684 (rdfint_2n[12], rgrint_2n, df_0n[12]);
  AND2 I685 (rdfint_2n[13], rgrint_2n, df_0n[13]);
  AND2 I686 (rdfint_2n[14], rgrint_2n, df_0n[14]);
  AND2 I687 (rdfint_2n[15], rgrint_2n, df_0n[15]);
  AND2 I688 (rdfint_2n[16], rgrint_2n, df_0n[16]);
  AND2 I689 (rdfint_2n[17], rgrint_2n, df_0n[17]);
  AND2 I690 (rdfint_2n[18], rgrint_2n, df_0n[18]);
  AND2 I691 (rdfint_2n[19], rgrint_2n, df_0n[19]);
  AND2 I692 (rdfint_2n[20], rgrint_2n, df_0n[20]);
  AND2 I693 (rdfint_2n[21], rgrint_2n, df_0n[21]);
  AND2 I694 (rdfint_2n[22], rgrint_2n, df_0n[22]);
  AND2 I695 (rdfint_2n[23], rgrint_2n, df_0n[23]);
  AND2 I696 (rdfint_2n[24], rgrint_2n, df_0n[24]);
  AND2 I697 (rdfint_2n[25], rgrint_2n, df_0n[25]);
  AND2 I698 (rdfint_2n[26], rgrint_2n, df_0n[26]);
  AND2 I699 (rdfint_2n[27], rgrint_2n, df_0n[27]);
  AND2 I700 (rdfint_2n[28], rgrint_2n, df_0n[28]);
  AND2 I701 (rdfint_2n[29], rgrint_2n, df_0n[29]);
  AND2 I702 (rdfint_2n[30], rgrint_2n, df_0n[30]);
  AND2 I703 (rdfint_2n[31], rgrint_2n, df_0n[31]);
  AND2 I704 (rdfint_2n[32], rgrint_2n, df_0n[32]);
  AND2 I705 (rdfint_1n[0], rgrint_1n, df_0n[0]);
  AND2 I706 (rdfint_1n[1], rgrint_1n, df_0n[1]);
  AND2 I707 (rdfint_1n[2], rgrint_1n, df_0n[2]);
  AND2 I708 (rdfint_1n[3], rgrint_1n, df_0n[3]);
  AND2 I709 (rdfint_1n[4], rgrint_1n, df_0n[4]);
  AND2 I710 (rdfint_1n[5], rgrint_1n, df_0n[5]);
  AND2 I711 (rdfint_1n[6], rgrint_1n, df_0n[6]);
  AND2 I712 (rdfint_1n[7], rgrint_1n, df_0n[7]);
  AND2 I713 (rdfint_1n[8], rgrint_1n, df_0n[8]);
  AND2 I714 (rdfint_1n[9], rgrint_1n, df_0n[9]);
  AND2 I715 (rdfint_1n[10], rgrint_1n, df_0n[10]);
  AND2 I716 (rdfint_1n[11], rgrint_1n, df_0n[11]);
  AND2 I717 (rdfint_1n[12], rgrint_1n, df_0n[12]);
  AND2 I718 (rdfint_1n[13], rgrint_1n, df_0n[13]);
  AND2 I719 (rdfint_1n[14], rgrint_1n, df_0n[14]);
  AND2 I720 (rdfint_1n[15], rgrint_1n, df_0n[15]);
  AND2 I721 (rdfint_1n[16], rgrint_1n, df_0n[16]);
  AND2 I722 (rdfint_1n[17], rgrint_1n, df_0n[17]);
  AND2 I723 (rdfint_1n[18], rgrint_1n, df_0n[18]);
  AND2 I724 (rdfint_1n[19], rgrint_1n, df_0n[19]);
  AND2 I725 (rdfint_1n[20], rgrint_1n, df_0n[20]);
  AND2 I726 (rdfint_1n[21], rgrint_1n, df_0n[21]);
  AND2 I727 (rdfint_1n[22], rgrint_1n, df_0n[22]);
  AND2 I728 (rdfint_1n[23], rgrint_1n, df_0n[23]);
  AND2 I729 (rdfint_1n[24], rgrint_1n, df_0n[24]);
  AND2 I730 (rdfint_1n[25], rgrint_1n, df_0n[25]);
  AND2 I731 (rdfint_1n[26], rgrint_1n, df_0n[26]);
  AND2 I732 (rdfint_1n[27], rgrint_1n, df_0n[27]);
  AND2 I733 (rdfint_1n[28], rgrint_1n, df_0n[28]);
  AND2 I734 (rdfint_1n[29], rgrint_1n, df_0n[29]);
  AND2 I735 (rdfint_1n[30], rgrint_1n, df_0n[30]);
  AND2 I736 (rdfint_1n[31], rgrint_1n, df_0n[31]);
  AND2 I737 (rdfint_1n[32], rgrint_1n, df_0n[32]);
  AND2 I738 (rdfint_1n[33], rgrint_1n, df_0n[33]);
  AND2 I739 (rdfint_0n[0], rgrint_0n, df_0n[0]);
  AND2 I740 (rdfint_0n[1], rgrint_0n, df_0n[1]);
  AND2 I741 (rdfint_0n[2], rgrint_0n, df_0n[2]);
  AND2 I742 (rdfint_0n[3], rgrint_0n, df_0n[3]);
  AND2 I743 (rdfint_0n[4], rgrint_0n, df_0n[4]);
  AND2 I744 (rdfint_0n[5], rgrint_0n, df_0n[5]);
  AND2 I745 (rdfint_0n[6], rgrint_0n, df_0n[6]);
  AND2 I746 (rdfint_0n[7], rgrint_0n, df_0n[7]);
  AND2 I747 (rdfint_0n[8], rgrint_0n, df_0n[8]);
  AND2 I748 (rdfint_0n[9], rgrint_0n, df_0n[9]);
  AND2 I749 (rdfint_0n[10], rgrint_0n, df_0n[10]);
  AND2 I750 (rdfint_0n[11], rgrint_0n, df_0n[11]);
  AND2 I751 (rdfint_0n[12], rgrint_0n, df_0n[12]);
  AND2 I752 (rdfint_0n[13], rgrint_0n, df_0n[13]);
  AND2 I753 (rdfint_0n[14], rgrint_0n, df_0n[14]);
  AND2 I754 (rdfint_0n[15], rgrint_0n, df_0n[15]);
  AND2 I755 (rdfint_0n[16], rgrint_0n, df_0n[16]);
  AND2 I756 (rdfint_0n[17], rgrint_0n, df_0n[17]);
  AND2 I757 (rdfint_0n[18], rgrint_0n, df_0n[18]);
  AND2 I758 (rdfint_0n[19], rgrint_0n, df_0n[19]);
  AND2 I759 (rdfint_0n[20], rgrint_0n, df_0n[20]);
  AND2 I760 (rdfint_0n[21], rgrint_0n, df_0n[21]);
  AND2 I761 (rdfint_0n[22], rgrint_0n, df_0n[22]);
  AND2 I762 (rdfint_0n[23], rgrint_0n, df_0n[23]);
  AND2 I763 (rdfint_0n[24], rgrint_0n, df_0n[24]);
  AND2 I764 (rdfint_0n[25], rgrint_0n, df_0n[25]);
  AND2 I765 (rdfint_0n[26], rgrint_0n, df_0n[26]);
  AND2 I766 (rdfint_0n[27], rgrint_0n, df_0n[27]);
  AND2 I767 (rdfint_0n[28], rgrint_0n, df_0n[28]);
  AND2 I768 (rdfint_0n[29], rgrint_0n, df_0n[29]);
  AND2 I769 (rdfint_0n[30], rgrint_0n, df_0n[30]);
  AND2 I770 (rdfint_0n[31], rgrint_0n, df_0n[31]);
  AND2 I771 (rdfint_0n[32], rgrint_0n, df_0n[32]);
  AND2 I772 (rdfint_0n[33], rgrint_0n, df_0n[33]);
  AND2 I773 (rdfint_0n[34], rgrint_0n, df_0n[34]);
  C3 I774 (internal_0n[7], wc_0n, wacks_0n[34], wacks_0n[33]);
  C3 I775 (internal_0n[8], wacks_0n[32], wacks_0n[31], wacks_0n[30]);
  C3 I776 (internal_0n[9], wacks_0n[29], wacks_0n[28], wacks_0n[27]);
  C3 I777 (internal_0n[10], wacks_0n[26], wacks_0n[25], wacks_0n[24]);
  C3 I778 (internal_0n[11], wacks_0n[23], wacks_0n[22], wacks_0n[21]);
  C3 I779 (internal_0n[12], wacks_0n[20], wacks_0n[19], wacks_0n[18]);
  C3 I780 (internal_0n[13], wacks_0n[17], wacks_0n[16], wacks_0n[15]);
  C3 I781 (internal_0n[14], wacks_0n[14], wacks_0n[13], wacks_0n[12]);
  C3 I782 (internal_0n[15], wacks_0n[11], wacks_0n[10], wacks_0n[9]);
  C3 I783 (internal_0n[16], wacks_0n[8], wacks_0n[7], wacks_0n[6]);
  C3 I784 (internal_0n[17], wacks_0n[5], wacks_0n[4], wacks_0n[3]);
  C3 I785 (internal_0n[18], wacks_0n[2], wacks_0n[1], wacks_0n[0]);
  C3 I786 (internal_0n[19], internal_0n[7], internal_0n[8], internal_0n[9]);
  C3 I787 (internal_0n[20], internal_0n[10], internal_0n[11], internal_0n[12]);
  C3 I788 (internal_0n[21], internal_0n[13], internal_0n[14], internal_0n[15]);
  C3 I789 (internal_0n[22], internal_0n[16], internal_0n[17], internal_0n[18]);
  C2 I790 (internal_0n[23], internal_0n[19], internal_0n[20]);
  C2 I791 (internal_0n[24], internal_0n[21], internal_0n[22]);
  C2 I792 (wdrint_0n, internal_0n[23], internal_0n[24]);
  assign wen_0n[34] = wc_0n;
  assign wen_0n[33] = wc_0n;
  assign wen_0n[32] = wc_0n;
  assign wen_0n[31] = wc_0n;
  assign wen_0n[30] = wc_0n;
  assign wen_0n[29] = wc_0n;
  assign wen_0n[28] = wc_0n;
  assign wen_0n[27] = wc_0n;
  assign wen_0n[26] = wc_0n;
  assign wen_0n[25] = wc_0n;
  assign wen_0n[24] = wc_0n;
  assign wen_0n[23] = wc_0n;
  assign wen_0n[22] = wc_0n;
  assign wen_0n[21] = wc_0n;
  assign wen_0n[20] = wc_0n;
  assign wen_0n[19] = wc_0n;
  assign wen_0n[18] = wc_0n;
  assign wen_0n[17] = wc_0n;
  assign wen_0n[16] = wc_0n;
  assign wen_0n[15] = wc_0n;
  assign wen_0n[14] = wc_0n;
  assign wen_0n[13] = wc_0n;
  assign wen_0n[12] = wc_0n;
  assign wen_0n[11] = wc_0n;
  assign wen_0n[10] = wc_0n;
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[34] = git_0n[34];
  assign wt_0n[33] = git_0n[33];
  assign wt_0n[32] = git_0n[32];
  assign wt_0n[31] = git_0n[31];
  assign wt_0n[30] = git_0n[30];
  assign wt_0n[29] = git_0n[29];
  assign wt_0n[28] = git_0n[28];
  assign wt_0n[27] = git_0n[27];
  assign wt_0n[26] = git_0n[26];
  assign wt_0n[25] = git_0n[25];
  assign wt_0n[24] = git_0n[24];
  assign wt_0n[23] = git_0n[23];
  assign wt_0n[22] = git_0n[22];
  assign wt_0n[21] = git_0n[21];
  assign wt_0n[20] = git_0n[20];
  assign wt_0n[19] = git_0n[19];
  assign wt_0n[18] = git_0n[18];
  assign wt_0n[17] = git_0n[17];
  assign wt_0n[16] = git_0n[16];
  assign wt_0n[15] = git_0n[15];
  assign wt_0n[14] = git_0n[14];
  assign wt_0n[13] = git_0n[13];
  assign wt_0n[12] = git_0n[12];
  assign wt_0n[11] = git_0n[11];
  assign wt_0n[10] = git_0n[10];
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[34] = gif_0n[34];
  assign wf_0n[33] = gif_0n[33];
  assign wf_0n[32] = gif_0n[32];
  assign wf_0n[31] = gif_0n[31];
  assign wf_0n[30] = gif_0n[30];
  assign wf_0n[29] = gif_0n[29];
  assign wf_0n[28] = gif_0n[28];
  assign wf_0n[27] = gif_0n[27];
  assign wf_0n[26] = gif_0n[26];
  assign wf_0n[25] = gif_0n[25];
  assign wf_0n[24] = gif_0n[24];
  assign wf_0n[23] = gif_0n[23];
  assign wf_0n[22] = gif_0n[22];
  assign wf_0n[21] = gif_0n[21];
  assign wf_0n[20] = gif_0n[20];
  assign wf_0n[19] = gif_0n[19];
  assign wf_0n[18] = gif_0n[18];
  assign wf_0n[17] = gif_0n[17];
  assign wf_0n[16] = gif_0n[16];
  assign wf_0n[15] = gif_0n[15];
  assign wf_0n[14] = gif_0n[14];
  assign wf_0n[13] = gif_0n[13];
  assign wf_0n[12] = gif_0n[12];
  assign wf_0n[11] = gif_0n[11];
  assign wf_0n[10] = gif_0n[10];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I898 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I900 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I901 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I902 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I903 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I904 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I905 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I906 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I907 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I908 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I909 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I910 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I911 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I912 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I913 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I914 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I915 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I916 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I917 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I918 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I919 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I920 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I921 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I922 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I923 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I924 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I925 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I926 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I927 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I928 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I929 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I930 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I931 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I932 (git_0n[32], wgtint_0n[32], ig_0n);
  AND2 I933 (git_0n[33], wgtint_0n[33], ig_0n);
  AND2 I934 (git_0n[34], wgtint_0n[34], ig_0n);
  AND2 I935 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I936 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I937 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I938 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I939 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I940 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I941 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I942 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I943 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I944 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I945 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I946 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I947 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I948 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I949 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I950 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I951 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I952 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I953 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I954 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I955 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I956 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I957 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I958 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I959 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I960 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I961 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I962 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I963 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I964 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I965 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I966 (gif_0n[31], wgfint_0n[31], ig_0n);
  AND2 I967 (gif_0n[32], wgfint_0n[32], ig_0n);
  AND2 I968 (gif_0n[33], wgfint_0n[33], ig_0n);
  AND2 I969 (gif_0n[34], wgfint_0n[34], ig_0n);
  C3 I970 (internal_0n[25], complete1451_0n[0], complete1451_0n[1], complete1451_0n[2]);
  C3 I971 (internal_0n[26], complete1451_0n[3], complete1451_0n[4], complete1451_0n[5]);
  C3 I972 (internal_0n[27], complete1451_0n[6], complete1451_0n[7], complete1451_0n[8]);
  C3 I973 (internal_0n[28], complete1451_0n[9], complete1451_0n[10], complete1451_0n[11]);
  C3 I974 (internal_0n[29], complete1451_0n[12], complete1451_0n[13], complete1451_0n[14]);
  C3 I975 (internal_0n[30], complete1451_0n[15], complete1451_0n[16], complete1451_0n[17]);
  C3 I976 (internal_0n[31], complete1451_0n[18], complete1451_0n[19], complete1451_0n[20]);
  C3 I977 (internal_0n[32], complete1451_0n[21], complete1451_0n[22], complete1451_0n[23]);
  C3 I978 (internal_0n[33], complete1451_0n[24], complete1451_0n[25], complete1451_0n[26]);
  C3 I979 (internal_0n[34], complete1451_0n[27], complete1451_0n[28], complete1451_0n[29]);
  C3 I980 (internal_0n[35], complete1451_0n[30], complete1451_0n[31], complete1451_0n[32]);
  C2 I981 (internal_0n[36], complete1451_0n[33], complete1451_0n[34]);
  C3 I982 (internal_0n[37], internal_0n[25], internal_0n[26], internal_0n[27]);
  C3 I983 (internal_0n[38], internal_0n[28], internal_0n[29], internal_0n[30]);
  C3 I984 (internal_0n[39], internal_0n[31], internal_0n[32], internal_0n[33]);
  C3 I985 (internal_0n[40], internal_0n[34], internal_0n[35], internal_0n[36]);
  C2 I986 (internal_0n[41], internal_0n[37], internal_0n[38]);
  C2 I987 (internal_0n[42], internal_0n[39], internal_0n[40]);
  C2 I988 (wc_0n, internal_0n[41], internal_0n[42]);
  OR2 I989 (complete1451_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I990 (complete1451_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I991 (complete1451_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I992 (complete1451_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I993 (complete1451_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I994 (complete1451_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I995 (complete1451_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I996 (complete1451_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I997 (complete1451_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I998 (complete1451_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I999 (complete1451_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I1000 (complete1451_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I1001 (complete1451_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I1002 (complete1451_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I1003 (complete1451_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I1004 (complete1451_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I1005 (complete1451_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I1006 (complete1451_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I1007 (complete1451_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I1008 (complete1451_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I1009 (complete1451_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I1010 (complete1451_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I1011 (complete1451_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I1012 (complete1451_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I1013 (complete1451_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I1014 (complete1451_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I1015 (complete1451_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I1016 (complete1451_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I1017 (complete1451_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I1018 (complete1451_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I1019 (complete1451_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I1020 (complete1451_0n[31], wgfint_0n[31], wgtint_0n[31]);
  OR2 I1021 (complete1451_0n[32], wgfint_0n[32], wgtint_0n[32]);
  OR2 I1022 (complete1451_0n[33], wgfint_0n[33], wgtint_0n[33]);
  OR2 I1023 (complete1451_0n[34], wgfint_0n[34], wgtint_0n[34]);
  AO22 I1024 (wacks_0n[34], gf1449_0n[34], df_0n[34], gt1450_0n[34], dt_0n[34]);
  NOR2 I1025 (dt_0n[34], df_0n[34], gf1449_0n[34]);
  NOR3 I1026 (df_0n[34], dt_0n[34], gt1450_0n[34], init_0n);
  AND2 I1027 (gt1450_0n[34], wt_0n[34], wen_0n[34]);
  AND2 I1028 (gf1449_0n[34], wf_0n[34], wen_0n[34]);
  AO22 I1029 (wacks_0n[33], gf1449_0n[33], df_0n[33], gt1450_0n[33], dt_0n[33]);
  NOR2 I1030 (dt_0n[33], df_0n[33], gf1449_0n[33]);
  NOR3 I1031 (df_0n[33], dt_0n[33], gt1450_0n[33], init_0n);
  AND2 I1032 (gt1450_0n[33], wt_0n[33], wen_0n[33]);
  AND2 I1033 (gf1449_0n[33], wf_0n[33], wen_0n[33]);
  AO22 I1034 (wacks_0n[32], gf1449_0n[32], df_0n[32], gt1450_0n[32], dt_0n[32]);
  NOR2 I1035 (dt_0n[32], df_0n[32], gf1449_0n[32]);
  NOR3 I1036 (df_0n[32], dt_0n[32], gt1450_0n[32], init_0n);
  AND2 I1037 (gt1450_0n[32], wt_0n[32], wen_0n[32]);
  AND2 I1038 (gf1449_0n[32], wf_0n[32], wen_0n[32]);
  AO22 I1039 (wacks_0n[31], gf1449_0n[31], df_0n[31], gt1450_0n[31], dt_0n[31]);
  NOR2 I1040 (dt_0n[31], df_0n[31], gf1449_0n[31]);
  NOR3 I1041 (df_0n[31], dt_0n[31], gt1450_0n[31], init_0n);
  AND2 I1042 (gt1450_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I1043 (gf1449_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I1044 (wacks_0n[30], gf1449_0n[30], df_0n[30], gt1450_0n[30], dt_0n[30]);
  NOR2 I1045 (dt_0n[30], df_0n[30], gf1449_0n[30]);
  NOR3 I1046 (df_0n[30], dt_0n[30], gt1450_0n[30], init_0n);
  AND2 I1047 (gt1450_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I1048 (gf1449_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I1049 (wacks_0n[29], gf1449_0n[29], df_0n[29], gt1450_0n[29], dt_0n[29]);
  NOR2 I1050 (dt_0n[29], df_0n[29], gf1449_0n[29]);
  NOR3 I1051 (df_0n[29], dt_0n[29], gt1450_0n[29], init_0n);
  AND2 I1052 (gt1450_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I1053 (gf1449_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I1054 (wacks_0n[28], gf1449_0n[28], df_0n[28], gt1450_0n[28], dt_0n[28]);
  NOR2 I1055 (dt_0n[28], df_0n[28], gf1449_0n[28]);
  NOR3 I1056 (df_0n[28], dt_0n[28], gt1450_0n[28], init_0n);
  AND2 I1057 (gt1450_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I1058 (gf1449_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I1059 (wacks_0n[27], gf1449_0n[27], df_0n[27], gt1450_0n[27], dt_0n[27]);
  NOR2 I1060 (dt_0n[27], df_0n[27], gf1449_0n[27]);
  NOR3 I1061 (df_0n[27], dt_0n[27], gt1450_0n[27], init_0n);
  AND2 I1062 (gt1450_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I1063 (gf1449_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I1064 (wacks_0n[26], gf1449_0n[26], df_0n[26], gt1450_0n[26], dt_0n[26]);
  NOR2 I1065 (dt_0n[26], df_0n[26], gf1449_0n[26]);
  NOR3 I1066 (df_0n[26], dt_0n[26], gt1450_0n[26], init_0n);
  AND2 I1067 (gt1450_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I1068 (gf1449_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I1069 (wacks_0n[25], gf1449_0n[25], df_0n[25], gt1450_0n[25], dt_0n[25]);
  NOR2 I1070 (dt_0n[25], df_0n[25], gf1449_0n[25]);
  NOR3 I1071 (df_0n[25], dt_0n[25], gt1450_0n[25], init_0n);
  AND2 I1072 (gt1450_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I1073 (gf1449_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I1074 (wacks_0n[24], gf1449_0n[24], df_0n[24], gt1450_0n[24], dt_0n[24]);
  NOR2 I1075 (dt_0n[24], df_0n[24], gf1449_0n[24]);
  NOR3 I1076 (df_0n[24], dt_0n[24], gt1450_0n[24], init_0n);
  AND2 I1077 (gt1450_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I1078 (gf1449_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I1079 (wacks_0n[23], gf1449_0n[23], df_0n[23], gt1450_0n[23], dt_0n[23]);
  NOR2 I1080 (dt_0n[23], df_0n[23], gf1449_0n[23]);
  NOR3 I1081 (df_0n[23], dt_0n[23], gt1450_0n[23], init_0n);
  AND2 I1082 (gt1450_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I1083 (gf1449_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I1084 (wacks_0n[22], gf1449_0n[22], df_0n[22], gt1450_0n[22], dt_0n[22]);
  NOR2 I1085 (dt_0n[22], df_0n[22], gf1449_0n[22]);
  NOR3 I1086 (df_0n[22], dt_0n[22], gt1450_0n[22], init_0n);
  AND2 I1087 (gt1450_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I1088 (gf1449_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I1089 (wacks_0n[21], gf1449_0n[21], df_0n[21], gt1450_0n[21], dt_0n[21]);
  NOR2 I1090 (dt_0n[21], df_0n[21], gf1449_0n[21]);
  NOR3 I1091 (df_0n[21], dt_0n[21], gt1450_0n[21], init_0n);
  AND2 I1092 (gt1450_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I1093 (gf1449_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I1094 (wacks_0n[20], gf1449_0n[20], df_0n[20], gt1450_0n[20], dt_0n[20]);
  NOR2 I1095 (dt_0n[20], df_0n[20], gf1449_0n[20]);
  NOR3 I1096 (df_0n[20], dt_0n[20], gt1450_0n[20], init_0n);
  AND2 I1097 (gt1450_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I1098 (gf1449_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I1099 (wacks_0n[19], gf1449_0n[19], df_0n[19], gt1450_0n[19], dt_0n[19]);
  NOR2 I1100 (dt_0n[19], df_0n[19], gf1449_0n[19]);
  NOR3 I1101 (df_0n[19], dt_0n[19], gt1450_0n[19], init_0n);
  AND2 I1102 (gt1450_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I1103 (gf1449_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I1104 (wacks_0n[18], gf1449_0n[18], df_0n[18], gt1450_0n[18], dt_0n[18]);
  NOR2 I1105 (dt_0n[18], df_0n[18], gf1449_0n[18]);
  NOR3 I1106 (df_0n[18], dt_0n[18], gt1450_0n[18], init_0n);
  AND2 I1107 (gt1450_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I1108 (gf1449_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I1109 (wacks_0n[17], gf1449_0n[17], df_0n[17], gt1450_0n[17], dt_0n[17]);
  NOR2 I1110 (dt_0n[17], df_0n[17], gf1449_0n[17]);
  NOR3 I1111 (df_0n[17], dt_0n[17], gt1450_0n[17], init_0n);
  AND2 I1112 (gt1450_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I1113 (gf1449_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I1114 (wacks_0n[16], gf1449_0n[16], df_0n[16], gt1450_0n[16], dt_0n[16]);
  NOR2 I1115 (dt_0n[16], df_0n[16], gf1449_0n[16]);
  NOR3 I1116 (df_0n[16], dt_0n[16], gt1450_0n[16], init_0n);
  AND2 I1117 (gt1450_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I1118 (gf1449_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I1119 (wacks_0n[15], gf1449_0n[15], df_0n[15], gt1450_0n[15], dt_0n[15]);
  NOR2 I1120 (dt_0n[15], df_0n[15], gf1449_0n[15]);
  NOR3 I1121 (df_0n[15], dt_0n[15], gt1450_0n[15], init_0n);
  AND2 I1122 (gt1450_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I1123 (gf1449_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I1124 (wacks_0n[14], gf1449_0n[14], df_0n[14], gt1450_0n[14], dt_0n[14]);
  NOR2 I1125 (dt_0n[14], df_0n[14], gf1449_0n[14]);
  NOR3 I1126 (df_0n[14], dt_0n[14], gt1450_0n[14], init_0n);
  AND2 I1127 (gt1450_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I1128 (gf1449_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I1129 (wacks_0n[13], gf1449_0n[13], df_0n[13], gt1450_0n[13], dt_0n[13]);
  NOR2 I1130 (dt_0n[13], df_0n[13], gf1449_0n[13]);
  NOR3 I1131 (df_0n[13], dt_0n[13], gt1450_0n[13], init_0n);
  AND2 I1132 (gt1450_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I1133 (gf1449_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I1134 (wacks_0n[12], gf1449_0n[12], df_0n[12], gt1450_0n[12], dt_0n[12]);
  NOR2 I1135 (dt_0n[12], df_0n[12], gf1449_0n[12]);
  NOR3 I1136 (df_0n[12], dt_0n[12], gt1450_0n[12], init_0n);
  AND2 I1137 (gt1450_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I1138 (gf1449_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I1139 (wacks_0n[11], gf1449_0n[11], df_0n[11], gt1450_0n[11], dt_0n[11]);
  NOR2 I1140 (dt_0n[11], df_0n[11], gf1449_0n[11]);
  NOR3 I1141 (df_0n[11], dt_0n[11], gt1450_0n[11], init_0n);
  AND2 I1142 (gt1450_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I1143 (gf1449_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I1144 (wacks_0n[10], gf1449_0n[10], df_0n[10], gt1450_0n[10], dt_0n[10]);
  NOR2 I1145 (dt_0n[10], df_0n[10], gf1449_0n[10]);
  NOR3 I1146 (df_0n[10], dt_0n[10], gt1450_0n[10], init_0n);
  AND2 I1147 (gt1450_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I1148 (gf1449_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I1149 (wacks_0n[9], gf1449_0n[9], df_0n[9], gt1450_0n[9], dt_0n[9]);
  NOR2 I1150 (dt_0n[9], df_0n[9], gf1449_0n[9]);
  NOR3 I1151 (df_0n[9], dt_0n[9], gt1450_0n[9], init_0n);
  AND2 I1152 (gt1450_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I1153 (gf1449_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I1154 (wacks_0n[8], gf1449_0n[8], df_0n[8], gt1450_0n[8], dt_0n[8]);
  NOR2 I1155 (dt_0n[8], df_0n[8], gf1449_0n[8]);
  NOR3 I1156 (df_0n[8], dt_0n[8], gt1450_0n[8], init_0n);
  AND2 I1157 (gt1450_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I1158 (gf1449_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I1159 (wacks_0n[7], gf1449_0n[7], df_0n[7], gt1450_0n[7], dt_0n[7]);
  NOR2 I1160 (dt_0n[7], df_0n[7], gf1449_0n[7]);
  NOR3 I1161 (df_0n[7], dt_0n[7], gt1450_0n[7], init_0n);
  AND2 I1162 (gt1450_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I1163 (gf1449_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I1164 (wacks_0n[6], gf1449_0n[6], df_0n[6], gt1450_0n[6], dt_0n[6]);
  NOR2 I1165 (dt_0n[6], df_0n[6], gf1449_0n[6]);
  NOR3 I1166 (df_0n[6], dt_0n[6], gt1450_0n[6], init_0n);
  AND2 I1167 (gt1450_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I1168 (gf1449_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I1169 (wacks_0n[5], gf1449_0n[5], df_0n[5], gt1450_0n[5], dt_0n[5]);
  NOR2 I1170 (dt_0n[5], df_0n[5], gf1449_0n[5]);
  NOR3 I1171 (df_0n[5], dt_0n[5], gt1450_0n[5], init_0n);
  AND2 I1172 (gt1450_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I1173 (gf1449_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I1174 (wacks_0n[4], gf1449_0n[4], df_0n[4], gt1450_0n[4], dt_0n[4]);
  NOR2 I1175 (dt_0n[4], df_0n[4], gf1449_0n[4]);
  NOR3 I1176 (df_0n[4], dt_0n[4], gt1450_0n[4], init_0n);
  AND2 I1177 (gt1450_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I1178 (gf1449_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I1179 (wacks_0n[3], gf1449_0n[3], df_0n[3], gt1450_0n[3], dt_0n[3]);
  NOR2 I1180 (dt_0n[3], df_0n[3], gf1449_0n[3]);
  NOR3 I1181 (df_0n[3], dt_0n[3], gt1450_0n[3], init_0n);
  AND2 I1182 (gt1450_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I1183 (gf1449_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I1184 (wacks_0n[2], gf1449_0n[2], df_0n[2], gt1450_0n[2], dt_0n[2]);
  NOR2 I1185 (dt_0n[2], df_0n[2], gf1449_0n[2]);
  NOR3 I1186 (df_0n[2], dt_0n[2], gt1450_0n[2], init_0n);
  AND2 I1187 (gt1450_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I1188 (gf1449_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I1189 (wacks_0n[1], gf1449_0n[1], df_0n[1], gt1450_0n[1], dt_0n[1]);
  NOR2 I1190 (dt_0n[1], df_0n[1], gf1449_0n[1]);
  NOR3 I1191 (df_0n[1], dt_0n[1], gt1450_0n[1], init_0n);
  AND2 I1192 (gt1450_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I1193 (gf1449_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I1194 (wacks_0n[0], gf1449_0n[0], df_0n[0], gt1450_0n[0], dt_0n[0]);
  NOR2 I1195 (dt_0n[0], df_0n[0], gf1449_0n[0]);
  NOR3 I1196 (df_0n[0], dt_0n[0], gt1450_0n[0], init_0n);
  AND2 I1197 (gt1450_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I1198 (gf1449_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I1199 (init_0n, initialise);
endmodule

module BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m90m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  initialise
);
  input [34:0] wg_0r0d;
  input [34:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [34:0] rd_0r0d;
  output [34:0] rd_0r1d;
  input rd_0a;
  output [34:0] rd_1r0d;
  output [34:0] rd_1r1d;
  input rd_1a;
  input initialise;
  wire [37:0] internal_0n;
  wire [34:0] wf_0n;
  wire [34:0] wt_0n;
  wire [34:0] df_0n;
  wire [34:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire wc_0n;
  wire [34:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [34:0] wgfint_0n;
  wire [34:0] wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire [34:0] rdfint_0n;
  wire [34:0] rdfint_1n;
  wire [34:0] rdtint_0n;
  wire [34:0] rdtint_1n;
  wire [34:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [34:0] gif_0n;
  wire [34:0] git_0n;
  wire [34:0] complete1486_0n;
  wire [34:0] gt1485_0n;
  wire [34:0] gf1484_0n;
  assign rgaint_1n = rd_1a;
  assign rd_1r0d[0] = rdfint_1n[0];
  assign rd_1r0d[1] = rdfint_1n[1];
  assign rd_1r0d[2] = rdfint_1n[2];
  assign rd_1r0d[3] = rdfint_1n[3];
  assign rd_1r0d[4] = rdfint_1n[4];
  assign rd_1r0d[5] = rdfint_1n[5];
  assign rd_1r0d[6] = rdfint_1n[6];
  assign rd_1r0d[7] = rdfint_1n[7];
  assign rd_1r0d[8] = rdfint_1n[8];
  assign rd_1r0d[9] = rdfint_1n[9];
  assign rd_1r0d[10] = rdfint_1n[10];
  assign rd_1r0d[11] = rdfint_1n[11];
  assign rd_1r0d[12] = rdfint_1n[12];
  assign rd_1r0d[13] = rdfint_1n[13];
  assign rd_1r0d[14] = rdfint_1n[14];
  assign rd_1r0d[15] = rdfint_1n[15];
  assign rd_1r0d[16] = rdfint_1n[16];
  assign rd_1r0d[17] = rdfint_1n[17];
  assign rd_1r0d[18] = rdfint_1n[18];
  assign rd_1r0d[19] = rdfint_1n[19];
  assign rd_1r0d[20] = rdfint_1n[20];
  assign rd_1r0d[21] = rdfint_1n[21];
  assign rd_1r0d[22] = rdfint_1n[22];
  assign rd_1r0d[23] = rdfint_1n[23];
  assign rd_1r0d[24] = rdfint_1n[24];
  assign rd_1r0d[25] = rdfint_1n[25];
  assign rd_1r0d[26] = rdfint_1n[26];
  assign rd_1r0d[27] = rdfint_1n[27];
  assign rd_1r0d[28] = rdfint_1n[28];
  assign rd_1r0d[29] = rdfint_1n[29];
  assign rd_1r0d[30] = rdfint_1n[30];
  assign rd_1r0d[31] = rdfint_1n[31];
  assign rd_1r0d[32] = rdfint_1n[32];
  assign rd_1r0d[33] = rdfint_1n[33];
  assign rd_1r0d[34] = rdfint_1n[34];
  assign rd_1r1d[0] = rdtint_1n[0];
  assign rd_1r1d[1] = rdtint_1n[1];
  assign rd_1r1d[2] = rdtint_1n[2];
  assign rd_1r1d[3] = rdtint_1n[3];
  assign rd_1r1d[4] = rdtint_1n[4];
  assign rd_1r1d[5] = rdtint_1n[5];
  assign rd_1r1d[6] = rdtint_1n[6];
  assign rd_1r1d[7] = rdtint_1n[7];
  assign rd_1r1d[8] = rdtint_1n[8];
  assign rd_1r1d[9] = rdtint_1n[9];
  assign rd_1r1d[10] = rdtint_1n[10];
  assign rd_1r1d[11] = rdtint_1n[11];
  assign rd_1r1d[12] = rdtint_1n[12];
  assign rd_1r1d[13] = rdtint_1n[13];
  assign rd_1r1d[14] = rdtint_1n[14];
  assign rd_1r1d[15] = rdtint_1n[15];
  assign rd_1r1d[16] = rdtint_1n[16];
  assign rd_1r1d[17] = rdtint_1n[17];
  assign rd_1r1d[18] = rdtint_1n[18];
  assign rd_1r1d[19] = rdtint_1n[19];
  assign rd_1r1d[20] = rdtint_1n[20];
  assign rd_1r1d[21] = rdtint_1n[21];
  assign rd_1r1d[22] = rdtint_1n[22];
  assign rd_1r1d[23] = rdtint_1n[23];
  assign rd_1r1d[24] = rdtint_1n[24];
  assign rd_1r1d[25] = rdtint_1n[25];
  assign rd_1r1d[26] = rdtint_1n[26];
  assign rd_1r1d[27] = rdtint_1n[27];
  assign rd_1r1d[28] = rdtint_1n[28];
  assign rd_1r1d[29] = rdtint_1n[29];
  assign rd_1r1d[30] = rdtint_1n[30];
  assign rd_1r1d[31] = rdtint_1n[31];
  assign rd_1r1d[32] = rdtint_1n[32];
  assign rd_1r1d[33] = rdtint_1n[33];
  assign rd_1r1d[34] = rdtint_1n[34];
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r0d[10] = rdfint_0n[10];
  assign rd_0r0d[11] = rdfint_0n[11];
  assign rd_0r0d[12] = rdfint_0n[12];
  assign rd_0r0d[13] = rdfint_0n[13];
  assign rd_0r0d[14] = rdfint_0n[14];
  assign rd_0r0d[15] = rdfint_0n[15];
  assign rd_0r0d[16] = rdfint_0n[16];
  assign rd_0r0d[17] = rdfint_0n[17];
  assign rd_0r0d[18] = rdfint_0n[18];
  assign rd_0r0d[19] = rdfint_0n[19];
  assign rd_0r0d[20] = rdfint_0n[20];
  assign rd_0r0d[21] = rdfint_0n[21];
  assign rd_0r0d[22] = rdfint_0n[22];
  assign rd_0r0d[23] = rdfint_0n[23];
  assign rd_0r0d[24] = rdfint_0n[24];
  assign rd_0r0d[25] = rdfint_0n[25];
  assign rd_0r0d[26] = rdfint_0n[26];
  assign rd_0r0d[27] = rdfint_0n[27];
  assign rd_0r0d[28] = rdfint_0n[28];
  assign rd_0r0d[29] = rdfint_0n[29];
  assign rd_0r0d[30] = rdfint_0n[30];
  assign rd_0r0d[31] = rdfint_0n[31];
  assign rd_0r0d[32] = rdfint_0n[32];
  assign rd_0r0d[33] = rdfint_0n[33];
  assign rd_0r0d[34] = rdfint_0n[34];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign rd_0r1d[10] = rdtint_0n[10];
  assign rd_0r1d[11] = rdtint_0n[11];
  assign rd_0r1d[12] = rdtint_0n[12];
  assign rd_0r1d[13] = rdtint_0n[13];
  assign rd_0r1d[14] = rdtint_0n[14];
  assign rd_0r1d[15] = rdtint_0n[15];
  assign rd_0r1d[16] = rdtint_0n[16];
  assign rd_0r1d[17] = rdtint_0n[17];
  assign rd_0r1d[18] = rdtint_0n[18];
  assign rd_0r1d[19] = rdtint_0n[19];
  assign rd_0r1d[20] = rdtint_0n[20];
  assign rd_0r1d[21] = rdtint_0n[21];
  assign rd_0r1d[22] = rdtint_0n[22];
  assign rd_0r1d[23] = rdtint_0n[23];
  assign rd_0r1d[24] = rdtint_0n[24];
  assign rd_0r1d[25] = rdtint_0n[25];
  assign rd_0r1d[26] = rdtint_0n[26];
  assign rd_0r1d[27] = rdtint_0n[27];
  assign rd_0r1d[28] = rdtint_0n[28];
  assign rd_0r1d[29] = rdtint_0n[29];
  assign rd_0r1d[30] = rdtint_0n[30];
  assign rd_0r1d[31] = rdtint_0n[31];
  assign rd_0r1d[32] = rdtint_0n[32];
  assign rd_0r1d[33] = rdtint_0n[33];
  assign rd_0r1d[34] = rdtint_0n[34];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgfint_0n[32] = wg_0r0d[32];
  assign wgfint_0n[33] = wg_0r0d[33];
  assign wgfint_0n[34] = wg_0r0d[34];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign wgtint_0n[32] = wg_0r1d[32];
  assign wgtint_0n[33] = wg_0r1d[33];
  assign wgtint_0n[34] = wg_0r1d[34];
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I219 (internal_0n[0], rgrint_0n, rgrint_1n);
  NOR2 I220 (internal_0n[1], rgaint_0n, rgaint_1n);
  AND2 I221 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I222 (rdtint_1n[0], rgrint_1n, dt_0n[0]);
  AND2 I223 (rdtint_1n[1], rgrint_1n, dt_0n[1]);
  AND2 I224 (rdtint_1n[2], rgrint_1n, dt_0n[2]);
  AND2 I225 (rdtint_1n[3], rgrint_1n, dt_0n[3]);
  AND2 I226 (rdtint_1n[4], rgrint_1n, dt_0n[4]);
  AND2 I227 (rdtint_1n[5], rgrint_1n, dt_0n[5]);
  AND2 I228 (rdtint_1n[6], rgrint_1n, dt_0n[6]);
  AND2 I229 (rdtint_1n[7], rgrint_1n, dt_0n[7]);
  AND2 I230 (rdtint_1n[8], rgrint_1n, dt_0n[8]);
  AND2 I231 (rdtint_1n[9], rgrint_1n, dt_0n[9]);
  AND2 I232 (rdtint_1n[10], rgrint_1n, dt_0n[10]);
  AND2 I233 (rdtint_1n[11], rgrint_1n, dt_0n[11]);
  AND2 I234 (rdtint_1n[12], rgrint_1n, dt_0n[12]);
  AND2 I235 (rdtint_1n[13], rgrint_1n, dt_0n[13]);
  AND2 I236 (rdtint_1n[14], rgrint_1n, dt_0n[14]);
  AND2 I237 (rdtint_1n[15], rgrint_1n, dt_0n[15]);
  AND2 I238 (rdtint_1n[16], rgrint_1n, dt_0n[16]);
  AND2 I239 (rdtint_1n[17], rgrint_1n, dt_0n[17]);
  AND2 I240 (rdtint_1n[18], rgrint_1n, dt_0n[18]);
  AND2 I241 (rdtint_1n[19], rgrint_1n, dt_0n[19]);
  AND2 I242 (rdtint_1n[20], rgrint_1n, dt_0n[20]);
  AND2 I243 (rdtint_1n[21], rgrint_1n, dt_0n[21]);
  AND2 I244 (rdtint_1n[22], rgrint_1n, dt_0n[22]);
  AND2 I245 (rdtint_1n[23], rgrint_1n, dt_0n[23]);
  AND2 I246 (rdtint_1n[24], rgrint_1n, dt_0n[24]);
  AND2 I247 (rdtint_1n[25], rgrint_1n, dt_0n[25]);
  AND2 I248 (rdtint_1n[26], rgrint_1n, dt_0n[26]);
  AND2 I249 (rdtint_1n[27], rgrint_1n, dt_0n[27]);
  AND2 I250 (rdtint_1n[28], rgrint_1n, dt_0n[28]);
  AND2 I251 (rdtint_1n[29], rgrint_1n, dt_0n[29]);
  AND2 I252 (rdtint_1n[30], rgrint_1n, dt_0n[30]);
  AND2 I253 (rdtint_1n[31], rgrint_1n, dt_0n[31]);
  AND2 I254 (rdtint_1n[32], rgrint_1n, dt_0n[32]);
  AND2 I255 (rdtint_1n[33], rgrint_1n, dt_0n[33]);
  AND2 I256 (rdtint_1n[34], rgrint_1n, dt_0n[34]);
  AND2 I257 (rdtint_0n[0], rgrint_0n, dt_0n[0]);
  AND2 I258 (rdtint_0n[1], rgrint_0n, dt_0n[1]);
  AND2 I259 (rdtint_0n[2], rgrint_0n, dt_0n[2]);
  AND2 I260 (rdtint_0n[3], rgrint_0n, dt_0n[3]);
  AND2 I261 (rdtint_0n[4], rgrint_0n, dt_0n[4]);
  AND2 I262 (rdtint_0n[5], rgrint_0n, dt_0n[5]);
  AND2 I263 (rdtint_0n[6], rgrint_0n, dt_0n[6]);
  AND2 I264 (rdtint_0n[7], rgrint_0n, dt_0n[7]);
  AND2 I265 (rdtint_0n[8], rgrint_0n, dt_0n[8]);
  AND2 I266 (rdtint_0n[9], rgrint_0n, dt_0n[9]);
  AND2 I267 (rdtint_0n[10], rgrint_0n, dt_0n[10]);
  AND2 I268 (rdtint_0n[11], rgrint_0n, dt_0n[11]);
  AND2 I269 (rdtint_0n[12], rgrint_0n, dt_0n[12]);
  AND2 I270 (rdtint_0n[13], rgrint_0n, dt_0n[13]);
  AND2 I271 (rdtint_0n[14], rgrint_0n, dt_0n[14]);
  AND2 I272 (rdtint_0n[15], rgrint_0n, dt_0n[15]);
  AND2 I273 (rdtint_0n[16], rgrint_0n, dt_0n[16]);
  AND2 I274 (rdtint_0n[17], rgrint_0n, dt_0n[17]);
  AND2 I275 (rdtint_0n[18], rgrint_0n, dt_0n[18]);
  AND2 I276 (rdtint_0n[19], rgrint_0n, dt_0n[19]);
  AND2 I277 (rdtint_0n[20], rgrint_0n, dt_0n[20]);
  AND2 I278 (rdtint_0n[21], rgrint_0n, dt_0n[21]);
  AND2 I279 (rdtint_0n[22], rgrint_0n, dt_0n[22]);
  AND2 I280 (rdtint_0n[23], rgrint_0n, dt_0n[23]);
  AND2 I281 (rdtint_0n[24], rgrint_0n, dt_0n[24]);
  AND2 I282 (rdtint_0n[25], rgrint_0n, dt_0n[25]);
  AND2 I283 (rdtint_0n[26], rgrint_0n, dt_0n[26]);
  AND2 I284 (rdtint_0n[27], rgrint_0n, dt_0n[27]);
  AND2 I285 (rdtint_0n[28], rgrint_0n, dt_0n[28]);
  AND2 I286 (rdtint_0n[29], rgrint_0n, dt_0n[29]);
  AND2 I287 (rdtint_0n[30], rgrint_0n, dt_0n[30]);
  AND2 I288 (rdtint_0n[31], rgrint_0n, dt_0n[31]);
  AND2 I289 (rdtint_0n[32], rgrint_0n, dt_0n[32]);
  AND2 I290 (rdtint_0n[33], rgrint_0n, dt_0n[33]);
  AND2 I291 (rdtint_0n[34], rgrint_0n, dt_0n[34]);
  AND2 I292 (rdfint_1n[0], rgrint_1n, df_0n[0]);
  AND2 I293 (rdfint_1n[1], rgrint_1n, df_0n[1]);
  AND2 I294 (rdfint_1n[2], rgrint_1n, df_0n[2]);
  AND2 I295 (rdfint_1n[3], rgrint_1n, df_0n[3]);
  AND2 I296 (rdfint_1n[4], rgrint_1n, df_0n[4]);
  AND2 I297 (rdfint_1n[5], rgrint_1n, df_0n[5]);
  AND2 I298 (rdfint_1n[6], rgrint_1n, df_0n[6]);
  AND2 I299 (rdfint_1n[7], rgrint_1n, df_0n[7]);
  AND2 I300 (rdfint_1n[8], rgrint_1n, df_0n[8]);
  AND2 I301 (rdfint_1n[9], rgrint_1n, df_0n[9]);
  AND2 I302 (rdfint_1n[10], rgrint_1n, df_0n[10]);
  AND2 I303 (rdfint_1n[11], rgrint_1n, df_0n[11]);
  AND2 I304 (rdfint_1n[12], rgrint_1n, df_0n[12]);
  AND2 I305 (rdfint_1n[13], rgrint_1n, df_0n[13]);
  AND2 I306 (rdfint_1n[14], rgrint_1n, df_0n[14]);
  AND2 I307 (rdfint_1n[15], rgrint_1n, df_0n[15]);
  AND2 I308 (rdfint_1n[16], rgrint_1n, df_0n[16]);
  AND2 I309 (rdfint_1n[17], rgrint_1n, df_0n[17]);
  AND2 I310 (rdfint_1n[18], rgrint_1n, df_0n[18]);
  AND2 I311 (rdfint_1n[19], rgrint_1n, df_0n[19]);
  AND2 I312 (rdfint_1n[20], rgrint_1n, df_0n[20]);
  AND2 I313 (rdfint_1n[21], rgrint_1n, df_0n[21]);
  AND2 I314 (rdfint_1n[22], rgrint_1n, df_0n[22]);
  AND2 I315 (rdfint_1n[23], rgrint_1n, df_0n[23]);
  AND2 I316 (rdfint_1n[24], rgrint_1n, df_0n[24]);
  AND2 I317 (rdfint_1n[25], rgrint_1n, df_0n[25]);
  AND2 I318 (rdfint_1n[26], rgrint_1n, df_0n[26]);
  AND2 I319 (rdfint_1n[27], rgrint_1n, df_0n[27]);
  AND2 I320 (rdfint_1n[28], rgrint_1n, df_0n[28]);
  AND2 I321 (rdfint_1n[29], rgrint_1n, df_0n[29]);
  AND2 I322 (rdfint_1n[30], rgrint_1n, df_0n[30]);
  AND2 I323 (rdfint_1n[31], rgrint_1n, df_0n[31]);
  AND2 I324 (rdfint_1n[32], rgrint_1n, df_0n[32]);
  AND2 I325 (rdfint_1n[33], rgrint_1n, df_0n[33]);
  AND2 I326 (rdfint_1n[34], rgrint_1n, df_0n[34]);
  AND2 I327 (rdfint_0n[0], rgrint_0n, df_0n[0]);
  AND2 I328 (rdfint_0n[1], rgrint_0n, df_0n[1]);
  AND2 I329 (rdfint_0n[2], rgrint_0n, df_0n[2]);
  AND2 I330 (rdfint_0n[3], rgrint_0n, df_0n[3]);
  AND2 I331 (rdfint_0n[4], rgrint_0n, df_0n[4]);
  AND2 I332 (rdfint_0n[5], rgrint_0n, df_0n[5]);
  AND2 I333 (rdfint_0n[6], rgrint_0n, df_0n[6]);
  AND2 I334 (rdfint_0n[7], rgrint_0n, df_0n[7]);
  AND2 I335 (rdfint_0n[8], rgrint_0n, df_0n[8]);
  AND2 I336 (rdfint_0n[9], rgrint_0n, df_0n[9]);
  AND2 I337 (rdfint_0n[10], rgrint_0n, df_0n[10]);
  AND2 I338 (rdfint_0n[11], rgrint_0n, df_0n[11]);
  AND2 I339 (rdfint_0n[12], rgrint_0n, df_0n[12]);
  AND2 I340 (rdfint_0n[13], rgrint_0n, df_0n[13]);
  AND2 I341 (rdfint_0n[14], rgrint_0n, df_0n[14]);
  AND2 I342 (rdfint_0n[15], rgrint_0n, df_0n[15]);
  AND2 I343 (rdfint_0n[16], rgrint_0n, df_0n[16]);
  AND2 I344 (rdfint_0n[17], rgrint_0n, df_0n[17]);
  AND2 I345 (rdfint_0n[18], rgrint_0n, df_0n[18]);
  AND2 I346 (rdfint_0n[19], rgrint_0n, df_0n[19]);
  AND2 I347 (rdfint_0n[20], rgrint_0n, df_0n[20]);
  AND2 I348 (rdfint_0n[21], rgrint_0n, df_0n[21]);
  AND2 I349 (rdfint_0n[22], rgrint_0n, df_0n[22]);
  AND2 I350 (rdfint_0n[23], rgrint_0n, df_0n[23]);
  AND2 I351 (rdfint_0n[24], rgrint_0n, df_0n[24]);
  AND2 I352 (rdfint_0n[25], rgrint_0n, df_0n[25]);
  AND2 I353 (rdfint_0n[26], rgrint_0n, df_0n[26]);
  AND2 I354 (rdfint_0n[27], rgrint_0n, df_0n[27]);
  AND2 I355 (rdfint_0n[28], rgrint_0n, df_0n[28]);
  AND2 I356 (rdfint_0n[29], rgrint_0n, df_0n[29]);
  AND2 I357 (rdfint_0n[30], rgrint_0n, df_0n[30]);
  AND2 I358 (rdfint_0n[31], rgrint_0n, df_0n[31]);
  AND2 I359 (rdfint_0n[32], rgrint_0n, df_0n[32]);
  AND2 I360 (rdfint_0n[33], rgrint_0n, df_0n[33]);
  AND2 I361 (rdfint_0n[34], rgrint_0n, df_0n[34]);
  C3 I362 (internal_0n[2], wc_0n, wacks_0n[34], wacks_0n[33]);
  C3 I363 (internal_0n[3], wacks_0n[32], wacks_0n[31], wacks_0n[30]);
  C3 I364 (internal_0n[4], wacks_0n[29], wacks_0n[28], wacks_0n[27]);
  C3 I365 (internal_0n[5], wacks_0n[26], wacks_0n[25], wacks_0n[24]);
  C3 I366 (internal_0n[6], wacks_0n[23], wacks_0n[22], wacks_0n[21]);
  C3 I367 (internal_0n[7], wacks_0n[20], wacks_0n[19], wacks_0n[18]);
  C3 I368 (internal_0n[8], wacks_0n[17], wacks_0n[16], wacks_0n[15]);
  C3 I369 (internal_0n[9], wacks_0n[14], wacks_0n[13], wacks_0n[12]);
  C3 I370 (internal_0n[10], wacks_0n[11], wacks_0n[10], wacks_0n[9]);
  C3 I371 (internal_0n[11], wacks_0n[8], wacks_0n[7], wacks_0n[6]);
  C3 I372 (internal_0n[12], wacks_0n[5], wacks_0n[4], wacks_0n[3]);
  C3 I373 (internal_0n[13], wacks_0n[2], wacks_0n[1], wacks_0n[0]);
  C3 I374 (internal_0n[14], internal_0n[2], internal_0n[3], internal_0n[4]);
  C3 I375 (internal_0n[15], internal_0n[5], internal_0n[6], internal_0n[7]);
  C3 I376 (internal_0n[16], internal_0n[8], internal_0n[9], internal_0n[10]);
  C3 I377 (internal_0n[17], internal_0n[11], internal_0n[12], internal_0n[13]);
  C2 I378 (internal_0n[18], internal_0n[14], internal_0n[15]);
  C2 I379 (internal_0n[19], internal_0n[16], internal_0n[17]);
  C2 I380 (wdrint_0n, internal_0n[18], internal_0n[19]);
  assign wen_0n[34] = wc_0n;
  assign wen_0n[33] = wc_0n;
  assign wen_0n[32] = wc_0n;
  assign wen_0n[31] = wc_0n;
  assign wen_0n[30] = wc_0n;
  assign wen_0n[29] = wc_0n;
  assign wen_0n[28] = wc_0n;
  assign wen_0n[27] = wc_0n;
  assign wen_0n[26] = wc_0n;
  assign wen_0n[25] = wc_0n;
  assign wen_0n[24] = wc_0n;
  assign wen_0n[23] = wc_0n;
  assign wen_0n[22] = wc_0n;
  assign wen_0n[21] = wc_0n;
  assign wen_0n[20] = wc_0n;
  assign wen_0n[19] = wc_0n;
  assign wen_0n[18] = wc_0n;
  assign wen_0n[17] = wc_0n;
  assign wen_0n[16] = wc_0n;
  assign wen_0n[15] = wc_0n;
  assign wen_0n[14] = wc_0n;
  assign wen_0n[13] = wc_0n;
  assign wen_0n[12] = wc_0n;
  assign wen_0n[11] = wc_0n;
  assign wen_0n[10] = wc_0n;
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[34] = git_0n[34];
  assign wt_0n[33] = git_0n[33];
  assign wt_0n[32] = git_0n[32];
  assign wt_0n[31] = git_0n[31];
  assign wt_0n[30] = git_0n[30];
  assign wt_0n[29] = git_0n[29];
  assign wt_0n[28] = git_0n[28];
  assign wt_0n[27] = git_0n[27];
  assign wt_0n[26] = git_0n[26];
  assign wt_0n[25] = git_0n[25];
  assign wt_0n[24] = git_0n[24];
  assign wt_0n[23] = git_0n[23];
  assign wt_0n[22] = git_0n[22];
  assign wt_0n[21] = git_0n[21];
  assign wt_0n[20] = git_0n[20];
  assign wt_0n[19] = git_0n[19];
  assign wt_0n[18] = git_0n[18];
  assign wt_0n[17] = git_0n[17];
  assign wt_0n[16] = git_0n[16];
  assign wt_0n[15] = git_0n[15];
  assign wt_0n[14] = git_0n[14];
  assign wt_0n[13] = git_0n[13];
  assign wt_0n[12] = git_0n[12];
  assign wt_0n[11] = git_0n[11];
  assign wt_0n[10] = git_0n[10];
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[34] = gif_0n[34];
  assign wf_0n[33] = gif_0n[33];
  assign wf_0n[32] = gif_0n[32];
  assign wf_0n[31] = gif_0n[31];
  assign wf_0n[30] = gif_0n[30];
  assign wf_0n[29] = gif_0n[29];
  assign wf_0n[28] = gif_0n[28];
  assign wf_0n[27] = gif_0n[27];
  assign wf_0n[26] = gif_0n[26];
  assign wf_0n[25] = gif_0n[25];
  assign wf_0n[24] = gif_0n[24];
  assign wf_0n[23] = gif_0n[23];
  assign wf_0n[22] = gif_0n[22];
  assign wf_0n[21] = gif_0n[21];
  assign wf_0n[20] = gif_0n[20];
  assign wf_0n[19] = gif_0n[19];
  assign wf_0n[18] = gif_0n[18];
  assign wf_0n[17] = gif_0n[17];
  assign wf_0n[16] = gif_0n[16];
  assign wf_0n[15] = gif_0n[15];
  assign wf_0n[14] = gif_0n[14];
  assign wf_0n[13] = gif_0n[13];
  assign wf_0n[12] = gif_0n[12];
  assign wf_0n[11] = gif_0n[11];
  assign wf_0n[10] = gif_0n[10];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I486 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I488 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I489 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I490 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I491 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I492 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I493 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I494 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I495 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I496 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I497 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I498 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I499 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I500 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I501 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I502 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I503 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I504 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I505 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I506 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I507 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I508 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I509 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I510 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I511 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I512 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I513 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I514 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I515 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I516 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I517 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I518 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I519 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I520 (git_0n[32], wgtint_0n[32], ig_0n);
  AND2 I521 (git_0n[33], wgtint_0n[33], ig_0n);
  AND2 I522 (git_0n[34], wgtint_0n[34], ig_0n);
  AND2 I523 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I524 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I525 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I526 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I527 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I528 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I529 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I530 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I531 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I532 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I533 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I534 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I535 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I536 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I537 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I538 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I539 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I540 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I541 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I542 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I543 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I544 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I545 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I546 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I547 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I548 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I549 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I550 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I551 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I552 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I553 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I554 (gif_0n[31], wgfint_0n[31], ig_0n);
  AND2 I555 (gif_0n[32], wgfint_0n[32], ig_0n);
  AND2 I556 (gif_0n[33], wgfint_0n[33], ig_0n);
  AND2 I557 (gif_0n[34], wgfint_0n[34], ig_0n);
  C3 I558 (internal_0n[20], complete1486_0n[0], complete1486_0n[1], complete1486_0n[2]);
  C3 I559 (internal_0n[21], complete1486_0n[3], complete1486_0n[4], complete1486_0n[5]);
  C3 I560 (internal_0n[22], complete1486_0n[6], complete1486_0n[7], complete1486_0n[8]);
  C3 I561 (internal_0n[23], complete1486_0n[9], complete1486_0n[10], complete1486_0n[11]);
  C3 I562 (internal_0n[24], complete1486_0n[12], complete1486_0n[13], complete1486_0n[14]);
  C3 I563 (internal_0n[25], complete1486_0n[15], complete1486_0n[16], complete1486_0n[17]);
  C3 I564 (internal_0n[26], complete1486_0n[18], complete1486_0n[19], complete1486_0n[20]);
  C3 I565 (internal_0n[27], complete1486_0n[21], complete1486_0n[22], complete1486_0n[23]);
  C3 I566 (internal_0n[28], complete1486_0n[24], complete1486_0n[25], complete1486_0n[26]);
  C3 I567 (internal_0n[29], complete1486_0n[27], complete1486_0n[28], complete1486_0n[29]);
  C3 I568 (internal_0n[30], complete1486_0n[30], complete1486_0n[31], complete1486_0n[32]);
  C2 I569 (internal_0n[31], complete1486_0n[33], complete1486_0n[34]);
  C3 I570 (internal_0n[32], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I571 (internal_0n[33], internal_0n[23], internal_0n[24], internal_0n[25]);
  C3 I572 (internal_0n[34], internal_0n[26], internal_0n[27], internal_0n[28]);
  C3 I573 (internal_0n[35], internal_0n[29], internal_0n[30], internal_0n[31]);
  C2 I574 (internal_0n[36], internal_0n[32], internal_0n[33]);
  C2 I575 (internal_0n[37], internal_0n[34], internal_0n[35]);
  C2 I576 (wc_0n, internal_0n[36], internal_0n[37]);
  OR2 I577 (complete1486_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I578 (complete1486_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I579 (complete1486_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I580 (complete1486_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I581 (complete1486_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I582 (complete1486_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I583 (complete1486_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I584 (complete1486_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I585 (complete1486_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I586 (complete1486_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I587 (complete1486_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I588 (complete1486_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I589 (complete1486_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I590 (complete1486_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I591 (complete1486_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I592 (complete1486_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I593 (complete1486_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I594 (complete1486_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I595 (complete1486_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I596 (complete1486_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I597 (complete1486_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I598 (complete1486_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I599 (complete1486_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I600 (complete1486_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I601 (complete1486_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I602 (complete1486_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I603 (complete1486_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I604 (complete1486_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I605 (complete1486_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I606 (complete1486_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I607 (complete1486_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I608 (complete1486_0n[31], wgfint_0n[31], wgtint_0n[31]);
  OR2 I609 (complete1486_0n[32], wgfint_0n[32], wgtint_0n[32]);
  OR2 I610 (complete1486_0n[33], wgfint_0n[33], wgtint_0n[33]);
  OR2 I611 (complete1486_0n[34], wgfint_0n[34], wgtint_0n[34]);
  AO22 I612 (wacks_0n[34], gf1484_0n[34], df_0n[34], gt1485_0n[34], dt_0n[34]);
  NOR2 I613 (dt_0n[34], df_0n[34], gf1484_0n[34]);
  NOR3 I614 (df_0n[34], dt_0n[34], gt1485_0n[34], init_0n);
  AND2 I615 (gt1485_0n[34], wt_0n[34], wen_0n[34]);
  AND2 I616 (gf1484_0n[34], wf_0n[34], wen_0n[34]);
  AO22 I617 (wacks_0n[33], gf1484_0n[33], df_0n[33], gt1485_0n[33], dt_0n[33]);
  NOR2 I618 (dt_0n[33], df_0n[33], gf1484_0n[33]);
  NOR3 I619 (df_0n[33], dt_0n[33], gt1485_0n[33], init_0n);
  AND2 I620 (gt1485_0n[33], wt_0n[33], wen_0n[33]);
  AND2 I621 (gf1484_0n[33], wf_0n[33], wen_0n[33]);
  AO22 I622 (wacks_0n[32], gf1484_0n[32], df_0n[32], gt1485_0n[32], dt_0n[32]);
  NOR2 I623 (dt_0n[32], df_0n[32], gf1484_0n[32]);
  NOR3 I624 (df_0n[32], dt_0n[32], gt1485_0n[32], init_0n);
  AND2 I625 (gt1485_0n[32], wt_0n[32], wen_0n[32]);
  AND2 I626 (gf1484_0n[32], wf_0n[32], wen_0n[32]);
  AO22 I627 (wacks_0n[31], gf1484_0n[31], df_0n[31], gt1485_0n[31], dt_0n[31]);
  NOR2 I628 (dt_0n[31], df_0n[31], gf1484_0n[31]);
  NOR3 I629 (df_0n[31], dt_0n[31], gt1485_0n[31], init_0n);
  AND2 I630 (gt1485_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I631 (gf1484_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I632 (wacks_0n[30], gf1484_0n[30], df_0n[30], gt1485_0n[30], dt_0n[30]);
  NOR2 I633 (dt_0n[30], df_0n[30], gf1484_0n[30]);
  NOR3 I634 (df_0n[30], dt_0n[30], gt1485_0n[30], init_0n);
  AND2 I635 (gt1485_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I636 (gf1484_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I637 (wacks_0n[29], gf1484_0n[29], df_0n[29], gt1485_0n[29], dt_0n[29]);
  NOR2 I638 (dt_0n[29], df_0n[29], gf1484_0n[29]);
  NOR3 I639 (df_0n[29], dt_0n[29], gt1485_0n[29], init_0n);
  AND2 I640 (gt1485_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I641 (gf1484_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I642 (wacks_0n[28], gf1484_0n[28], df_0n[28], gt1485_0n[28], dt_0n[28]);
  NOR2 I643 (dt_0n[28], df_0n[28], gf1484_0n[28]);
  NOR3 I644 (df_0n[28], dt_0n[28], gt1485_0n[28], init_0n);
  AND2 I645 (gt1485_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I646 (gf1484_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I647 (wacks_0n[27], gf1484_0n[27], df_0n[27], gt1485_0n[27], dt_0n[27]);
  NOR2 I648 (dt_0n[27], df_0n[27], gf1484_0n[27]);
  NOR3 I649 (df_0n[27], dt_0n[27], gt1485_0n[27], init_0n);
  AND2 I650 (gt1485_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I651 (gf1484_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I652 (wacks_0n[26], gf1484_0n[26], df_0n[26], gt1485_0n[26], dt_0n[26]);
  NOR2 I653 (dt_0n[26], df_0n[26], gf1484_0n[26]);
  NOR3 I654 (df_0n[26], dt_0n[26], gt1485_0n[26], init_0n);
  AND2 I655 (gt1485_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I656 (gf1484_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I657 (wacks_0n[25], gf1484_0n[25], df_0n[25], gt1485_0n[25], dt_0n[25]);
  NOR2 I658 (dt_0n[25], df_0n[25], gf1484_0n[25]);
  NOR3 I659 (df_0n[25], dt_0n[25], gt1485_0n[25], init_0n);
  AND2 I660 (gt1485_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I661 (gf1484_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I662 (wacks_0n[24], gf1484_0n[24], df_0n[24], gt1485_0n[24], dt_0n[24]);
  NOR2 I663 (dt_0n[24], df_0n[24], gf1484_0n[24]);
  NOR3 I664 (df_0n[24], dt_0n[24], gt1485_0n[24], init_0n);
  AND2 I665 (gt1485_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I666 (gf1484_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I667 (wacks_0n[23], gf1484_0n[23], df_0n[23], gt1485_0n[23], dt_0n[23]);
  NOR2 I668 (dt_0n[23], df_0n[23], gf1484_0n[23]);
  NOR3 I669 (df_0n[23], dt_0n[23], gt1485_0n[23], init_0n);
  AND2 I670 (gt1485_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I671 (gf1484_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I672 (wacks_0n[22], gf1484_0n[22], df_0n[22], gt1485_0n[22], dt_0n[22]);
  NOR2 I673 (dt_0n[22], df_0n[22], gf1484_0n[22]);
  NOR3 I674 (df_0n[22], dt_0n[22], gt1485_0n[22], init_0n);
  AND2 I675 (gt1485_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I676 (gf1484_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I677 (wacks_0n[21], gf1484_0n[21], df_0n[21], gt1485_0n[21], dt_0n[21]);
  NOR2 I678 (dt_0n[21], df_0n[21], gf1484_0n[21]);
  NOR3 I679 (df_0n[21], dt_0n[21], gt1485_0n[21], init_0n);
  AND2 I680 (gt1485_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I681 (gf1484_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I682 (wacks_0n[20], gf1484_0n[20], df_0n[20], gt1485_0n[20], dt_0n[20]);
  NOR2 I683 (dt_0n[20], df_0n[20], gf1484_0n[20]);
  NOR3 I684 (df_0n[20], dt_0n[20], gt1485_0n[20], init_0n);
  AND2 I685 (gt1485_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I686 (gf1484_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I687 (wacks_0n[19], gf1484_0n[19], df_0n[19], gt1485_0n[19], dt_0n[19]);
  NOR2 I688 (dt_0n[19], df_0n[19], gf1484_0n[19]);
  NOR3 I689 (df_0n[19], dt_0n[19], gt1485_0n[19], init_0n);
  AND2 I690 (gt1485_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I691 (gf1484_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I692 (wacks_0n[18], gf1484_0n[18], df_0n[18], gt1485_0n[18], dt_0n[18]);
  NOR2 I693 (dt_0n[18], df_0n[18], gf1484_0n[18]);
  NOR3 I694 (df_0n[18], dt_0n[18], gt1485_0n[18], init_0n);
  AND2 I695 (gt1485_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I696 (gf1484_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I697 (wacks_0n[17], gf1484_0n[17], df_0n[17], gt1485_0n[17], dt_0n[17]);
  NOR2 I698 (dt_0n[17], df_0n[17], gf1484_0n[17]);
  NOR3 I699 (df_0n[17], dt_0n[17], gt1485_0n[17], init_0n);
  AND2 I700 (gt1485_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I701 (gf1484_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I702 (wacks_0n[16], gf1484_0n[16], df_0n[16], gt1485_0n[16], dt_0n[16]);
  NOR2 I703 (dt_0n[16], df_0n[16], gf1484_0n[16]);
  NOR3 I704 (df_0n[16], dt_0n[16], gt1485_0n[16], init_0n);
  AND2 I705 (gt1485_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I706 (gf1484_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I707 (wacks_0n[15], gf1484_0n[15], df_0n[15], gt1485_0n[15], dt_0n[15]);
  NOR2 I708 (dt_0n[15], df_0n[15], gf1484_0n[15]);
  NOR3 I709 (df_0n[15], dt_0n[15], gt1485_0n[15], init_0n);
  AND2 I710 (gt1485_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I711 (gf1484_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I712 (wacks_0n[14], gf1484_0n[14], df_0n[14], gt1485_0n[14], dt_0n[14]);
  NOR2 I713 (dt_0n[14], df_0n[14], gf1484_0n[14]);
  NOR3 I714 (df_0n[14], dt_0n[14], gt1485_0n[14], init_0n);
  AND2 I715 (gt1485_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I716 (gf1484_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I717 (wacks_0n[13], gf1484_0n[13], df_0n[13], gt1485_0n[13], dt_0n[13]);
  NOR2 I718 (dt_0n[13], df_0n[13], gf1484_0n[13]);
  NOR3 I719 (df_0n[13], dt_0n[13], gt1485_0n[13], init_0n);
  AND2 I720 (gt1485_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I721 (gf1484_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I722 (wacks_0n[12], gf1484_0n[12], df_0n[12], gt1485_0n[12], dt_0n[12]);
  NOR2 I723 (dt_0n[12], df_0n[12], gf1484_0n[12]);
  NOR3 I724 (df_0n[12], dt_0n[12], gt1485_0n[12], init_0n);
  AND2 I725 (gt1485_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I726 (gf1484_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I727 (wacks_0n[11], gf1484_0n[11], df_0n[11], gt1485_0n[11], dt_0n[11]);
  NOR2 I728 (dt_0n[11], df_0n[11], gf1484_0n[11]);
  NOR3 I729 (df_0n[11], dt_0n[11], gt1485_0n[11], init_0n);
  AND2 I730 (gt1485_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I731 (gf1484_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I732 (wacks_0n[10], gf1484_0n[10], df_0n[10], gt1485_0n[10], dt_0n[10]);
  NOR2 I733 (dt_0n[10], df_0n[10], gf1484_0n[10]);
  NOR3 I734 (df_0n[10], dt_0n[10], gt1485_0n[10], init_0n);
  AND2 I735 (gt1485_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I736 (gf1484_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I737 (wacks_0n[9], gf1484_0n[9], df_0n[9], gt1485_0n[9], dt_0n[9]);
  NOR2 I738 (dt_0n[9], df_0n[9], gf1484_0n[9]);
  NOR3 I739 (df_0n[9], dt_0n[9], gt1485_0n[9], init_0n);
  AND2 I740 (gt1485_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I741 (gf1484_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I742 (wacks_0n[8], gf1484_0n[8], df_0n[8], gt1485_0n[8], dt_0n[8]);
  NOR2 I743 (dt_0n[8], df_0n[8], gf1484_0n[8]);
  NOR3 I744 (df_0n[8], dt_0n[8], gt1485_0n[8], init_0n);
  AND2 I745 (gt1485_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I746 (gf1484_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I747 (wacks_0n[7], gf1484_0n[7], df_0n[7], gt1485_0n[7], dt_0n[7]);
  NOR2 I748 (dt_0n[7], df_0n[7], gf1484_0n[7]);
  NOR3 I749 (df_0n[7], dt_0n[7], gt1485_0n[7], init_0n);
  AND2 I750 (gt1485_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I751 (gf1484_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I752 (wacks_0n[6], gf1484_0n[6], df_0n[6], gt1485_0n[6], dt_0n[6]);
  NOR2 I753 (dt_0n[6], df_0n[6], gf1484_0n[6]);
  NOR3 I754 (df_0n[6], dt_0n[6], gt1485_0n[6], init_0n);
  AND2 I755 (gt1485_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I756 (gf1484_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I757 (wacks_0n[5], gf1484_0n[5], df_0n[5], gt1485_0n[5], dt_0n[5]);
  NOR2 I758 (dt_0n[5], df_0n[5], gf1484_0n[5]);
  NOR3 I759 (df_0n[5], dt_0n[5], gt1485_0n[5], init_0n);
  AND2 I760 (gt1485_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I761 (gf1484_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I762 (wacks_0n[4], gf1484_0n[4], df_0n[4], gt1485_0n[4], dt_0n[4]);
  NOR2 I763 (dt_0n[4], df_0n[4], gf1484_0n[4]);
  NOR3 I764 (df_0n[4], dt_0n[4], gt1485_0n[4], init_0n);
  AND2 I765 (gt1485_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I766 (gf1484_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I767 (wacks_0n[3], gf1484_0n[3], df_0n[3], gt1485_0n[3], dt_0n[3]);
  NOR2 I768 (dt_0n[3], df_0n[3], gf1484_0n[3]);
  NOR3 I769 (df_0n[3], dt_0n[3], gt1485_0n[3], init_0n);
  AND2 I770 (gt1485_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I771 (gf1484_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I772 (wacks_0n[2], gf1484_0n[2], df_0n[2], gt1485_0n[2], dt_0n[2]);
  NOR2 I773 (dt_0n[2], df_0n[2], gf1484_0n[2]);
  NOR3 I774 (df_0n[2], dt_0n[2], gt1485_0n[2], init_0n);
  AND2 I775 (gt1485_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I776 (gf1484_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I777 (wacks_0n[1], gf1484_0n[1], df_0n[1], gt1485_0n[1], dt_0n[1]);
  NOR2 I778 (dt_0n[1], df_0n[1], gf1484_0n[1]);
  NOR3 I779 (df_0n[1], dt_0n[1], gt1485_0n[1], init_0n);
  AND2 I780 (gt1485_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I781 (gf1484_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I782 (wacks_0n[0], gf1484_0n[0], df_0n[0], gt1485_0n[0], dt_0n[0]);
  NOR2 I783 (dt_0n[0], df_0n[0], gf1484_0n[0]);
  NOR3 I784 (df_0n[0], dt_0n[0], gt1485_0n[0], init_0n);
  AND2 I785 (gt1485_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I786 (gf1484_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I787 (init_0n, initialise);
endmodule

module BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m91m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rg_2r, rg_2a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  rd_2r0d, rd_2r1d, rd_2a,
  initialise
);
  input [34:0] wg_0r0d;
  input [34:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [34:0] rd_0r0d;
  output [34:0] rd_0r1d;
  input rd_0a;
  output [34:0] rd_1r0d;
  output [34:0] rd_1r1d;
  input rd_1a;
  output [34:0] rd_2r0d;
  output [34:0] rd_2r1d;
  input rd_2a;
  input initialise;
  wire [37:0] internal_0n;
  wire [34:0] wf_0n;
  wire [34:0] wt_0n;
  wire [34:0] df_0n;
  wire [34:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire rgrint_2n;
  wire wc_0n;
  wire [34:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [34:0] wgfint_0n;
  wire [34:0] wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire rgaint_2n;
  wire [34:0] rdfint_0n;
  wire [34:0] rdfint_1n;
  wire [34:0] rdfint_2n;
  wire [34:0] rdtint_0n;
  wire [34:0] rdtint_1n;
  wire [34:0] rdtint_2n;
  wire [34:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [34:0] gif_0n;
  wire [34:0] git_0n;
  wire [34:0] complete1501_0n;
  wire [34:0] gt1500_0n;
  wire [34:0] gf1499_0n;
  assign rgaint_2n = rd_2a;
  assign rd_2r0d[0] = rdfint_2n[0];
  assign rd_2r0d[1] = rdfint_2n[1];
  assign rd_2r0d[2] = rdfint_2n[2];
  assign rd_2r0d[3] = rdfint_2n[3];
  assign rd_2r0d[4] = rdfint_2n[4];
  assign rd_2r0d[5] = rdfint_2n[5];
  assign rd_2r0d[6] = rdfint_2n[6];
  assign rd_2r0d[7] = rdfint_2n[7];
  assign rd_2r0d[8] = rdfint_2n[8];
  assign rd_2r0d[9] = rdfint_2n[9];
  assign rd_2r0d[10] = rdfint_2n[10];
  assign rd_2r0d[11] = rdfint_2n[11];
  assign rd_2r0d[12] = rdfint_2n[12];
  assign rd_2r0d[13] = rdfint_2n[13];
  assign rd_2r0d[14] = rdfint_2n[14];
  assign rd_2r0d[15] = rdfint_2n[15];
  assign rd_2r0d[16] = rdfint_2n[16];
  assign rd_2r0d[17] = rdfint_2n[17];
  assign rd_2r0d[18] = rdfint_2n[18];
  assign rd_2r0d[19] = rdfint_2n[19];
  assign rd_2r0d[20] = rdfint_2n[20];
  assign rd_2r0d[21] = rdfint_2n[21];
  assign rd_2r0d[22] = rdfint_2n[22];
  assign rd_2r0d[23] = rdfint_2n[23];
  assign rd_2r0d[24] = rdfint_2n[24];
  assign rd_2r0d[25] = rdfint_2n[25];
  assign rd_2r0d[26] = rdfint_2n[26];
  assign rd_2r0d[27] = rdfint_2n[27];
  assign rd_2r0d[28] = rdfint_2n[28];
  assign rd_2r0d[29] = rdfint_2n[29];
  assign rd_2r0d[30] = rdfint_2n[30];
  assign rd_2r0d[31] = rdfint_2n[31];
  assign rd_2r0d[32] = rdfint_2n[32];
  assign rd_2r0d[33] = rdfint_2n[33];
  assign rd_2r0d[34] = rdfint_2n[34];
  assign rd_2r1d[0] = rdtint_2n[0];
  assign rd_2r1d[1] = rdtint_2n[1];
  assign rd_2r1d[2] = rdtint_2n[2];
  assign rd_2r1d[3] = rdtint_2n[3];
  assign rd_2r1d[4] = rdtint_2n[4];
  assign rd_2r1d[5] = rdtint_2n[5];
  assign rd_2r1d[6] = rdtint_2n[6];
  assign rd_2r1d[7] = rdtint_2n[7];
  assign rd_2r1d[8] = rdtint_2n[8];
  assign rd_2r1d[9] = rdtint_2n[9];
  assign rd_2r1d[10] = rdtint_2n[10];
  assign rd_2r1d[11] = rdtint_2n[11];
  assign rd_2r1d[12] = rdtint_2n[12];
  assign rd_2r1d[13] = rdtint_2n[13];
  assign rd_2r1d[14] = rdtint_2n[14];
  assign rd_2r1d[15] = rdtint_2n[15];
  assign rd_2r1d[16] = rdtint_2n[16];
  assign rd_2r1d[17] = rdtint_2n[17];
  assign rd_2r1d[18] = rdtint_2n[18];
  assign rd_2r1d[19] = rdtint_2n[19];
  assign rd_2r1d[20] = rdtint_2n[20];
  assign rd_2r1d[21] = rdtint_2n[21];
  assign rd_2r1d[22] = rdtint_2n[22];
  assign rd_2r1d[23] = rdtint_2n[23];
  assign rd_2r1d[24] = rdtint_2n[24];
  assign rd_2r1d[25] = rdtint_2n[25];
  assign rd_2r1d[26] = rdtint_2n[26];
  assign rd_2r1d[27] = rdtint_2n[27];
  assign rd_2r1d[28] = rdtint_2n[28];
  assign rd_2r1d[29] = rdtint_2n[29];
  assign rd_2r1d[30] = rdtint_2n[30];
  assign rd_2r1d[31] = rdtint_2n[31];
  assign rd_2r1d[32] = rdtint_2n[32];
  assign rd_2r1d[33] = rdtint_2n[33];
  assign rd_2r1d[34] = rdtint_2n[34];
  assign rgaint_1n = rd_1a;
  assign rd_1r0d[0] = rdfint_1n[0];
  assign rd_1r0d[1] = rdfint_1n[1];
  assign rd_1r0d[2] = rdfint_1n[2];
  assign rd_1r0d[3] = rdfint_1n[3];
  assign rd_1r0d[4] = rdfint_1n[4];
  assign rd_1r0d[5] = rdfint_1n[5];
  assign rd_1r0d[6] = rdfint_1n[6];
  assign rd_1r0d[7] = rdfint_1n[7];
  assign rd_1r0d[8] = rdfint_1n[8];
  assign rd_1r0d[9] = rdfint_1n[9];
  assign rd_1r0d[10] = rdfint_1n[10];
  assign rd_1r0d[11] = rdfint_1n[11];
  assign rd_1r0d[12] = rdfint_1n[12];
  assign rd_1r0d[13] = rdfint_1n[13];
  assign rd_1r0d[14] = rdfint_1n[14];
  assign rd_1r0d[15] = rdfint_1n[15];
  assign rd_1r0d[16] = rdfint_1n[16];
  assign rd_1r0d[17] = rdfint_1n[17];
  assign rd_1r0d[18] = rdfint_1n[18];
  assign rd_1r0d[19] = rdfint_1n[19];
  assign rd_1r0d[20] = rdfint_1n[20];
  assign rd_1r0d[21] = rdfint_1n[21];
  assign rd_1r0d[22] = rdfint_1n[22];
  assign rd_1r0d[23] = rdfint_1n[23];
  assign rd_1r0d[24] = rdfint_1n[24];
  assign rd_1r0d[25] = rdfint_1n[25];
  assign rd_1r0d[26] = rdfint_1n[26];
  assign rd_1r0d[27] = rdfint_1n[27];
  assign rd_1r0d[28] = rdfint_1n[28];
  assign rd_1r0d[29] = rdfint_1n[29];
  assign rd_1r0d[30] = rdfint_1n[30];
  assign rd_1r0d[31] = rdfint_1n[31];
  assign rd_1r0d[32] = rdfint_1n[32];
  assign rd_1r0d[33] = rdfint_1n[33];
  assign rd_1r0d[34] = rdfint_1n[34];
  assign rd_1r1d[0] = rdtint_1n[0];
  assign rd_1r1d[1] = rdtint_1n[1];
  assign rd_1r1d[2] = rdtint_1n[2];
  assign rd_1r1d[3] = rdtint_1n[3];
  assign rd_1r1d[4] = rdtint_1n[4];
  assign rd_1r1d[5] = rdtint_1n[5];
  assign rd_1r1d[6] = rdtint_1n[6];
  assign rd_1r1d[7] = rdtint_1n[7];
  assign rd_1r1d[8] = rdtint_1n[8];
  assign rd_1r1d[9] = rdtint_1n[9];
  assign rd_1r1d[10] = rdtint_1n[10];
  assign rd_1r1d[11] = rdtint_1n[11];
  assign rd_1r1d[12] = rdtint_1n[12];
  assign rd_1r1d[13] = rdtint_1n[13];
  assign rd_1r1d[14] = rdtint_1n[14];
  assign rd_1r1d[15] = rdtint_1n[15];
  assign rd_1r1d[16] = rdtint_1n[16];
  assign rd_1r1d[17] = rdtint_1n[17];
  assign rd_1r1d[18] = rdtint_1n[18];
  assign rd_1r1d[19] = rdtint_1n[19];
  assign rd_1r1d[20] = rdtint_1n[20];
  assign rd_1r1d[21] = rdtint_1n[21];
  assign rd_1r1d[22] = rdtint_1n[22];
  assign rd_1r1d[23] = rdtint_1n[23];
  assign rd_1r1d[24] = rdtint_1n[24];
  assign rd_1r1d[25] = rdtint_1n[25];
  assign rd_1r1d[26] = rdtint_1n[26];
  assign rd_1r1d[27] = rdtint_1n[27];
  assign rd_1r1d[28] = rdtint_1n[28];
  assign rd_1r1d[29] = rdtint_1n[29];
  assign rd_1r1d[30] = rdtint_1n[30];
  assign rd_1r1d[31] = rdtint_1n[31];
  assign rd_1r1d[32] = rdtint_1n[32];
  assign rd_1r1d[33] = rdtint_1n[33];
  assign rd_1r1d[34] = rdtint_1n[34];
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r0d[10] = rdfint_0n[10];
  assign rd_0r0d[11] = rdfint_0n[11];
  assign rd_0r0d[12] = rdfint_0n[12];
  assign rd_0r0d[13] = rdfint_0n[13];
  assign rd_0r0d[14] = rdfint_0n[14];
  assign rd_0r0d[15] = rdfint_0n[15];
  assign rd_0r0d[16] = rdfint_0n[16];
  assign rd_0r0d[17] = rdfint_0n[17];
  assign rd_0r0d[18] = rdfint_0n[18];
  assign rd_0r0d[19] = rdfint_0n[19];
  assign rd_0r0d[20] = rdfint_0n[20];
  assign rd_0r0d[21] = rdfint_0n[21];
  assign rd_0r0d[22] = rdfint_0n[22];
  assign rd_0r0d[23] = rdfint_0n[23];
  assign rd_0r0d[24] = rdfint_0n[24];
  assign rd_0r0d[25] = rdfint_0n[25];
  assign rd_0r0d[26] = rdfint_0n[26];
  assign rd_0r0d[27] = rdfint_0n[27];
  assign rd_0r0d[28] = rdfint_0n[28];
  assign rd_0r0d[29] = rdfint_0n[29];
  assign rd_0r0d[30] = rdfint_0n[30];
  assign rd_0r0d[31] = rdfint_0n[31];
  assign rd_0r0d[32] = rdfint_0n[32];
  assign rd_0r0d[33] = rdfint_0n[33];
  assign rd_0r0d[34] = rdfint_0n[34];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign rd_0r1d[10] = rdtint_0n[10];
  assign rd_0r1d[11] = rdtint_0n[11];
  assign rd_0r1d[12] = rdtint_0n[12];
  assign rd_0r1d[13] = rdtint_0n[13];
  assign rd_0r1d[14] = rdtint_0n[14];
  assign rd_0r1d[15] = rdtint_0n[15];
  assign rd_0r1d[16] = rdtint_0n[16];
  assign rd_0r1d[17] = rdtint_0n[17];
  assign rd_0r1d[18] = rdtint_0n[18];
  assign rd_0r1d[19] = rdtint_0n[19];
  assign rd_0r1d[20] = rdtint_0n[20];
  assign rd_0r1d[21] = rdtint_0n[21];
  assign rd_0r1d[22] = rdtint_0n[22];
  assign rd_0r1d[23] = rdtint_0n[23];
  assign rd_0r1d[24] = rdtint_0n[24];
  assign rd_0r1d[25] = rdtint_0n[25];
  assign rd_0r1d[26] = rdtint_0n[26];
  assign rd_0r1d[27] = rdtint_0n[27];
  assign rd_0r1d[28] = rdtint_0n[28];
  assign rd_0r1d[29] = rdtint_0n[29];
  assign rd_0r1d[30] = rdtint_0n[30];
  assign rd_0r1d[31] = rdtint_0n[31];
  assign rd_0r1d[32] = rdtint_0n[32];
  assign rd_0r1d[33] = rdtint_0n[33];
  assign rd_0r1d[34] = rdtint_0n[34];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgfint_0n[32] = wg_0r0d[32];
  assign wgfint_0n[33] = wg_0r0d[33];
  assign wgfint_0n[34] = wg_0r0d[34];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign wgtint_0n[32] = wg_0r1d[32];
  assign wgtint_0n[33] = wg_0r1d[33];
  assign wgtint_0n[34] = wg_0r1d[34];
  assign rg_2a = rgaint_2n;
  assign rgrint_2n = rg_2r;
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR3 I292 (internal_0n[0], rgrint_0n, rgrint_1n, rgrint_2n);
  NOR3 I293 (internal_0n[1], rgaint_0n, rgaint_1n, rgaint_2n);
  AND2 I294 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I295 (rdtint_2n[0], rgrint_2n, dt_0n[0]);
  AND2 I296 (rdtint_2n[1], rgrint_2n, dt_0n[1]);
  AND2 I297 (rdtint_2n[2], rgrint_2n, dt_0n[2]);
  AND2 I298 (rdtint_2n[3], rgrint_2n, dt_0n[3]);
  AND2 I299 (rdtint_2n[4], rgrint_2n, dt_0n[4]);
  AND2 I300 (rdtint_2n[5], rgrint_2n, dt_0n[5]);
  AND2 I301 (rdtint_2n[6], rgrint_2n, dt_0n[6]);
  AND2 I302 (rdtint_2n[7], rgrint_2n, dt_0n[7]);
  AND2 I303 (rdtint_2n[8], rgrint_2n, dt_0n[8]);
  AND2 I304 (rdtint_2n[9], rgrint_2n, dt_0n[9]);
  AND2 I305 (rdtint_2n[10], rgrint_2n, dt_0n[10]);
  AND2 I306 (rdtint_2n[11], rgrint_2n, dt_0n[11]);
  AND2 I307 (rdtint_2n[12], rgrint_2n, dt_0n[12]);
  AND2 I308 (rdtint_2n[13], rgrint_2n, dt_0n[13]);
  AND2 I309 (rdtint_2n[14], rgrint_2n, dt_0n[14]);
  AND2 I310 (rdtint_2n[15], rgrint_2n, dt_0n[15]);
  AND2 I311 (rdtint_2n[16], rgrint_2n, dt_0n[16]);
  AND2 I312 (rdtint_2n[17], rgrint_2n, dt_0n[17]);
  AND2 I313 (rdtint_2n[18], rgrint_2n, dt_0n[18]);
  AND2 I314 (rdtint_2n[19], rgrint_2n, dt_0n[19]);
  AND2 I315 (rdtint_2n[20], rgrint_2n, dt_0n[20]);
  AND2 I316 (rdtint_2n[21], rgrint_2n, dt_0n[21]);
  AND2 I317 (rdtint_2n[22], rgrint_2n, dt_0n[22]);
  AND2 I318 (rdtint_2n[23], rgrint_2n, dt_0n[23]);
  AND2 I319 (rdtint_2n[24], rgrint_2n, dt_0n[24]);
  AND2 I320 (rdtint_2n[25], rgrint_2n, dt_0n[25]);
  AND2 I321 (rdtint_2n[26], rgrint_2n, dt_0n[26]);
  AND2 I322 (rdtint_2n[27], rgrint_2n, dt_0n[27]);
  AND2 I323 (rdtint_2n[28], rgrint_2n, dt_0n[28]);
  AND2 I324 (rdtint_2n[29], rgrint_2n, dt_0n[29]);
  AND2 I325 (rdtint_2n[30], rgrint_2n, dt_0n[30]);
  AND2 I326 (rdtint_2n[31], rgrint_2n, dt_0n[31]);
  AND2 I327 (rdtint_2n[32], rgrint_2n, dt_0n[32]);
  AND2 I328 (rdtint_2n[33], rgrint_2n, dt_0n[33]);
  AND2 I329 (rdtint_2n[34], rgrint_2n, dt_0n[34]);
  AND2 I330 (rdtint_1n[0], rgrint_1n, dt_0n[0]);
  AND2 I331 (rdtint_1n[1], rgrint_1n, dt_0n[1]);
  AND2 I332 (rdtint_1n[2], rgrint_1n, dt_0n[2]);
  AND2 I333 (rdtint_1n[3], rgrint_1n, dt_0n[3]);
  AND2 I334 (rdtint_1n[4], rgrint_1n, dt_0n[4]);
  AND2 I335 (rdtint_1n[5], rgrint_1n, dt_0n[5]);
  AND2 I336 (rdtint_1n[6], rgrint_1n, dt_0n[6]);
  AND2 I337 (rdtint_1n[7], rgrint_1n, dt_0n[7]);
  AND2 I338 (rdtint_1n[8], rgrint_1n, dt_0n[8]);
  AND2 I339 (rdtint_1n[9], rgrint_1n, dt_0n[9]);
  AND2 I340 (rdtint_1n[10], rgrint_1n, dt_0n[10]);
  AND2 I341 (rdtint_1n[11], rgrint_1n, dt_0n[11]);
  AND2 I342 (rdtint_1n[12], rgrint_1n, dt_0n[12]);
  AND2 I343 (rdtint_1n[13], rgrint_1n, dt_0n[13]);
  AND2 I344 (rdtint_1n[14], rgrint_1n, dt_0n[14]);
  AND2 I345 (rdtint_1n[15], rgrint_1n, dt_0n[15]);
  AND2 I346 (rdtint_1n[16], rgrint_1n, dt_0n[16]);
  AND2 I347 (rdtint_1n[17], rgrint_1n, dt_0n[17]);
  AND2 I348 (rdtint_1n[18], rgrint_1n, dt_0n[18]);
  AND2 I349 (rdtint_1n[19], rgrint_1n, dt_0n[19]);
  AND2 I350 (rdtint_1n[20], rgrint_1n, dt_0n[20]);
  AND2 I351 (rdtint_1n[21], rgrint_1n, dt_0n[21]);
  AND2 I352 (rdtint_1n[22], rgrint_1n, dt_0n[22]);
  AND2 I353 (rdtint_1n[23], rgrint_1n, dt_0n[23]);
  AND2 I354 (rdtint_1n[24], rgrint_1n, dt_0n[24]);
  AND2 I355 (rdtint_1n[25], rgrint_1n, dt_0n[25]);
  AND2 I356 (rdtint_1n[26], rgrint_1n, dt_0n[26]);
  AND2 I357 (rdtint_1n[27], rgrint_1n, dt_0n[27]);
  AND2 I358 (rdtint_1n[28], rgrint_1n, dt_0n[28]);
  AND2 I359 (rdtint_1n[29], rgrint_1n, dt_0n[29]);
  AND2 I360 (rdtint_1n[30], rgrint_1n, dt_0n[30]);
  AND2 I361 (rdtint_1n[31], rgrint_1n, dt_0n[31]);
  AND2 I362 (rdtint_1n[32], rgrint_1n, dt_0n[32]);
  AND2 I363 (rdtint_1n[33], rgrint_1n, dt_0n[33]);
  AND2 I364 (rdtint_1n[34], rgrint_1n, dt_0n[34]);
  AND2 I365 (rdtint_0n[0], rgrint_0n, dt_0n[0]);
  AND2 I366 (rdtint_0n[1], rgrint_0n, dt_0n[1]);
  AND2 I367 (rdtint_0n[2], rgrint_0n, dt_0n[2]);
  AND2 I368 (rdtint_0n[3], rgrint_0n, dt_0n[3]);
  AND2 I369 (rdtint_0n[4], rgrint_0n, dt_0n[4]);
  AND2 I370 (rdtint_0n[5], rgrint_0n, dt_0n[5]);
  AND2 I371 (rdtint_0n[6], rgrint_0n, dt_0n[6]);
  AND2 I372 (rdtint_0n[7], rgrint_0n, dt_0n[7]);
  AND2 I373 (rdtint_0n[8], rgrint_0n, dt_0n[8]);
  AND2 I374 (rdtint_0n[9], rgrint_0n, dt_0n[9]);
  AND2 I375 (rdtint_0n[10], rgrint_0n, dt_0n[10]);
  AND2 I376 (rdtint_0n[11], rgrint_0n, dt_0n[11]);
  AND2 I377 (rdtint_0n[12], rgrint_0n, dt_0n[12]);
  AND2 I378 (rdtint_0n[13], rgrint_0n, dt_0n[13]);
  AND2 I379 (rdtint_0n[14], rgrint_0n, dt_0n[14]);
  AND2 I380 (rdtint_0n[15], rgrint_0n, dt_0n[15]);
  AND2 I381 (rdtint_0n[16], rgrint_0n, dt_0n[16]);
  AND2 I382 (rdtint_0n[17], rgrint_0n, dt_0n[17]);
  AND2 I383 (rdtint_0n[18], rgrint_0n, dt_0n[18]);
  AND2 I384 (rdtint_0n[19], rgrint_0n, dt_0n[19]);
  AND2 I385 (rdtint_0n[20], rgrint_0n, dt_0n[20]);
  AND2 I386 (rdtint_0n[21], rgrint_0n, dt_0n[21]);
  AND2 I387 (rdtint_0n[22], rgrint_0n, dt_0n[22]);
  AND2 I388 (rdtint_0n[23], rgrint_0n, dt_0n[23]);
  AND2 I389 (rdtint_0n[24], rgrint_0n, dt_0n[24]);
  AND2 I390 (rdtint_0n[25], rgrint_0n, dt_0n[25]);
  AND2 I391 (rdtint_0n[26], rgrint_0n, dt_0n[26]);
  AND2 I392 (rdtint_0n[27], rgrint_0n, dt_0n[27]);
  AND2 I393 (rdtint_0n[28], rgrint_0n, dt_0n[28]);
  AND2 I394 (rdtint_0n[29], rgrint_0n, dt_0n[29]);
  AND2 I395 (rdtint_0n[30], rgrint_0n, dt_0n[30]);
  AND2 I396 (rdtint_0n[31], rgrint_0n, dt_0n[31]);
  AND2 I397 (rdtint_0n[32], rgrint_0n, dt_0n[32]);
  AND2 I398 (rdtint_0n[33], rgrint_0n, dt_0n[33]);
  AND2 I399 (rdtint_0n[34], rgrint_0n, dt_0n[34]);
  AND2 I400 (rdfint_2n[0], rgrint_2n, df_0n[0]);
  AND2 I401 (rdfint_2n[1], rgrint_2n, df_0n[1]);
  AND2 I402 (rdfint_2n[2], rgrint_2n, df_0n[2]);
  AND2 I403 (rdfint_2n[3], rgrint_2n, df_0n[3]);
  AND2 I404 (rdfint_2n[4], rgrint_2n, df_0n[4]);
  AND2 I405 (rdfint_2n[5], rgrint_2n, df_0n[5]);
  AND2 I406 (rdfint_2n[6], rgrint_2n, df_0n[6]);
  AND2 I407 (rdfint_2n[7], rgrint_2n, df_0n[7]);
  AND2 I408 (rdfint_2n[8], rgrint_2n, df_0n[8]);
  AND2 I409 (rdfint_2n[9], rgrint_2n, df_0n[9]);
  AND2 I410 (rdfint_2n[10], rgrint_2n, df_0n[10]);
  AND2 I411 (rdfint_2n[11], rgrint_2n, df_0n[11]);
  AND2 I412 (rdfint_2n[12], rgrint_2n, df_0n[12]);
  AND2 I413 (rdfint_2n[13], rgrint_2n, df_0n[13]);
  AND2 I414 (rdfint_2n[14], rgrint_2n, df_0n[14]);
  AND2 I415 (rdfint_2n[15], rgrint_2n, df_0n[15]);
  AND2 I416 (rdfint_2n[16], rgrint_2n, df_0n[16]);
  AND2 I417 (rdfint_2n[17], rgrint_2n, df_0n[17]);
  AND2 I418 (rdfint_2n[18], rgrint_2n, df_0n[18]);
  AND2 I419 (rdfint_2n[19], rgrint_2n, df_0n[19]);
  AND2 I420 (rdfint_2n[20], rgrint_2n, df_0n[20]);
  AND2 I421 (rdfint_2n[21], rgrint_2n, df_0n[21]);
  AND2 I422 (rdfint_2n[22], rgrint_2n, df_0n[22]);
  AND2 I423 (rdfint_2n[23], rgrint_2n, df_0n[23]);
  AND2 I424 (rdfint_2n[24], rgrint_2n, df_0n[24]);
  AND2 I425 (rdfint_2n[25], rgrint_2n, df_0n[25]);
  AND2 I426 (rdfint_2n[26], rgrint_2n, df_0n[26]);
  AND2 I427 (rdfint_2n[27], rgrint_2n, df_0n[27]);
  AND2 I428 (rdfint_2n[28], rgrint_2n, df_0n[28]);
  AND2 I429 (rdfint_2n[29], rgrint_2n, df_0n[29]);
  AND2 I430 (rdfint_2n[30], rgrint_2n, df_0n[30]);
  AND2 I431 (rdfint_2n[31], rgrint_2n, df_0n[31]);
  AND2 I432 (rdfint_2n[32], rgrint_2n, df_0n[32]);
  AND2 I433 (rdfint_2n[33], rgrint_2n, df_0n[33]);
  AND2 I434 (rdfint_2n[34], rgrint_2n, df_0n[34]);
  AND2 I435 (rdfint_1n[0], rgrint_1n, df_0n[0]);
  AND2 I436 (rdfint_1n[1], rgrint_1n, df_0n[1]);
  AND2 I437 (rdfint_1n[2], rgrint_1n, df_0n[2]);
  AND2 I438 (rdfint_1n[3], rgrint_1n, df_0n[3]);
  AND2 I439 (rdfint_1n[4], rgrint_1n, df_0n[4]);
  AND2 I440 (rdfint_1n[5], rgrint_1n, df_0n[5]);
  AND2 I441 (rdfint_1n[6], rgrint_1n, df_0n[6]);
  AND2 I442 (rdfint_1n[7], rgrint_1n, df_0n[7]);
  AND2 I443 (rdfint_1n[8], rgrint_1n, df_0n[8]);
  AND2 I444 (rdfint_1n[9], rgrint_1n, df_0n[9]);
  AND2 I445 (rdfint_1n[10], rgrint_1n, df_0n[10]);
  AND2 I446 (rdfint_1n[11], rgrint_1n, df_0n[11]);
  AND2 I447 (rdfint_1n[12], rgrint_1n, df_0n[12]);
  AND2 I448 (rdfint_1n[13], rgrint_1n, df_0n[13]);
  AND2 I449 (rdfint_1n[14], rgrint_1n, df_0n[14]);
  AND2 I450 (rdfint_1n[15], rgrint_1n, df_0n[15]);
  AND2 I451 (rdfint_1n[16], rgrint_1n, df_0n[16]);
  AND2 I452 (rdfint_1n[17], rgrint_1n, df_0n[17]);
  AND2 I453 (rdfint_1n[18], rgrint_1n, df_0n[18]);
  AND2 I454 (rdfint_1n[19], rgrint_1n, df_0n[19]);
  AND2 I455 (rdfint_1n[20], rgrint_1n, df_0n[20]);
  AND2 I456 (rdfint_1n[21], rgrint_1n, df_0n[21]);
  AND2 I457 (rdfint_1n[22], rgrint_1n, df_0n[22]);
  AND2 I458 (rdfint_1n[23], rgrint_1n, df_0n[23]);
  AND2 I459 (rdfint_1n[24], rgrint_1n, df_0n[24]);
  AND2 I460 (rdfint_1n[25], rgrint_1n, df_0n[25]);
  AND2 I461 (rdfint_1n[26], rgrint_1n, df_0n[26]);
  AND2 I462 (rdfint_1n[27], rgrint_1n, df_0n[27]);
  AND2 I463 (rdfint_1n[28], rgrint_1n, df_0n[28]);
  AND2 I464 (rdfint_1n[29], rgrint_1n, df_0n[29]);
  AND2 I465 (rdfint_1n[30], rgrint_1n, df_0n[30]);
  AND2 I466 (rdfint_1n[31], rgrint_1n, df_0n[31]);
  AND2 I467 (rdfint_1n[32], rgrint_1n, df_0n[32]);
  AND2 I468 (rdfint_1n[33], rgrint_1n, df_0n[33]);
  AND2 I469 (rdfint_1n[34], rgrint_1n, df_0n[34]);
  AND2 I470 (rdfint_0n[0], rgrint_0n, df_0n[0]);
  AND2 I471 (rdfint_0n[1], rgrint_0n, df_0n[1]);
  AND2 I472 (rdfint_0n[2], rgrint_0n, df_0n[2]);
  AND2 I473 (rdfint_0n[3], rgrint_0n, df_0n[3]);
  AND2 I474 (rdfint_0n[4], rgrint_0n, df_0n[4]);
  AND2 I475 (rdfint_0n[5], rgrint_0n, df_0n[5]);
  AND2 I476 (rdfint_0n[6], rgrint_0n, df_0n[6]);
  AND2 I477 (rdfint_0n[7], rgrint_0n, df_0n[7]);
  AND2 I478 (rdfint_0n[8], rgrint_0n, df_0n[8]);
  AND2 I479 (rdfint_0n[9], rgrint_0n, df_0n[9]);
  AND2 I480 (rdfint_0n[10], rgrint_0n, df_0n[10]);
  AND2 I481 (rdfint_0n[11], rgrint_0n, df_0n[11]);
  AND2 I482 (rdfint_0n[12], rgrint_0n, df_0n[12]);
  AND2 I483 (rdfint_0n[13], rgrint_0n, df_0n[13]);
  AND2 I484 (rdfint_0n[14], rgrint_0n, df_0n[14]);
  AND2 I485 (rdfint_0n[15], rgrint_0n, df_0n[15]);
  AND2 I486 (rdfint_0n[16], rgrint_0n, df_0n[16]);
  AND2 I487 (rdfint_0n[17], rgrint_0n, df_0n[17]);
  AND2 I488 (rdfint_0n[18], rgrint_0n, df_0n[18]);
  AND2 I489 (rdfint_0n[19], rgrint_0n, df_0n[19]);
  AND2 I490 (rdfint_0n[20], rgrint_0n, df_0n[20]);
  AND2 I491 (rdfint_0n[21], rgrint_0n, df_0n[21]);
  AND2 I492 (rdfint_0n[22], rgrint_0n, df_0n[22]);
  AND2 I493 (rdfint_0n[23], rgrint_0n, df_0n[23]);
  AND2 I494 (rdfint_0n[24], rgrint_0n, df_0n[24]);
  AND2 I495 (rdfint_0n[25], rgrint_0n, df_0n[25]);
  AND2 I496 (rdfint_0n[26], rgrint_0n, df_0n[26]);
  AND2 I497 (rdfint_0n[27], rgrint_0n, df_0n[27]);
  AND2 I498 (rdfint_0n[28], rgrint_0n, df_0n[28]);
  AND2 I499 (rdfint_0n[29], rgrint_0n, df_0n[29]);
  AND2 I500 (rdfint_0n[30], rgrint_0n, df_0n[30]);
  AND2 I501 (rdfint_0n[31], rgrint_0n, df_0n[31]);
  AND2 I502 (rdfint_0n[32], rgrint_0n, df_0n[32]);
  AND2 I503 (rdfint_0n[33], rgrint_0n, df_0n[33]);
  AND2 I504 (rdfint_0n[34], rgrint_0n, df_0n[34]);
  C3 I505 (internal_0n[2], wc_0n, wacks_0n[34], wacks_0n[33]);
  C3 I506 (internal_0n[3], wacks_0n[32], wacks_0n[31], wacks_0n[30]);
  C3 I507 (internal_0n[4], wacks_0n[29], wacks_0n[28], wacks_0n[27]);
  C3 I508 (internal_0n[5], wacks_0n[26], wacks_0n[25], wacks_0n[24]);
  C3 I509 (internal_0n[6], wacks_0n[23], wacks_0n[22], wacks_0n[21]);
  C3 I510 (internal_0n[7], wacks_0n[20], wacks_0n[19], wacks_0n[18]);
  C3 I511 (internal_0n[8], wacks_0n[17], wacks_0n[16], wacks_0n[15]);
  C3 I512 (internal_0n[9], wacks_0n[14], wacks_0n[13], wacks_0n[12]);
  C3 I513 (internal_0n[10], wacks_0n[11], wacks_0n[10], wacks_0n[9]);
  C3 I514 (internal_0n[11], wacks_0n[8], wacks_0n[7], wacks_0n[6]);
  C3 I515 (internal_0n[12], wacks_0n[5], wacks_0n[4], wacks_0n[3]);
  C3 I516 (internal_0n[13], wacks_0n[2], wacks_0n[1], wacks_0n[0]);
  C3 I517 (internal_0n[14], internal_0n[2], internal_0n[3], internal_0n[4]);
  C3 I518 (internal_0n[15], internal_0n[5], internal_0n[6], internal_0n[7]);
  C3 I519 (internal_0n[16], internal_0n[8], internal_0n[9], internal_0n[10]);
  C3 I520 (internal_0n[17], internal_0n[11], internal_0n[12], internal_0n[13]);
  C2 I521 (internal_0n[18], internal_0n[14], internal_0n[15]);
  C2 I522 (internal_0n[19], internal_0n[16], internal_0n[17]);
  C2 I523 (wdrint_0n, internal_0n[18], internal_0n[19]);
  assign wen_0n[34] = wc_0n;
  assign wen_0n[33] = wc_0n;
  assign wen_0n[32] = wc_0n;
  assign wen_0n[31] = wc_0n;
  assign wen_0n[30] = wc_0n;
  assign wen_0n[29] = wc_0n;
  assign wen_0n[28] = wc_0n;
  assign wen_0n[27] = wc_0n;
  assign wen_0n[26] = wc_0n;
  assign wen_0n[25] = wc_0n;
  assign wen_0n[24] = wc_0n;
  assign wen_0n[23] = wc_0n;
  assign wen_0n[22] = wc_0n;
  assign wen_0n[21] = wc_0n;
  assign wen_0n[20] = wc_0n;
  assign wen_0n[19] = wc_0n;
  assign wen_0n[18] = wc_0n;
  assign wen_0n[17] = wc_0n;
  assign wen_0n[16] = wc_0n;
  assign wen_0n[15] = wc_0n;
  assign wen_0n[14] = wc_0n;
  assign wen_0n[13] = wc_0n;
  assign wen_0n[12] = wc_0n;
  assign wen_0n[11] = wc_0n;
  assign wen_0n[10] = wc_0n;
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[34] = git_0n[34];
  assign wt_0n[33] = git_0n[33];
  assign wt_0n[32] = git_0n[32];
  assign wt_0n[31] = git_0n[31];
  assign wt_0n[30] = git_0n[30];
  assign wt_0n[29] = git_0n[29];
  assign wt_0n[28] = git_0n[28];
  assign wt_0n[27] = git_0n[27];
  assign wt_0n[26] = git_0n[26];
  assign wt_0n[25] = git_0n[25];
  assign wt_0n[24] = git_0n[24];
  assign wt_0n[23] = git_0n[23];
  assign wt_0n[22] = git_0n[22];
  assign wt_0n[21] = git_0n[21];
  assign wt_0n[20] = git_0n[20];
  assign wt_0n[19] = git_0n[19];
  assign wt_0n[18] = git_0n[18];
  assign wt_0n[17] = git_0n[17];
  assign wt_0n[16] = git_0n[16];
  assign wt_0n[15] = git_0n[15];
  assign wt_0n[14] = git_0n[14];
  assign wt_0n[13] = git_0n[13];
  assign wt_0n[12] = git_0n[12];
  assign wt_0n[11] = git_0n[11];
  assign wt_0n[10] = git_0n[10];
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[34] = gif_0n[34];
  assign wf_0n[33] = gif_0n[33];
  assign wf_0n[32] = gif_0n[32];
  assign wf_0n[31] = gif_0n[31];
  assign wf_0n[30] = gif_0n[30];
  assign wf_0n[29] = gif_0n[29];
  assign wf_0n[28] = gif_0n[28];
  assign wf_0n[27] = gif_0n[27];
  assign wf_0n[26] = gif_0n[26];
  assign wf_0n[25] = gif_0n[25];
  assign wf_0n[24] = gif_0n[24];
  assign wf_0n[23] = gif_0n[23];
  assign wf_0n[22] = gif_0n[22];
  assign wf_0n[21] = gif_0n[21];
  assign wf_0n[20] = gif_0n[20];
  assign wf_0n[19] = gif_0n[19];
  assign wf_0n[18] = gif_0n[18];
  assign wf_0n[17] = gif_0n[17];
  assign wf_0n[16] = gif_0n[16];
  assign wf_0n[15] = gif_0n[15];
  assign wf_0n[14] = gif_0n[14];
  assign wf_0n[13] = gif_0n[13];
  assign wf_0n[12] = gif_0n[12];
  assign wf_0n[11] = gif_0n[11];
  assign wf_0n[10] = gif_0n[10];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I629 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I631 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I632 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I633 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I634 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I635 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I636 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I637 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I638 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I639 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I640 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I641 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I642 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I643 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I644 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I645 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I646 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I647 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I648 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I649 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I650 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I651 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I652 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I653 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I654 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I655 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I656 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I657 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I658 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I659 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I660 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I661 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I662 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I663 (git_0n[32], wgtint_0n[32], ig_0n);
  AND2 I664 (git_0n[33], wgtint_0n[33], ig_0n);
  AND2 I665 (git_0n[34], wgtint_0n[34], ig_0n);
  AND2 I666 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I667 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I668 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I669 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I670 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I671 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I672 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I673 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I674 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I675 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I676 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I677 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I678 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I679 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I680 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I681 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I682 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I683 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I684 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I685 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I686 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I687 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I688 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I689 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I690 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I691 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I692 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I693 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I694 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I695 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I696 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I697 (gif_0n[31], wgfint_0n[31], ig_0n);
  AND2 I698 (gif_0n[32], wgfint_0n[32], ig_0n);
  AND2 I699 (gif_0n[33], wgfint_0n[33], ig_0n);
  AND2 I700 (gif_0n[34], wgfint_0n[34], ig_0n);
  C3 I701 (internal_0n[20], complete1501_0n[0], complete1501_0n[1], complete1501_0n[2]);
  C3 I702 (internal_0n[21], complete1501_0n[3], complete1501_0n[4], complete1501_0n[5]);
  C3 I703 (internal_0n[22], complete1501_0n[6], complete1501_0n[7], complete1501_0n[8]);
  C3 I704 (internal_0n[23], complete1501_0n[9], complete1501_0n[10], complete1501_0n[11]);
  C3 I705 (internal_0n[24], complete1501_0n[12], complete1501_0n[13], complete1501_0n[14]);
  C3 I706 (internal_0n[25], complete1501_0n[15], complete1501_0n[16], complete1501_0n[17]);
  C3 I707 (internal_0n[26], complete1501_0n[18], complete1501_0n[19], complete1501_0n[20]);
  C3 I708 (internal_0n[27], complete1501_0n[21], complete1501_0n[22], complete1501_0n[23]);
  C3 I709 (internal_0n[28], complete1501_0n[24], complete1501_0n[25], complete1501_0n[26]);
  C3 I710 (internal_0n[29], complete1501_0n[27], complete1501_0n[28], complete1501_0n[29]);
  C3 I711 (internal_0n[30], complete1501_0n[30], complete1501_0n[31], complete1501_0n[32]);
  C2 I712 (internal_0n[31], complete1501_0n[33], complete1501_0n[34]);
  C3 I713 (internal_0n[32], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I714 (internal_0n[33], internal_0n[23], internal_0n[24], internal_0n[25]);
  C3 I715 (internal_0n[34], internal_0n[26], internal_0n[27], internal_0n[28]);
  C3 I716 (internal_0n[35], internal_0n[29], internal_0n[30], internal_0n[31]);
  C2 I717 (internal_0n[36], internal_0n[32], internal_0n[33]);
  C2 I718 (internal_0n[37], internal_0n[34], internal_0n[35]);
  C2 I719 (wc_0n, internal_0n[36], internal_0n[37]);
  OR2 I720 (complete1501_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I721 (complete1501_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I722 (complete1501_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I723 (complete1501_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I724 (complete1501_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I725 (complete1501_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I726 (complete1501_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I727 (complete1501_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I728 (complete1501_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I729 (complete1501_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I730 (complete1501_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I731 (complete1501_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I732 (complete1501_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I733 (complete1501_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I734 (complete1501_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I735 (complete1501_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I736 (complete1501_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I737 (complete1501_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I738 (complete1501_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I739 (complete1501_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I740 (complete1501_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I741 (complete1501_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I742 (complete1501_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I743 (complete1501_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I744 (complete1501_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I745 (complete1501_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I746 (complete1501_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I747 (complete1501_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I748 (complete1501_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I749 (complete1501_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I750 (complete1501_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I751 (complete1501_0n[31], wgfint_0n[31], wgtint_0n[31]);
  OR2 I752 (complete1501_0n[32], wgfint_0n[32], wgtint_0n[32]);
  OR2 I753 (complete1501_0n[33], wgfint_0n[33], wgtint_0n[33]);
  OR2 I754 (complete1501_0n[34], wgfint_0n[34], wgtint_0n[34]);
  AO22 I755 (wacks_0n[34], gf1499_0n[34], df_0n[34], gt1500_0n[34], dt_0n[34]);
  NOR2 I756 (dt_0n[34], df_0n[34], gf1499_0n[34]);
  NOR3 I757 (df_0n[34], dt_0n[34], gt1500_0n[34], init_0n);
  AND2 I758 (gt1500_0n[34], wt_0n[34], wen_0n[34]);
  AND2 I759 (gf1499_0n[34], wf_0n[34], wen_0n[34]);
  AO22 I760 (wacks_0n[33], gf1499_0n[33], df_0n[33], gt1500_0n[33], dt_0n[33]);
  NOR2 I761 (dt_0n[33], df_0n[33], gf1499_0n[33]);
  NOR3 I762 (df_0n[33], dt_0n[33], gt1500_0n[33], init_0n);
  AND2 I763 (gt1500_0n[33], wt_0n[33], wen_0n[33]);
  AND2 I764 (gf1499_0n[33], wf_0n[33], wen_0n[33]);
  AO22 I765 (wacks_0n[32], gf1499_0n[32], df_0n[32], gt1500_0n[32], dt_0n[32]);
  NOR2 I766 (dt_0n[32], df_0n[32], gf1499_0n[32]);
  NOR3 I767 (df_0n[32], dt_0n[32], gt1500_0n[32], init_0n);
  AND2 I768 (gt1500_0n[32], wt_0n[32], wen_0n[32]);
  AND2 I769 (gf1499_0n[32], wf_0n[32], wen_0n[32]);
  AO22 I770 (wacks_0n[31], gf1499_0n[31], df_0n[31], gt1500_0n[31], dt_0n[31]);
  NOR2 I771 (dt_0n[31], df_0n[31], gf1499_0n[31]);
  NOR3 I772 (df_0n[31], dt_0n[31], gt1500_0n[31], init_0n);
  AND2 I773 (gt1500_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I774 (gf1499_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I775 (wacks_0n[30], gf1499_0n[30], df_0n[30], gt1500_0n[30], dt_0n[30]);
  NOR2 I776 (dt_0n[30], df_0n[30], gf1499_0n[30]);
  NOR3 I777 (df_0n[30], dt_0n[30], gt1500_0n[30], init_0n);
  AND2 I778 (gt1500_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I779 (gf1499_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I780 (wacks_0n[29], gf1499_0n[29], df_0n[29], gt1500_0n[29], dt_0n[29]);
  NOR2 I781 (dt_0n[29], df_0n[29], gf1499_0n[29]);
  NOR3 I782 (df_0n[29], dt_0n[29], gt1500_0n[29], init_0n);
  AND2 I783 (gt1500_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I784 (gf1499_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I785 (wacks_0n[28], gf1499_0n[28], df_0n[28], gt1500_0n[28], dt_0n[28]);
  NOR2 I786 (dt_0n[28], df_0n[28], gf1499_0n[28]);
  NOR3 I787 (df_0n[28], dt_0n[28], gt1500_0n[28], init_0n);
  AND2 I788 (gt1500_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I789 (gf1499_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I790 (wacks_0n[27], gf1499_0n[27], df_0n[27], gt1500_0n[27], dt_0n[27]);
  NOR2 I791 (dt_0n[27], df_0n[27], gf1499_0n[27]);
  NOR3 I792 (df_0n[27], dt_0n[27], gt1500_0n[27], init_0n);
  AND2 I793 (gt1500_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I794 (gf1499_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I795 (wacks_0n[26], gf1499_0n[26], df_0n[26], gt1500_0n[26], dt_0n[26]);
  NOR2 I796 (dt_0n[26], df_0n[26], gf1499_0n[26]);
  NOR3 I797 (df_0n[26], dt_0n[26], gt1500_0n[26], init_0n);
  AND2 I798 (gt1500_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I799 (gf1499_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I800 (wacks_0n[25], gf1499_0n[25], df_0n[25], gt1500_0n[25], dt_0n[25]);
  NOR2 I801 (dt_0n[25], df_0n[25], gf1499_0n[25]);
  NOR3 I802 (df_0n[25], dt_0n[25], gt1500_0n[25], init_0n);
  AND2 I803 (gt1500_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I804 (gf1499_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I805 (wacks_0n[24], gf1499_0n[24], df_0n[24], gt1500_0n[24], dt_0n[24]);
  NOR2 I806 (dt_0n[24], df_0n[24], gf1499_0n[24]);
  NOR3 I807 (df_0n[24], dt_0n[24], gt1500_0n[24], init_0n);
  AND2 I808 (gt1500_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I809 (gf1499_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I810 (wacks_0n[23], gf1499_0n[23], df_0n[23], gt1500_0n[23], dt_0n[23]);
  NOR2 I811 (dt_0n[23], df_0n[23], gf1499_0n[23]);
  NOR3 I812 (df_0n[23], dt_0n[23], gt1500_0n[23], init_0n);
  AND2 I813 (gt1500_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I814 (gf1499_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I815 (wacks_0n[22], gf1499_0n[22], df_0n[22], gt1500_0n[22], dt_0n[22]);
  NOR2 I816 (dt_0n[22], df_0n[22], gf1499_0n[22]);
  NOR3 I817 (df_0n[22], dt_0n[22], gt1500_0n[22], init_0n);
  AND2 I818 (gt1500_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I819 (gf1499_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I820 (wacks_0n[21], gf1499_0n[21], df_0n[21], gt1500_0n[21], dt_0n[21]);
  NOR2 I821 (dt_0n[21], df_0n[21], gf1499_0n[21]);
  NOR3 I822 (df_0n[21], dt_0n[21], gt1500_0n[21], init_0n);
  AND2 I823 (gt1500_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I824 (gf1499_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I825 (wacks_0n[20], gf1499_0n[20], df_0n[20], gt1500_0n[20], dt_0n[20]);
  NOR2 I826 (dt_0n[20], df_0n[20], gf1499_0n[20]);
  NOR3 I827 (df_0n[20], dt_0n[20], gt1500_0n[20], init_0n);
  AND2 I828 (gt1500_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I829 (gf1499_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I830 (wacks_0n[19], gf1499_0n[19], df_0n[19], gt1500_0n[19], dt_0n[19]);
  NOR2 I831 (dt_0n[19], df_0n[19], gf1499_0n[19]);
  NOR3 I832 (df_0n[19], dt_0n[19], gt1500_0n[19], init_0n);
  AND2 I833 (gt1500_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I834 (gf1499_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I835 (wacks_0n[18], gf1499_0n[18], df_0n[18], gt1500_0n[18], dt_0n[18]);
  NOR2 I836 (dt_0n[18], df_0n[18], gf1499_0n[18]);
  NOR3 I837 (df_0n[18], dt_0n[18], gt1500_0n[18], init_0n);
  AND2 I838 (gt1500_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I839 (gf1499_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I840 (wacks_0n[17], gf1499_0n[17], df_0n[17], gt1500_0n[17], dt_0n[17]);
  NOR2 I841 (dt_0n[17], df_0n[17], gf1499_0n[17]);
  NOR3 I842 (df_0n[17], dt_0n[17], gt1500_0n[17], init_0n);
  AND2 I843 (gt1500_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I844 (gf1499_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I845 (wacks_0n[16], gf1499_0n[16], df_0n[16], gt1500_0n[16], dt_0n[16]);
  NOR2 I846 (dt_0n[16], df_0n[16], gf1499_0n[16]);
  NOR3 I847 (df_0n[16], dt_0n[16], gt1500_0n[16], init_0n);
  AND2 I848 (gt1500_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I849 (gf1499_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I850 (wacks_0n[15], gf1499_0n[15], df_0n[15], gt1500_0n[15], dt_0n[15]);
  NOR2 I851 (dt_0n[15], df_0n[15], gf1499_0n[15]);
  NOR3 I852 (df_0n[15], dt_0n[15], gt1500_0n[15], init_0n);
  AND2 I853 (gt1500_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I854 (gf1499_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I855 (wacks_0n[14], gf1499_0n[14], df_0n[14], gt1500_0n[14], dt_0n[14]);
  NOR2 I856 (dt_0n[14], df_0n[14], gf1499_0n[14]);
  NOR3 I857 (df_0n[14], dt_0n[14], gt1500_0n[14], init_0n);
  AND2 I858 (gt1500_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I859 (gf1499_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I860 (wacks_0n[13], gf1499_0n[13], df_0n[13], gt1500_0n[13], dt_0n[13]);
  NOR2 I861 (dt_0n[13], df_0n[13], gf1499_0n[13]);
  NOR3 I862 (df_0n[13], dt_0n[13], gt1500_0n[13], init_0n);
  AND2 I863 (gt1500_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I864 (gf1499_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I865 (wacks_0n[12], gf1499_0n[12], df_0n[12], gt1500_0n[12], dt_0n[12]);
  NOR2 I866 (dt_0n[12], df_0n[12], gf1499_0n[12]);
  NOR3 I867 (df_0n[12], dt_0n[12], gt1500_0n[12], init_0n);
  AND2 I868 (gt1500_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I869 (gf1499_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I870 (wacks_0n[11], gf1499_0n[11], df_0n[11], gt1500_0n[11], dt_0n[11]);
  NOR2 I871 (dt_0n[11], df_0n[11], gf1499_0n[11]);
  NOR3 I872 (df_0n[11], dt_0n[11], gt1500_0n[11], init_0n);
  AND2 I873 (gt1500_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I874 (gf1499_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I875 (wacks_0n[10], gf1499_0n[10], df_0n[10], gt1500_0n[10], dt_0n[10]);
  NOR2 I876 (dt_0n[10], df_0n[10], gf1499_0n[10]);
  NOR3 I877 (df_0n[10], dt_0n[10], gt1500_0n[10], init_0n);
  AND2 I878 (gt1500_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I879 (gf1499_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I880 (wacks_0n[9], gf1499_0n[9], df_0n[9], gt1500_0n[9], dt_0n[9]);
  NOR2 I881 (dt_0n[9], df_0n[9], gf1499_0n[9]);
  NOR3 I882 (df_0n[9], dt_0n[9], gt1500_0n[9], init_0n);
  AND2 I883 (gt1500_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I884 (gf1499_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I885 (wacks_0n[8], gf1499_0n[8], df_0n[8], gt1500_0n[8], dt_0n[8]);
  NOR2 I886 (dt_0n[8], df_0n[8], gf1499_0n[8]);
  NOR3 I887 (df_0n[8], dt_0n[8], gt1500_0n[8], init_0n);
  AND2 I888 (gt1500_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I889 (gf1499_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I890 (wacks_0n[7], gf1499_0n[7], df_0n[7], gt1500_0n[7], dt_0n[7]);
  NOR2 I891 (dt_0n[7], df_0n[7], gf1499_0n[7]);
  NOR3 I892 (df_0n[7], dt_0n[7], gt1500_0n[7], init_0n);
  AND2 I893 (gt1500_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I894 (gf1499_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I895 (wacks_0n[6], gf1499_0n[6], df_0n[6], gt1500_0n[6], dt_0n[6]);
  NOR2 I896 (dt_0n[6], df_0n[6], gf1499_0n[6]);
  NOR3 I897 (df_0n[6], dt_0n[6], gt1500_0n[6], init_0n);
  AND2 I898 (gt1500_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I899 (gf1499_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I900 (wacks_0n[5], gf1499_0n[5], df_0n[5], gt1500_0n[5], dt_0n[5]);
  NOR2 I901 (dt_0n[5], df_0n[5], gf1499_0n[5]);
  NOR3 I902 (df_0n[5], dt_0n[5], gt1500_0n[5], init_0n);
  AND2 I903 (gt1500_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I904 (gf1499_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I905 (wacks_0n[4], gf1499_0n[4], df_0n[4], gt1500_0n[4], dt_0n[4]);
  NOR2 I906 (dt_0n[4], df_0n[4], gf1499_0n[4]);
  NOR3 I907 (df_0n[4], dt_0n[4], gt1500_0n[4], init_0n);
  AND2 I908 (gt1500_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I909 (gf1499_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I910 (wacks_0n[3], gf1499_0n[3], df_0n[3], gt1500_0n[3], dt_0n[3]);
  NOR2 I911 (dt_0n[3], df_0n[3], gf1499_0n[3]);
  NOR3 I912 (df_0n[3], dt_0n[3], gt1500_0n[3], init_0n);
  AND2 I913 (gt1500_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I914 (gf1499_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I915 (wacks_0n[2], gf1499_0n[2], df_0n[2], gt1500_0n[2], dt_0n[2]);
  NOR2 I916 (dt_0n[2], df_0n[2], gf1499_0n[2]);
  NOR3 I917 (df_0n[2], dt_0n[2], gt1500_0n[2], init_0n);
  AND2 I918 (gt1500_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I919 (gf1499_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I920 (wacks_0n[1], gf1499_0n[1], df_0n[1], gt1500_0n[1], dt_0n[1]);
  NOR2 I921 (dt_0n[1], df_0n[1], gf1499_0n[1]);
  NOR3 I922 (df_0n[1], dt_0n[1], gt1500_0n[1], init_0n);
  AND2 I923 (gt1500_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I924 (gf1499_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I925 (wacks_0n[0], gf1499_0n[0], df_0n[0], gt1500_0n[0], dt_0n[0]);
  NOR2 I926 (dt_0n[0], df_0n[0], gf1499_0n[0]);
  NOR3 I927 (df_0n[0], dt_0n[0], gt1500_0n[0], init_0n);
  AND2 I928 (gt1500_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I929 (gf1499_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I930 (init_0n, initialise);
endmodule

module BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m92m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rg_2r, rg_2a,
  rg_3r, rg_3a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  rd_2r0d, rd_2r1d, rd_2a,
  rd_3r0d, rd_3r1d, rd_3a,
  initialise
);
  input [34:0] wg_0r0d;
  input [34:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  output [31:0] rd_0r0d;
  output [31:0] rd_0r1d;
  input rd_0a;
  output rd_1r0d;
  output rd_1r1d;
  input rd_1a;
  output rd_2r0d;
  output rd_2r1d;
  input rd_2a;
  output [32:0] rd_3r0d;
  output [32:0] rd_3r1d;
  input rd_3a;
  input initialise;
  wire [38:0] internal_0n;
  wire [34:0] wf_0n;
  wire [34:0] wt_0n;
  wire [34:0] df_0n;
  wire [34:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire rgrint_2n;
  wire rgrint_3n;
  wire wc_0n;
  wire [34:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [34:0] wgfint_0n;
  wire [34:0] wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire rgaint_2n;
  wire rgaint_3n;
  wire [31:0] rdfint_0n;
  wire rdfint_1n;
  wire rdfint_2n;
  wire [32:0] rdfint_3n;
  wire [31:0] rdtint_0n;
  wire rdtint_1n;
  wire rdtint_2n;
  wire [32:0] rdtint_3n;
  wire [34:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [34:0] gif_0n;
  wire [34:0] git_0n;
  wire [34:0] complete1520_0n;
  wire [34:0] gt1519_0n;
  wire [34:0] gf1518_0n;
  assign rgaint_3n = rd_3a;
  assign rd_3r0d[0] = rdfint_3n[0];
  assign rd_3r0d[1] = rdfint_3n[1];
  assign rd_3r0d[2] = rdfint_3n[2];
  assign rd_3r0d[3] = rdfint_3n[3];
  assign rd_3r0d[4] = rdfint_3n[4];
  assign rd_3r0d[5] = rdfint_3n[5];
  assign rd_3r0d[6] = rdfint_3n[6];
  assign rd_3r0d[7] = rdfint_3n[7];
  assign rd_3r0d[8] = rdfint_3n[8];
  assign rd_3r0d[9] = rdfint_3n[9];
  assign rd_3r0d[10] = rdfint_3n[10];
  assign rd_3r0d[11] = rdfint_3n[11];
  assign rd_3r0d[12] = rdfint_3n[12];
  assign rd_3r0d[13] = rdfint_3n[13];
  assign rd_3r0d[14] = rdfint_3n[14];
  assign rd_3r0d[15] = rdfint_3n[15];
  assign rd_3r0d[16] = rdfint_3n[16];
  assign rd_3r0d[17] = rdfint_3n[17];
  assign rd_3r0d[18] = rdfint_3n[18];
  assign rd_3r0d[19] = rdfint_3n[19];
  assign rd_3r0d[20] = rdfint_3n[20];
  assign rd_3r0d[21] = rdfint_3n[21];
  assign rd_3r0d[22] = rdfint_3n[22];
  assign rd_3r0d[23] = rdfint_3n[23];
  assign rd_3r0d[24] = rdfint_3n[24];
  assign rd_3r0d[25] = rdfint_3n[25];
  assign rd_3r0d[26] = rdfint_3n[26];
  assign rd_3r0d[27] = rdfint_3n[27];
  assign rd_3r0d[28] = rdfint_3n[28];
  assign rd_3r0d[29] = rdfint_3n[29];
  assign rd_3r0d[30] = rdfint_3n[30];
  assign rd_3r0d[31] = rdfint_3n[31];
  assign rd_3r0d[32] = rdfint_3n[32];
  assign rd_3r1d[0] = rdtint_3n[0];
  assign rd_3r1d[1] = rdtint_3n[1];
  assign rd_3r1d[2] = rdtint_3n[2];
  assign rd_3r1d[3] = rdtint_3n[3];
  assign rd_3r1d[4] = rdtint_3n[4];
  assign rd_3r1d[5] = rdtint_3n[5];
  assign rd_3r1d[6] = rdtint_3n[6];
  assign rd_3r1d[7] = rdtint_3n[7];
  assign rd_3r1d[8] = rdtint_3n[8];
  assign rd_3r1d[9] = rdtint_3n[9];
  assign rd_3r1d[10] = rdtint_3n[10];
  assign rd_3r1d[11] = rdtint_3n[11];
  assign rd_3r1d[12] = rdtint_3n[12];
  assign rd_3r1d[13] = rdtint_3n[13];
  assign rd_3r1d[14] = rdtint_3n[14];
  assign rd_3r1d[15] = rdtint_3n[15];
  assign rd_3r1d[16] = rdtint_3n[16];
  assign rd_3r1d[17] = rdtint_3n[17];
  assign rd_3r1d[18] = rdtint_3n[18];
  assign rd_3r1d[19] = rdtint_3n[19];
  assign rd_3r1d[20] = rdtint_3n[20];
  assign rd_3r1d[21] = rdtint_3n[21];
  assign rd_3r1d[22] = rdtint_3n[22];
  assign rd_3r1d[23] = rdtint_3n[23];
  assign rd_3r1d[24] = rdtint_3n[24];
  assign rd_3r1d[25] = rdtint_3n[25];
  assign rd_3r1d[26] = rdtint_3n[26];
  assign rd_3r1d[27] = rdtint_3n[27];
  assign rd_3r1d[28] = rdtint_3n[28];
  assign rd_3r1d[29] = rdtint_3n[29];
  assign rd_3r1d[30] = rdtint_3n[30];
  assign rd_3r1d[31] = rdtint_3n[31];
  assign rd_3r1d[32] = rdtint_3n[32];
  assign rgaint_2n = rd_2a;
  assign rd_2r0d = rdfint_2n;
  assign rd_2r1d = rdtint_2n;
  assign rgaint_1n = rd_1a;
  assign rd_1r0d = rdfint_1n;
  assign rd_1r1d = rdtint_1n;
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r0d[10] = rdfint_0n[10];
  assign rd_0r0d[11] = rdfint_0n[11];
  assign rd_0r0d[12] = rdfint_0n[12];
  assign rd_0r0d[13] = rdfint_0n[13];
  assign rd_0r0d[14] = rdfint_0n[14];
  assign rd_0r0d[15] = rdfint_0n[15];
  assign rd_0r0d[16] = rdfint_0n[16];
  assign rd_0r0d[17] = rdfint_0n[17];
  assign rd_0r0d[18] = rdfint_0n[18];
  assign rd_0r0d[19] = rdfint_0n[19];
  assign rd_0r0d[20] = rdfint_0n[20];
  assign rd_0r0d[21] = rdfint_0n[21];
  assign rd_0r0d[22] = rdfint_0n[22];
  assign rd_0r0d[23] = rdfint_0n[23];
  assign rd_0r0d[24] = rdfint_0n[24];
  assign rd_0r0d[25] = rdfint_0n[25];
  assign rd_0r0d[26] = rdfint_0n[26];
  assign rd_0r0d[27] = rdfint_0n[27];
  assign rd_0r0d[28] = rdfint_0n[28];
  assign rd_0r0d[29] = rdfint_0n[29];
  assign rd_0r0d[30] = rdfint_0n[30];
  assign rd_0r0d[31] = rdfint_0n[31];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign rd_0r1d[10] = rdtint_0n[10];
  assign rd_0r1d[11] = rdtint_0n[11];
  assign rd_0r1d[12] = rdtint_0n[12];
  assign rd_0r1d[13] = rdtint_0n[13];
  assign rd_0r1d[14] = rdtint_0n[14];
  assign rd_0r1d[15] = rdtint_0n[15];
  assign rd_0r1d[16] = rdtint_0n[16];
  assign rd_0r1d[17] = rdtint_0n[17];
  assign rd_0r1d[18] = rdtint_0n[18];
  assign rd_0r1d[19] = rdtint_0n[19];
  assign rd_0r1d[20] = rdtint_0n[20];
  assign rd_0r1d[21] = rdtint_0n[21];
  assign rd_0r1d[22] = rdtint_0n[22];
  assign rd_0r1d[23] = rdtint_0n[23];
  assign rd_0r1d[24] = rdtint_0n[24];
  assign rd_0r1d[25] = rdtint_0n[25];
  assign rd_0r1d[26] = rdtint_0n[26];
  assign rd_0r1d[27] = rdtint_0n[27];
  assign rd_0r1d[28] = rdtint_0n[28];
  assign rd_0r1d[29] = rdtint_0n[29];
  assign rd_0r1d[30] = rdtint_0n[30];
  assign rd_0r1d[31] = rdtint_0n[31];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgfint_0n[32] = wg_0r0d[32];
  assign wgfint_0n[33] = wg_0r0d[33];
  assign wgfint_0n[34] = wg_0r0d[34];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign wgtint_0n[32] = wg_0r1d[32];
  assign wgtint_0n[33] = wg_0r1d[33];
  assign wgtint_0n[34] = wg_0r1d[34];
  assign rg_3a = rgaint_3n;
  assign rgrint_3n = rg_3r;
  assign rg_2a = rgaint_2n;
  assign rgrint_2n = rg_2r;
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR3 I219 (internal_0n[0], rgrint_0n, rgrint_1n, rgrint_2n);
  NOR3 I220 (internal_0n[1], rgrint_3n, rgaint_0n, rgaint_1n);
  NOR2 I221 (internal_0n[2], rgaint_2n, rgaint_3n);
  AND3 I222 (nanyread_0n, internal_0n[0], internal_0n[1], internal_0n[2]);
  AND2 I223 (rdtint_3n[0], rgrint_3n, dt_0n[2]);
  AND2 I224 (rdtint_3n[1], rgrint_3n, dt_0n[3]);
  AND2 I225 (rdtint_3n[2], rgrint_3n, dt_0n[4]);
  AND2 I226 (rdtint_3n[3], rgrint_3n, dt_0n[5]);
  AND2 I227 (rdtint_3n[4], rgrint_3n, dt_0n[6]);
  AND2 I228 (rdtint_3n[5], rgrint_3n, dt_0n[7]);
  AND2 I229 (rdtint_3n[6], rgrint_3n, dt_0n[8]);
  AND2 I230 (rdtint_3n[7], rgrint_3n, dt_0n[9]);
  AND2 I231 (rdtint_3n[8], rgrint_3n, dt_0n[10]);
  AND2 I232 (rdtint_3n[9], rgrint_3n, dt_0n[11]);
  AND2 I233 (rdtint_3n[10], rgrint_3n, dt_0n[12]);
  AND2 I234 (rdtint_3n[11], rgrint_3n, dt_0n[13]);
  AND2 I235 (rdtint_3n[12], rgrint_3n, dt_0n[14]);
  AND2 I236 (rdtint_3n[13], rgrint_3n, dt_0n[15]);
  AND2 I237 (rdtint_3n[14], rgrint_3n, dt_0n[16]);
  AND2 I238 (rdtint_3n[15], rgrint_3n, dt_0n[17]);
  AND2 I239 (rdtint_3n[16], rgrint_3n, dt_0n[18]);
  AND2 I240 (rdtint_3n[17], rgrint_3n, dt_0n[19]);
  AND2 I241 (rdtint_3n[18], rgrint_3n, dt_0n[20]);
  AND2 I242 (rdtint_3n[19], rgrint_3n, dt_0n[21]);
  AND2 I243 (rdtint_3n[20], rgrint_3n, dt_0n[22]);
  AND2 I244 (rdtint_3n[21], rgrint_3n, dt_0n[23]);
  AND2 I245 (rdtint_3n[22], rgrint_3n, dt_0n[24]);
  AND2 I246 (rdtint_3n[23], rgrint_3n, dt_0n[25]);
  AND2 I247 (rdtint_3n[24], rgrint_3n, dt_0n[26]);
  AND2 I248 (rdtint_3n[25], rgrint_3n, dt_0n[27]);
  AND2 I249 (rdtint_3n[26], rgrint_3n, dt_0n[28]);
  AND2 I250 (rdtint_3n[27], rgrint_3n, dt_0n[29]);
  AND2 I251 (rdtint_3n[28], rgrint_3n, dt_0n[30]);
  AND2 I252 (rdtint_3n[29], rgrint_3n, dt_0n[31]);
  AND2 I253 (rdtint_3n[30], rgrint_3n, dt_0n[32]);
  AND2 I254 (rdtint_3n[31], rgrint_3n, dt_0n[33]);
  AND2 I255 (rdtint_3n[32], rgrint_3n, dt_0n[34]);
  AND2 I256 (rdtint_2n, rgrint_2n, dt_0n[34]);
  AND2 I257 (rdtint_1n, rgrint_1n, dt_0n[34]);
  AND2 I258 (rdtint_0n[0], rgrint_0n, dt_0n[1]);
  AND2 I259 (rdtint_0n[1], rgrint_0n, dt_0n[2]);
  AND2 I260 (rdtint_0n[2], rgrint_0n, dt_0n[3]);
  AND2 I261 (rdtint_0n[3], rgrint_0n, dt_0n[4]);
  AND2 I262 (rdtint_0n[4], rgrint_0n, dt_0n[5]);
  AND2 I263 (rdtint_0n[5], rgrint_0n, dt_0n[6]);
  AND2 I264 (rdtint_0n[6], rgrint_0n, dt_0n[7]);
  AND2 I265 (rdtint_0n[7], rgrint_0n, dt_0n[8]);
  AND2 I266 (rdtint_0n[8], rgrint_0n, dt_0n[9]);
  AND2 I267 (rdtint_0n[9], rgrint_0n, dt_0n[10]);
  AND2 I268 (rdtint_0n[10], rgrint_0n, dt_0n[11]);
  AND2 I269 (rdtint_0n[11], rgrint_0n, dt_0n[12]);
  AND2 I270 (rdtint_0n[12], rgrint_0n, dt_0n[13]);
  AND2 I271 (rdtint_0n[13], rgrint_0n, dt_0n[14]);
  AND2 I272 (rdtint_0n[14], rgrint_0n, dt_0n[15]);
  AND2 I273 (rdtint_0n[15], rgrint_0n, dt_0n[16]);
  AND2 I274 (rdtint_0n[16], rgrint_0n, dt_0n[17]);
  AND2 I275 (rdtint_0n[17], rgrint_0n, dt_0n[18]);
  AND2 I276 (rdtint_0n[18], rgrint_0n, dt_0n[19]);
  AND2 I277 (rdtint_0n[19], rgrint_0n, dt_0n[20]);
  AND2 I278 (rdtint_0n[20], rgrint_0n, dt_0n[21]);
  AND2 I279 (rdtint_0n[21], rgrint_0n, dt_0n[22]);
  AND2 I280 (rdtint_0n[22], rgrint_0n, dt_0n[23]);
  AND2 I281 (rdtint_0n[23], rgrint_0n, dt_0n[24]);
  AND2 I282 (rdtint_0n[24], rgrint_0n, dt_0n[25]);
  AND2 I283 (rdtint_0n[25], rgrint_0n, dt_0n[26]);
  AND2 I284 (rdtint_0n[26], rgrint_0n, dt_0n[27]);
  AND2 I285 (rdtint_0n[27], rgrint_0n, dt_0n[28]);
  AND2 I286 (rdtint_0n[28], rgrint_0n, dt_0n[29]);
  AND2 I287 (rdtint_0n[29], rgrint_0n, dt_0n[30]);
  AND2 I288 (rdtint_0n[30], rgrint_0n, dt_0n[31]);
  AND2 I289 (rdtint_0n[31], rgrint_0n, dt_0n[32]);
  AND2 I290 (rdfint_3n[0], rgrint_3n, df_0n[2]);
  AND2 I291 (rdfint_3n[1], rgrint_3n, df_0n[3]);
  AND2 I292 (rdfint_3n[2], rgrint_3n, df_0n[4]);
  AND2 I293 (rdfint_3n[3], rgrint_3n, df_0n[5]);
  AND2 I294 (rdfint_3n[4], rgrint_3n, df_0n[6]);
  AND2 I295 (rdfint_3n[5], rgrint_3n, df_0n[7]);
  AND2 I296 (rdfint_3n[6], rgrint_3n, df_0n[8]);
  AND2 I297 (rdfint_3n[7], rgrint_3n, df_0n[9]);
  AND2 I298 (rdfint_3n[8], rgrint_3n, df_0n[10]);
  AND2 I299 (rdfint_3n[9], rgrint_3n, df_0n[11]);
  AND2 I300 (rdfint_3n[10], rgrint_3n, df_0n[12]);
  AND2 I301 (rdfint_3n[11], rgrint_3n, df_0n[13]);
  AND2 I302 (rdfint_3n[12], rgrint_3n, df_0n[14]);
  AND2 I303 (rdfint_3n[13], rgrint_3n, df_0n[15]);
  AND2 I304 (rdfint_3n[14], rgrint_3n, df_0n[16]);
  AND2 I305 (rdfint_3n[15], rgrint_3n, df_0n[17]);
  AND2 I306 (rdfint_3n[16], rgrint_3n, df_0n[18]);
  AND2 I307 (rdfint_3n[17], rgrint_3n, df_0n[19]);
  AND2 I308 (rdfint_3n[18], rgrint_3n, df_0n[20]);
  AND2 I309 (rdfint_3n[19], rgrint_3n, df_0n[21]);
  AND2 I310 (rdfint_3n[20], rgrint_3n, df_0n[22]);
  AND2 I311 (rdfint_3n[21], rgrint_3n, df_0n[23]);
  AND2 I312 (rdfint_3n[22], rgrint_3n, df_0n[24]);
  AND2 I313 (rdfint_3n[23], rgrint_3n, df_0n[25]);
  AND2 I314 (rdfint_3n[24], rgrint_3n, df_0n[26]);
  AND2 I315 (rdfint_3n[25], rgrint_3n, df_0n[27]);
  AND2 I316 (rdfint_3n[26], rgrint_3n, df_0n[28]);
  AND2 I317 (rdfint_3n[27], rgrint_3n, df_0n[29]);
  AND2 I318 (rdfint_3n[28], rgrint_3n, df_0n[30]);
  AND2 I319 (rdfint_3n[29], rgrint_3n, df_0n[31]);
  AND2 I320 (rdfint_3n[30], rgrint_3n, df_0n[32]);
  AND2 I321 (rdfint_3n[31], rgrint_3n, df_0n[33]);
  AND2 I322 (rdfint_3n[32], rgrint_3n, df_0n[34]);
  AND2 I323 (rdfint_2n, rgrint_2n, df_0n[34]);
  AND2 I324 (rdfint_1n, rgrint_1n, df_0n[34]);
  AND2 I325 (rdfint_0n[0], rgrint_0n, df_0n[1]);
  AND2 I326 (rdfint_0n[1], rgrint_0n, df_0n[2]);
  AND2 I327 (rdfint_0n[2], rgrint_0n, df_0n[3]);
  AND2 I328 (rdfint_0n[3], rgrint_0n, df_0n[4]);
  AND2 I329 (rdfint_0n[4], rgrint_0n, df_0n[5]);
  AND2 I330 (rdfint_0n[5], rgrint_0n, df_0n[6]);
  AND2 I331 (rdfint_0n[6], rgrint_0n, df_0n[7]);
  AND2 I332 (rdfint_0n[7], rgrint_0n, df_0n[8]);
  AND2 I333 (rdfint_0n[8], rgrint_0n, df_0n[9]);
  AND2 I334 (rdfint_0n[9], rgrint_0n, df_0n[10]);
  AND2 I335 (rdfint_0n[10], rgrint_0n, df_0n[11]);
  AND2 I336 (rdfint_0n[11], rgrint_0n, df_0n[12]);
  AND2 I337 (rdfint_0n[12], rgrint_0n, df_0n[13]);
  AND2 I338 (rdfint_0n[13], rgrint_0n, df_0n[14]);
  AND2 I339 (rdfint_0n[14], rgrint_0n, df_0n[15]);
  AND2 I340 (rdfint_0n[15], rgrint_0n, df_0n[16]);
  AND2 I341 (rdfint_0n[16], rgrint_0n, df_0n[17]);
  AND2 I342 (rdfint_0n[17], rgrint_0n, df_0n[18]);
  AND2 I343 (rdfint_0n[18], rgrint_0n, df_0n[19]);
  AND2 I344 (rdfint_0n[19], rgrint_0n, df_0n[20]);
  AND2 I345 (rdfint_0n[20], rgrint_0n, df_0n[21]);
  AND2 I346 (rdfint_0n[21], rgrint_0n, df_0n[22]);
  AND2 I347 (rdfint_0n[22], rgrint_0n, df_0n[23]);
  AND2 I348 (rdfint_0n[23], rgrint_0n, df_0n[24]);
  AND2 I349 (rdfint_0n[24], rgrint_0n, df_0n[25]);
  AND2 I350 (rdfint_0n[25], rgrint_0n, df_0n[26]);
  AND2 I351 (rdfint_0n[26], rgrint_0n, df_0n[27]);
  AND2 I352 (rdfint_0n[27], rgrint_0n, df_0n[28]);
  AND2 I353 (rdfint_0n[28], rgrint_0n, df_0n[29]);
  AND2 I354 (rdfint_0n[29], rgrint_0n, df_0n[30]);
  AND2 I355 (rdfint_0n[30], rgrint_0n, df_0n[31]);
  AND2 I356 (rdfint_0n[31], rgrint_0n, df_0n[32]);
  C3 I357 (internal_0n[3], wc_0n, wacks_0n[34], wacks_0n[33]);
  C3 I358 (internal_0n[4], wacks_0n[32], wacks_0n[31], wacks_0n[30]);
  C3 I359 (internal_0n[5], wacks_0n[29], wacks_0n[28], wacks_0n[27]);
  C3 I360 (internal_0n[6], wacks_0n[26], wacks_0n[25], wacks_0n[24]);
  C3 I361 (internal_0n[7], wacks_0n[23], wacks_0n[22], wacks_0n[21]);
  C3 I362 (internal_0n[8], wacks_0n[20], wacks_0n[19], wacks_0n[18]);
  C3 I363 (internal_0n[9], wacks_0n[17], wacks_0n[16], wacks_0n[15]);
  C3 I364 (internal_0n[10], wacks_0n[14], wacks_0n[13], wacks_0n[12]);
  C3 I365 (internal_0n[11], wacks_0n[11], wacks_0n[10], wacks_0n[9]);
  C3 I366 (internal_0n[12], wacks_0n[8], wacks_0n[7], wacks_0n[6]);
  C3 I367 (internal_0n[13], wacks_0n[5], wacks_0n[4], wacks_0n[3]);
  C3 I368 (internal_0n[14], wacks_0n[2], wacks_0n[1], wacks_0n[0]);
  C3 I369 (internal_0n[15], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I370 (internal_0n[16], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I371 (internal_0n[17], internal_0n[9], internal_0n[10], internal_0n[11]);
  C3 I372 (internal_0n[18], internal_0n[12], internal_0n[13], internal_0n[14]);
  C2 I373 (internal_0n[19], internal_0n[15], internal_0n[16]);
  C2 I374 (internal_0n[20], internal_0n[17], internal_0n[18]);
  C2 I375 (wdrint_0n, internal_0n[19], internal_0n[20]);
  assign wen_0n[34] = wc_0n;
  assign wen_0n[33] = wc_0n;
  assign wen_0n[32] = wc_0n;
  assign wen_0n[31] = wc_0n;
  assign wen_0n[30] = wc_0n;
  assign wen_0n[29] = wc_0n;
  assign wen_0n[28] = wc_0n;
  assign wen_0n[27] = wc_0n;
  assign wen_0n[26] = wc_0n;
  assign wen_0n[25] = wc_0n;
  assign wen_0n[24] = wc_0n;
  assign wen_0n[23] = wc_0n;
  assign wen_0n[22] = wc_0n;
  assign wen_0n[21] = wc_0n;
  assign wen_0n[20] = wc_0n;
  assign wen_0n[19] = wc_0n;
  assign wen_0n[18] = wc_0n;
  assign wen_0n[17] = wc_0n;
  assign wen_0n[16] = wc_0n;
  assign wen_0n[15] = wc_0n;
  assign wen_0n[14] = wc_0n;
  assign wen_0n[13] = wc_0n;
  assign wen_0n[12] = wc_0n;
  assign wen_0n[11] = wc_0n;
  assign wen_0n[10] = wc_0n;
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[34] = git_0n[34];
  assign wt_0n[33] = git_0n[33];
  assign wt_0n[32] = git_0n[32];
  assign wt_0n[31] = git_0n[31];
  assign wt_0n[30] = git_0n[30];
  assign wt_0n[29] = git_0n[29];
  assign wt_0n[28] = git_0n[28];
  assign wt_0n[27] = git_0n[27];
  assign wt_0n[26] = git_0n[26];
  assign wt_0n[25] = git_0n[25];
  assign wt_0n[24] = git_0n[24];
  assign wt_0n[23] = git_0n[23];
  assign wt_0n[22] = git_0n[22];
  assign wt_0n[21] = git_0n[21];
  assign wt_0n[20] = git_0n[20];
  assign wt_0n[19] = git_0n[19];
  assign wt_0n[18] = git_0n[18];
  assign wt_0n[17] = git_0n[17];
  assign wt_0n[16] = git_0n[16];
  assign wt_0n[15] = git_0n[15];
  assign wt_0n[14] = git_0n[14];
  assign wt_0n[13] = git_0n[13];
  assign wt_0n[12] = git_0n[12];
  assign wt_0n[11] = git_0n[11];
  assign wt_0n[10] = git_0n[10];
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[34] = gif_0n[34];
  assign wf_0n[33] = gif_0n[33];
  assign wf_0n[32] = gif_0n[32];
  assign wf_0n[31] = gif_0n[31];
  assign wf_0n[30] = gif_0n[30];
  assign wf_0n[29] = gif_0n[29];
  assign wf_0n[28] = gif_0n[28];
  assign wf_0n[27] = gif_0n[27];
  assign wf_0n[26] = gif_0n[26];
  assign wf_0n[25] = gif_0n[25];
  assign wf_0n[24] = gif_0n[24];
  assign wf_0n[23] = gif_0n[23];
  assign wf_0n[22] = gif_0n[22];
  assign wf_0n[21] = gif_0n[21];
  assign wf_0n[20] = gif_0n[20];
  assign wf_0n[19] = gif_0n[19];
  assign wf_0n[18] = gif_0n[18];
  assign wf_0n[17] = gif_0n[17];
  assign wf_0n[16] = gif_0n[16];
  assign wf_0n[15] = gif_0n[15];
  assign wf_0n[14] = gif_0n[14];
  assign wf_0n[13] = gif_0n[13];
  assign wf_0n[12] = gif_0n[12];
  assign wf_0n[11] = gif_0n[11];
  assign wf_0n[10] = gif_0n[10];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I481 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I483 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I484 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I485 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I486 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I487 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I488 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I489 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I490 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I491 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I492 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I493 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I494 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I495 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I496 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I497 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I498 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I499 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I500 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I501 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I502 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I503 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I504 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I505 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I506 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I507 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I508 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I509 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I510 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I511 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I512 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I513 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I514 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I515 (git_0n[32], wgtint_0n[32], ig_0n);
  AND2 I516 (git_0n[33], wgtint_0n[33], ig_0n);
  AND2 I517 (git_0n[34], wgtint_0n[34], ig_0n);
  AND2 I518 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I519 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I520 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I521 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I522 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I523 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I524 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I525 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I526 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I527 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I528 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I529 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I530 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I531 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I532 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I533 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I534 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I535 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I536 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I537 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I538 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I539 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I540 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I541 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I542 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I543 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I544 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I545 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I546 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I547 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I548 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I549 (gif_0n[31], wgfint_0n[31], ig_0n);
  AND2 I550 (gif_0n[32], wgfint_0n[32], ig_0n);
  AND2 I551 (gif_0n[33], wgfint_0n[33], ig_0n);
  AND2 I552 (gif_0n[34], wgfint_0n[34], ig_0n);
  C3 I553 (internal_0n[21], complete1520_0n[0], complete1520_0n[1], complete1520_0n[2]);
  C3 I554 (internal_0n[22], complete1520_0n[3], complete1520_0n[4], complete1520_0n[5]);
  C3 I555 (internal_0n[23], complete1520_0n[6], complete1520_0n[7], complete1520_0n[8]);
  C3 I556 (internal_0n[24], complete1520_0n[9], complete1520_0n[10], complete1520_0n[11]);
  C3 I557 (internal_0n[25], complete1520_0n[12], complete1520_0n[13], complete1520_0n[14]);
  C3 I558 (internal_0n[26], complete1520_0n[15], complete1520_0n[16], complete1520_0n[17]);
  C3 I559 (internal_0n[27], complete1520_0n[18], complete1520_0n[19], complete1520_0n[20]);
  C3 I560 (internal_0n[28], complete1520_0n[21], complete1520_0n[22], complete1520_0n[23]);
  C3 I561 (internal_0n[29], complete1520_0n[24], complete1520_0n[25], complete1520_0n[26]);
  C3 I562 (internal_0n[30], complete1520_0n[27], complete1520_0n[28], complete1520_0n[29]);
  C3 I563 (internal_0n[31], complete1520_0n[30], complete1520_0n[31], complete1520_0n[32]);
  C2 I564 (internal_0n[32], complete1520_0n[33], complete1520_0n[34]);
  C3 I565 (internal_0n[33], internal_0n[21], internal_0n[22], internal_0n[23]);
  C3 I566 (internal_0n[34], internal_0n[24], internal_0n[25], internal_0n[26]);
  C3 I567 (internal_0n[35], internal_0n[27], internal_0n[28], internal_0n[29]);
  C3 I568 (internal_0n[36], internal_0n[30], internal_0n[31], internal_0n[32]);
  C2 I569 (internal_0n[37], internal_0n[33], internal_0n[34]);
  C2 I570 (internal_0n[38], internal_0n[35], internal_0n[36]);
  C2 I571 (wc_0n, internal_0n[37], internal_0n[38]);
  OR2 I572 (complete1520_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I573 (complete1520_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I574 (complete1520_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I575 (complete1520_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I576 (complete1520_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I577 (complete1520_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I578 (complete1520_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I579 (complete1520_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I580 (complete1520_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I581 (complete1520_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I582 (complete1520_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I583 (complete1520_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I584 (complete1520_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I585 (complete1520_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I586 (complete1520_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I587 (complete1520_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I588 (complete1520_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I589 (complete1520_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I590 (complete1520_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I591 (complete1520_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I592 (complete1520_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I593 (complete1520_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I594 (complete1520_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I595 (complete1520_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I596 (complete1520_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I597 (complete1520_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I598 (complete1520_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I599 (complete1520_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I600 (complete1520_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I601 (complete1520_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I602 (complete1520_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I603 (complete1520_0n[31], wgfint_0n[31], wgtint_0n[31]);
  OR2 I604 (complete1520_0n[32], wgfint_0n[32], wgtint_0n[32]);
  OR2 I605 (complete1520_0n[33], wgfint_0n[33], wgtint_0n[33]);
  OR2 I606 (complete1520_0n[34], wgfint_0n[34], wgtint_0n[34]);
  AO22 I607 (wacks_0n[34], gf1518_0n[34], df_0n[34], gt1519_0n[34], dt_0n[34]);
  NOR2 I608 (dt_0n[34], df_0n[34], gf1518_0n[34]);
  NOR3 I609 (df_0n[34], dt_0n[34], gt1519_0n[34], init_0n);
  AND2 I610 (gt1519_0n[34], wt_0n[34], wen_0n[34]);
  AND2 I611 (gf1518_0n[34], wf_0n[34], wen_0n[34]);
  AO22 I612 (wacks_0n[33], gf1518_0n[33], df_0n[33], gt1519_0n[33], dt_0n[33]);
  NOR2 I613 (dt_0n[33], df_0n[33], gf1518_0n[33]);
  NOR3 I614 (df_0n[33], dt_0n[33], gt1519_0n[33], init_0n);
  AND2 I615 (gt1519_0n[33], wt_0n[33], wen_0n[33]);
  AND2 I616 (gf1518_0n[33], wf_0n[33], wen_0n[33]);
  AO22 I617 (wacks_0n[32], gf1518_0n[32], df_0n[32], gt1519_0n[32], dt_0n[32]);
  NOR2 I618 (dt_0n[32], df_0n[32], gf1518_0n[32]);
  NOR3 I619 (df_0n[32], dt_0n[32], gt1519_0n[32], init_0n);
  AND2 I620 (gt1519_0n[32], wt_0n[32], wen_0n[32]);
  AND2 I621 (gf1518_0n[32], wf_0n[32], wen_0n[32]);
  AO22 I622 (wacks_0n[31], gf1518_0n[31], df_0n[31], gt1519_0n[31], dt_0n[31]);
  NOR2 I623 (dt_0n[31], df_0n[31], gf1518_0n[31]);
  NOR3 I624 (df_0n[31], dt_0n[31], gt1519_0n[31], init_0n);
  AND2 I625 (gt1519_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I626 (gf1518_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I627 (wacks_0n[30], gf1518_0n[30], df_0n[30], gt1519_0n[30], dt_0n[30]);
  NOR2 I628 (dt_0n[30], df_0n[30], gf1518_0n[30]);
  NOR3 I629 (df_0n[30], dt_0n[30], gt1519_0n[30], init_0n);
  AND2 I630 (gt1519_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I631 (gf1518_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I632 (wacks_0n[29], gf1518_0n[29], df_0n[29], gt1519_0n[29], dt_0n[29]);
  NOR2 I633 (dt_0n[29], df_0n[29], gf1518_0n[29]);
  NOR3 I634 (df_0n[29], dt_0n[29], gt1519_0n[29], init_0n);
  AND2 I635 (gt1519_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I636 (gf1518_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I637 (wacks_0n[28], gf1518_0n[28], df_0n[28], gt1519_0n[28], dt_0n[28]);
  NOR2 I638 (dt_0n[28], df_0n[28], gf1518_0n[28]);
  NOR3 I639 (df_0n[28], dt_0n[28], gt1519_0n[28], init_0n);
  AND2 I640 (gt1519_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I641 (gf1518_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I642 (wacks_0n[27], gf1518_0n[27], df_0n[27], gt1519_0n[27], dt_0n[27]);
  NOR2 I643 (dt_0n[27], df_0n[27], gf1518_0n[27]);
  NOR3 I644 (df_0n[27], dt_0n[27], gt1519_0n[27], init_0n);
  AND2 I645 (gt1519_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I646 (gf1518_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I647 (wacks_0n[26], gf1518_0n[26], df_0n[26], gt1519_0n[26], dt_0n[26]);
  NOR2 I648 (dt_0n[26], df_0n[26], gf1518_0n[26]);
  NOR3 I649 (df_0n[26], dt_0n[26], gt1519_0n[26], init_0n);
  AND2 I650 (gt1519_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I651 (gf1518_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I652 (wacks_0n[25], gf1518_0n[25], df_0n[25], gt1519_0n[25], dt_0n[25]);
  NOR2 I653 (dt_0n[25], df_0n[25], gf1518_0n[25]);
  NOR3 I654 (df_0n[25], dt_0n[25], gt1519_0n[25], init_0n);
  AND2 I655 (gt1519_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I656 (gf1518_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I657 (wacks_0n[24], gf1518_0n[24], df_0n[24], gt1519_0n[24], dt_0n[24]);
  NOR2 I658 (dt_0n[24], df_0n[24], gf1518_0n[24]);
  NOR3 I659 (df_0n[24], dt_0n[24], gt1519_0n[24], init_0n);
  AND2 I660 (gt1519_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I661 (gf1518_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I662 (wacks_0n[23], gf1518_0n[23], df_0n[23], gt1519_0n[23], dt_0n[23]);
  NOR2 I663 (dt_0n[23], df_0n[23], gf1518_0n[23]);
  NOR3 I664 (df_0n[23], dt_0n[23], gt1519_0n[23], init_0n);
  AND2 I665 (gt1519_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I666 (gf1518_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I667 (wacks_0n[22], gf1518_0n[22], df_0n[22], gt1519_0n[22], dt_0n[22]);
  NOR2 I668 (dt_0n[22], df_0n[22], gf1518_0n[22]);
  NOR3 I669 (df_0n[22], dt_0n[22], gt1519_0n[22], init_0n);
  AND2 I670 (gt1519_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I671 (gf1518_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I672 (wacks_0n[21], gf1518_0n[21], df_0n[21], gt1519_0n[21], dt_0n[21]);
  NOR2 I673 (dt_0n[21], df_0n[21], gf1518_0n[21]);
  NOR3 I674 (df_0n[21], dt_0n[21], gt1519_0n[21], init_0n);
  AND2 I675 (gt1519_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I676 (gf1518_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I677 (wacks_0n[20], gf1518_0n[20], df_0n[20], gt1519_0n[20], dt_0n[20]);
  NOR2 I678 (dt_0n[20], df_0n[20], gf1518_0n[20]);
  NOR3 I679 (df_0n[20], dt_0n[20], gt1519_0n[20], init_0n);
  AND2 I680 (gt1519_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I681 (gf1518_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I682 (wacks_0n[19], gf1518_0n[19], df_0n[19], gt1519_0n[19], dt_0n[19]);
  NOR2 I683 (dt_0n[19], df_0n[19], gf1518_0n[19]);
  NOR3 I684 (df_0n[19], dt_0n[19], gt1519_0n[19], init_0n);
  AND2 I685 (gt1519_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I686 (gf1518_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I687 (wacks_0n[18], gf1518_0n[18], df_0n[18], gt1519_0n[18], dt_0n[18]);
  NOR2 I688 (dt_0n[18], df_0n[18], gf1518_0n[18]);
  NOR3 I689 (df_0n[18], dt_0n[18], gt1519_0n[18], init_0n);
  AND2 I690 (gt1519_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I691 (gf1518_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I692 (wacks_0n[17], gf1518_0n[17], df_0n[17], gt1519_0n[17], dt_0n[17]);
  NOR2 I693 (dt_0n[17], df_0n[17], gf1518_0n[17]);
  NOR3 I694 (df_0n[17], dt_0n[17], gt1519_0n[17], init_0n);
  AND2 I695 (gt1519_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I696 (gf1518_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I697 (wacks_0n[16], gf1518_0n[16], df_0n[16], gt1519_0n[16], dt_0n[16]);
  NOR2 I698 (dt_0n[16], df_0n[16], gf1518_0n[16]);
  NOR3 I699 (df_0n[16], dt_0n[16], gt1519_0n[16], init_0n);
  AND2 I700 (gt1519_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I701 (gf1518_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I702 (wacks_0n[15], gf1518_0n[15], df_0n[15], gt1519_0n[15], dt_0n[15]);
  NOR2 I703 (dt_0n[15], df_0n[15], gf1518_0n[15]);
  NOR3 I704 (df_0n[15], dt_0n[15], gt1519_0n[15], init_0n);
  AND2 I705 (gt1519_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I706 (gf1518_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I707 (wacks_0n[14], gf1518_0n[14], df_0n[14], gt1519_0n[14], dt_0n[14]);
  NOR2 I708 (dt_0n[14], df_0n[14], gf1518_0n[14]);
  NOR3 I709 (df_0n[14], dt_0n[14], gt1519_0n[14], init_0n);
  AND2 I710 (gt1519_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I711 (gf1518_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I712 (wacks_0n[13], gf1518_0n[13], df_0n[13], gt1519_0n[13], dt_0n[13]);
  NOR2 I713 (dt_0n[13], df_0n[13], gf1518_0n[13]);
  NOR3 I714 (df_0n[13], dt_0n[13], gt1519_0n[13], init_0n);
  AND2 I715 (gt1519_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I716 (gf1518_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I717 (wacks_0n[12], gf1518_0n[12], df_0n[12], gt1519_0n[12], dt_0n[12]);
  NOR2 I718 (dt_0n[12], df_0n[12], gf1518_0n[12]);
  NOR3 I719 (df_0n[12], dt_0n[12], gt1519_0n[12], init_0n);
  AND2 I720 (gt1519_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I721 (gf1518_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I722 (wacks_0n[11], gf1518_0n[11], df_0n[11], gt1519_0n[11], dt_0n[11]);
  NOR2 I723 (dt_0n[11], df_0n[11], gf1518_0n[11]);
  NOR3 I724 (df_0n[11], dt_0n[11], gt1519_0n[11], init_0n);
  AND2 I725 (gt1519_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I726 (gf1518_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I727 (wacks_0n[10], gf1518_0n[10], df_0n[10], gt1519_0n[10], dt_0n[10]);
  NOR2 I728 (dt_0n[10], df_0n[10], gf1518_0n[10]);
  NOR3 I729 (df_0n[10], dt_0n[10], gt1519_0n[10], init_0n);
  AND2 I730 (gt1519_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I731 (gf1518_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I732 (wacks_0n[9], gf1518_0n[9], df_0n[9], gt1519_0n[9], dt_0n[9]);
  NOR2 I733 (dt_0n[9], df_0n[9], gf1518_0n[9]);
  NOR3 I734 (df_0n[9], dt_0n[9], gt1519_0n[9], init_0n);
  AND2 I735 (gt1519_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I736 (gf1518_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I737 (wacks_0n[8], gf1518_0n[8], df_0n[8], gt1519_0n[8], dt_0n[8]);
  NOR2 I738 (dt_0n[8], df_0n[8], gf1518_0n[8]);
  NOR3 I739 (df_0n[8], dt_0n[8], gt1519_0n[8], init_0n);
  AND2 I740 (gt1519_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I741 (gf1518_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I742 (wacks_0n[7], gf1518_0n[7], df_0n[7], gt1519_0n[7], dt_0n[7]);
  NOR2 I743 (dt_0n[7], df_0n[7], gf1518_0n[7]);
  NOR3 I744 (df_0n[7], dt_0n[7], gt1519_0n[7], init_0n);
  AND2 I745 (gt1519_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I746 (gf1518_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I747 (wacks_0n[6], gf1518_0n[6], df_0n[6], gt1519_0n[6], dt_0n[6]);
  NOR2 I748 (dt_0n[6], df_0n[6], gf1518_0n[6]);
  NOR3 I749 (df_0n[6], dt_0n[6], gt1519_0n[6], init_0n);
  AND2 I750 (gt1519_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I751 (gf1518_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I752 (wacks_0n[5], gf1518_0n[5], df_0n[5], gt1519_0n[5], dt_0n[5]);
  NOR2 I753 (dt_0n[5], df_0n[5], gf1518_0n[5]);
  NOR3 I754 (df_0n[5], dt_0n[5], gt1519_0n[5], init_0n);
  AND2 I755 (gt1519_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I756 (gf1518_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I757 (wacks_0n[4], gf1518_0n[4], df_0n[4], gt1519_0n[4], dt_0n[4]);
  NOR2 I758 (dt_0n[4], df_0n[4], gf1518_0n[4]);
  NOR3 I759 (df_0n[4], dt_0n[4], gt1519_0n[4], init_0n);
  AND2 I760 (gt1519_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I761 (gf1518_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I762 (wacks_0n[3], gf1518_0n[3], df_0n[3], gt1519_0n[3], dt_0n[3]);
  NOR2 I763 (dt_0n[3], df_0n[3], gf1518_0n[3]);
  NOR3 I764 (df_0n[3], dt_0n[3], gt1519_0n[3], init_0n);
  AND2 I765 (gt1519_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I766 (gf1518_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I767 (wacks_0n[2], gf1518_0n[2], df_0n[2], gt1519_0n[2], dt_0n[2]);
  NOR2 I768 (dt_0n[2], df_0n[2], gf1518_0n[2]);
  NOR3 I769 (df_0n[2], dt_0n[2], gt1519_0n[2], init_0n);
  AND2 I770 (gt1519_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I771 (gf1518_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I772 (wacks_0n[1], gf1518_0n[1], df_0n[1], gt1519_0n[1], dt_0n[1]);
  NOR2 I773 (dt_0n[1], df_0n[1], gf1518_0n[1]);
  NOR3 I774 (df_0n[1], dt_0n[1], gt1519_0n[1], init_0n);
  AND2 I775 (gt1519_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I776 (gf1518_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I777 (wacks_0n[0], gf1518_0n[0], df_0n[0], gt1519_0n[0], dt_0n[0]);
  NOR2 I778 (dt_0n[0], df_0n[0], gf1518_0n[0]);
  NOR3 I779 (df_0n[0], dt_0n[0], gt1519_0n[0], init_0n);
  AND2 I780 (gt1519_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I781 (gf1518_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I782 (init_0n, initialise);
endmodule

module BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m93m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  initialise
);
  input [34:0] wg_0r0d;
  input [34:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [31:0] rd_0r0d;
  output [31:0] rd_0r1d;
  input rd_0a;
  output [2:0] rd_1r0d;
  output [2:0] rd_1r1d;
  input rd_1a;
  input initialise;
  wire [37:0] internal_0n;
  wire [34:0] wf_0n;
  wire [34:0] wt_0n;
  wire [34:0] df_0n;
  wire [34:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire wc_0n;
  wire [34:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [34:0] wgfint_0n;
  wire [34:0] wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire [31:0] rdfint_0n;
  wire [2:0] rdfint_1n;
  wire [31:0] rdtint_0n;
  wire [2:0] rdtint_1n;
  wire [34:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [34:0] gif_0n;
  wire [34:0] git_0n;
  wire [34:0] complete1543_0n;
  wire [34:0] gt1542_0n;
  wire [34:0] gf1541_0n;
  assign rgaint_1n = rd_1a;
  assign rd_1r0d[0] = rdfint_1n[0];
  assign rd_1r0d[1] = rdfint_1n[1];
  assign rd_1r0d[2] = rdfint_1n[2];
  assign rd_1r1d[0] = rdtint_1n[0];
  assign rd_1r1d[1] = rdtint_1n[1];
  assign rd_1r1d[2] = rdtint_1n[2];
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r0d[10] = rdfint_0n[10];
  assign rd_0r0d[11] = rdfint_0n[11];
  assign rd_0r0d[12] = rdfint_0n[12];
  assign rd_0r0d[13] = rdfint_0n[13];
  assign rd_0r0d[14] = rdfint_0n[14];
  assign rd_0r0d[15] = rdfint_0n[15];
  assign rd_0r0d[16] = rdfint_0n[16];
  assign rd_0r0d[17] = rdfint_0n[17];
  assign rd_0r0d[18] = rdfint_0n[18];
  assign rd_0r0d[19] = rdfint_0n[19];
  assign rd_0r0d[20] = rdfint_0n[20];
  assign rd_0r0d[21] = rdfint_0n[21];
  assign rd_0r0d[22] = rdfint_0n[22];
  assign rd_0r0d[23] = rdfint_0n[23];
  assign rd_0r0d[24] = rdfint_0n[24];
  assign rd_0r0d[25] = rdfint_0n[25];
  assign rd_0r0d[26] = rdfint_0n[26];
  assign rd_0r0d[27] = rdfint_0n[27];
  assign rd_0r0d[28] = rdfint_0n[28];
  assign rd_0r0d[29] = rdfint_0n[29];
  assign rd_0r0d[30] = rdfint_0n[30];
  assign rd_0r0d[31] = rdfint_0n[31];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign rd_0r1d[10] = rdtint_0n[10];
  assign rd_0r1d[11] = rdtint_0n[11];
  assign rd_0r1d[12] = rdtint_0n[12];
  assign rd_0r1d[13] = rdtint_0n[13];
  assign rd_0r1d[14] = rdtint_0n[14];
  assign rd_0r1d[15] = rdtint_0n[15];
  assign rd_0r1d[16] = rdtint_0n[16];
  assign rd_0r1d[17] = rdtint_0n[17];
  assign rd_0r1d[18] = rdtint_0n[18];
  assign rd_0r1d[19] = rdtint_0n[19];
  assign rd_0r1d[20] = rdtint_0n[20];
  assign rd_0r1d[21] = rdtint_0n[21];
  assign rd_0r1d[22] = rdtint_0n[22];
  assign rd_0r1d[23] = rdtint_0n[23];
  assign rd_0r1d[24] = rdtint_0n[24];
  assign rd_0r1d[25] = rdtint_0n[25];
  assign rd_0r1d[26] = rdtint_0n[26];
  assign rd_0r1d[27] = rdtint_0n[27];
  assign rd_0r1d[28] = rdtint_0n[28];
  assign rd_0r1d[29] = rdtint_0n[29];
  assign rd_0r1d[30] = rdtint_0n[30];
  assign rd_0r1d[31] = rdtint_0n[31];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgfint_0n[32] = wg_0r0d[32];
  assign wgfint_0n[33] = wg_0r0d[33];
  assign wgfint_0n[34] = wg_0r0d[34];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign wgtint_0n[32] = wg_0r1d[32];
  assign wgtint_0n[33] = wg_0r1d[33];
  assign wgtint_0n[34] = wg_0r1d[34];
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I149 (internal_0n[0], rgrint_0n, rgrint_1n);
  NOR2 I150 (internal_0n[1], rgaint_0n, rgaint_1n);
  AND2 I151 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I152 (rdtint_1n[0], rgrint_1n, dt_0n[0]);
  AND2 I153 (rdtint_1n[1], rgrint_1n, dt_0n[1]);
  AND2 I154 (rdtint_1n[2], rgrint_1n, dt_0n[2]);
  AND2 I155 (rdtint_0n[0], rgrint_0n, dt_0n[3]);
  AND2 I156 (rdtint_0n[1], rgrint_0n, dt_0n[4]);
  AND2 I157 (rdtint_0n[2], rgrint_0n, dt_0n[5]);
  AND2 I158 (rdtint_0n[3], rgrint_0n, dt_0n[6]);
  AND2 I159 (rdtint_0n[4], rgrint_0n, dt_0n[7]);
  AND2 I160 (rdtint_0n[5], rgrint_0n, dt_0n[8]);
  AND2 I161 (rdtint_0n[6], rgrint_0n, dt_0n[9]);
  AND2 I162 (rdtint_0n[7], rgrint_0n, dt_0n[10]);
  AND2 I163 (rdtint_0n[8], rgrint_0n, dt_0n[11]);
  AND2 I164 (rdtint_0n[9], rgrint_0n, dt_0n[12]);
  AND2 I165 (rdtint_0n[10], rgrint_0n, dt_0n[13]);
  AND2 I166 (rdtint_0n[11], rgrint_0n, dt_0n[14]);
  AND2 I167 (rdtint_0n[12], rgrint_0n, dt_0n[15]);
  AND2 I168 (rdtint_0n[13], rgrint_0n, dt_0n[16]);
  AND2 I169 (rdtint_0n[14], rgrint_0n, dt_0n[17]);
  AND2 I170 (rdtint_0n[15], rgrint_0n, dt_0n[18]);
  AND2 I171 (rdtint_0n[16], rgrint_0n, dt_0n[19]);
  AND2 I172 (rdtint_0n[17], rgrint_0n, dt_0n[20]);
  AND2 I173 (rdtint_0n[18], rgrint_0n, dt_0n[21]);
  AND2 I174 (rdtint_0n[19], rgrint_0n, dt_0n[22]);
  AND2 I175 (rdtint_0n[20], rgrint_0n, dt_0n[23]);
  AND2 I176 (rdtint_0n[21], rgrint_0n, dt_0n[24]);
  AND2 I177 (rdtint_0n[22], rgrint_0n, dt_0n[25]);
  AND2 I178 (rdtint_0n[23], rgrint_0n, dt_0n[26]);
  AND2 I179 (rdtint_0n[24], rgrint_0n, dt_0n[27]);
  AND2 I180 (rdtint_0n[25], rgrint_0n, dt_0n[28]);
  AND2 I181 (rdtint_0n[26], rgrint_0n, dt_0n[29]);
  AND2 I182 (rdtint_0n[27], rgrint_0n, dt_0n[30]);
  AND2 I183 (rdtint_0n[28], rgrint_0n, dt_0n[31]);
  AND2 I184 (rdtint_0n[29], rgrint_0n, dt_0n[32]);
  AND2 I185 (rdtint_0n[30], rgrint_0n, dt_0n[33]);
  AND2 I186 (rdtint_0n[31], rgrint_0n, dt_0n[34]);
  AND2 I187 (rdfint_1n[0], rgrint_1n, df_0n[0]);
  AND2 I188 (rdfint_1n[1], rgrint_1n, df_0n[1]);
  AND2 I189 (rdfint_1n[2], rgrint_1n, df_0n[2]);
  AND2 I190 (rdfint_0n[0], rgrint_0n, df_0n[3]);
  AND2 I191 (rdfint_0n[1], rgrint_0n, df_0n[4]);
  AND2 I192 (rdfint_0n[2], rgrint_0n, df_0n[5]);
  AND2 I193 (rdfint_0n[3], rgrint_0n, df_0n[6]);
  AND2 I194 (rdfint_0n[4], rgrint_0n, df_0n[7]);
  AND2 I195 (rdfint_0n[5], rgrint_0n, df_0n[8]);
  AND2 I196 (rdfint_0n[6], rgrint_0n, df_0n[9]);
  AND2 I197 (rdfint_0n[7], rgrint_0n, df_0n[10]);
  AND2 I198 (rdfint_0n[8], rgrint_0n, df_0n[11]);
  AND2 I199 (rdfint_0n[9], rgrint_0n, df_0n[12]);
  AND2 I200 (rdfint_0n[10], rgrint_0n, df_0n[13]);
  AND2 I201 (rdfint_0n[11], rgrint_0n, df_0n[14]);
  AND2 I202 (rdfint_0n[12], rgrint_0n, df_0n[15]);
  AND2 I203 (rdfint_0n[13], rgrint_0n, df_0n[16]);
  AND2 I204 (rdfint_0n[14], rgrint_0n, df_0n[17]);
  AND2 I205 (rdfint_0n[15], rgrint_0n, df_0n[18]);
  AND2 I206 (rdfint_0n[16], rgrint_0n, df_0n[19]);
  AND2 I207 (rdfint_0n[17], rgrint_0n, df_0n[20]);
  AND2 I208 (rdfint_0n[18], rgrint_0n, df_0n[21]);
  AND2 I209 (rdfint_0n[19], rgrint_0n, df_0n[22]);
  AND2 I210 (rdfint_0n[20], rgrint_0n, df_0n[23]);
  AND2 I211 (rdfint_0n[21], rgrint_0n, df_0n[24]);
  AND2 I212 (rdfint_0n[22], rgrint_0n, df_0n[25]);
  AND2 I213 (rdfint_0n[23], rgrint_0n, df_0n[26]);
  AND2 I214 (rdfint_0n[24], rgrint_0n, df_0n[27]);
  AND2 I215 (rdfint_0n[25], rgrint_0n, df_0n[28]);
  AND2 I216 (rdfint_0n[26], rgrint_0n, df_0n[29]);
  AND2 I217 (rdfint_0n[27], rgrint_0n, df_0n[30]);
  AND2 I218 (rdfint_0n[28], rgrint_0n, df_0n[31]);
  AND2 I219 (rdfint_0n[29], rgrint_0n, df_0n[32]);
  AND2 I220 (rdfint_0n[30], rgrint_0n, df_0n[33]);
  AND2 I221 (rdfint_0n[31], rgrint_0n, df_0n[34]);
  C3 I222 (internal_0n[2], wc_0n, wacks_0n[34], wacks_0n[33]);
  C3 I223 (internal_0n[3], wacks_0n[32], wacks_0n[31], wacks_0n[30]);
  C3 I224 (internal_0n[4], wacks_0n[29], wacks_0n[28], wacks_0n[27]);
  C3 I225 (internal_0n[5], wacks_0n[26], wacks_0n[25], wacks_0n[24]);
  C3 I226 (internal_0n[6], wacks_0n[23], wacks_0n[22], wacks_0n[21]);
  C3 I227 (internal_0n[7], wacks_0n[20], wacks_0n[19], wacks_0n[18]);
  C3 I228 (internal_0n[8], wacks_0n[17], wacks_0n[16], wacks_0n[15]);
  C3 I229 (internal_0n[9], wacks_0n[14], wacks_0n[13], wacks_0n[12]);
  C3 I230 (internal_0n[10], wacks_0n[11], wacks_0n[10], wacks_0n[9]);
  C3 I231 (internal_0n[11], wacks_0n[8], wacks_0n[7], wacks_0n[6]);
  C3 I232 (internal_0n[12], wacks_0n[5], wacks_0n[4], wacks_0n[3]);
  C3 I233 (internal_0n[13], wacks_0n[2], wacks_0n[1], wacks_0n[0]);
  C3 I234 (internal_0n[14], internal_0n[2], internal_0n[3], internal_0n[4]);
  C3 I235 (internal_0n[15], internal_0n[5], internal_0n[6], internal_0n[7]);
  C3 I236 (internal_0n[16], internal_0n[8], internal_0n[9], internal_0n[10]);
  C3 I237 (internal_0n[17], internal_0n[11], internal_0n[12], internal_0n[13]);
  C2 I238 (internal_0n[18], internal_0n[14], internal_0n[15]);
  C2 I239 (internal_0n[19], internal_0n[16], internal_0n[17]);
  C2 I240 (wdrint_0n, internal_0n[18], internal_0n[19]);
  assign wen_0n[34] = wc_0n;
  assign wen_0n[33] = wc_0n;
  assign wen_0n[32] = wc_0n;
  assign wen_0n[31] = wc_0n;
  assign wen_0n[30] = wc_0n;
  assign wen_0n[29] = wc_0n;
  assign wen_0n[28] = wc_0n;
  assign wen_0n[27] = wc_0n;
  assign wen_0n[26] = wc_0n;
  assign wen_0n[25] = wc_0n;
  assign wen_0n[24] = wc_0n;
  assign wen_0n[23] = wc_0n;
  assign wen_0n[22] = wc_0n;
  assign wen_0n[21] = wc_0n;
  assign wen_0n[20] = wc_0n;
  assign wen_0n[19] = wc_0n;
  assign wen_0n[18] = wc_0n;
  assign wen_0n[17] = wc_0n;
  assign wen_0n[16] = wc_0n;
  assign wen_0n[15] = wc_0n;
  assign wen_0n[14] = wc_0n;
  assign wen_0n[13] = wc_0n;
  assign wen_0n[12] = wc_0n;
  assign wen_0n[11] = wc_0n;
  assign wen_0n[10] = wc_0n;
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[34] = git_0n[34];
  assign wt_0n[33] = git_0n[33];
  assign wt_0n[32] = git_0n[32];
  assign wt_0n[31] = git_0n[31];
  assign wt_0n[30] = git_0n[30];
  assign wt_0n[29] = git_0n[29];
  assign wt_0n[28] = git_0n[28];
  assign wt_0n[27] = git_0n[27];
  assign wt_0n[26] = git_0n[26];
  assign wt_0n[25] = git_0n[25];
  assign wt_0n[24] = git_0n[24];
  assign wt_0n[23] = git_0n[23];
  assign wt_0n[22] = git_0n[22];
  assign wt_0n[21] = git_0n[21];
  assign wt_0n[20] = git_0n[20];
  assign wt_0n[19] = git_0n[19];
  assign wt_0n[18] = git_0n[18];
  assign wt_0n[17] = git_0n[17];
  assign wt_0n[16] = git_0n[16];
  assign wt_0n[15] = git_0n[15];
  assign wt_0n[14] = git_0n[14];
  assign wt_0n[13] = git_0n[13];
  assign wt_0n[12] = git_0n[12];
  assign wt_0n[11] = git_0n[11];
  assign wt_0n[10] = git_0n[10];
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[34] = gif_0n[34];
  assign wf_0n[33] = gif_0n[33];
  assign wf_0n[32] = gif_0n[32];
  assign wf_0n[31] = gif_0n[31];
  assign wf_0n[30] = gif_0n[30];
  assign wf_0n[29] = gif_0n[29];
  assign wf_0n[28] = gif_0n[28];
  assign wf_0n[27] = gif_0n[27];
  assign wf_0n[26] = gif_0n[26];
  assign wf_0n[25] = gif_0n[25];
  assign wf_0n[24] = gif_0n[24];
  assign wf_0n[23] = gif_0n[23];
  assign wf_0n[22] = gif_0n[22];
  assign wf_0n[21] = gif_0n[21];
  assign wf_0n[20] = gif_0n[20];
  assign wf_0n[19] = gif_0n[19];
  assign wf_0n[18] = gif_0n[18];
  assign wf_0n[17] = gif_0n[17];
  assign wf_0n[16] = gif_0n[16];
  assign wf_0n[15] = gif_0n[15];
  assign wf_0n[14] = gif_0n[14];
  assign wf_0n[13] = gif_0n[13];
  assign wf_0n[12] = gif_0n[12];
  assign wf_0n[11] = gif_0n[11];
  assign wf_0n[10] = gif_0n[10];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I346 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I348 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I349 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I350 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I351 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I352 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I353 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I354 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I355 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I356 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I357 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I358 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I359 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I360 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I361 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I362 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I363 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I364 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I365 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I366 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I367 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I368 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I369 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I370 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I371 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I372 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I373 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I374 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I375 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I376 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I377 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I378 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I379 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I380 (git_0n[32], wgtint_0n[32], ig_0n);
  AND2 I381 (git_0n[33], wgtint_0n[33], ig_0n);
  AND2 I382 (git_0n[34], wgtint_0n[34], ig_0n);
  AND2 I383 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I384 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I385 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I386 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I387 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I388 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I389 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I390 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I391 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I392 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I393 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I394 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I395 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I396 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I397 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I398 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I399 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I400 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I401 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I402 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I403 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I404 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I405 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I406 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I407 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I408 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I409 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I410 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I411 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I412 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I413 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I414 (gif_0n[31], wgfint_0n[31], ig_0n);
  AND2 I415 (gif_0n[32], wgfint_0n[32], ig_0n);
  AND2 I416 (gif_0n[33], wgfint_0n[33], ig_0n);
  AND2 I417 (gif_0n[34], wgfint_0n[34], ig_0n);
  C3 I418 (internal_0n[20], complete1543_0n[0], complete1543_0n[1], complete1543_0n[2]);
  C3 I419 (internal_0n[21], complete1543_0n[3], complete1543_0n[4], complete1543_0n[5]);
  C3 I420 (internal_0n[22], complete1543_0n[6], complete1543_0n[7], complete1543_0n[8]);
  C3 I421 (internal_0n[23], complete1543_0n[9], complete1543_0n[10], complete1543_0n[11]);
  C3 I422 (internal_0n[24], complete1543_0n[12], complete1543_0n[13], complete1543_0n[14]);
  C3 I423 (internal_0n[25], complete1543_0n[15], complete1543_0n[16], complete1543_0n[17]);
  C3 I424 (internal_0n[26], complete1543_0n[18], complete1543_0n[19], complete1543_0n[20]);
  C3 I425 (internal_0n[27], complete1543_0n[21], complete1543_0n[22], complete1543_0n[23]);
  C3 I426 (internal_0n[28], complete1543_0n[24], complete1543_0n[25], complete1543_0n[26]);
  C3 I427 (internal_0n[29], complete1543_0n[27], complete1543_0n[28], complete1543_0n[29]);
  C3 I428 (internal_0n[30], complete1543_0n[30], complete1543_0n[31], complete1543_0n[32]);
  C2 I429 (internal_0n[31], complete1543_0n[33], complete1543_0n[34]);
  C3 I430 (internal_0n[32], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I431 (internal_0n[33], internal_0n[23], internal_0n[24], internal_0n[25]);
  C3 I432 (internal_0n[34], internal_0n[26], internal_0n[27], internal_0n[28]);
  C3 I433 (internal_0n[35], internal_0n[29], internal_0n[30], internal_0n[31]);
  C2 I434 (internal_0n[36], internal_0n[32], internal_0n[33]);
  C2 I435 (internal_0n[37], internal_0n[34], internal_0n[35]);
  C2 I436 (wc_0n, internal_0n[36], internal_0n[37]);
  OR2 I437 (complete1543_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I438 (complete1543_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I439 (complete1543_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I440 (complete1543_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I441 (complete1543_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I442 (complete1543_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I443 (complete1543_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I444 (complete1543_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I445 (complete1543_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I446 (complete1543_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I447 (complete1543_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I448 (complete1543_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I449 (complete1543_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I450 (complete1543_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I451 (complete1543_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I452 (complete1543_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I453 (complete1543_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I454 (complete1543_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I455 (complete1543_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I456 (complete1543_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I457 (complete1543_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I458 (complete1543_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I459 (complete1543_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I460 (complete1543_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I461 (complete1543_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I462 (complete1543_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I463 (complete1543_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I464 (complete1543_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I465 (complete1543_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I466 (complete1543_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I467 (complete1543_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I468 (complete1543_0n[31], wgfint_0n[31], wgtint_0n[31]);
  OR2 I469 (complete1543_0n[32], wgfint_0n[32], wgtint_0n[32]);
  OR2 I470 (complete1543_0n[33], wgfint_0n[33], wgtint_0n[33]);
  OR2 I471 (complete1543_0n[34], wgfint_0n[34], wgtint_0n[34]);
  AO22 I472 (wacks_0n[34], gf1541_0n[34], df_0n[34], gt1542_0n[34], dt_0n[34]);
  NOR2 I473 (dt_0n[34], df_0n[34], gf1541_0n[34]);
  NOR3 I474 (df_0n[34], dt_0n[34], gt1542_0n[34], init_0n);
  AND2 I475 (gt1542_0n[34], wt_0n[34], wen_0n[34]);
  AND2 I476 (gf1541_0n[34], wf_0n[34], wen_0n[34]);
  AO22 I477 (wacks_0n[33], gf1541_0n[33], df_0n[33], gt1542_0n[33], dt_0n[33]);
  NOR2 I478 (dt_0n[33], df_0n[33], gf1541_0n[33]);
  NOR3 I479 (df_0n[33], dt_0n[33], gt1542_0n[33], init_0n);
  AND2 I480 (gt1542_0n[33], wt_0n[33], wen_0n[33]);
  AND2 I481 (gf1541_0n[33], wf_0n[33], wen_0n[33]);
  AO22 I482 (wacks_0n[32], gf1541_0n[32], df_0n[32], gt1542_0n[32], dt_0n[32]);
  NOR2 I483 (dt_0n[32], df_0n[32], gf1541_0n[32]);
  NOR3 I484 (df_0n[32], dt_0n[32], gt1542_0n[32], init_0n);
  AND2 I485 (gt1542_0n[32], wt_0n[32], wen_0n[32]);
  AND2 I486 (gf1541_0n[32], wf_0n[32], wen_0n[32]);
  AO22 I487 (wacks_0n[31], gf1541_0n[31], df_0n[31], gt1542_0n[31], dt_0n[31]);
  NOR2 I488 (dt_0n[31], df_0n[31], gf1541_0n[31]);
  NOR3 I489 (df_0n[31], dt_0n[31], gt1542_0n[31], init_0n);
  AND2 I490 (gt1542_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I491 (gf1541_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I492 (wacks_0n[30], gf1541_0n[30], df_0n[30], gt1542_0n[30], dt_0n[30]);
  NOR2 I493 (dt_0n[30], df_0n[30], gf1541_0n[30]);
  NOR3 I494 (df_0n[30], dt_0n[30], gt1542_0n[30], init_0n);
  AND2 I495 (gt1542_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I496 (gf1541_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I497 (wacks_0n[29], gf1541_0n[29], df_0n[29], gt1542_0n[29], dt_0n[29]);
  NOR2 I498 (dt_0n[29], df_0n[29], gf1541_0n[29]);
  NOR3 I499 (df_0n[29], dt_0n[29], gt1542_0n[29], init_0n);
  AND2 I500 (gt1542_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I501 (gf1541_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I502 (wacks_0n[28], gf1541_0n[28], df_0n[28], gt1542_0n[28], dt_0n[28]);
  NOR2 I503 (dt_0n[28], df_0n[28], gf1541_0n[28]);
  NOR3 I504 (df_0n[28], dt_0n[28], gt1542_0n[28], init_0n);
  AND2 I505 (gt1542_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I506 (gf1541_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I507 (wacks_0n[27], gf1541_0n[27], df_0n[27], gt1542_0n[27], dt_0n[27]);
  NOR2 I508 (dt_0n[27], df_0n[27], gf1541_0n[27]);
  NOR3 I509 (df_0n[27], dt_0n[27], gt1542_0n[27], init_0n);
  AND2 I510 (gt1542_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I511 (gf1541_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I512 (wacks_0n[26], gf1541_0n[26], df_0n[26], gt1542_0n[26], dt_0n[26]);
  NOR2 I513 (dt_0n[26], df_0n[26], gf1541_0n[26]);
  NOR3 I514 (df_0n[26], dt_0n[26], gt1542_0n[26], init_0n);
  AND2 I515 (gt1542_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I516 (gf1541_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I517 (wacks_0n[25], gf1541_0n[25], df_0n[25], gt1542_0n[25], dt_0n[25]);
  NOR2 I518 (dt_0n[25], df_0n[25], gf1541_0n[25]);
  NOR3 I519 (df_0n[25], dt_0n[25], gt1542_0n[25], init_0n);
  AND2 I520 (gt1542_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I521 (gf1541_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I522 (wacks_0n[24], gf1541_0n[24], df_0n[24], gt1542_0n[24], dt_0n[24]);
  NOR2 I523 (dt_0n[24], df_0n[24], gf1541_0n[24]);
  NOR3 I524 (df_0n[24], dt_0n[24], gt1542_0n[24], init_0n);
  AND2 I525 (gt1542_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I526 (gf1541_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I527 (wacks_0n[23], gf1541_0n[23], df_0n[23], gt1542_0n[23], dt_0n[23]);
  NOR2 I528 (dt_0n[23], df_0n[23], gf1541_0n[23]);
  NOR3 I529 (df_0n[23], dt_0n[23], gt1542_0n[23], init_0n);
  AND2 I530 (gt1542_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I531 (gf1541_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I532 (wacks_0n[22], gf1541_0n[22], df_0n[22], gt1542_0n[22], dt_0n[22]);
  NOR2 I533 (dt_0n[22], df_0n[22], gf1541_0n[22]);
  NOR3 I534 (df_0n[22], dt_0n[22], gt1542_0n[22], init_0n);
  AND2 I535 (gt1542_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I536 (gf1541_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I537 (wacks_0n[21], gf1541_0n[21], df_0n[21], gt1542_0n[21], dt_0n[21]);
  NOR2 I538 (dt_0n[21], df_0n[21], gf1541_0n[21]);
  NOR3 I539 (df_0n[21], dt_0n[21], gt1542_0n[21], init_0n);
  AND2 I540 (gt1542_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I541 (gf1541_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I542 (wacks_0n[20], gf1541_0n[20], df_0n[20], gt1542_0n[20], dt_0n[20]);
  NOR2 I543 (dt_0n[20], df_0n[20], gf1541_0n[20]);
  NOR3 I544 (df_0n[20], dt_0n[20], gt1542_0n[20], init_0n);
  AND2 I545 (gt1542_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I546 (gf1541_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I547 (wacks_0n[19], gf1541_0n[19], df_0n[19], gt1542_0n[19], dt_0n[19]);
  NOR2 I548 (dt_0n[19], df_0n[19], gf1541_0n[19]);
  NOR3 I549 (df_0n[19], dt_0n[19], gt1542_0n[19], init_0n);
  AND2 I550 (gt1542_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I551 (gf1541_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I552 (wacks_0n[18], gf1541_0n[18], df_0n[18], gt1542_0n[18], dt_0n[18]);
  NOR2 I553 (dt_0n[18], df_0n[18], gf1541_0n[18]);
  NOR3 I554 (df_0n[18], dt_0n[18], gt1542_0n[18], init_0n);
  AND2 I555 (gt1542_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I556 (gf1541_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I557 (wacks_0n[17], gf1541_0n[17], df_0n[17], gt1542_0n[17], dt_0n[17]);
  NOR2 I558 (dt_0n[17], df_0n[17], gf1541_0n[17]);
  NOR3 I559 (df_0n[17], dt_0n[17], gt1542_0n[17], init_0n);
  AND2 I560 (gt1542_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I561 (gf1541_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I562 (wacks_0n[16], gf1541_0n[16], df_0n[16], gt1542_0n[16], dt_0n[16]);
  NOR2 I563 (dt_0n[16], df_0n[16], gf1541_0n[16]);
  NOR3 I564 (df_0n[16], dt_0n[16], gt1542_0n[16], init_0n);
  AND2 I565 (gt1542_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I566 (gf1541_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I567 (wacks_0n[15], gf1541_0n[15], df_0n[15], gt1542_0n[15], dt_0n[15]);
  NOR2 I568 (dt_0n[15], df_0n[15], gf1541_0n[15]);
  NOR3 I569 (df_0n[15], dt_0n[15], gt1542_0n[15], init_0n);
  AND2 I570 (gt1542_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I571 (gf1541_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I572 (wacks_0n[14], gf1541_0n[14], df_0n[14], gt1542_0n[14], dt_0n[14]);
  NOR2 I573 (dt_0n[14], df_0n[14], gf1541_0n[14]);
  NOR3 I574 (df_0n[14], dt_0n[14], gt1542_0n[14], init_0n);
  AND2 I575 (gt1542_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I576 (gf1541_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I577 (wacks_0n[13], gf1541_0n[13], df_0n[13], gt1542_0n[13], dt_0n[13]);
  NOR2 I578 (dt_0n[13], df_0n[13], gf1541_0n[13]);
  NOR3 I579 (df_0n[13], dt_0n[13], gt1542_0n[13], init_0n);
  AND2 I580 (gt1542_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I581 (gf1541_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I582 (wacks_0n[12], gf1541_0n[12], df_0n[12], gt1542_0n[12], dt_0n[12]);
  NOR2 I583 (dt_0n[12], df_0n[12], gf1541_0n[12]);
  NOR3 I584 (df_0n[12], dt_0n[12], gt1542_0n[12], init_0n);
  AND2 I585 (gt1542_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I586 (gf1541_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I587 (wacks_0n[11], gf1541_0n[11], df_0n[11], gt1542_0n[11], dt_0n[11]);
  NOR2 I588 (dt_0n[11], df_0n[11], gf1541_0n[11]);
  NOR3 I589 (df_0n[11], dt_0n[11], gt1542_0n[11], init_0n);
  AND2 I590 (gt1542_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I591 (gf1541_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I592 (wacks_0n[10], gf1541_0n[10], df_0n[10], gt1542_0n[10], dt_0n[10]);
  NOR2 I593 (dt_0n[10], df_0n[10], gf1541_0n[10]);
  NOR3 I594 (df_0n[10], dt_0n[10], gt1542_0n[10], init_0n);
  AND2 I595 (gt1542_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I596 (gf1541_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I597 (wacks_0n[9], gf1541_0n[9], df_0n[9], gt1542_0n[9], dt_0n[9]);
  NOR2 I598 (dt_0n[9], df_0n[9], gf1541_0n[9]);
  NOR3 I599 (df_0n[9], dt_0n[9], gt1542_0n[9], init_0n);
  AND2 I600 (gt1542_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I601 (gf1541_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I602 (wacks_0n[8], gf1541_0n[8], df_0n[8], gt1542_0n[8], dt_0n[8]);
  NOR2 I603 (dt_0n[8], df_0n[8], gf1541_0n[8]);
  NOR3 I604 (df_0n[8], dt_0n[8], gt1542_0n[8], init_0n);
  AND2 I605 (gt1542_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I606 (gf1541_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I607 (wacks_0n[7], gf1541_0n[7], df_0n[7], gt1542_0n[7], dt_0n[7]);
  NOR2 I608 (dt_0n[7], df_0n[7], gf1541_0n[7]);
  NOR3 I609 (df_0n[7], dt_0n[7], gt1542_0n[7], init_0n);
  AND2 I610 (gt1542_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I611 (gf1541_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I612 (wacks_0n[6], gf1541_0n[6], df_0n[6], gt1542_0n[6], dt_0n[6]);
  NOR2 I613 (dt_0n[6], df_0n[6], gf1541_0n[6]);
  NOR3 I614 (df_0n[6], dt_0n[6], gt1542_0n[6], init_0n);
  AND2 I615 (gt1542_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I616 (gf1541_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I617 (wacks_0n[5], gf1541_0n[5], df_0n[5], gt1542_0n[5], dt_0n[5]);
  NOR2 I618 (dt_0n[5], df_0n[5], gf1541_0n[5]);
  NOR3 I619 (df_0n[5], dt_0n[5], gt1542_0n[5], init_0n);
  AND2 I620 (gt1542_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I621 (gf1541_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I622 (wacks_0n[4], gf1541_0n[4], df_0n[4], gt1542_0n[4], dt_0n[4]);
  NOR2 I623 (dt_0n[4], df_0n[4], gf1541_0n[4]);
  NOR3 I624 (df_0n[4], dt_0n[4], gt1542_0n[4], init_0n);
  AND2 I625 (gt1542_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I626 (gf1541_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I627 (wacks_0n[3], gf1541_0n[3], df_0n[3], gt1542_0n[3], dt_0n[3]);
  NOR2 I628 (dt_0n[3], df_0n[3], gf1541_0n[3]);
  NOR3 I629 (df_0n[3], dt_0n[3], gt1542_0n[3], init_0n);
  AND2 I630 (gt1542_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I631 (gf1541_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I632 (wacks_0n[2], gf1541_0n[2], df_0n[2], gt1542_0n[2], dt_0n[2]);
  NOR2 I633 (dt_0n[2], df_0n[2], gf1541_0n[2]);
  NOR3 I634 (df_0n[2], dt_0n[2], gt1542_0n[2], init_0n);
  AND2 I635 (gt1542_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I636 (gf1541_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I637 (wacks_0n[1], gf1541_0n[1], df_0n[1], gt1542_0n[1], dt_0n[1]);
  NOR2 I638 (dt_0n[1], df_0n[1], gf1541_0n[1]);
  NOR3 I639 (df_0n[1], dt_0n[1], gt1542_0n[1], init_0n);
  AND2 I640 (gt1542_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I641 (gf1541_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I642 (wacks_0n[0], gf1541_0n[0], df_0n[0], gt1542_0n[0], dt_0n[0]);
  NOR2 I643 (dt_0n[0], df_0n[0], gf1541_0n[0]);
  NOR3 I644 (df_0n[0], dt_0n[0], gt1542_0n[0], init_0n);
  AND2 I645 (gt1542_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I646 (gf1541_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I647 (init_0n, initialise);
endmodule

module BrzV_35_l6__28_29_l45__28_28_280_2035_29_2_m94m (
  wg_0r0d, wg_0r1d, wg_0a,
  wg_1r0d, wg_1r1d, wg_1a,
  wd_0r, wd_0a,
  wd_1r, wd_1a,
  rg_0r, rg_0a,
  rd_0r0d, rd_0r1d, rd_0a,
  initialise
);
  input [34:0] wg_0r0d;
  input [34:0] wg_0r1d;
  output wg_0a;
  input [34:0] wg_1r0d;
  input [34:0] wg_1r1d;
  output wg_1a;
  output wd_0r;
  input wd_0a;
  output wd_1r;
  input wd_1a;
  input rg_0r;
  output rg_0a;
  output [34:0] rd_0r0d;
  output [34:0] rd_0r1d;
  input rd_0a;
  input initialise;
  wire [71:0] internal_0n;
  wire [34:0] wf_0n;
  wire [34:0] wt_0n;
  wire [34:0] df_0n;
  wire [34:0] dt_0n;
  wire rgrint_0n;
  wire wc_0n;
  wire wc_1n;
  wire [34:0] wacks_0n;
  wire wdrint_0n;
  wire wdrint_1n;
  wire wgaint_0n;
  wire wgaint_1n;
  wire [34:0] wgfint_0n;
  wire [34:0] wgfint_1n;
  wire [34:0] wgtint_0n;
  wire [34:0] wgtint_1n;
  wire rgaint_0n;
  wire [34:0] rdfint_0n;
  wire [34:0] rdtint_0n;
  wire [34:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire igc_1n;
  wire ig_0n;
  wire ig_1n;
  wire [34:0] gif_0n;
  wire [34:0] gif_1n;
  wire [34:0] git_0n;
  wire [34:0] git_1n;
  wire [34:0] complete1559_0n;
  wire [34:0] complete1558_0n;
  wire [34:0] gt1557_0n;
  wire [34:0] gf1556_0n;
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r0d[10] = rdfint_0n[10];
  assign rd_0r0d[11] = rdfint_0n[11];
  assign rd_0r0d[12] = rdfint_0n[12];
  assign rd_0r0d[13] = rdfint_0n[13];
  assign rd_0r0d[14] = rdfint_0n[14];
  assign rd_0r0d[15] = rdfint_0n[15];
  assign rd_0r0d[16] = rdfint_0n[16];
  assign rd_0r0d[17] = rdfint_0n[17];
  assign rd_0r0d[18] = rdfint_0n[18];
  assign rd_0r0d[19] = rdfint_0n[19];
  assign rd_0r0d[20] = rdfint_0n[20];
  assign rd_0r0d[21] = rdfint_0n[21];
  assign rd_0r0d[22] = rdfint_0n[22];
  assign rd_0r0d[23] = rdfint_0n[23];
  assign rd_0r0d[24] = rdfint_0n[24];
  assign rd_0r0d[25] = rdfint_0n[25];
  assign rd_0r0d[26] = rdfint_0n[26];
  assign rd_0r0d[27] = rdfint_0n[27];
  assign rd_0r0d[28] = rdfint_0n[28];
  assign rd_0r0d[29] = rdfint_0n[29];
  assign rd_0r0d[30] = rdfint_0n[30];
  assign rd_0r0d[31] = rdfint_0n[31];
  assign rd_0r0d[32] = rdfint_0n[32];
  assign rd_0r0d[33] = rdfint_0n[33];
  assign rd_0r0d[34] = rdfint_0n[34];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign rd_0r1d[10] = rdtint_0n[10];
  assign rd_0r1d[11] = rdtint_0n[11];
  assign rd_0r1d[12] = rdtint_0n[12];
  assign rd_0r1d[13] = rdtint_0n[13];
  assign rd_0r1d[14] = rdtint_0n[14];
  assign rd_0r1d[15] = rdtint_0n[15];
  assign rd_0r1d[16] = rdtint_0n[16];
  assign rd_0r1d[17] = rdtint_0n[17];
  assign rd_0r1d[18] = rdtint_0n[18];
  assign rd_0r1d[19] = rdtint_0n[19];
  assign rd_0r1d[20] = rdtint_0n[20];
  assign rd_0r1d[21] = rdtint_0n[21];
  assign rd_0r1d[22] = rdtint_0n[22];
  assign rd_0r1d[23] = rdtint_0n[23];
  assign rd_0r1d[24] = rdtint_0n[24];
  assign rd_0r1d[25] = rdtint_0n[25];
  assign rd_0r1d[26] = rdtint_0n[26];
  assign rd_0r1d[27] = rdtint_0n[27];
  assign rd_0r1d[28] = rdtint_0n[28];
  assign rd_0r1d[29] = rdtint_0n[29];
  assign rd_0r1d[30] = rdtint_0n[30];
  assign rd_0r1d[31] = rdtint_0n[31];
  assign rd_0r1d[32] = rdtint_0n[32];
  assign rd_0r1d[33] = rdtint_0n[33];
  assign rd_0r1d[34] = rdtint_0n[34];
  assign wg_1a = wgaint_1n;
  assign wgfint_1n[0] = wg_1r0d[0];
  assign wgfint_1n[1] = wg_1r0d[1];
  assign wgfint_1n[2] = wg_1r0d[2];
  assign wgfint_1n[3] = wg_1r0d[3];
  assign wgfint_1n[4] = wg_1r0d[4];
  assign wgfint_1n[5] = wg_1r0d[5];
  assign wgfint_1n[6] = wg_1r0d[6];
  assign wgfint_1n[7] = wg_1r0d[7];
  assign wgfint_1n[8] = wg_1r0d[8];
  assign wgfint_1n[9] = wg_1r0d[9];
  assign wgfint_1n[10] = wg_1r0d[10];
  assign wgfint_1n[11] = wg_1r0d[11];
  assign wgfint_1n[12] = wg_1r0d[12];
  assign wgfint_1n[13] = wg_1r0d[13];
  assign wgfint_1n[14] = wg_1r0d[14];
  assign wgfint_1n[15] = wg_1r0d[15];
  assign wgfint_1n[16] = wg_1r0d[16];
  assign wgfint_1n[17] = wg_1r0d[17];
  assign wgfint_1n[18] = wg_1r0d[18];
  assign wgfint_1n[19] = wg_1r0d[19];
  assign wgfint_1n[20] = wg_1r0d[20];
  assign wgfint_1n[21] = wg_1r0d[21];
  assign wgfint_1n[22] = wg_1r0d[22];
  assign wgfint_1n[23] = wg_1r0d[23];
  assign wgfint_1n[24] = wg_1r0d[24];
  assign wgfint_1n[25] = wg_1r0d[25];
  assign wgfint_1n[26] = wg_1r0d[26];
  assign wgfint_1n[27] = wg_1r0d[27];
  assign wgfint_1n[28] = wg_1r0d[28];
  assign wgfint_1n[29] = wg_1r0d[29];
  assign wgfint_1n[30] = wg_1r0d[30];
  assign wgfint_1n[31] = wg_1r0d[31];
  assign wgfint_1n[32] = wg_1r0d[32];
  assign wgfint_1n[33] = wg_1r0d[33];
  assign wgfint_1n[34] = wg_1r0d[34];
  assign wgtint_1n[0] = wg_1r1d[0];
  assign wgtint_1n[1] = wg_1r1d[1];
  assign wgtint_1n[2] = wg_1r1d[2];
  assign wgtint_1n[3] = wg_1r1d[3];
  assign wgtint_1n[4] = wg_1r1d[4];
  assign wgtint_1n[5] = wg_1r1d[5];
  assign wgtint_1n[6] = wg_1r1d[6];
  assign wgtint_1n[7] = wg_1r1d[7];
  assign wgtint_1n[8] = wg_1r1d[8];
  assign wgtint_1n[9] = wg_1r1d[9];
  assign wgtint_1n[10] = wg_1r1d[10];
  assign wgtint_1n[11] = wg_1r1d[11];
  assign wgtint_1n[12] = wg_1r1d[12];
  assign wgtint_1n[13] = wg_1r1d[13];
  assign wgtint_1n[14] = wg_1r1d[14];
  assign wgtint_1n[15] = wg_1r1d[15];
  assign wgtint_1n[16] = wg_1r1d[16];
  assign wgtint_1n[17] = wg_1r1d[17];
  assign wgtint_1n[18] = wg_1r1d[18];
  assign wgtint_1n[19] = wg_1r1d[19];
  assign wgtint_1n[20] = wg_1r1d[20];
  assign wgtint_1n[21] = wg_1r1d[21];
  assign wgtint_1n[22] = wg_1r1d[22];
  assign wgtint_1n[23] = wg_1r1d[23];
  assign wgtint_1n[24] = wg_1r1d[24];
  assign wgtint_1n[25] = wg_1r1d[25];
  assign wgtint_1n[26] = wg_1r1d[26];
  assign wgtint_1n[27] = wg_1r1d[27];
  assign wgtint_1n[28] = wg_1r1d[28];
  assign wgtint_1n[29] = wg_1r1d[29];
  assign wgtint_1n[30] = wg_1r1d[30];
  assign wgtint_1n[31] = wg_1r1d[31];
  assign wgtint_1n[32] = wg_1r1d[32];
  assign wgtint_1n[33] = wg_1r1d[33];
  assign wgtint_1n[34] = wg_1r1d[34];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgfint_0n[32] = wg_0r0d[32];
  assign wgfint_0n[33] = wg_0r0d[33];
  assign wgfint_0n[34] = wg_0r0d[34];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign wgtint_0n[32] = wg_0r1d[32];
  assign wgtint_0n[33] = wg_0r1d[33];
  assign wgtint_0n[34] = wg_0r1d[34];
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_1n = wd_1a;
  assign wd_1r = wdrint_1n;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I219 (nanyread_0n, rgrint_0n, rgaint_0n);
  AND2 I220 (rdtint_0n[0], rgrint_0n, dt_0n[0]);
  AND2 I221 (rdtint_0n[1], rgrint_0n, dt_0n[1]);
  AND2 I222 (rdtint_0n[2], rgrint_0n, dt_0n[2]);
  AND2 I223 (rdtint_0n[3], rgrint_0n, dt_0n[3]);
  AND2 I224 (rdtint_0n[4], rgrint_0n, dt_0n[4]);
  AND2 I225 (rdtint_0n[5], rgrint_0n, dt_0n[5]);
  AND2 I226 (rdtint_0n[6], rgrint_0n, dt_0n[6]);
  AND2 I227 (rdtint_0n[7], rgrint_0n, dt_0n[7]);
  AND2 I228 (rdtint_0n[8], rgrint_0n, dt_0n[8]);
  AND2 I229 (rdtint_0n[9], rgrint_0n, dt_0n[9]);
  AND2 I230 (rdtint_0n[10], rgrint_0n, dt_0n[10]);
  AND2 I231 (rdtint_0n[11], rgrint_0n, dt_0n[11]);
  AND2 I232 (rdtint_0n[12], rgrint_0n, dt_0n[12]);
  AND2 I233 (rdtint_0n[13], rgrint_0n, dt_0n[13]);
  AND2 I234 (rdtint_0n[14], rgrint_0n, dt_0n[14]);
  AND2 I235 (rdtint_0n[15], rgrint_0n, dt_0n[15]);
  AND2 I236 (rdtint_0n[16], rgrint_0n, dt_0n[16]);
  AND2 I237 (rdtint_0n[17], rgrint_0n, dt_0n[17]);
  AND2 I238 (rdtint_0n[18], rgrint_0n, dt_0n[18]);
  AND2 I239 (rdtint_0n[19], rgrint_0n, dt_0n[19]);
  AND2 I240 (rdtint_0n[20], rgrint_0n, dt_0n[20]);
  AND2 I241 (rdtint_0n[21], rgrint_0n, dt_0n[21]);
  AND2 I242 (rdtint_0n[22], rgrint_0n, dt_0n[22]);
  AND2 I243 (rdtint_0n[23], rgrint_0n, dt_0n[23]);
  AND2 I244 (rdtint_0n[24], rgrint_0n, dt_0n[24]);
  AND2 I245 (rdtint_0n[25], rgrint_0n, dt_0n[25]);
  AND2 I246 (rdtint_0n[26], rgrint_0n, dt_0n[26]);
  AND2 I247 (rdtint_0n[27], rgrint_0n, dt_0n[27]);
  AND2 I248 (rdtint_0n[28], rgrint_0n, dt_0n[28]);
  AND2 I249 (rdtint_0n[29], rgrint_0n, dt_0n[29]);
  AND2 I250 (rdtint_0n[30], rgrint_0n, dt_0n[30]);
  AND2 I251 (rdtint_0n[31], rgrint_0n, dt_0n[31]);
  AND2 I252 (rdtint_0n[32], rgrint_0n, dt_0n[32]);
  AND2 I253 (rdtint_0n[33], rgrint_0n, dt_0n[33]);
  AND2 I254 (rdtint_0n[34], rgrint_0n, dt_0n[34]);
  AND2 I255 (rdfint_0n[0], rgrint_0n, df_0n[0]);
  AND2 I256 (rdfint_0n[1], rgrint_0n, df_0n[1]);
  AND2 I257 (rdfint_0n[2], rgrint_0n, df_0n[2]);
  AND2 I258 (rdfint_0n[3], rgrint_0n, df_0n[3]);
  AND2 I259 (rdfint_0n[4], rgrint_0n, df_0n[4]);
  AND2 I260 (rdfint_0n[5], rgrint_0n, df_0n[5]);
  AND2 I261 (rdfint_0n[6], rgrint_0n, df_0n[6]);
  AND2 I262 (rdfint_0n[7], rgrint_0n, df_0n[7]);
  AND2 I263 (rdfint_0n[8], rgrint_0n, df_0n[8]);
  AND2 I264 (rdfint_0n[9], rgrint_0n, df_0n[9]);
  AND2 I265 (rdfint_0n[10], rgrint_0n, df_0n[10]);
  AND2 I266 (rdfint_0n[11], rgrint_0n, df_0n[11]);
  AND2 I267 (rdfint_0n[12], rgrint_0n, df_0n[12]);
  AND2 I268 (rdfint_0n[13], rgrint_0n, df_0n[13]);
  AND2 I269 (rdfint_0n[14], rgrint_0n, df_0n[14]);
  AND2 I270 (rdfint_0n[15], rgrint_0n, df_0n[15]);
  AND2 I271 (rdfint_0n[16], rgrint_0n, df_0n[16]);
  AND2 I272 (rdfint_0n[17], rgrint_0n, df_0n[17]);
  AND2 I273 (rdfint_0n[18], rgrint_0n, df_0n[18]);
  AND2 I274 (rdfint_0n[19], rgrint_0n, df_0n[19]);
  AND2 I275 (rdfint_0n[20], rgrint_0n, df_0n[20]);
  AND2 I276 (rdfint_0n[21], rgrint_0n, df_0n[21]);
  AND2 I277 (rdfint_0n[22], rgrint_0n, df_0n[22]);
  AND2 I278 (rdfint_0n[23], rgrint_0n, df_0n[23]);
  AND2 I279 (rdfint_0n[24], rgrint_0n, df_0n[24]);
  AND2 I280 (rdfint_0n[25], rgrint_0n, df_0n[25]);
  AND2 I281 (rdfint_0n[26], rgrint_0n, df_0n[26]);
  AND2 I282 (rdfint_0n[27], rgrint_0n, df_0n[27]);
  AND2 I283 (rdfint_0n[28], rgrint_0n, df_0n[28]);
  AND2 I284 (rdfint_0n[29], rgrint_0n, df_0n[29]);
  AND2 I285 (rdfint_0n[30], rgrint_0n, df_0n[30]);
  AND2 I286 (rdfint_0n[31], rgrint_0n, df_0n[31]);
  AND2 I287 (rdfint_0n[32], rgrint_0n, df_0n[32]);
  AND2 I288 (rdfint_0n[33], rgrint_0n, df_0n[33]);
  AND2 I289 (rdfint_0n[34], rgrint_0n, df_0n[34]);
  C3 I290 (internal_0n[0], wc_1n, wacks_0n[34], wacks_0n[33]);
  C3 I291 (internal_0n[1], wacks_0n[32], wacks_0n[31], wacks_0n[30]);
  C3 I292 (internal_0n[2], wacks_0n[29], wacks_0n[28], wacks_0n[27]);
  C3 I293 (internal_0n[3], wacks_0n[26], wacks_0n[25], wacks_0n[24]);
  C3 I294 (internal_0n[4], wacks_0n[23], wacks_0n[22], wacks_0n[21]);
  C3 I295 (internal_0n[5], wacks_0n[20], wacks_0n[19], wacks_0n[18]);
  C3 I296 (internal_0n[6], wacks_0n[17], wacks_0n[16], wacks_0n[15]);
  C3 I297 (internal_0n[7], wacks_0n[14], wacks_0n[13], wacks_0n[12]);
  C3 I298 (internal_0n[8], wacks_0n[11], wacks_0n[10], wacks_0n[9]);
  C3 I299 (internal_0n[9], wacks_0n[8], wacks_0n[7], wacks_0n[6]);
  C3 I300 (internal_0n[10], wacks_0n[5], wacks_0n[4], wacks_0n[3]);
  C3 I301 (internal_0n[11], wacks_0n[2], wacks_0n[1], wacks_0n[0]);
  C3 I302 (internal_0n[12], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I303 (internal_0n[13], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I304 (internal_0n[14], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I305 (internal_0n[15], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I306 (internal_0n[16], internal_0n[12], internal_0n[13]);
  C2 I307 (internal_0n[17], internal_0n[14], internal_0n[15]);
  C2 I308 (wdrint_1n, internal_0n[16], internal_0n[17]);
  C3 I309 (internal_0n[18], wc_0n, wacks_0n[34], wacks_0n[33]);
  C3 I310 (internal_0n[19], wacks_0n[32], wacks_0n[31], wacks_0n[30]);
  C3 I311 (internal_0n[20], wacks_0n[29], wacks_0n[28], wacks_0n[27]);
  C3 I312 (internal_0n[21], wacks_0n[26], wacks_0n[25], wacks_0n[24]);
  C3 I313 (internal_0n[22], wacks_0n[23], wacks_0n[22], wacks_0n[21]);
  C3 I314 (internal_0n[23], wacks_0n[20], wacks_0n[19], wacks_0n[18]);
  C3 I315 (internal_0n[24], wacks_0n[17], wacks_0n[16], wacks_0n[15]);
  C3 I316 (internal_0n[25], wacks_0n[14], wacks_0n[13], wacks_0n[12]);
  C3 I317 (internal_0n[26], wacks_0n[11], wacks_0n[10], wacks_0n[9]);
  C3 I318 (internal_0n[27], wacks_0n[8], wacks_0n[7], wacks_0n[6]);
  C3 I319 (internal_0n[28], wacks_0n[5], wacks_0n[4], wacks_0n[3]);
  C3 I320 (internal_0n[29], wacks_0n[2], wacks_0n[1], wacks_0n[0]);
  C3 I321 (internal_0n[30], internal_0n[18], internal_0n[19], internal_0n[20]);
  C3 I322 (internal_0n[31], internal_0n[21], internal_0n[22], internal_0n[23]);
  C3 I323 (internal_0n[32], internal_0n[24], internal_0n[25], internal_0n[26]);
  C3 I324 (internal_0n[33], internal_0n[27], internal_0n[28], internal_0n[29]);
  C2 I325 (internal_0n[34], internal_0n[30], internal_0n[31]);
  C2 I326 (internal_0n[35], internal_0n[32], internal_0n[33]);
  C2 I327 (wdrint_0n, internal_0n[34], internal_0n[35]);
  OR2 I328 (wen_0n[34], wc_1n, wc_0n);
  OR2 I329 (wen_0n[33], wc_1n, wc_0n);
  OR2 I330 (wen_0n[32], wc_1n, wc_0n);
  OR2 I331 (wen_0n[31], wc_1n, wc_0n);
  OR2 I332 (wen_0n[30], wc_1n, wc_0n);
  OR2 I333 (wen_0n[29], wc_1n, wc_0n);
  OR2 I334 (wen_0n[28], wc_1n, wc_0n);
  OR2 I335 (wen_0n[27], wc_1n, wc_0n);
  OR2 I336 (wen_0n[26], wc_1n, wc_0n);
  OR2 I337 (wen_0n[25], wc_1n, wc_0n);
  OR2 I338 (wen_0n[24], wc_1n, wc_0n);
  OR2 I339 (wen_0n[23], wc_1n, wc_0n);
  OR2 I340 (wen_0n[22], wc_1n, wc_0n);
  OR2 I341 (wen_0n[21], wc_1n, wc_0n);
  OR2 I342 (wen_0n[20], wc_1n, wc_0n);
  OR2 I343 (wen_0n[19], wc_1n, wc_0n);
  OR2 I344 (wen_0n[18], wc_1n, wc_0n);
  OR2 I345 (wen_0n[17], wc_1n, wc_0n);
  OR2 I346 (wen_0n[16], wc_1n, wc_0n);
  OR2 I347 (wen_0n[15], wc_1n, wc_0n);
  OR2 I348 (wen_0n[14], wc_1n, wc_0n);
  OR2 I349 (wen_0n[13], wc_1n, wc_0n);
  OR2 I350 (wen_0n[12], wc_1n, wc_0n);
  OR2 I351 (wen_0n[11], wc_1n, wc_0n);
  OR2 I352 (wen_0n[10], wc_1n, wc_0n);
  OR2 I353 (wen_0n[9], wc_1n, wc_0n);
  OR2 I354 (wen_0n[8], wc_1n, wc_0n);
  OR2 I355 (wen_0n[7], wc_1n, wc_0n);
  OR2 I356 (wen_0n[6], wc_1n, wc_0n);
  OR2 I357 (wen_0n[5], wc_1n, wc_0n);
  OR2 I358 (wen_0n[4], wc_1n, wc_0n);
  OR2 I359 (wen_0n[3], wc_1n, wc_0n);
  OR2 I360 (wen_0n[2], wc_1n, wc_0n);
  OR2 I361 (wen_0n[1], wc_1n, wc_0n);
  OR2 I362 (wen_0n[0], wc_1n, wc_0n);
  OR2 I363 (wt_0n[34], git_1n[34], git_0n[34]);
  OR2 I364 (wt_0n[33], git_1n[33], git_0n[33]);
  OR2 I365 (wt_0n[32], git_1n[32], git_0n[32]);
  OR2 I366 (wt_0n[31], git_1n[31], git_0n[31]);
  OR2 I367 (wt_0n[30], git_1n[30], git_0n[30]);
  OR2 I368 (wt_0n[29], git_1n[29], git_0n[29]);
  OR2 I369 (wt_0n[28], git_1n[28], git_0n[28]);
  OR2 I370 (wt_0n[27], git_1n[27], git_0n[27]);
  OR2 I371 (wt_0n[26], git_1n[26], git_0n[26]);
  OR2 I372 (wt_0n[25], git_1n[25], git_0n[25]);
  OR2 I373 (wt_0n[24], git_1n[24], git_0n[24]);
  OR2 I374 (wt_0n[23], git_1n[23], git_0n[23]);
  OR2 I375 (wt_0n[22], git_1n[22], git_0n[22]);
  OR2 I376 (wt_0n[21], git_1n[21], git_0n[21]);
  OR2 I377 (wt_0n[20], git_1n[20], git_0n[20]);
  OR2 I378 (wt_0n[19], git_1n[19], git_0n[19]);
  OR2 I379 (wt_0n[18], git_1n[18], git_0n[18]);
  OR2 I380 (wt_0n[17], git_1n[17], git_0n[17]);
  OR2 I381 (wt_0n[16], git_1n[16], git_0n[16]);
  OR2 I382 (wt_0n[15], git_1n[15], git_0n[15]);
  OR2 I383 (wt_0n[14], git_1n[14], git_0n[14]);
  OR2 I384 (wt_0n[13], git_1n[13], git_0n[13]);
  OR2 I385 (wt_0n[12], git_1n[12], git_0n[12]);
  OR2 I386 (wt_0n[11], git_1n[11], git_0n[11]);
  OR2 I387 (wt_0n[10], git_1n[10], git_0n[10]);
  OR2 I388 (wt_0n[9], git_1n[9], git_0n[9]);
  OR2 I389 (wt_0n[8], git_1n[8], git_0n[8]);
  OR2 I390 (wt_0n[7], git_1n[7], git_0n[7]);
  OR2 I391 (wt_0n[6], git_1n[6], git_0n[6]);
  OR2 I392 (wt_0n[5], git_1n[5], git_0n[5]);
  OR2 I393 (wt_0n[4], git_1n[4], git_0n[4]);
  OR2 I394 (wt_0n[3], git_1n[3], git_0n[3]);
  OR2 I395 (wt_0n[2], git_1n[2], git_0n[2]);
  OR2 I396 (wt_0n[1], git_1n[1], git_0n[1]);
  OR2 I397 (wt_0n[0], git_1n[0], git_0n[0]);
  OR2 I398 (wf_0n[34], gif_1n[34], gif_0n[34]);
  OR2 I399 (wf_0n[33], gif_1n[33], gif_0n[33]);
  OR2 I400 (wf_0n[32], gif_1n[32], gif_0n[32]);
  OR2 I401 (wf_0n[31], gif_1n[31], gif_0n[31]);
  OR2 I402 (wf_0n[30], gif_1n[30], gif_0n[30]);
  OR2 I403 (wf_0n[29], gif_1n[29], gif_0n[29]);
  OR2 I404 (wf_0n[28], gif_1n[28], gif_0n[28]);
  OR2 I405 (wf_0n[27], gif_1n[27], gif_0n[27]);
  OR2 I406 (wf_0n[26], gif_1n[26], gif_0n[26]);
  OR2 I407 (wf_0n[25], gif_1n[25], gif_0n[25]);
  OR2 I408 (wf_0n[24], gif_1n[24], gif_0n[24]);
  OR2 I409 (wf_0n[23], gif_1n[23], gif_0n[23]);
  OR2 I410 (wf_0n[22], gif_1n[22], gif_0n[22]);
  OR2 I411 (wf_0n[21], gif_1n[21], gif_0n[21]);
  OR2 I412 (wf_0n[20], gif_1n[20], gif_0n[20]);
  OR2 I413 (wf_0n[19], gif_1n[19], gif_0n[19]);
  OR2 I414 (wf_0n[18], gif_1n[18], gif_0n[18]);
  OR2 I415 (wf_0n[17], gif_1n[17], gif_0n[17]);
  OR2 I416 (wf_0n[16], gif_1n[16], gif_0n[16]);
  OR2 I417 (wf_0n[15], gif_1n[15], gif_0n[15]);
  OR2 I418 (wf_0n[14], gif_1n[14], gif_0n[14]);
  OR2 I419 (wf_0n[13], gif_1n[13], gif_0n[13]);
  OR2 I420 (wf_0n[12], gif_1n[12], gif_0n[12]);
  OR2 I421 (wf_0n[11], gif_1n[11], gif_0n[11]);
  OR2 I422 (wf_0n[10], gif_1n[10], gif_0n[10]);
  OR2 I423 (wf_0n[9], gif_1n[9], gif_0n[9]);
  OR2 I424 (wf_0n[8], gif_1n[8], gif_0n[8]);
  OR2 I425 (wf_0n[7], gif_1n[7], gif_0n[7]);
  OR2 I426 (wf_0n[6], gif_1n[6], gif_0n[6]);
  OR2 I427 (wf_0n[5], gif_1n[5], gif_0n[5]);
  OR2 I428 (wf_0n[4], gif_1n[4], gif_0n[4]);
  OR2 I429 (wf_0n[3], gif_1n[3], gif_0n[3]);
  OR2 I430 (wf_0n[2], gif_1n[2], gif_0n[2]);
  OR2 I431 (wf_0n[1], gif_1n[1], gif_0n[1]);
  OR2 I432 (wf_0n[0], gif_1n[0], gif_0n[0]);
  AC2 I433 (ig_0n, igc_0n, nanyread_0n);
  AC2 I434 (ig_1n, igc_1n, nanyread_0n);
  assign igc_0n = wc_0n;
  assign igc_1n = wc_1n;
  AND2 I437 (git_1n[0], wgtint_1n[0], ig_1n);
  AND2 I438 (git_1n[1], wgtint_1n[1], ig_1n);
  AND2 I439 (git_1n[2], wgtint_1n[2], ig_1n);
  AND2 I440 (git_1n[3], wgtint_1n[3], ig_1n);
  AND2 I441 (git_1n[4], wgtint_1n[4], ig_1n);
  AND2 I442 (git_1n[5], wgtint_1n[5], ig_1n);
  AND2 I443 (git_1n[6], wgtint_1n[6], ig_1n);
  AND2 I444 (git_1n[7], wgtint_1n[7], ig_1n);
  AND2 I445 (git_1n[8], wgtint_1n[8], ig_1n);
  AND2 I446 (git_1n[9], wgtint_1n[9], ig_1n);
  AND2 I447 (git_1n[10], wgtint_1n[10], ig_1n);
  AND2 I448 (git_1n[11], wgtint_1n[11], ig_1n);
  AND2 I449 (git_1n[12], wgtint_1n[12], ig_1n);
  AND2 I450 (git_1n[13], wgtint_1n[13], ig_1n);
  AND2 I451 (git_1n[14], wgtint_1n[14], ig_1n);
  AND2 I452 (git_1n[15], wgtint_1n[15], ig_1n);
  AND2 I453 (git_1n[16], wgtint_1n[16], ig_1n);
  AND2 I454 (git_1n[17], wgtint_1n[17], ig_1n);
  AND2 I455 (git_1n[18], wgtint_1n[18], ig_1n);
  AND2 I456 (git_1n[19], wgtint_1n[19], ig_1n);
  AND2 I457 (git_1n[20], wgtint_1n[20], ig_1n);
  AND2 I458 (git_1n[21], wgtint_1n[21], ig_1n);
  AND2 I459 (git_1n[22], wgtint_1n[22], ig_1n);
  AND2 I460 (git_1n[23], wgtint_1n[23], ig_1n);
  AND2 I461 (git_1n[24], wgtint_1n[24], ig_1n);
  AND2 I462 (git_1n[25], wgtint_1n[25], ig_1n);
  AND2 I463 (git_1n[26], wgtint_1n[26], ig_1n);
  AND2 I464 (git_1n[27], wgtint_1n[27], ig_1n);
  AND2 I465 (git_1n[28], wgtint_1n[28], ig_1n);
  AND2 I466 (git_1n[29], wgtint_1n[29], ig_1n);
  AND2 I467 (git_1n[30], wgtint_1n[30], ig_1n);
  AND2 I468 (git_1n[31], wgtint_1n[31], ig_1n);
  AND2 I469 (git_1n[32], wgtint_1n[32], ig_1n);
  AND2 I470 (git_1n[33], wgtint_1n[33], ig_1n);
  AND2 I471 (git_1n[34], wgtint_1n[34], ig_1n);
  AND2 I472 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I473 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I474 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I475 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I476 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I477 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I478 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I479 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I480 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I481 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I482 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I483 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I484 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I485 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I486 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I487 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I488 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I489 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I490 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I491 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I492 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I493 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I494 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I495 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I496 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I497 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I498 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I499 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I500 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I501 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I502 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I503 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I504 (git_0n[32], wgtint_0n[32], ig_0n);
  AND2 I505 (git_0n[33], wgtint_0n[33], ig_0n);
  AND2 I506 (git_0n[34], wgtint_0n[34], ig_0n);
  AND2 I507 (gif_1n[0], wgfint_1n[0], ig_1n);
  AND2 I508 (gif_1n[1], wgfint_1n[1], ig_1n);
  AND2 I509 (gif_1n[2], wgfint_1n[2], ig_1n);
  AND2 I510 (gif_1n[3], wgfint_1n[3], ig_1n);
  AND2 I511 (gif_1n[4], wgfint_1n[4], ig_1n);
  AND2 I512 (gif_1n[5], wgfint_1n[5], ig_1n);
  AND2 I513 (gif_1n[6], wgfint_1n[6], ig_1n);
  AND2 I514 (gif_1n[7], wgfint_1n[7], ig_1n);
  AND2 I515 (gif_1n[8], wgfint_1n[8], ig_1n);
  AND2 I516 (gif_1n[9], wgfint_1n[9], ig_1n);
  AND2 I517 (gif_1n[10], wgfint_1n[10], ig_1n);
  AND2 I518 (gif_1n[11], wgfint_1n[11], ig_1n);
  AND2 I519 (gif_1n[12], wgfint_1n[12], ig_1n);
  AND2 I520 (gif_1n[13], wgfint_1n[13], ig_1n);
  AND2 I521 (gif_1n[14], wgfint_1n[14], ig_1n);
  AND2 I522 (gif_1n[15], wgfint_1n[15], ig_1n);
  AND2 I523 (gif_1n[16], wgfint_1n[16], ig_1n);
  AND2 I524 (gif_1n[17], wgfint_1n[17], ig_1n);
  AND2 I525 (gif_1n[18], wgfint_1n[18], ig_1n);
  AND2 I526 (gif_1n[19], wgfint_1n[19], ig_1n);
  AND2 I527 (gif_1n[20], wgfint_1n[20], ig_1n);
  AND2 I528 (gif_1n[21], wgfint_1n[21], ig_1n);
  AND2 I529 (gif_1n[22], wgfint_1n[22], ig_1n);
  AND2 I530 (gif_1n[23], wgfint_1n[23], ig_1n);
  AND2 I531 (gif_1n[24], wgfint_1n[24], ig_1n);
  AND2 I532 (gif_1n[25], wgfint_1n[25], ig_1n);
  AND2 I533 (gif_1n[26], wgfint_1n[26], ig_1n);
  AND2 I534 (gif_1n[27], wgfint_1n[27], ig_1n);
  AND2 I535 (gif_1n[28], wgfint_1n[28], ig_1n);
  AND2 I536 (gif_1n[29], wgfint_1n[29], ig_1n);
  AND2 I537 (gif_1n[30], wgfint_1n[30], ig_1n);
  AND2 I538 (gif_1n[31], wgfint_1n[31], ig_1n);
  AND2 I539 (gif_1n[32], wgfint_1n[32], ig_1n);
  AND2 I540 (gif_1n[33], wgfint_1n[33], ig_1n);
  AND2 I541 (gif_1n[34], wgfint_1n[34], ig_1n);
  AND2 I542 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I543 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I544 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I545 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I546 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I547 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I548 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I549 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I550 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I551 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I552 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I553 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I554 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I555 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I556 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I557 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I558 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I559 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I560 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I561 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I562 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I563 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I564 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I565 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I566 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I567 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I568 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I569 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I570 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I571 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I572 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I573 (gif_0n[31], wgfint_0n[31], ig_0n);
  AND2 I574 (gif_0n[32], wgfint_0n[32], ig_0n);
  AND2 I575 (gif_0n[33], wgfint_0n[33], ig_0n);
  AND2 I576 (gif_0n[34], wgfint_0n[34], ig_0n);
  C3 I577 (internal_0n[36], complete1559_0n[0], complete1559_0n[1], complete1559_0n[2]);
  C3 I578 (internal_0n[37], complete1559_0n[3], complete1559_0n[4], complete1559_0n[5]);
  C3 I579 (internal_0n[38], complete1559_0n[6], complete1559_0n[7], complete1559_0n[8]);
  C3 I580 (internal_0n[39], complete1559_0n[9], complete1559_0n[10], complete1559_0n[11]);
  C3 I581 (internal_0n[40], complete1559_0n[12], complete1559_0n[13], complete1559_0n[14]);
  C3 I582 (internal_0n[41], complete1559_0n[15], complete1559_0n[16], complete1559_0n[17]);
  C3 I583 (internal_0n[42], complete1559_0n[18], complete1559_0n[19], complete1559_0n[20]);
  C3 I584 (internal_0n[43], complete1559_0n[21], complete1559_0n[22], complete1559_0n[23]);
  C3 I585 (internal_0n[44], complete1559_0n[24], complete1559_0n[25], complete1559_0n[26]);
  C3 I586 (internal_0n[45], complete1559_0n[27], complete1559_0n[28], complete1559_0n[29]);
  C3 I587 (internal_0n[46], complete1559_0n[30], complete1559_0n[31], complete1559_0n[32]);
  C2 I588 (internal_0n[47], complete1559_0n[33], complete1559_0n[34]);
  C3 I589 (internal_0n[48], internal_0n[36], internal_0n[37], internal_0n[38]);
  C3 I590 (internal_0n[49], internal_0n[39], internal_0n[40], internal_0n[41]);
  C3 I591 (internal_0n[50], internal_0n[42], internal_0n[43], internal_0n[44]);
  C3 I592 (internal_0n[51], internal_0n[45], internal_0n[46], internal_0n[47]);
  C2 I593 (internal_0n[52], internal_0n[48], internal_0n[49]);
  C2 I594 (internal_0n[53], internal_0n[50], internal_0n[51]);
  C2 I595 (wc_1n, internal_0n[52], internal_0n[53]);
  OR2 I596 (complete1559_0n[0], wgfint_1n[0], wgtint_1n[0]);
  OR2 I597 (complete1559_0n[1], wgfint_1n[1], wgtint_1n[1]);
  OR2 I598 (complete1559_0n[2], wgfint_1n[2], wgtint_1n[2]);
  OR2 I599 (complete1559_0n[3], wgfint_1n[3], wgtint_1n[3]);
  OR2 I600 (complete1559_0n[4], wgfint_1n[4], wgtint_1n[4]);
  OR2 I601 (complete1559_0n[5], wgfint_1n[5], wgtint_1n[5]);
  OR2 I602 (complete1559_0n[6], wgfint_1n[6], wgtint_1n[6]);
  OR2 I603 (complete1559_0n[7], wgfint_1n[7], wgtint_1n[7]);
  OR2 I604 (complete1559_0n[8], wgfint_1n[8], wgtint_1n[8]);
  OR2 I605 (complete1559_0n[9], wgfint_1n[9], wgtint_1n[9]);
  OR2 I606 (complete1559_0n[10], wgfint_1n[10], wgtint_1n[10]);
  OR2 I607 (complete1559_0n[11], wgfint_1n[11], wgtint_1n[11]);
  OR2 I608 (complete1559_0n[12], wgfint_1n[12], wgtint_1n[12]);
  OR2 I609 (complete1559_0n[13], wgfint_1n[13], wgtint_1n[13]);
  OR2 I610 (complete1559_0n[14], wgfint_1n[14], wgtint_1n[14]);
  OR2 I611 (complete1559_0n[15], wgfint_1n[15], wgtint_1n[15]);
  OR2 I612 (complete1559_0n[16], wgfint_1n[16], wgtint_1n[16]);
  OR2 I613 (complete1559_0n[17], wgfint_1n[17], wgtint_1n[17]);
  OR2 I614 (complete1559_0n[18], wgfint_1n[18], wgtint_1n[18]);
  OR2 I615 (complete1559_0n[19], wgfint_1n[19], wgtint_1n[19]);
  OR2 I616 (complete1559_0n[20], wgfint_1n[20], wgtint_1n[20]);
  OR2 I617 (complete1559_0n[21], wgfint_1n[21], wgtint_1n[21]);
  OR2 I618 (complete1559_0n[22], wgfint_1n[22], wgtint_1n[22]);
  OR2 I619 (complete1559_0n[23], wgfint_1n[23], wgtint_1n[23]);
  OR2 I620 (complete1559_0n[24], wgfint_1n[24], wgtint_1n[24]);
  OR2 I621 (complete1559_0n[25], wgfint_1n[25], wgtint_1n[25]);
  OR2 I622 (complete1559_0n[26], wgfint_1n[26], wgtint_1n[26]);
  OR2 I623 (complete1559_0n[27], wgfint_1n[27], wgtint_1n[27]);
  OR2 I624 (complete1559_0n[28], wgfint_1n[28], wgtint_1n[28]);
  OR2 I625 (complete1559_0n[29], wgfint_1n[29], wgtint_1n[29]);
  OR2 I626 (complete1559_0n[30], wgfint_1n[30], wgtint_1n[30]);
  OR2 I627 (complete1559_0n[31], wgfint_1n[31], wgtint_1n[31]);
  OR2 I628 (complete1559_0n[32], wgfint_1n[32], wgtint_1n[32]);
  OR2 I629 (complete1559_0n[33], wgfint_1n[33], wgtint_1n[33]);
  OR2 I630 (complete1559_0n[34], wgfint_1n[34], wgtint_1n[34]);
  C3 I631 (internal_0n[54], complete1558_0n[0], complete1558_0n[1], complete1558_0n[2]);
  C3 I632 (internal_0n[55], complete1558_0n[3], complete1558_0n[4], complete1558_0n[5]);
  C3 I633 (internal_0n[56], complete1558_0n[6], complete1558_0n[7], complete1558_0n[8]);
  C3 I634 (internal_0n[57], complete1558_0n[9], complete1558_0n[10], complete1558_0n[11]);
  C3 I635 (internal_0n[58], complete1558_0n[12], complete1558_0n[13], complete1558_0n[14]);
  C3 I636 (internal_0n[59], complete1558_0n[15], complete1558_0n[16], complete1558_0n[17]);
  C3 I637 (internal_0n[60], complete1558_0n[18], complete1558_0n[19], complete1558_0n[20]);
  C3 I638 (internal_0n[61], complete1558_0n[21], complete1558_0n[22], complete1558_0n[23]);
  C3 I639 (internal_0n[62], complete1558_0n[24], complete1558_0n[25], complete1558_0n[26]);
  C3 I640 (internal_0n[63], complete1558_0n[27], complete1558_0n[28], complete1558_0n[29]);
  C3 I641 (internal_0n[64], complete1558_0n[30], complete1558_0n[31], complete1558_0n[32]);
  C2 I642 (internal_0n[65], complete1558_0n[33], complete1558_0n[34]);
  C3 I643 (internal_0n[66], internal_0n[54], internal_0n[55], internal_0n[56]);
  C3 I644 (internal_0n[67], internal_0n[57], internal_0n[58], internal_0n[59]);
  C3 I645 (internal_0n[68], internal_0n[60], internal_0n[61], internal_0n[62]);
  C3 I646 (internal_0n[69], internal_0n[63], internal_0n[64], internal_0n[65]);
  C2 I647 (internal_0n[70], internal_0n[66], internal_0n[67]);
  C2 I648 (internal_0n[71], internal_0n[68], internal_0n[69]);
  C2 I649 (wc_0n, internal_0n[70], internal_0n[71]);
  OR2 I650 (complete1558_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I651 (complete1558_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I652 (complete1558_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I653 (complete1558_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I654 (complete1558_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I655 (complete1558_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I656 (complete1558_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I657 (complete1558_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I658 (complete1558_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I659 (complete1558_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I660 (complete1558_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I661 (complete1558_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I662 (complete1558_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I663 (complete1558_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I664 (complete1558_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I665 (complete1558_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I666 (complete1558_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I667 (complete1558_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I668 (complete1558_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I669 (complete1558_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I670 (complete1558_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I671 (complete1558_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I672 (complete1558_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I673 (complete1558_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I674 (complete1558_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I675 (complete1558_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I676 (complete1558_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I677 (complete1558_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I678 (complete1558_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I679 (complete1558_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I680 (complete1558_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I681 (complete1558_0n[31], wgfint_0n[31], wgtint_0n[31]);
  OR2 I682 (complete1558_0n[32], wgfint_0n[32], wgtint_0n[32]);
  OR2 I683 (complete1558_0n[33], wgfint_0n[33], wgtint_0n[33]);
  OR2 I684 (complete1558_0n[34], wgfint_0n[34], wgtint_0n[34]);
  AO22 I685 (wacks_0n[34], gf1556_0n[34], df_0n[34], gt1557_0n[34], dt_0n[34]);
  NOR2 I686 (dt_0n[34], df_0n[34], gf1556_0n[34]);
  NOR3 I687 (df_0n[34], dt_0n[34], gt1557_0n[34], init_0n);
  AND2 I688 (gt1557_0n[34], wt_0n[34], wen_0n[34]);
  AND2 I689 (gf1556_0n[34], wf_0n[34], wen_0n[34]);
  AO22 I690 (wacks_0n[33], gf1556_0n[33], df_0n[33], gt1557_0n[33], dt_0n[33]);
  NOR2 I691 (dt_0n[33], df_0n[33], gf1556_0n[33]);
  NOR3 I692 (df_0n[33], dt_0n[33], gt1557_0n[33], init_0n);
  AND2 I693 (gt1557_0n[33], wt_0n[33], wen_0n[33]);
  AND2 I694 (gf1556_0n[33], wf_0n[33], wen_0n[33]);
  AO22 I695 (wacks_0n[32], gf1556_0n[32], df_0n[32], gt1557_0n[32], dt_0n[32]);
  NOR2 I696 (dt_0n[32], df_0n[32], gf1556_0n[32]);
  NOR3 I697 (df_0n[32], dt_0n[32], gt1557_0n[32], init_0n);
  AND2 I698 (gt1557_0n[32], wt_0n[32], wen_0n[32]);
  AND2 I699 (gf1556_0n[32], wf_0n[32], wen_0n[32]);
  AO22 I700 (wacks_0n[31], gf1556_0n[31], df_0n[31], gt1557_0n[31], dt_0n[31]);
  NOR2 I701 (dt_0n[31], df_0n[31], gf1556_0n[31]);
  NOR3 I702 (df_0n[31], dt_0n[31], gt1557_0n[31], init_0n);
  AND2 I703 (gt1557_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I704 (gf1556_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I705 (wacks_0n[30], gf1556_0n[30], df_0n[30], gt1557_0n[30], dt_0n[30]);
  NOR2 I706 (dt_0n[30], df_0n[30], gf1556_0n[30]);
  NOR3 I707 (df_0n[30], dt_0n[30], gt1557_0n[30], init_0n);
  AND2 I708 (gt1557_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I709 (gf1556_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I710 (wacks_0n[29], gf1556_0n[29], df_0n[29], gt1557_0n[29], dt_0n[29]);
  NOR2 I711 (dt_0n[29], df_0n[29], gf1556_0n[29]);
  NOR3 I712 (df_0n[29], dt_0n[29], gt1557_0n[29], init_0n);
  AND2 I713 (gt1557_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I714 (gf1556_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I715 (wacks_0n[28], gf1556_0n[28], df_0n[28], gt1557_0n[28], dt_0n[28]);
  NOR2 I716 (dt_0n[28], df_0n[28], gf1556_0n[28]);
  NOR3 I717 (df_0n[28], dt_0n[28], gt1557_0n[28], init_0n);
  AND2 I718 (gt1557_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I719 (gf1556_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I720 (wacks_0n[27], gf1556_0n[27], df_0n[27], gt1557_0n[27], dt_0n[27]);
  NOR2 I721 (dt_0n[27], df_0n[27], gf1556_0n[27]);
  NOR3 I722 (df_0n[27], dt_0n[27], gt1557_0n[27], init_0n);
  AND2 I723 (gt1557_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I724 (gf1556_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I725 (wacks_0n[26], gf1556_0n[26], df_0n[26], gt1557_0n[26], dt_0n[26]);
  NOR2 I726 (dt_0n[26], df_0n[26], gf1556_0n[26]);
  NOR3 I727 (df_0n[26], dt_0n[26], gt1557_0n[26], init_0n);
  AND2 I728 (gt1557_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I729 (gf1556_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I730 (wacks_0n[25], gf1556_0n[25], df_0n[25], gt1557_0n[25], dt_0n[25]);
  NOR2 I731 (dt_0n[25], df_0n[25], gf1556_0n[25]);
  NOR3 I732 (df_0n[25], dt_0n[25], gt1557_0n[25], init_0n);
  AND2 I733 (gt1557_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I734 (gf1556_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I735 (wacks_0n[24], gf1556_0n[24], df_0n[24], gt1557_0n[24], dt_0n[24]);
  NOR2 I736 (dt_0n[24], df_0n[24], gf1556_0n[24]);
  NOR3 I737 (df_0n[24], dt_0n[24], gt1557_0n[24], init_0n);
  AND2 I738 (gt1557_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I739 (gf1556_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I740 (wacks_0n[23], gf1556_0n[23], df_0n[23], gt1557_0n[23], dt_0n[23]);
  NOR2 I741 (dt_0n[23], df_0n[23], gf1556_0n[23]);
  NOR3 I742 (df_0n[23], dt_0n[23], gt1557_0n[23], init_0n);
  AND2 I743 (gt1557_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I744 (gf1556_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I745 (wacks_0n[22], gf1556_0n[22], df_0n[22], gt1557_0n[22], dt_0n[22]);
  NOR2 I746 (dt_0n[22], df_0n[22], gf1556_0n[22]);
  NOR3 I747 (df_0n[22], dt_0n[22], gt1557_0n[22], init_0n);
  AND2 I748 (gt1557_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I749 (gf1556_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I750 (wacks_0n[21], gf1556_0n[21], df_0n[21], gt1557_0n[21], dt_0n[21]);
  NOR2 I751 (dt_0n[21], df_0n[21], gf1556_0n[21]);
  NOR3 I752 (df_0n[21], dt_0n[21], gt1557_0n[21], init_0n);
  AND2 I753 (gt1557_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I754 (gf1556_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I755 (wacks_0n[20], gf1556_0n[20], df_0n[20], gt1557_0n[20], dt_0n[20]);
  NOR2 I756 (dt_0n[20], df_0n[20], gf1556_0n[20]);
  NOR3 I757 (df_0n[20], dt_0n[20], gt1557_0n[20], init_0n);
  AND2 I758 (gt1557_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I759 (gf1556_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I760 (wacks_0n[19], gf1556_0n[19], df_0n[19], gt1557_0n[19], dt_0n[19]);
  NOR2 I761 (dt_0n[19], df_0n[19], gf1556_0n[19]);
  NOR3 I762 (df_0n[19], dt_0n[19], gt1557_0n[19], init_0n);
  AND2 I763 (gt1557_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I764 (gf1556_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I765 (wacks_0n[18], gf1556_0n[18], df_0n[18], gt1557_0n[18], dt_0n[18]);
  NOR2 I766 (dt_0n[18], df_0n[18], gf1556_0n[18]);
  NOR3 I767 (df_0n[18], dt_0n[18], gt1557_0n[18], init_0n);
  AND2 I768 (gt1557_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I769 (gf1556_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I770 (wacks_0n[17], gf1556_0n[17], df_0n[17], gt1557_0n[17], dt_0n[17]);
  NOR2 I771 (dt_0n[17], df_0n[17], gf1556_0n[17]);
  NOR3 I772 (df_0n[17], dt_0n[17], gt1557_0n[17], init_0n);
  AND2 I773 (gt1557_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I774 (gf1556_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I775 (wacks_0n[16], gf1556_0n[16], df_0n[16], gt1557_0n[16], dt_0n[16]);
  NOR2 I776 (dt_0n[16], df_0n[16], gf1556_0n[16]);
  NOR3 I777 (df_0n[16], dt_0n[16], gt1557_0n[16], init_0n);
  AND2 I778 (gt1557_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I779 (gf1556_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I780 (wacks_0n[15], gf1556_0n[15], df_0n[15], gt1557_0n[15], dt_0n[15]);
  NOR2 I781 (dt_0n[15], df_0n[15], gf1556_0n[15]);
  NOR3 I782 (df_0n[15], dt_0n[15], gt1557_0n[15], init_0n);
  AND2 I783 (gt1557_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I784 (gf1556_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I785 (wacks_0n[14], gf1556_0n[14], df_0n[14], gt1557_0n[14], dt_0n[14]);
  NOR2 I786 (dt_0n[14], df_0n[14], gf1556_0n[14]);
  NOR3 I787 (df_0n[14], dt_0n[14], gt1557_0n[14], init_0n);
  AND2 I788 (gt1557_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I789 (gf1556_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I790 (wacks_0n[13], gf1556_0n[13], df_0n[13], gt1557_0n[13], dt_0n[13]);
  NOR2 I791 (dt_0n[13], df_0n[13], gf1556_0n[13]);
  NOR3 I792 (df_0n[13], dt_0n[13], gt1557_0n[13], init_0n);
  AND2 I793 (gt1557_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I794 (gf1556_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I795 (wacks_0n[12], gf1556_0n[12], df_0n[12], gt1557_0n[12], dt_0n[12]);
  NOR2 I796 (dt_0n[12], df_0n[12], gf1556_0n[12]);
  NOR3 I797 (df_0n[12], dt_0n[12], gt1557_0n[12], init_0n);
  AND2 I798 (gt1557_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I799 (gf1556_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I800 (wacks_0n[11], gf1556_0n[11], df_0n[11], gt1557_0n[11], dt_0n[11]);
  NOR2 I801 (dt_0n[11], df_0n[11], gf1556_0n[11]);
  NOR3 I802 (df_0n[11], dt_0n[11], gt1557_0n[11], init_0n);
  AND2 I803 (gt1557_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I804 (gf1556_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I805 (wacks_0n[10], gf1556_0n[10], df_0n[10], gt1557_0n[10], dt_0n[10]);
  NOR2 I806 (dt_0n[10], df_0n[10], gf1556_0n[10]);
  NOR3 I807 (df_0n[10], dt_0n[10], gt1557_0n[10], init_0n);
  AND2 I808 (gt1557_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I809 (gf1556_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I810 (wacks_0n[9], gf1556_0n[9], df_0n[9], gt1557_0n[9], dt_0n[9]);
  NOR2 I811 (dt_0n[9], df_0n[9], gf1556_0n[9]);
  NOR3 I812 (df_0n[9], dt_0n[9], gt1557_0n[9], init_0n);
  AND2 I813 (gt1557_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I814 (gf1556_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I815 (wacks_0n[8], gf1556_0n[8], df_0n[8], gt1557_0n[8], dt_0n[8]);
  NOR2 I816 (dt_0n[8], df_0n[8], gf1556_0n[8]);
  NOR3 I817 (df_0n[8], dt_0n[8], gt1557_0n[8], init_0n);
  AND2 I818 (gt1557_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I819 (gf1556_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I820 (wacks_0n[7], gf1556_0n[7], df_0n[7], gt1557_0n[7], dt_0n[7]);
  NOR2 I821 (dt_0n[7], df_0n[7], gf1556_0n[7]);
  NOR3 I822 (df_0n[7], dt_0n[7], gt1557_0n[7], init_0n);
  AND2 I823 (gt1557_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I824 (gf1556_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I825 (wacks_0n[6], gf1556_0n[6], df_0n[6], gt1557_0n[6], dt_0n[6]);
  NOR2 I826 (dt_0n[6], df_0n[6], gf1556_0n[6]);
  NOR3 I827 (df_0n[6], dt_0n[6], gt1557_0n[6], init_0n);
  AND2 I828 (gt1557_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I829 (gf1556_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I830 (wacks_0n[5], gf1556_0n[5], df_0n[5], gt1557_0n[5], dt_0n[5]);
  NOR2 I831 (dt_0n[5], df_0n[5], gf1556_0n[5]);
  NOR3 I832 (df_0n[5], dt_0n[5], gt1557_0n[5], init_0n);
  AND2 I833 (gt1557_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I834 (gf1556_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I835 (wacks_0n[4], gf1556_0n[4], df_0n[4], gt1557_0n[4], dt_0n[4]);
  NOR2 I836 (dt_0n[4], df_0n[4], gf1556_0n[4]);
  NOR3 I837 (df_0n[4], dt_0n[4], gt1557_0n[4], init_0n);
  AND2 I838 (gt1557_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I839 (gf1556_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I840 (wacks_0n[3], gf1556_0n[3], df_0n[3], gt1557_0n[3], dt_0n[3]);
  NOR2 I841 (dt_0n[3], df_0n[3], gf1556_0n[3]);
  NOR3 I842 (df_0n[3], dt_0n[3], gt1557_0n[3], init_0n);
  AND2 I843 (gt1557_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I844 (gf1556_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I845 (wacks_0n[2], gf1556_0n[2], df_0n[2], gt1557_0n[2], dt_0n[2]);
  NOR2 I846 (dt_0n[2], df_0n[2], gf1556_0n[2]);
  NOR3 I847 (df_0n[2], dt_0n[2], gt1557_0n[2], init_0n);
  AND2 I848 (gt1557_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I849 (gf1556_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I850 (wacks_0n[1], gf1556_0n[1], df_0n[1], gt1557_0n[1], dt_0n[1]);
  NOR2 I851 (dt_0n[1], df_0n[1], gf1556_0n[1]);
  NOR3 I852 (df_0n[1], dt_0n[1], gt1557_0n[1], init_0n);
  AND2 I853 (gt1557_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I854 (gf1556_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I855 (wacks_0n[0], gf1556_0n[0], df_0n[0], gt1557_0n[0], dt_0n[0]);
  NOR2 I856 (dt_0n[0], df_0n[0], gf1556_0n[0]);
  NOR3 I857 (df_0n[0], dt_0n[0], gt1557_0n[0], init_0n);
  AND2 I858 (gt1557_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I859 (gf1556_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I860 (init_0n, initialise);
endmodule

module BrzV_36_l6__28_29_l24__28_28_280_2036_29_2_m95m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  initialise
);
  input [35:0] wg_0r0d;
  input [35:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [35:0] rd_0r0d;
  output [35:0] rd_0r1d;
  input rd_0a;
  output [3:0] rd_1r0d;
  output [3:0] rd_1r1d;
  input rd_1a;
  input initialise;
  wire [39:0] internal_0n;
  wire [35:0] wf_0n;
  wire [35:0] wt_0n;
  wire [35:0] df_0n;
  wire [35:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire wc_0n;
  wire [35:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [35:0] wgfint_0n;
  wire [35:0] wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire [35:0] rdfint_0n;
  wire [3:0] rdfint_1n;
  wire [35:0] rdtint_0n;
  wire [3:0] rdtint_1n;
  wire [35:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [35:0] gif_0n;
  wire [35:0] git_0n;
  wire [35:0] complete1574_0n;
  wire [35:0] gt1573_0n;
  wire [35:0] gf1572_0n;
  assign rgaint_1n = rd_1a;
  assign rd_1r0d[0] = rdfint_1n[0];
  assign rd_1r0d[1] = rdfint_1n[1];
  assign rd_1r0d[2] = rdfint_1n[2];
  assign rd_1r0d[3] = rdfint_1n[3];
  assign rd_1r1d[0] = rdtint_1n[0];
  assign rd_1r1d[1] = rdtint_1n[1];
  assign rd_1r1d[2] = rdtint_1n[2];
  assign rd_1r1d[3] = rdtint_1n[3];
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r0d[10] = rdfint_0n[10];
  assign rd_0r0d[11] = rdfint_0n[11];
  assign rd_0r0d[12] = rdfint_0n[12];
  assign rd_0r0d[13] = rdfint_0n[13];
  assign rd_0r0d[14] = rdfint_0n[14];
  assign rd_0r0d[15] = rdfint_0n[15];
  assign rd_0r0d[16] = rdfint_0n[16];
  assign rd_0r0d[17] = rdfint_0n[17];
  assign rd_0r0d[18] = rdfint_0n[18];
  assign rd_0r0d[19] = rdfint_0n[19];
  assign rd_0r0d[20] = rdfint_0n[20];
  assign rd_0r0d[21] = rdfint_0n[21];
  assign rd_0r0d[22] = rdfint_0n[22];
  assign rd_0r0d[23] = rdfint_0n[23];
  assign rd_0r0d[24] = rdfint_0n[24];
  assign rd_0r0d[25] = rdfint_0n[25];
  assign rd_0r0d[26] = rdfint_0n[26];
  assign rd_0r0d[27] = rdfint_0n[27];
  assign rd_0r0d[28] = rdfint_0n[28];
  assign rd_0r0d[29] = rdfint_0n[29];
  assign rd_0r0d[30] = rdfint_0n[30];
  assign rd_0r0d[31] = rdfint_0n[31];
  assign rd_0r0d[32] = rdfint_0n[32];
  assign rd_0r0d[33] = rdfint_0n[33];
  assign rd_0r0d[34] = rdfint_0n[34];
  assign rd_0r0d[35] = rdfint_0n[35];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign rd_0r1d[10] = rdtint_0n[10];
  assign rd_0r1d[11] = rdtint_0n[11];
  assign rd_0r1d[12] = rdtint_0n[12];
  assign rd_0r1d[13] = rdtint_0n[13];
  assign rd_0r1d[14] = rdtint_0n[14];
  assign rd_0r1d[15] = rdtint_0n[15];
  assign rd_0r1d[16] = rdtint_0n[16];
  assign rd_0r1d[17] = rdtint_0n[17];
  assign rd_0r1d[18] = rdtint_0n[18];
  assign rd_0r1d[19] = rdtint_0n[19];
  assign rd_0r1d[20] = rdtint_0n[20];
  assign rd_0r1d[21] = rdtint_0n[21];
  assign rd_0r1d[22] = rdtint_0n[22];
  assign rd_0r1d[23] = rdtint_0n[23];
  assign rd_0r1d[24] = rdtint_0n[24];
  assign rd_0r1d[25] = rdtint_0n[25];
  assign rd_0r1d[26] = rdtint_0n[26];
  assign rd_0r1d[27] = rdtint_0n[27];
  assign rd_0r1d[28] = rdtint_0n[28];
  assign rd_0r1d[29] = rdtint_0n[29];
  assign rd_0r1d[30] = rdtint_0n[30];
  assign rd_0r1d[31] = rdtint_0n[31];
  assign rd_0r1d[32] = rdtint_0n[32];
  assign rd_0r1d[33] = rdtint_0n[33];
  assign rd_0r1d[34] = rdtint_0n[34];
  assign rd_0r1d[35] = rdtint_0n[35];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgfint_0n[32] = wg_0r0d[32];
  assign wgfint_0n[33] = wg_0r0d[33];
  assign wgfint_0n[34] = wg_0r0d[34];
  assign wgfint_0n[35] = wg_0r0d[35];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign wgtint_0n[32] = wg_0r1d[32];
  assign wgtint_0n[33] = wg_0r1d[33];
  assign wgtint_0n[34] = wg_0r1d[34];
  assign wgtint_0n[35] = wg_0r1d[35];
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I161 (internal_0n[0], rgrint_0n, rgrint_1n);
  NOR2 I162 (internal_0n[1], rgaint_0n, rgaint_1n);
  AND2 I163 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I164 (rdtint_1n[0], rgrint_1n, dt_0n[0]);
  AND2 I165 (rdtint_1n[1], rgrint_1n, dt_0n[1]);
  AND2 I166 (rdtint_1n[2], rgrint_1n, dt_0n[2]);
  AND2 I167 (rdtint_1n[3], rgrint_1n, dt_0n[3]);
  AND2 I168 (rdtint_0n[0], rgrint_0n, dt_0n[0]);
  AND2 I169 (rdtint_0n[1], rgrint_0n, dt_0n[1]);
  AND2 I170 (rdtint_0n[2], rgrint_0n, dt_0n[2]);
  AND2 I171 (rdtint_0n[3], rgrint_0n, dt_0n[3]);
  AND2 I172 (rdtint_0n[4], rgrint_0n, dt_0n[4]);
  AND2 I173 (rdtint_0n[5], rgrint_0n, dt_0n[5]);
  AND2 I174 (rdtint_0n[6], rgrint_0n, dt_0n[6]);
  AND2 I175 (rdtint_0n[7], rgrint_0n, dt_0n[7]);
  AND2 I176 (rdtint_0n[8], rgrint_0n, dt_0n[8]);
  AND2 I177 (rdtint_0n[9], rgrint_0n, dt_0n[9]);
  AND2 I178 (rdtint_0n[10], rgrint_0n, dt_0n[10]);
  AND2 I179 (rdtint_0n[11], rgrint_0n, dt_0n[11]);
  AND2 I180 (rdtint_0n[12], rgrint_0n, dt_0n[12]);
  AND2 I181 (rdtint_0n[13], rgrint_0n, dt_0n[13]);
  AND2 I182 (rdtint_0n[14], rgrint_0n, dt_0n[14]);
  AND2 I183 (rdtint_0n[15], rgrint_0n, dt_0n[15]);
  AND2 I184 (rdtint_0n[16], rgrint_0n, dt_0n[16]);
  AND2 I185 (rdtint_0n[17], rgrint_0n, dt_0n[17]);
  AND2 I186 (rdtint_0n[18], rgrint_0n, dt_0n[18]);
  AND2 I187 (rdtint_0n[19], rgrint_0n, dt_0n[19]);
  AND2 I188 (rdtint_0n[20], rgrint_0n, dt_0n[20]);
  AND2 I189 (rdtint_0n[21], rgrint_0n, dt_0n[21]);
  AND2 I190 (rdtint_0n[22], rgrint_0n, dt_0n[22]);
  AND2 I191 (rdtint_0n[23], rgrint_0n, dt_0n[23]);
  AND2 I192 (rdtint_0n[24], rgrint_0n, dt_0n[24]);
  AND2 I193 (rdtint_0n[25], rgrint_0n, dt_0n[25]);
  AND2 I194 (rdtint_0n[26], rgrint_0n, dt_0n[26]);
  AND2 I195 (rdtint_0n[27], rgrint_0n, dt_0n[27]);
  AND2 I196 (rdtint_0n[28], rgrint_0n, dt_0n[28]);
  AND2 I197 (rdtint_0n[29], rgrint_0n, dt_0n[29]);
  AND2 I198 (rdtint_0n[30], rgrint_0n, dt_0n[30]);
  AND2 I199 (rdtint_0n[31], rgrint_0n, dt_0n[31]);
  AND2 I200 (rdtint_0n[32], rgrint_0n, dt_0n[32]);
  AND2 I201 (rdtint_0n[33], rgrint_0n, dt_0n[33]);
  AND2 I202 (rdtint_0n[34], rgrint_0n, dt_0n[34]);
  AND2 I203 (rdtint_0n[35], rgrint_0n, dt_0n[35]);
  AND2 I204 (rdfint_1n[0], rgrint_1n, df_0n[0]);
  AND2 I205 (rdfint_1n[1], rgrint_1n, df_0n[1]);
  AND2 I206 (rdfint_1n[2], rgrint_1n, df_0n[2]);
  AND2 I207 (rdfint_1n[3], rgrint_1n, df_0n[3]);
  AND2 I208 (rdfint_0n[0], rgrint_0n, df_0n[0]);
  AND2 I209 (rdfint_0n[1], rgrint_0n, df_0n[1]);
  AND2 I210 (rdfint_0n[2], rgrint_0n, df_0n[2]);
  AND2 I211 (rdfint_0n[3], rgrint_0n, df_0n[3]);
  AND2 I212 (rdfint_0n[4], rgrint_0n, df_0n[4]);
  AND2 I213 (rdfint_0n[5], rgrint_0n, df_0n[5]);
  AND2 I214 (rdfint_0n[6], rgrint_0n, df_0n[6]);
  AND2 I215 (rdfint_0n[7], rgrint_0n, df_0n[7]);
  AND2 I216 (rdfint_0n[8], rgrint_0n, df_0n[8]);
  AND2 I217 (rdfint_0n[9], rgrint_0n, df_0n[9]);
  AND2 I218 (rdfint_0n[10], rgrint_0n, df_0n[10]);
  AND2 I219 (rdfint_0n[11], rgrint_0n, df_0n[11]);
  AND2 I220 (rdfint_0n[12], rgrint_0n, df_0n[12]);
  AND2 I221 (rdfint_0n[13], rgrint_0n, df_0n[13]);
  AND2 I222 (rdfint_0n[14], rgrint_0n, df_0n[14]);
  AND2 I223 (rdfint_0n[15], rgrint_0n, df_0n[15]);
  AND2 I224 (rdfint_0n[16], rgrint_0n, df_0n[16]);
  AND2 I225 (rdfint_0n[17], rgrint_0n, df_0n[17]);
  AND2 I226 (rdfint_0n[18], rgrint_0n, df_0n[18]);
  AND2 I227 (rdfint_0n[19], rgrint_0n, df_0n[19]);
  AND2 I228 (rdfint_0n[20], rgrint_0n, df_0n[20]);
  AND2 I229 (rdfint_0n[21], rgrint_0n, df_0n[21]);
  AND2 I230 (rdfint_0n[22], rgrint_0n, df_0n[22]);
  AND2 I231 (rdfint_0n[23], rgrint_0n, df_0n[23]);
  AND2 I232 (rdfint_0n[24], rgrint_0n, df_0n[24]);
  AND2 I233 (rdfint_0n[25], rgrint_0n, df_0n[25]);
  AND2 I234 (rdfint_0n[26], rgrint_0n, df_0n[26]);
  AND2 I235 (rdfint_0n[27], rgrint_0n, df_0n[27]);
  AND2 I236 (rdfint_0n[28], rgrint_0n, df_0n[28]);
  AND2 I237 (rdfint_0n[29], rgrint_0n, df_0n[29]);
  AND2 I238 (rdfint_0n[30], rgrint_0n, df_0n[30]);
  AND2 I239 (rdfint_0n[31], rgrint_0n, df_0n[31]);
  AND2 I240 (rdfint_0n[32], rgrint_0n, df_0n[32]);
  AND2 I241 (rdfint_0n[33], rgrint_0n, df_0n[33]);
  AND2 I242 (rdfint_0n[34], rgrint_0n, df_0n[34]);
  AND2 I243 (rdfint_0n[35], rgrint_0n, df_0n[35]);
  C3 I244 (internal_0n[2], wc_0n, wacks_0n[35], wacks_0n[34]);
  C3 I245 (internal_0n[3], wacks_0n[33], wacks_0n[32], wacks_0n[31]);
  C3 I246 (internal_0n[4], wacks_0n[30], wacks_0n[29], wacks_0n[28]);
  C3 I247 (internal_0n[5], wacks_0n[27], wacks_0n[26], wacks_0n[25]);
  C3 I248 (internal_0n[6], wacks_0n[24], wacks_0n[23], wacks_0n[22]);
  C3 I249 (internal_0n[7], wacks_0n[21], wacks_0n[20], wacks_0n[19]);
  C3 I250 (internal_0n[8], wacks_0n[18], wacks_0n[17], wacks_0n[16]);
  C3 I251 (internal_0n[9], wacks_0n[15], wacks_0n[14], wacks_0n[13]);
  C3 I252 (internal_0n[10], wacks_0n[12], wacks_0n[11], wacks_0n[10]);
  C3 I253 (internal_0n[11], wacks_0n[9], wacks_0n[8], wacks_0n[7]);
  C3 I254 (internal_0n[12], wacks_0n[6], wacks_0n[5], wacks_0n[4]);
  C2 I255 (internal_0n[13], wacks_0n[3], wacks_0n[2]);
  C2 I256 (internal_0n[14], wacks_0n[1], wacks_0n[0]);
  C3 I257 (internal_0n[15], internal_0n[2], internal_0n[3], internal_0n[4]);
  C3 I258 (internal_0n[16], internal_0n[5], internal_0n[6], internal_0n[7]);
  C3 I259 (internal_0n[17], internal_0n[8], internal_0n[9], internal_0n[10]);
  C2 I260 (internal_0n[18], internal_0n[11], internal_0n[12]);
  C2 I261 (internal_0n[19], internal_0n[13], internal_0n[14]);
  C3 I262 (internal_0n[20], internal_0n[15], internal_0n[16], internal_0n[17]);
  C2 I263 (internal_0n[21], internal_0n[18], internal_0n[19]);
  C2 I264 (wdrint_0n, internal_0n[20], internal_0n[21]);
  assign wen_0n[35] = wc_0n;
  assign wen_0n[34] = wc_0n;
  assign wen_0n[33] = wc_0n;
  assign wen_0n[32] = wc_0n;
  assign wen_0n[31] = wc_0n;
  assign wen_0n[30] = wc_0n;
  assign wen_0n[29] = wc_0n;
  assign wen_0n[28] = wc_0n;
  assign wen_0n[27] = wc_0n;
  assign wen_0n[26] = wc_0n;
  assign wen_0n[25] = wc_0n;
  assign wen_0n[24] = wc_0n;
  assign wen_0n[23] = wc_0n;
  assign wen_0n[22] = wc_0n;
  assign wen_0n[21] = wc_0n;
  assign wen_0n[20] = wc_0n;
  assign wen_0n[19] = wc_0n;
  assign wen_0n[18] = wc_0n;
  assign wen_0n[17] = wc_0n;
  assign wen_0n[16] = wc_0n;
  assign wen_0n[15] = wc_0n;
  assign wen_0n[14] = wc_0n;
  assign wen_0n[13] = wc_0n;
  assign wen_0n[12] = wc_0n;
  assign wen_0n[11] = wc_0n;
  assign wen_0n[10] = wc_0n;
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[35] = git_0n[35];
  assign wt_0n[34] = git_0n[34];
  assign wt_0n[33] = git_0n[33];
  assign wt_0n[32] = git_0n[32];
  assign wt_0n[31] = git_0n[31];
  assign wt_0n[30] = git_0n[30];
  assign wt_0n[29] = git_0n[29];
  assign wt_0n[28] = git_0n[28];
  assign wt_0n[27] = git_0n[27];
  assign wt_0n[26] = git_0n[26];
  assign wt_0n[25] = git_0n[25];
  assign wt_0n[24] = git_0n[24];
  assign wt_0n[23] = git_0n[23];
  assign wt_0n[22] = git_0n[22];
  assign wt_0n[21] = git_0n[21];
  assign wt_0n[20] = git_0n[20];
  assign wt_0n[19] = git_0n[19];
  assign wt_0n[18] = git_0n[18];
  assign wt_0n[17] = git_0n[17];
  assign wt_0n[16] = git_0n[16];
  assign wt_0n[15] = git_0n[15];
  assign wt_0n[14] = git_0n[14];
  assign wt_0n[13] = git_0n[13];
  assign wt_0n[12] = git_0n[12];
  assign wt_0n[11] = git_0n[11];
  assign wt_0n[10] = git_0n[10];
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[35] = gif_0n[35];
  assign wf_0n[34] = gif_0n[34];
  assign wf_0n[33] = gif_0n[33];
  assign wf_0n[32] = gif_0n[32];
  assign wf_0n[31] = gif_0n[31];
  assign wf_0n[30] = gif_0n[30];
  assign wf_0n[29] = gif_0n[29];
  assign wf_0n[28] = gif_0n[28];
  assign wf_0n[27] = gif_0n[27];
  assign wf_0n[26] = gif_0n[26];
  assign wf_0n[25] = gif_0n[25];
  assign wf_0n[24] = gif_0n[24];
  assign wf_0n[23] = gif_0n[23];
  assign wf_0n[22] = gif_0n[22];
  assign wf_0n[21] = gif_0n[21];
  assign wf_0n[20] = gif_0n[20];
  assign wf_0n[19] = gif_0n[19];
  assign wf_0n[18] = gif_0n[18];
  assign wf_0n[17] = gif_0n[17];
  assign wf_0n[16] = gif_0n[16];
  assign wf_0n[15] = gif_0n[15];
  assign wf_0n[14] = gif_0n[14];
  assign wf_0n[13] = gif_0n[13];
  assign wf_0n[12] = gif_0n[12];
  assign wf_0n[11] = gif_0n[11];
  assign wf_0n[10] = gif_0n[10];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I373 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I375 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I376 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I377 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I378 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I379 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I380 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I381 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I382 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I383 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I384 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I385 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I386 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I387 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I388 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I389 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I390 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I391 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I392 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I393 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I394 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I395 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I396 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I397 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I398 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I399 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I400 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I401 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I402 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I403 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I404 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I405 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I406 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I407 (git_0n[32], wgtint_0n[32], ig_0n);
  AND2 I408 (git_0n[33], wgtint_0n[33], ig_0n);
  AND2 I409 (git_0n[34], wgtint_0n[34], ig_0n);
  AND2 I410 (git_0n[35], wgtint_0n[35], ig_0n);
  AND2 I411 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I412 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I413 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I414 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I415 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I416 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I417 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I418 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I419 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I420 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I421 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I422 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I423 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I424 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I425 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I426 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I427 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I428 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I429 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I430 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I431 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I432 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I433 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I434 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I435 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I436 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I437 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I438 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I439 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I440 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I441 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I442 (gif_0n[31], wgfint_0n[31], ig_0n);
  AND2 I443 (gif_0n[32], wgfint_0n[32], ig_0n);
  AND2 I444 (gif_0n[33], wgfint_0n[33], ig_0n);
  AND2 I445 (gif_0n[34], wgfint_0n[34], ig_0n);
  AND2 I446 (gif_0n[35], wgfint_0n[35], ig_0n);
  C3 I447 (internal_0n[22], complete1574_0n[0], complete1574_0n[1], complete1574_0n[2]);
  C3 I448 (internal_0n[23], complete1574_0n[3], complete1574_0n[4], complete1574_0n[5]);
  C3 I449 (internal_0n[24], complete1574_0n[6], complete1574_0n[7], complete1574_0n[8]);
  C3 I450 (internal_0n[25], complete1574_0n[9], complete1574_0n[10], complete1574_0n[11]);
  C3 I451 (internal_0n[26], complete1574_0n[12], complete1574_0n[13], complete1574_0n[14]);
  C3 I452 (internal_0n[27], complete1574_0n[15], complete1574_0n[16], complete1574_0n[17]);
  C3 I453 (internal_0n[28], complete1574_0n[18], complete1574_0n[19], complete1574_0n[20]);
  C3 I454 (internal_0n[29], complete1574_0n[21], complete1574_0n[22], complete1574_0n[23]);
  C3 I455 (internal_0n[30], complete1574_0n[24], complete1574_0n[25], complete1574_0n[26]);
  C3 I456 (internal_0n[31], complete1574_0n[27], complete1574_0n[28], complete1574_0n[29]);
  C3 I457 (internal_0n[32], complete1574_0n[30], complete1574_0n[31], complete1574_0n[32]);
  C3 I458 (internal_0n[33], complete1574_0n[33], complete1574_0n[34], complete1574_0n[35]);
  C3 I459 (internal_0n[34], internal_0n[22], internal_0n[23], internal_0n[24]);
  C3 I460 (internal_0n[35], internal_0n[25], internal_0n[26], internal_0n[27]);
  C3 I461 (internal_0n[36], internal_0n[28], internal_0n[29], internal_0n[30]);
  C3 I462 (internal_0n[37], internal_0n[31], internal_0n[32], internal_0n[33]);
  C2 I463 (internal_0n[38], internal_0n[34], internal_0n[35]);
  C2 I464 (internal_0n[39], internal_0n[36], internal_0n[37]);
  C2 I465 (wc_0n, internal_0n[38], internal_0n[39]);
  OR2 I466 (complete1574_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I467 (complete1574_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I468 (complete1574_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I469 (complete1574_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I470 (complete1574_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I471 (complete1574_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I472 (complete1574_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I473 (complete1574_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I474 (complete1574_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I475 (complete1574_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I476 (complete1574_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I477 (complete1574_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I478 (complete1574_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I479 (complete1574_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I480 (complete1574_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I481 (complete1574_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I482 (complete1574_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I483 (complete1574_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I484 (complete1574_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I485 (complete1574_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I486 (complete1574_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I487 (complete1574_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I488 (complete1574_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I489 (complete1574_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I490 (complete1574_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I491 (complete1574_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I492 (complete1574_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I493 (complete1574_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I494 (complete1574_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I495 (complete1574_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I496 (complete1574_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I497 (complete1574_0n[31], wgfint_0n[31], wgtint_0n[31]);
  OR2 I498 (complete1574_0n[32], wgfint_0n[32], wgtint_0n[32]);
  OR2 I499 (complete1574_0n[33], wgfint_0n[33], wgtint_0n[33]);
  OR2 I500 (complete1574_0n[34], wgfint_0n[34], wgtint_0n[34]);
  OR2 I501 (complete1574_0n[35], wgfint_0n[35], wgtint_0n[35]);
  AO22 I502 (wacks_0n[35], gf1572_0n[35], df_0n[35], gt1573_0n[35], dt_0n[35]);
  NOR2 I503 (dt_0n[35], df_0n[35], gf1572_0n[35]);
  NOR3 I504 (df_0n[35], dt_0n[35], gt1573_0n[35], init_0n);
  AND2 I505 (gt1573_0n[35], wt_0n[35], wen_0n[35]);
  AND2 I506 (gf1572_0n[35], wf_0n[35], wen_0n[35]);
  AO22 I507 (wacks_0n[34], gf1572_0n[34], df_0n[34], gt1573_0n[34], dt_0n[34]);
  NOR2 I508 (dt_0n[34], df_0n[34], gf1572_0n[34]);
  NOR3 I509 (df_0n[34], dt_0n[34], gt1573_0n[34], init_0n);
  AND2 I510 (gt1573_0n[34], wt_0n[34], wen_0n[34]);
  AND2 I511 (gf1572_0n[34], wf_0n[34], wen_0n[34]);
  AO22 I512 (wacks_0n[33], gf1572_0n[33], df_0n[33], gt1573_0n[33], dt_0n[33]);
  NOR2 I513 (dt_0n[33], df_0n[33], gf1572_0n[33]);
  NOR3 I514 (df_0n[33], dt_0n[33], gt1573_0n[33], init_0n);
  AND2 I515 (gt1573_0n[33], wt_0n[33], wen_0n[33]);
  AND2 I516 (gf1572_0n[33], wf_0n[33], wen_0n[33]);
  AO22 I517 (wacks_0n[32], gf1572_0n[32], df_0n[32], gt1573_0n[32], dt_0n[32]);
  NOR2 I518 (dt_0n[32], df_0n[32], gf1572_0n[32]);
  NOR3 I519 (df_0n[32], dt_0n[32], gt1573_0n[32], init_0n);
  AND2 I520 (gt1573_0n[32], wt_0n[32], wen_0n[32]);
  AND2 I521 (gf1572_0n[32], wf_0n[32], wen_0n[32]);
  AO22 I522 (wacks_0n[31], gf1572_0n[31], df_0n[31], gt1573_0n[31], dt_0n[31]);
  NOR2 I523 (dt_0n[31], df_0n[31], gf1572_0n[31]);
  NOR3 I524 (df_0n[31], dt_0n[31], gt1573_0n[31], init_0n);
  AND2 I525 (gt1573_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I526 (gf1572_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I527 (wacks_0n[30], gf1572_0n[30], df_0n[30], gt1573_0n[30], dt_0n[30]);
  NOR2 I528 (dt_0n[30], df_0n[30], gf1572_0n[30]);
  NOR3 I529 (df_0n[30], dt_0n[30], gt1573_0n[30], init_0n);
  AND2 I530 (gt1573_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I531 (gf1572_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I532 (wacks_0n[29], gf1572_0n[29], df_0n[29], gt1573_0n[29], dt_0n[29]);
  NOR2 I533 (dt_0n[29], df_0n[29], gf1572_0n[29]);
  NOR3 I534 (df_0n[29], dt_0n[29], gt1573_0n[29], init_0n);
  AND2 I535 (gt1573_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I536 (gf1572_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I537 (wacks_0n[28], gf1572_0n[28], df_0n[28], gt1573_0n[28], dt_0n[28]);
  NOR2 I538 (dt_0n[28], df_0n[28], gf1572_0n[28]);
  NOR3 I539 (df_0n[28], dt_0n[28], gt1573_0n[28], init_0n);
  AND2 I540 (gt1573_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I541 (gf1572_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I542 (wacks_0n[27], gf1572_0n[27], df_0n[27], gt1573_0n[27], dt_0n[27]);
  NOR2 I543 (dt_0n[27], df_0n[27], gf1572_0n[27]);
  NOR3 I544 (df_0n[27], dt_0n[27], gt1573_0n[27], init_0n);
  AND2 I545 (gt1573_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I546 (gf1572_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I547 (wacks_0n[26], gf1572_0n[26], df_0n[26], gt1573_0n[26], dt_0n[26]);
  NOR2 I548 (dt_0n[26], df_0n[26], gf1572_0n[26]);
  NOR3 I549 (df_0n[26], dt_0n[26], gt1573_0n[26], init_0n);
  AND2 I550 (gt1573_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I551 (gf1572_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I552 (wacks_0n[25], gf1572_0n[25], df_0n[25], gt1573_0n[25], dt_0n[25]);
  NOR2 I553 (dt_0n[25], df_0n[25], gf1572_0n[25]);
  NOR3 I554 (df_0n[25], dt_0n[25], gt1573_0n[25], init_0n);
  AND2 I555 (gt1573_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I556 (gf1572_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I557 (wacks_0n[24], gf1572_0n[24], df_0n[24], gt1573_0n[24], dt_0n[24]);
  NOR2 I558 (dt_0n[24], df_0n[24], gf1572_0n[24]);
  NOR3 I559 (df_0n[24], dt_0n[24], gt1573_0n[24], init_0n);
  AND2 I560 (gt1573_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I561 (gf1572_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I562 (wacks_0n[23], gf1572_0n[23], df_0n[23], gt1573_0n[23], dt_0n[23]);
  NOR2 I563 (dt_0n[23], df_0n[23], gf1572_0n[23]);
  NOR3 I564 (df_0n[23], dt_0n[23], gt1573_0n[23], init_0n);
  AND2 I565 (gt1573_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I566 (gf1572_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I567 (wacks_0n[22], gf1572_0n[22], df_0n[22], gt1573_0n[22], dt_0n[22]);
  NOR2 I568 (dt_0n[22], df_0n[22], gf1572_0n[22]);
  NOR3 I569 (df_0n[22], dt_0n[22], gt1573_0n[22], init_0n);
  AND2 I570 (gt1573_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I571 (gf1572_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I572 (wacks_0n[21], gf1572_0n[21], df_0n[21], gt1573_0n[21], dt_0n[21]);
  NOR2 I573 (dt_0n[21], df_0n[21], gf1572_0n[21]);
  NOR3 I574 (df_0n[21], dt_0n[21], gt1573_0n[21], init_0n);
  AND2 I575 (gt1573_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I576 (gf1572_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I577 (wacks_0n[20], gf1572_0n[20], df_0n[20], gt1573_0n[20], dt_0n[20]);
  NOR2 I578 (dt_0n[20], df_0n[20], gf1572_0n[20]);
  NOR3 I579 (df_0n[20], dt_0n[20], gt1573_0n[20], init_0n);
  AND2 I580 (gt1573_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I581 (gf1572_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I582 (wacks_0n[19], gf1572_0n[19], df_0n[19], gt1573_0n[19], dt_0n[19]);
  NOR2 I583 (dt_0n[19], df_0n[19], gf1572_0n[19]);
  NOR3 I584 (df_0n[19], dt_0n[19], gt1573_0n[19], init_0n);
  AND2 I585 (gt1573_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I586 (gf1572_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I587 (wacks_0n[18], gf1572_0n[18], df_0n[18], gt1573_0n[18], dt_0n[18]);
  NOR2 I588 (dt_0n[18], df_0n[18], gf1572_0n[18]);
  NOR3 I589 (df_0n[18], dt_0n[18], gt1573_0n[18], init_0n);
  AND2 I590 (gt1573_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I591 (gf1572_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I592 (wacks_0n[17], gf1572_0n[17], df_0n[17], gt1573_0n[17], dt_0n[17]);
  NOR2 I593 (dt_0n[17], df_0n[17], gf1572_0n[17]);
  NOR3 I594 (df_0n[17], dt_0n[17], gt1573_0n[17], init_0n);
  AND2 I595 (gt1573_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I596 (gf1572_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I597 (wacks_0n[16], gf1572_0n[16], df_0n[16], gt1573_0n[16], dt_0n[16]);
  NOR2 I598 (dt_0n[16], df_0n[16], gf1572_0n[16]);
  NOR3 I599 (df_0n[16], dt_0n[16], gt1573_0n[16], init_0n);
  AND2 I600 (gt1573_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I601 (gf1572_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I602 (wacks_0n[15], gf1572_0n[15], df_0n[15], gt1573_0n[15], dt_0n[15]);
  NOR2 I603 (dt_0n[15], df_0n[15], gf1572_0n[15]);
  NOR3 I604 (df_0n[15], dt_0n[15], gt1573_0n[15], init_0n);
  AND2 I605 (gt1573_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I606 (gf1572_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I607 (wacks_0n[14], gf1572_0n[14], df_0n[14], gt1573_0n[14], dt_0n[14]);
  NOR2 I608 (dt_0n[14], df_0n[14], gf1572_0n[14]);
  NOR3 I609 (df_0n[14], dt_0n[14], gt1573_0n[14], init_0n);
  AND2 I610 (gt1573_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I611 (gf1572_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I612 (wacks_0n[13], gf1572_0n[13], df_0n[13], gt1573_0n[13], dt_0n[13]);
  NOR2 I613 (dt_0n[13], df_0n[13], gf1572_0n[13]);
  NOR3 I614 (df_0n[13], dt_0n[13], gt1573_0n[13], init_0n);
  AND2 I615 (gt1573_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I616 (gf1572_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I617 (wacks_0n[12], gf1572_0n[12], df_0n[12], gt1573_0n[12], dt_0n[12]);
  NOR2 I618 (dt_0n[12], df_0n[12], gf1572_0n[12]);
  NOR3 I619 (df_0n[12], dt_0n[12], gt1573_0n[12], init_0n);
  AND2 I620 (gt1573_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I621 (gf1572_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I622 (wacks_0n[11], gf1572_0n[11], df_0n[11], gt1573_0n[11], dt_0n[11]);
  NOR2 I623 (dt_0n[11], df_0n[11], gf1572_0n[11]);
  NOR3 I624 (df_0n[11], dt_0n[11], gt1573_0n[11], init_0n);
  AND2 I625 (gt1573_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I626 (gf1572_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I627 (wacks_0n[10], gf1572_0n[10], df_0n[10], gt1573_0n[10], dt_0n[10]);
  NOR2 I628 (dt_0n[10], df_0n[10], gf1572_0n[10]);
  NOR3 I629 (df_0n[10], dt_0n[10], gt1573_0n[10], init_0n);
  AND2 I630 (gt1573_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I631 (gf1572_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I632 (wacks_0n[9], gf1572_0n[9], df_0n[9], gt1573_0n[9], dt_0n[9]);
  NOR2 I633 (dt_0n[9], df_0n[9], gf1572_0n[9]);
  NOR3 I634 (df_0n[9], dt_0n[9], gt1573_0n[9], init_0n);
  AND2 I635 (gt1573_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I636 (gf1572_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I637 (wacks_0n[8], gf1572_0n[8], df_0n[8], gt1573_0n[8], dt_0n[8]);
  NOR2 I638 (dt_0n[8], df_0n[8], gf1572_0n[8]);
  NOR3 I639 (df_0n[8], dt_0n[8], gt1573_0n[8], init_0n);
  AND2 I640 (gt1573_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I641 (gf1572_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I642 (wacks_0n[7], gf1572_0n[7], df_0n[7], gt1573_0n[7], dt_0n[7]);
  NOR2 I643 (dt_0n[7], df_0n[7], gf1572_0n[7]);
  NOR3 I644 (df_0n[7], dt_0n[7], gt1573_0n[7], init_0n);
  AND2 I645 (gt1573_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I646 (gf1572_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I647 (wacks_0n[6], gf1572_0n[6], df_0n[6], gt1573_0n[6], dt_0n[6]);
  NOR2 I648 (dt_0n[6], df_0n[6], gf1572_0n[6]);
  NOR3 I649 (df_0n[6], dt_0n[6], gt1573_0n[6], init_0n);
  AND2 I650 (gt1573_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I651 (gf1572_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I652 (wacks_0n[5], gf1572_0n[5], df_0n[5], gt1573_0n[5], dt_0n[5]);
  NOR2 I653 (dt_0n[5], df_0n[5], gf1572_0n[5]);
  NOR3 I654 (df_0n[5], dt_0n[5], gt1573_0n[5], init_0n);
  AND2 I655 (gt1573_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I656 (gf1572_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I657 (wacks_0n[4], gf1572_0n[4], df_0n[4], gt1573_0n[4], dt_0n[4]);
  NOR2 I658 (dt_0n[4], df_0n[4], gf1572_0n[4]);
  NOR3 I659 (df_0n[4], dt_0n[4], gt1573_0n[4], init_0n);
  AND2 I660 (gt1573_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I661 (gf1572_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I662 (wacks_0n[3], gf1572_0n[3], df_0n[3], gt1573_0n[3], dt_0n[3]);
  NOR2 I663 (dt_0n[3], df_0n[3], gf1572_0n[3]);
  NOR3 I664 (df_0n[3], dt_0n[3], gt1573_0n[3], init_0n);
  AND2 I665 (gt1573_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I666 (gf1572_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I667 (wacks_0n[2], gf1572_0n[2], df_0n[2], gt1573_0n[2], dt_0n[2]);
  NOR2 I668 (dt_0n[2], df_0n[2], gf1572_0n[2]);
  NOR3 I669 (df_0n[2], dt_0n[2], gt1573_0n[2], init_0n);
  AND2 I670 (gt1573_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I671 (gf1572_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I672 (wacks_0n[1], gf1572_0n[1], df_0n[1], gt1573_0n[1], dt_0n[1]);
  NOR2 I673 (dt_0n[1], df_0n[1], gf1572_0n[1]);
  NOR3 I674 (df_0n[1], dt_0n[1], gt1573_0n[1], init_0n);
  AND2 I675 (gt1573_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I676 (gf1572_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I677 (wacks_0n[0], gf1572_0n[0], df_0n[0], gt1573_0n[0], dt_0n[0]);
  NOR2 I678 (dt_0n[0], df_0n[0], gf1572_0n[0]);
  NOR3 I679 (df_0n[0], dt_0n[0], gt1573_0n[0], init_0n);
  AND2 I680 (gt1573_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I681 (gf1572_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I682 (init_0n, initialise);
endmodule

module BrzV_36_l6__28_29_l24__28_28_280_2036_29_2_m96m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  initialise
);
  input [35:0] wg_0r0d;
  input [35:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [31:0] rd_0r0d;
  output [31:0] rd_0r1d;
  input rd_0a;
  output [35:0] rd_1r0d;
  output [35:0] rd_1r1d;
  input rd_1a;
  input initialise;
  wire [39:0] internal_0n;
  wire [35:0] wf_0n;
  wire [35:0] wt_0n;
  wire [35:0] df_0n;
  wire [35:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire wc_0n;
  wire [35:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [35:0] wgfint_0n;
  wire [35:0] wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire [31:0] rdfint_0n;
  wire [35:0] rdfint_1n;
  wire [31:0] rdtint_0n;
  wire [35:0] rdtint_1n;
  wire [35:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [35:0] gif_0n;
  wire [35:0] git_0n;
  wire [35:0] complete1589_0n;
  wire [35:0] gt1588_0n;
  wire [35:0] gf1587_0n;
  assign rgaint_1n = rd_1a;
  assign rd_1r0d[0] = rdfint_1n[0];
  assign rd_1r0d[1] = rdfint_1n[1];
  assign rd_1r0d[2] = rdfint_1n[2];
  assign rd_1r0d[3] = rdfint_1n[3];
  assign rd_1r0d[4] = rdfint_1n[4];
  assign rd_1r0d[5] = rdfint_1n[5];
  assign rd_1r0d[6] = rdfint_1n[6];
  assign rd_1r0d[7] = rdfint_1n[7];
  assign rd_1r0d[8] = rdfint_1n[8];
  assign rd_1r0d[9] = rdfint_1n[9];
  assign rd_1r0d[10] = rdfint_1n[10];
  assign rd_1r0d[11] = rdfint_1n[11];
  assign rd_1r0d[12] = rdfint_1n[12];
  assign rd_1r0d[13] = rdfint_1n[13];
  assign rd_1r0d[14] = rdfint_1n[14];
  assign rd_1r0d[15] = rdfint_1n[15];
  assign rd_1r0d[16] = rdfint_1n[16];
  assign rd_1r0d[17] = rdfint_1n[17];
  assign rd_1r0d[18] = rdfint_1n[18];
  assign rd_1r0d[19] = rdfint_1n[19];
  assign rd_1r0d[20] = rdfint_1n[20];
  assign rd_1r0d[21] = rdfint_1n[21];
  assign rd_1r0d[22] = rdfint_1n[22];
  assign rd_1r0d[23] = rdfint_1n[23];
  assign rd_1r0d[24] = rdfint_1n[24];
  assign rd_1r0d[25] = rdfint_1n[25];
  assign rd_1r0d[26] = rdfint_1n[26];
  assign rd_1r0d[27] = rdfint_1n[27];
  assign rd_1r0d[28] = rdfint_1n[28];
  assign rd_1r0d[29] = rdfint_1n[29];
  assign rd_1r0d[30] = rdfint_1n[30];
  assign rd_1r0d[31] = rdfint_1n[31];
  assign rd_1r0d[32] = rdfint_1n[32];
  assign rd_1r0d[33] = rdfint_1n[33];
  assign rd_1r0d[34] = rdfint_1n[34];
  assign rd_1r0d[35] = rdfint_1n[35];
  assign rd_1r1d[0] = rdtint_1n[0];
  assign rd_1r1d[1] = rdtint_1n[1];
  assign rd_1r1d[2] = rdtint_1n[2];
  assign rd_1r1d[3] = rdtint_1n[3];
  assign rd_1r1d[4] = rdtint_1n[4];
  assign rd_1r1d[5] = rdtint_1n[5];
  assign rd_1r1d[6] = rdtint_1n[6];
  assign rd_1r1d[7] = rdtint_1n[7];
  assign rd_1r1d[8] = rdtint_1n[8];
  assign rd_1r1d[9] = rdtint_1n[9];
  assign rd_1r1d[10] = rdtint_1n[10];
  assign rd_1r1d[11] = rdtint_1n[11];
  assign rd_1r1d[12] = rdtint_1n[12];
  assign rd_1r1d[13] = rdtint_1n[13];
  assign rd_1r1d[14] = rdtint_1n[14];
  assign rd_1r1d[15] = rdtint_1n[15];
  assign rd_1r1d[16] = rdtint_1n[16];
  assign rd_1r1d[17] = rdtint_1n[17];
  assign rd_1r1d[18] = rdtint_1n[18];
  assign rd_1r1d[19] = rdtint_1n[19];
  assign rd_1r1d[20] = rdtint_1n[20];
  assign rd_1r1d[21] = rdtint_1n[21];
  assign rd_1r1d[22] = rdtint_1n[22];
  assign rd_1r1d[23] = rdtint_1n[23];
  assign rd_1r1d[24] = rdtint_1n[24];
  assign rd_1r1d[25] = rdtint_1n[25];
  assign rd_1r1d[26] = rdtint_1n[26];
  assign rd_1r1d[27] = rdtint_1n[27];
  assign rd_1r1d[28] = rdtint_1n[28];
  assign rd_1r1d[29] = rdtint_1n[29];
  assign rd_1r1d[30] = rdtint_1n[30];
  assign rd_1r1d[31] = rdtint_1n[31];
  assign rd_1r1d[32] = rdtint_1n[32];
  assign rd_1r1d[33] = rdtint_1n[33];
  assign rd_1r1d[34] = rdtint_1n[34];
  assign rd_1r1d[35] = rdtint_1n[35];
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r0d[10] = rdfint_0n[10];
  assign rd_0r0d[11] = rdfint_0n[11];
  assign rd_0r0d[12] = rdfint_0n[12];
  assign rd_0r0d[13] = rdfint_0n[13];
  assign rd_0r0d[14] = rdfint_0n[14];
  assign rd_0r0d[15] = rdfint_0n[15];
  assign rd_0r0d[16] = rdfint_0n[16];
  assign rd_0r0d[17] = rdfint_0n[17];
  assign rd_0r0d[18] = rdfint_0n[18];
  assign rd_0r0d[19] = rdfint_0n[19];
  assign rd_0r0d[20] = rdfint_0n[20];
  assign rd_0r0d[21] = rdfint_0n[21];
  assign rd_0r0d[22] = rdfint_0n[22];
  assign rd_0r0d[23] = rdfint_0n[23];
  assign rd_0r0d[24] = rdfint_0n[24];
  assign rd_0r0d[25] = rdfint_0n[25];
  assign rd_0r0d[26] = rdfint_0n[26];
  assign rd_0r0d[27] = rdfint_0n[27];
  assign rd_0r0d[28] = rdfint_0n[28];
  assign rd_0r0d[29] = rdfint_0n[29];
  assign rd_0r0d[30] = rdfint_0n[30];
  assign rd_0r0d[31] = rdfint_0n[31];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign rd_0r1d[10] = rdtint_0n[10];
  assign rd_0r1d[11] = rdtint_0n[11];
  assign rd_0r1d[12] = rdtint_0n[12];
  assign rd_0r1d[13] = rdtint_0n[13];
  assign rd_0r1d[14] = rdtint_0n[14];
  assign rd_0r1d[15] = rdtint_0n[15];
  assign rd_0r1d[16] = rdtint_0n[16];
  assign rd_0r1d[17] = rdtint_0n[17];
  assign rd_0r1d[18] = rdtint_0n[18];
  assign rd_0r1d[19] = rdtint_0n[19];
  assign rd_0r1d[20] = rdtint_0n[20];
  assign rd_0r1d[21] = rdtint_0n[21];
  assign rd_0r1d[22] = rdtint_0n[22];
  assign rd_0r1d[23] = rdtint_0n[23];
  assign rd_0r1d[24] = rdtint_0n[24];
  assign rd_0r1d[25] = rdtint_0n[25];
  assign rd_0r1d[26] = rdtint_0n[26];
  assign rd_0r1d[27] = rdtint_0n[27];
  assign rd_0r1d[28] = rdtint_0n[28];
  assign rd_0r1d[29] = rdtint_0n[29];
  assign rd_0r1d[30] = rdtint_0n[30];
  assign rd_0r1d[31] = rdtint_0n[31];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgfint_0n[32] = wg_0r0d[32];
  assign wgfint_0n[33] = wg_0r0d[33];
  assign wgfint_0n[34] = wg_0r0d[34];
  assign wgfint_0n[35] = wg_0r0d[35];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign wgtint_0n[32] = wg_0r1d[32];
  assign wgtint_0n[33] = wg_0r1d[33];
  assign wgtint_0n[34] = wg_0r1d[34];
  assign wgtint_0n[35] = wg_0r1d[35];
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I217 (internal_0n[0], rgrint_0n, rgrint_1n);
  NOR2 I218 (internal_0n[1], rgaint_0n, rgaint_1n);
  AND2 I219 (nanyread_0n, internal_0n[0], internal_0n[1]);
  AND2 I220 (rdtint_1n[0], rgrint_1n, dt_0n[0]);
  AND2 I221 (rdtint_1n[1], rgrint_1n, dt_0n[1]);
  AND2 I222 (rdtint_1n[2], rgrint_1n, dt_0n[2]);
  AND2 I223 (rdtint_1n[3], rgrint_1n, dt_0n[3]);
  AND2 I224 (rdtint_1n[4], rgrint_1n, dt_0n[4]);
  AND2 I225 (rdtint_1n[5], rgrint_1n, dt_0n[5]);
  AND2 I226 (rdtint_1n[6], rgrint_1n, dt_0n[6]);
  AND2 I227 (rdtint_1n[7], rgrint_1n, dt_0n[7]);
  AND2 I228 (rdtint_1n[8], rgrint_1n, dt_0n[8]);
  AND2 I229 (rdtint_1n[9], rgrint_1n, dt_0n[9]);
  AND2 I230 (rdtint_1n[10], rgrint_1n, dt_0n[10]);
  AND2 I231 (rdtint_1n[11], rgrint_1n, dt_0n[11]);
  AND2 I232 (rdtint_1n[12], rgrint_1n, dt_0n[12]);
  AND2 I233 (rdtint_1n[13], rgrint_1n, dt_0n[13]);
  AND2 I234 (rdtint_1n[14], rgrint_1n, dt_0n[14]);
  AND2 I235 (rdtint_1n[15], rgrint_1n, dt_0n[15]);
  AND2 I236 (rdtint_1n[16], rgrint_1n, dt_0n[16]);
  AND2 I237 (rdtint_1n[17], rgrint_1n, dt_0n[17]);
  AND2 I238 (rdtint_1n[18], rgrint_1n, dt_0n[18]);
  AND2 I239 (rdtint_1n[19], rgrint_1n, dt_0n[19]);
  AND2 I240 (rdtint_1n[20], rgrint_1n, dt_0n[20]);
  AND2 I241 (rdtint_1n[21], rgrint_1n, dt_0n[21]);
  AND2 I242 (rdtint_1n[22], rgrint_1n, dt_0n[22]);
  AND2 I243 (rdtint_1n[23], rgrint_1n, dt_0n[23]);
  AND2 I244 (rdtint_1n[24], rgrint_1n, dt_0n[24]);
  AND2 I245 (rdtint_1n[25], rgrint_1n, dt_0n[25]);
  AND2 I246 (rdtint_1n[26], rgrint_1n, dt_0n[26]);
  AND2 I247 (rdtint_1n[27], rgrint_1n, dt_0n[27]);
  AND2 I248 (rdtint_1n[28], rgrint_1n, dt_0n[28]);
  AND2 I249 (rdtint_1n[29], rgrint_1n, dt_0n[29]);
  AND2 I250 (rdtint_1n[30], rgrint_1n, dt_0n[30]);
  AND2 I251 (rdtint_1n[31], rgrint_1n, dt_0n[31]);
  AND2 I252 (rdtint_1n[32], rgrint_1n, dt_0n[32]);
  AND2 I253 (rdtint_1n[33], rgrint_1n, dt_0n[33]);
  AND2 I254 (rdtint_1n[34], rgrint_1n, dt_0n[34]);
  AND2 I255 (rdtint_1n[35], rgrint_1n, dt_0n[35]);
  AND2 I256 (rdtint_0n[0], rgrint_0n, dt_0n[2]);
  AND2 I257 (rdtint_0n[1], rgrint_0n, dt_0n[3]);
  AND2 I258 (rdtint_0n[2], rgrint_0n, dt_0n[4]);
  AND2 I259 (rdtint_0n[3], rgrint_0n, dt_0n[5]);
  AND2 I260 (rdtint_0n[4], rgrint_0n, dt_0n[6]);
  AND2 I261 (rdtint_0n[5], rgrint_0n, dt_0n[7]);
  AND2 I262 (rdtint_0n[6], rgrint_0n, dt_0n[8]);
  AND2 I263 (rdtint_0n[7], rgrint_0n, dt_0n[9]);
  AND2 I264 (rdtint_0n[8], rgrint_0n, dt_0n[10]);
  AND2 I265 (rdtint_0n[9], rgrint_0n, dt_0n[11]);
  AND2 I266 (rdtint_0n[10], rgrint_0n, dt_0n[12]);
  AND2 I267 (rdtint_0n[11], rgrint_0n, dt_0n[13]);
  AND2 I268 (rdtint_0n[12], rgrint_0n, dt_0n[14]);
  AND2 I269 (rdtint_0n[13], rgrint_0n, dt_0n[15]);
  AND2 I270 (rdtint_0n[14], rgrint_0n, dt_0n[16]);
  AND2 I271 (rdtint_0n[15], rgrint_0n, dt_0n[17]);
  AND2 I272 (rdtint_0n[16], rgrint_0n, dt_0n[18]);
  AND2 I273 (rdtint_0n[17], rgrint_0n, dt_0n[19]);
  AND2 I274 (rdtint_0n[18], rgrint_0n, dt_0n[20]);
  AND2 I275 (rdtint_0n[19], rgrint_0n, dt_0n[21]);
  AND2 I276 (rdtint_0n[20], rgrint_0n, dt_0n[22]);
  AND2 I277 (rdtint_0n[21], rgrint_0n, dt_0n[23]);
  AND2 I278 (rdtint_0n[22], rgrint_0n, dt_0n[24]);
  AND2 I279 (rdtint_0n[23], rgrint_0n, dt_0n[25]);
  AND2 I280 (rdtint_0n[24], rgrint_0n, dt_0n[26]);
  AND2 I281 (rdtint_0n[25], rgrint_0n, dt_0n[27]);
  AND2 I282 (rdtint_0n[26], rgrint_0n, dt_0n[28]);
  AND2 I283 (rdtint_0n[27], rgrint_0n, dt_0n[29]);
  AND2 I284 (rdtint_0n[28], rgrint_0n, dt_0n[30]);
  AND2 I285 (rdtint_0n[29], rgrint_0n, dt_0n[31]);
  AND2 I286 (rdtint_0n[30], rgrint_0n, dt_0n[32]);
  AND2 I287 (rdtint_0n[31], rgrint_0n, dt_0n[33]);
  AND2 I288 (rdfint_1n[0], rgrint_1n, df_0n[0]);
  AND2 I289 (rdfint_1n[1], rgrint_1n, df_0n[1]);
  AND2 I290 (rdfint_1n[2], rgrint_1n, df_0n[2]);
  AND2 I291 (rdfint_1n[3], rgrint_1n, df_0n[3]);
  AND2 I292 (rdfint_1n[4], rgrint_1n, df_0n[4]);
  AND2 I293 (rdfint_1n[5], rgrint_1n, df_0n[5]);
  AND2 I294 (rdfint_1n[6], rgrint_1n, df_0n[6]);
  AND2 I295 (rdfint_1n[7], rgrint_1n, df_0n[7]);
  AND2 I296 (rdfint_1n[8], rgrint_1n, df_0n[8]);
  AND2 I297 (rdfint_1n[9], rgrint_1n, df_0n[9]);
  AND2 I298 (rdfint_1n[10], rgrint_1n, df_0n[10]);
  AND2 I299 (rdfint_1n[11], rgrint_1n, df_0n[11]);
  AND2 I300 (rdfint_1n[12], rgrint_1n, df_0n[12]);
  AND2 I301 (rdfint_1n[13], rgrint_1n, df_0n[13]);
  AND2 I302 (rdfint_1n[14], rgrint_1n, df_0n[14]);
  AND2 I303 (rdfint_1n[15], rgrint_1n, df_0n[15]);
  AND2 I304 (rdfint_1n[16], rgrint_1n, df_0n[16]);
  AND2 I305 (rdfint_1n[17], rgrint_1n, df_0n[17]);
  AND2 I306 (rdfint_1n[18], rgrint_1n, df_0n[18]);
  AND2 I307 (rdfint_1n[19], rgrint_1n, df_0n[19]);
  AND2 I308 (rdfint_1n[20], rgrint_1n, df_0n[20]);
  AND2 I309 (rdfint_1n[21], rgrint_1n, df_0n[21]);
  AND2 I310 (rdfint_1n[22], rgrint_1n, df_0n[22]);
  AND2 I311 (rdfint_1n[23], rgrint_1n, df_0n[23]);
  AND2 I312 (rdfint_1n[24], rgrint_1n, df_0n[24]);
  AND2 I313 (rdfint_1n[25], rgrint_1n, df_0n[25]);
  AND2 I314 (rdfint_1n[26], rgrint_1n, df_0n[26]);
  AND2 I315 (rdfint_1n[27], rgrint_1n, df_0n[27]);
  AND2 I316 (rdfint_1n[28], rgrint_1n, df_0n[28]);
  AND2 I317 (rdfint_1n[29], rgrint_1n, df_0n[29]);
  AND2 I318 (rdfint_1n[30], rgrint_1n, df_0n[30]);
  AND2 I319 (rdfint_1n[31], rgrint_1n, df_0n[31]);
  AND2 I320 (rdfint_1n[32], rgrint_1n, df_0n[32]);
  AND2 I321 (rdfint_1n[33], rgrint_1n, df_0n[33]);
  AND2 I322 (rdfint_1n[34], rgrint_1n, df_0n[34]);
  AND2 I323 (rdfint_1n[35], rgrint_1n, df_0n[35]);
  AND2 I324 (rdfint_0n[0], rgrint_0n, df_0n[2]);
  AND2 I325 (rdfint_0n[1], rgrint_0n, df_0n[3]);
  AND2 I326 (rdfint_0n[2], rgrint_0n, df_0n[4]);
  AND2 I327 (rdfint_0n[3], rgrint_0n, df_0n[5]);
  AND2 I328 (rdfint_0n[4], rgrint_0n, df_0n[6]);
  AND2 I329 (rdfint_0n[5], rgrint_0n, df_0n[7]);
  AND2 I330 (rdfint_0n[6], rgrint_0n, df_0n[8]);
  AND2 I331 (rdfint_0n[7], rgrint_0n, df_0n[9]);
  AND2 I332 (rdfint_0n[8], rgrint_0n, df_0n[10]);
  AND2 I333 (rdfint_0n[9], rgrint_0n, df_0n[11]);
  AND2 I334 (rdfint_0n[10], rgrint_0n, df_0n[12]);
  AND2 I335 (rdfint_0n[11], rgrint_0n, df_0n[13]);
  AND2 I336 (rdfint_0n[12], rgrint_0n, df_0n[14]);
  AND2 I337 (rdfint_0n[13], rgrint_0n, df_0n[15]);
  AND2 I338 (rdfint_0n[14], rgrint_0n, df_0n[16]);
  AND2 I339 (rdfint_0n[15], rgrint_0n, df_0n[17]);
  AND2 I340 (rdfint_0n[16], rgrint_0n, df_0n[18]);
  AND2 I341 (rdfint_0n[17], rgrint_0n, df_0n[19]);
  AND2 I342 (rdfint_0n[18], rgrint_0n, df_0n[20]);
  AND2 I343 (rdfint_0n[19], rgrint_0n, df_0n[21]);
  AND2 I344 (rdfint_0n[20], rgrint_0n, df_0n[22]);
  AND2 I345 (rdfint_0n[21], rgrint_0n, df_0n[23]);
  AND2 I346 (rdfint_0n[22], rgrint_0n, df_0n[24]);
  AND2 I347 (rdfint_0n[23], rgrint_0n, df_0n[25]);
  AND2 I348 (rdfint_0n[24], rgrint_0n, df_0n[26]);
  AND2 I349 (rdfint_0n[25], rgrint_0n, df_0n[27]);
  AND2 I350 (rdfint_0n[26], rgrint_0n, df_0n[28]);
  AND2 I351 (rdfint_0n[27], rgrint_0n, df_0n[29]);
  AND2 I352 (rdfint_0n[28], rgrint_0n, df_0n[30]);
  AND2 I353 (rdfint_0n[29], rgrint_0n, df_0n[31]);
  AND2 I354 (rdfint_0n[30], rgrint_0n, df_0n[32]);
  AND2 I355 (rdfint_0n[31], rgrint_0n, df_0n[33]);
  C3 I356 (internal_0n[2], wc_0n, wacks_0n[35], wacks_0n[34]);
  C3 I357 (internal_0n[3], wacks_0n[33], wacks_0n[32], wacks_0n[31]);
  C3 I358 (internal_0n[4], wacks_0n[30], wacks_0n[29], wacks_0n[28]);
  C3 I359 (internal_0n[5], wacks_0n[27], wacks_0n[26], wacks_0n[25]);
  C3 I360 (internal_0n[6], wacks_0n[24], wacks_0n[23], wacks_0n[22]);
  C3 I361 (internal_0n[7], wacks_0n[21], wacks_0n[20], wacks_0n[19]);
  C3 I362 (internal_0n[8], wacks_0n[18], wacks_0n[17], wacks_0n[16]);
  C3 I363 (internal_0n[9], wacks_0n[15], wacks_0n[14], wacks_0n[13]);
  C3 I364 (internal_0n[10], wacks_0n[12], wacks_0n[11], wacks_0n[10]);
  C3 I365 (internal_0n[11], wacks_0n[9], wacks_0n[8], wacks_0n[7]);
  C3 I366 (internal_0n[12], wacks_0n[6], wacks_0n[5], wacks_0n[4]);
  C2 I367 (internal_0n[13], wacks_0n[3], wacks_0n[2]);
  C2 I368 (internal_0n[14], wacks_0n[1], wacks_0n[0]);
  C3 I369 (internal_0n[15], internal_0n[2], internal_0n[3], internal_0n[4]);
  C3 I370 (internal_0n[16], internal_0n[5], internal_0n[6], internal_0n[7]);
  C3 I371 (internal_0n[17], internal_0n[8], internal_0n[9], internal_0n[10]);
  C2 I372 (internal_0n[18], internal_0n[11], internal_0n[12]);
  C2 I373 (internal_0n[19], internal_0n[13], internal_0n[14]);
  C3 I374 (internal_0n[20], internal_0n[15], internal_0n[16], internal_0n[17]);
  C2 I375 (internal_0n[21], internal_0n[18], internal_0n[19]);
  C2 I376 (wdrint_0n, internal_0n[20], internal_0n[21]);
  assign wen_0n[35] = wc_0n;
  assign wen_0n[34] = wc_0n;
  assign wen_0n[33] = wc_0n;
  assign wen_0n[32] = wc_0n;
  assign wen_0n[31] = wc_0n;
  assign wen_0n[30] = wc_0n;
  assign wen_0n[29] = wc_0n;
  assign wen_0n[28] = wc_0n;
  assign wen_0n[27] = wc_0n;
  assign wen_0n[26] = wc_0n;
  assign wen_0n[25] = wc_0n;
  assign wen_0n[24] = wc_0n;
  assign wen_0n[23] = wc_0n;
  assign wen_0n[22] = wc_0n;
  assign wen_0n[21] = wc_0n;
  assign wen_0n[20] = wc_0n;
  assign wen_0n[19] = wc_0n;
  assign wen_0n[18] = wc_0n;
  assign wen_0n[17] = wc_0n;
  assign wen_0n[16] = wc_0n;
  assign wen_0n[15] = wc_0n;
  assign wen_0n[14] = wc_0n;
  assign wen_0n[13] = wc_0n;
  assign wen_0n[12] = wc_0n;
  assign wen_0n[11] = wc_0n;
  assign wen_0n[10] = wc_0n;
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[35] = git_0n[35];
  assign wt_0n[34] = git_0n[34];
  assign wt_0n[33] = git_0n[33];
  assign wt_0n[32] = git_0n[32];
  assign wt_0n[31] = git_0n[31];
  assign wt_0n[30] = git_0n[30];
  assign wt_0n[29] = git_0n[29];
  assign wt_0n[28] = git_0n[28];
  assign wt_0n[27] = git_0n[27];
  assign wt_0n[26] = git_0n[26];
  assign wt_0n[25] = git_0n[25];
  assign wt_0n[24] = git_0n[24];
  assign wt_0n[23] = git_0n[23];
  assign wt_0n[22] = git_0n[22];
  assign wt_0n[21] = git_0n[21];
  assign wt_0n[20] = git_0n[20];
  assign wt_0n[19] = git_0n[19];
  assign wt_0n[18] = git_0n[18];
  assign wt_0n[17] = git_0n[17];
  assign wt_0n[16] = git_0n[16];
  assign wt_0n[15] = git_0n[15];
  assign wt_0n[14] = git_0n[14];
  assign wt_0n[13] = git_0n[13];
  assign wt_0n[12] = git_0n[12];
  assign wt_0n[11] = git_0n[11];
  assign wt_0n[10] = git_0n[10];
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[35] = gif_0n[35];
  assign wf_0n[34] = gif_0n[34];
  assign wf_0n[33] = gif_0n[33];
  assign wf_0n[32] = gif_0n[32];
  assign wf_0n[31] = gif_0n[31];
  assign wf_0n[30] = gif_0n[30];
  assign wf_0n[29] = gif_0n[29];
  assign wf_0n[28] = gif_0n[28];
  assign wf_0n[27] = gif_0n[27];
  assign wf_0n[26] = gif_0n[26];
  assign wf_0n[25] = gif_0n[25];
  assign wf_0n[24] = gif_0n[24];
  assign wf_0n[23] = gif_0n[23];
  assign wf_0n[22] = gif_0n[22];
  assign wf_0n[21] = gif_0n[21];
  assign wf_0n[20] = gif_0n[20];
  assign wf_0n[19] = gif_0n[19];
  assign wf_0n[18] = gif_0n[18];
  assign wf_0n[17] = gif_0n[17];
  assign wf_0n[16] = gif_0n[16];
  assign wf_0n[15] = gif_0n[15];
  assign wf_0n[14] = gif_0n[14];
  assign wf_0n[13] = gif_0n[13];
  assign wf_0n[12] = gif_0n[12];
  assign wf_0n[11] = gif_0n[11];
  assign wf_0n[10] = gif_0n[10];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I485 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I487 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I488 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I489 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I490 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I491 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I492 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I493 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I494 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I495 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I496 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I497 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I498 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I499 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I500 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I501 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I502 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I503 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I504 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I505 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I506 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I507 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I508 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I509 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I510 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I511 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I512 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I513 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I514 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I515 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I516 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I517 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I518 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I519 (git_0n[32], wgtint_0n[32], ig_0n);
  AND2 I520 (git_0n[33], wgtint_0n[33], ig_0n);
  AND2 I521 (git_0n[34], wgtint_0n[34], ig_0n);
  AND2 I522 (git_0n[35], wgtint_0n[35], ig_0n);
  AND2 I523 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I524 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I525 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I526 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I527 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I528 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I529 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I530 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I531 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I532 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I533 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I534 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I535 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I536 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I537 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I538 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I539 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I540 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I541 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I542 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I543 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I544 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I545 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I546 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I547 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I548 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I549 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I550 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I551 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I552 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I553 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I554 (gif_0n[31], wgfint_0n[31], ig_0n);
  AND2 I555 (gif_0n[32], wgfint_0n[32], ig_0n);
  AND2 I556 (gif_0n[33], wgfint_0n[33], ig_0n);
  AND2 I557 (gif_0n[34], wgfint_0n[34], ig_0n);
  AND2 I558 (gif_0n[35], wgfint_0n[35], ig_0n);
  C3 I559 (internal_0n[22], complete1589_0n[0], complete1589_0n[1], complete1589_0n[2]);
  C3 I560 (internal_0n[23], complete1589_0n[3], complete1589_0n[4], complete1589_0n[5]);
  C3 I561 (internal_0n[24], complete1589_0n[6], complete1589_0n[7], complete1589_0n[8]);
  C3 I562 (internal_0n[25], complete1589_0n[9], complete1589_0n[10], complete1589_0n[11]);
  C3 I563 (internal_0n[26], complete1589_0n[12], complete1589_0n[13], complete1589_0n[14]);
  C3 I564 (internal_0n[27], complete1589_0n[15], complete1589_0n[16], complete1589_0n[17]);
  C3 I565 (internal_0n[28], complete1589_0n[18], complete1589_0n[19], complete1589_0n[20]);
  C3 I566 (internal_0n[29], complete1589_0n[21], complete1589_0n[22], complete1589_0n[23]);
  C3 I567 (internal_0n[30], complete1589_0n[24], complete1589_0n[25], complete1589_0n[26]);
  C3 I568 (internal_0n[31], complete1589_0n[27], complete1589_0n[28], complete1589_0n[29]);
  C3 I569 (internal_0n[32], complete1589_0n[30], complete1589_0n[31], complete1589_0n[32]);
  C3 I570 (internal_0n[33], complete1589_0n[33], complete1589_0n[34], complete1589_0n[35]);
  C3 I571 (internal_0n[34], internal_0n[22], internal_0n[23], internal_0n[24]);
  C3 I572 (internal_0n[35], internal_0n[25], internal_0n[26], internal_0n[27]);
  C3 I573 (internal_0n[36], internal_0n[28], internal_0n[29], internal_0n[30]);
  C3 I574 (internal_0n[37], internal_0n[31], internal_0n[32], internal_0n[33]);
  C2 I575 (internal_0n[38], internal_0n[34], internal_0n[35]);
  C2 I576 (internal_0n[39], internal_0n[36], internal_0n[37]);
  C2 I577 (wc_0n, internal_0n[38], internal_0n[39]);
  OR2 I578 (complete1589_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I579 (complete1589_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I580 (complete1589_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I581 (complete1589_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I582 (complete1589_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I583 (complete1589_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I584 (complete1589_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I585 (complete1589_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I586 (complete1589_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I587 (complete1589_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I588 (complete1589_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I589 (complete1589_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I590 (complete1589_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I591 (complete1589_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I592 (complete1589_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I593 (complete1589_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I594 (complete1589_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I595 (complete1589_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I596 (complete1589_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I597 (complete1589_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I598 (complete1589_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I599 (complete1589_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I600 (complete1589_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I601 (complete1589_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I602 (complete1589_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I603 (complete1589_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I604 (complete1589_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I605 (complete1589_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I606 (complete1589_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I607 (complete1589_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I608 (complete1589_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I609 (complete1589_0n[31], wgfint_0n[31], wgtint_0n[31]);
  OR2 I610 (complete1589_0n[32], wgfint_0n[32], wgtint_0n[32]);
  OR2 I611 (complete1589_0n[33], wgfint_0n[33], wgtint_0n[33]);
  OR2 I612 (complete1589_0n[34], wgfint_0n[34], wgtint_0n[34]);
  OR2 I613 (complete1589_0n[35], wgfint_0n[35], wgtint_0n[35]);
  AO22 I614 (wacks_0n[35], gf1587_0n[35], df_0n[35], gt1588_0n[35], dt_0n[35]);
  NOR2 I615 (dt_0n[35], df_0n[35], gf1587_0n[35]);
  NOR3 I616 (df_0n[35], dt_0n[35], gt1588_0n[35], init_0n);
  AND2 I617 (gt1588_0n[35], wt_0n[35], wen_0n[35]);
  AND2 I618 (gf1587_0n[35], wf_0n[35], wen_0n[35]);
  AO22 I619 (wacks_0n[34], gf1587_0n[34], df_0n[34], gt1588_0n[34], dt_0n[34]);
  NOR2 I620 (dt_0n[34], df_0n[34], gf1587_0n[34]);
  NOR3 I621 (df_0n[34], dt_0n[34], gt1588_0n[34], init_0n);
  AND2 I622 (gt1588_0n[34], wt_0n[34], wen_0n[34]);
  AND2 I623 (gf1587_0n[34], wf_0n[34], wen_0n[34]);
  AO22 I624 (wacks_0n[33], gf1587_0n[33], df_0n[33], gt1588_0n[33], dt_0n[33]);
  NOR2 I625 (dt_0n[33], df_0n[33], gf1587_0n[33]);
  NOR3 I626 (df_0n[33], dt_0n[33], gt1588_0n[33], init_0n);
  AND2 I627 (gt1588_0n[33], wt_0n[33], wen_0n[33]);
  AND2 I628 (gf1587_0n[33], wf_0n[33], wen_0n[33]);
  AO22 I629 (wacks_0n[32], gf1587_0n[32], df_0n[32], gt1588_0n[32], dt_0n[32]);
  NOR2 I630 (dt_0n[32], df_0n[32], gf1587_0n[32]);
  NOR3 I631 (df_0n[32], dt_0n[32], gt1588_0n[32], init_0n);
  AND2 I632 (gt1588_0n[32], wt_0n[32], wen_0n[32]);
  AND2 I633 (gf1587_0n[32], wf_0n[32], wen_0n[32]);
  AO22 I634 (wacks_0n[31], gf1587_0n[31], df_0n[31], gt1588_0n[31], dt_0n[31]);
  NOR2 I635 (dt_0n[31], df_0n[31], gf1587_0n[31]);
  NOR3 I636 (df_0n[31], dt_0n[31], gt1588_0n[31], init_0n);
  AND2 I637 (gt1588_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I638 (gf1587_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I639 (wacks_0n[30], gf1587_0n[30], df_0n[30], gt1588_0n[30], dt_0n[30]);
  NOR2 I640 (dt_0n[30], df_0n[30], gf1587_0n[30]);
  NOR3 I641 (df_0n[30], dt_0n[30], gt1588_0n[30], init_0n);
  AND2 I642 (gt1588_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I643 (gf1587_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I644 (wacks_0n[29], gf1587_0n[29], df_0n[29], gt1588_0n[29], dt_0n[29]);
  NOR2 I645 (dt_0n[29], df_0n[29], gf1587_0n[29]);
  NOR3 I646 (df_0n[29], dt_0n[29], gt1588_0n[29], init_0n);
  AND2 I647 (gt1588_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I648 (gf1587_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I649 (wacks_0n[28], gf1587_0n[28], df_0n[28], gt1588_0n[28], dt_0n[28]);
  NOR2 I650 (dt_0n[28], df_0n[28], gf1587_0n[28]);
  NOR3 I651 (df_0n[28], dt_0n[28], gt1588_0n[28], init_0n);
  AND2 I652 (gt1588_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I653 (gf1587_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I654 (wacks_0n[27], gf1587_0n[27], df_0n[27], gt1588_0n[27], dt_0n[27]);
  NOR2 I655 (dt_0n[27], df_0n[27], gf1587_0n[27]);
  NOR3 I656 (df_0n[27], dt_0n[27], gt1588_0n[27], init_0n);
  AND2 I657 (gt1588_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I658 (gf1587_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I659 (wacks_0n[26], gf1587_0n[26], df_0n[26], gt1588_0n[26], dt_0n[26]);
  NOR2 I660 (dt_0n[26], df_0n[26], gf1587_0n[26]);
  NOR3 I661 (df_0n[26], dt_0n[26], gt1588_0n[26], init_0n);
  AND2 I662 (gt1588_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I663 (gf1587_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I664 (wacks_0n[25], gf1587_0n[25], df_0n[25], gt1588_0n[25], dt_0n[25]);
  NOR2 I665 (dt_0n[25], df_0n[25], gf1587_0n[25]);
  NOR3 I666 (df_0n[25], dt_0n[25], gt1588_0n[25], init_0n);
  AND2 I667 (gt1588_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I668 (gf1587_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I669 (wacks_0n[24], gf1587_0n[24], df_0n[24], gt1588_0n[24], dt_0n[24]);
  NOR2 I670 (dt_0n[24], df_0n[24], gf1587_0n[24]);
  NOR3 I671 (df_0n[24], dt_0n[24], gt1588_0n[24], init_0n);
  AND2 I672 (gt1588_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I673 (gf1587_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I674 (wacks_0n[23], gf1587_0n[23], df_0n[23], gt1588_0n[23], dt_0n[23]);
  NOR2 I675 (dt_0n[23], df_0n[23], gf1587_0n[23]);
  NOR3 I676 (df_0n[23], dt_0n[23], gt1588_0n[23], init_0n);
  AND2 I677 (gt1588_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I678 (gf1587_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I679 (wacks_0n[22], gf1587_0n[22], df_0n[22], gt1588_0n[22], dt_0n[22]);
  NOR2 I680 (dt_0n[22], df_0n[22], gf1587_0n[22]);
  NOR3 I681 (df_0n[22], dt_0n[22], gt1588_0n[22], init_0n);
  AND2 I682 (gt1588_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I683 (gf1587_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I684 (wacks_0n[21], gf1587_0n[21], df_0n[21], gt1588_0n[21], dt_0n[21]);
  NOR2 I685 (dt_0n[21], df_0n[21], gf1587_0n[21]);
  NOR3 I686 (df_0n[21], dt_0n[21], gt1588_0n[21], init_0n);
  AND2 I687 (gt1588_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I688 (gf1587_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I689 (wacks_0n[20], gf1587_0n[20], df_0n[20], gt1588_0n[20], dt_0n[20]);
  NOR2 I690 (dt_0n[20], df_0n[20], gf1587_0n[20]);
  NOR3 I691 (df_0n[20], dt_0n[20], gt1588_0n[20], init_0n);
  AND2 I692 (gt1588_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I693 (gf1587_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I694 (wacks_0n[19], gf1587_0n[19], df_0n[19], gt1588_0n[19], dt_0n[19]);
  NOR2 I695 (dt_0n[19], df_0n[19], gf1587_0n[19]);
  NOR3 I696 (df_0n[19], dt_0n[19], gt1588_0n[19], init_0n);
  AND2 I697 (gt1588_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I698 (gf1587_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I699 (wacks_0n[18], gf1587_0n[18], df_0n[18], gt1588_0n[18], dt_0n[18]);
  NOR2 I700 (dt_0n[18], df_0n[18], gf1587_0n[18]);
  NOR3 I701 (df_0n[18], dt_0n[18], gt1588_0n[18], init_0n);
  AND2 I702 (gt1588_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I703 (gf1587_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I704 (wacks_0n[17], gf1587_0n[17], df_0n[17], gt1588_0n[17], dt_0n[17]);
  NOR2 I705 (dt_0n[17], df_0n[17], gf1587_0n[17]);
  NOR3 I706 (df_0n[17], dt_0n[17], gt1588_0n[17], init_0n);
  AND2 I707 (gt1588_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I708 (gf1587_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I709 (wacks_0n[16], gf1587_0n[16], df_0n[16], gt1588_0n[16], dt_0n[16]);
  NOR2 I710 (dt_0n[16], df_0n[16], gf1587_0n[16]);
  NOR3 I711 (df_0n[16], dt_0n[16], gt1588_0n[16], init_0n);
  AND2 I712 (gt1588_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I713 (gf1587_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I714 (wacks_0n[15], gf1587_0n[15], df_0n[15], gt1588_0n[15], dt_0n[15]);
  NOR2 I715 (dt_0n[15], df_0n[15], gf1587_0n[15]);
  NOR3 I716 (df_0n[15], dt_0n[15], gt1588_0n[15], init_0n);
  AND2 I717 (gt1588_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I718 (gf1587_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I719 (wacks_0n[14], gf1587_0n[14], df_0n[14], gt1588_0n[14], dt_0n[14]);
  NOR2 I720 (dt_0n[14], df_0n[14], gf1587_0n[14]);
  NOR3 I721 (df_0n[14], dt_0n[14], gt1588_0n[14], init_0n);
  AND2 I722 (gt1588_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I723 (gf1587_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I724 (wacks_0n[13], gf1587_0n[13], df_0n[13], gt1588_0n[13], dt_0n[13]);
  NOR2 I725 (dt_0n[13], df_0n[13], gf1587_0n[13]);
  NOR3 I726 (df_0n[13], dt_0n[13], gt1588_0n[13], init_0n);
  AND2 I727 (gt1588_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I728 (gf1587_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I729 (wacks_0n[12], gf1587_0n[12], df_0n[12], gt1588_0n[12], dt_0n[12]);
  NOR2 I730 (dt_0n[12], df_0n[12], gf1587_0n[12]);
  NOR3 I731 (df_0n[12], dt_0n[12], gt1588_0n[12], init_0n);
  AND2 I732 (gt1588_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I733 (gf1587_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I734 (wacks_0n[11], gf1587_0n[11], df_0n[11], gt1588_0n[11], dt_0n[11]);
  NOR2 I735 (dt_0n[11], df_0n[11], gf1587_0n[11]);
  NOR3 I736 (df_0n[11], dt_0n[11], gt1588_0n[11], init_0n);
  AND2 I737 (gt1588_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I738 (gf1587_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I739 (wacks_0n[10], gf1587_0n[10], df_0n[10], gt1588_0n[10], dt_0n[10]);
  NOR2 I740 (dt_0n[10], df_0n[10], gf1587_0n[10]);
  NOR3 I741 (df_0n[10], dt_0n[10], gt1588_0n[10], init_0n);
  AND2 I742 (gt1588_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I743 (gf1587_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I744 (wacks_0n[9], gf1587_0n[9], df_0n[9], gt1588_0n[9], dt_0n[9]);
  NOR2 I745 (dt_0n[9], df_0n[9], gf1587_0n[9]);
  NOR3 I746 (df_0n[9], dt_0n[9], gt1588_0n[9], init_0n);
  AND2 I747 (gt1588_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I748 (gf1587_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I749 (wacks_0n[8], gf1587_0n[8], df_0n[8], gt1588_0n[8], dt_0n[8]);
  NOR2 I750 (dt_0n[8], df_0n[8], gf1587_0n[8]);
  NOR3 I751 (df_0n[8], dt_0n[8], gt1588_0n[8], init_0n);
  AND2 I752 (gt1588_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I753 (gf1587_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I754 (wacks_0n[7], gf1587_0n[7], df_0n[7], gt1588_0n[7], dt_0n[7]);
  NOR2 I755 (dt_0n[7], df_0n[7], gf1587_0n[7]);
  NOR3 I756 (df_0n[7], dt_0n[7], gt1588_0n[7], init_0n);
  AND2 I757 (gt1588_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I758 (gf1587_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I759 (wacks_0n[6], gf1587_0n[6], df_0n[6], gt1588_0n[6], dt_0n[6]);
  NOR2 I760 (dt_0n[6], df_0n[6], gf1587_0n[6]);
  NOR3 I761 (df_0n[6], dt_0n[6], gt1588_0n[6], init_0n);
  AND2 I762 (gt1588_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I763 (gf1587_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I764 (wacks_0n[5], gf1587_0n[5], df_0n[5], gt1588_0n[5], dt_0n[5]);
  NOR2 I765 (dt_0n[5], df_0n[5], gf1587_0n[5]);
  NOR3 I766 (df_0n[5], dt_0n[5], gt1588_0n[5], init_0n);
  AND2 I767 (gt1588_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I768 (gf1587_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I769 (wacks_0n[4], gf1587_0n[4], df_0n[4], gt1588_0n[4], dt_0n[4]);
  NOR2 I770 (dt_0n[4], df_0n[4], gf1587_0n[4]);
  NOR3 I771 (df_0n[4], dt_0n[4], gt1588_0n[4], init_0n);
  AND2 I772 (gt1588_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I773 (gf1587_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I774 (wacks_0n[3], gf1587_0n[3], df_0n[3], gt1588_0n[3], dt_0n[3]);
  NOR2 I775 (dt_0n[3], df_0n[3], gf1587_0n[3]);
  NOR3 I776 (df_0n[3], dt_0n[3], gt1588_0n[3], init_0n);
  AND2 I777 (gt1588_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I778 (gf1587_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I779 (wacks_0n[2], gf1587_0n[2], df_0n[2], gt1588_0n[2], dt_0n[2]);
  NOR2 I780 (dt_0n[2], df_0n[2], gf1587_0n[2]);
  NOR3 I781 (df_0n[2], dt_0n[2], gt1588_0n[2], init_0n);
  AND2 I782 (gt1588_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I783 (gf1587_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I784 (wacks_0n[1], gf1587_0n[1], df_0n[1], gt1588_0n[1], dt_0n[1]);
  NOR2 I785 (dt_0n[1], df_0n[1], gf1587_0n[1]);
  NOR3 I786 (df_0n[1], dt_0n[1], gt1588_0n[1], init_0n);
  AND2 I787 (gt1588_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I788 (gf1587_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I789 (wacks_0n[0], gf1587_0n[0], df_0n[0], gt1588_0n[0], dt_0n[0]);
  NOR2 I790 (dt_0n[0], df_0n[0], gf1587_0n[0]);
  NOR3 I791 (df_0n[0], dt_0n[0], gt1588_0n[0], init_0n);
  AND2 I792 (gt1588_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I793 (gf1587_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I794 (init_0n, initialise);
endmodule

module BrzV_36_l6__28_29_l24__28_28_280_2036_29_2_m97m (
  wg_0r0d, wg_0r1d, wg_0a,
  wd_0r, wd_0a,
  rg_0r, rg_0a,
  rg_1r, rg_1a,
  rg_2r, rg_2a,
  rg_3r, rg_3a,
  rd_0r0d, rd_0r1d, rd_0a,
  rd_1r0d, rd_1r1d, rd_1a,
  rd_2r0d, rd_2r1d, rd_2a,
  rd_3r0d, rd_3r1d, rd_3a,
  initialise
);
  input [35:0] wg_0r0d;
  input [35:0] wg_0r1d;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  output rd_0r0d;
  output rd_0r1d;
  input rd_0a;
  output [31:0] rd_1r0d;
  output [31:0] rd_1r1d;
  input rd_1a;
  output [3:0] rd_2r0d;
  output [3:0] rd_2r1d;
  input rd_2a;
  output [35:0] rd_3r0d;
  output [35:0] rd_3r1d;
  input rd_3a;
  input initialise;
  wire [40:0] internal_0n;
  wire [35:0] wf_0n;
  wire [35:0] wt_0n;
  wire [35:0] df_0n;
  wire [35:0] dt_0n;
  wire rgrint_0n;
  wire rgrint_1n;
  wire rgrint_2n;
  wire rgrint_3n;
  wire wc_0n;
  wire [35:0] wacks_0n;
  wire wdrint_0n;
  wire wgaint_0n;
  wire [35:0] wgfint_0n;
  wire [35:0] wgtint_0n;
  wire rgaint_0n;
  wire rgaint_1n;
  wire rgaint_2n;
  wire rgaint_3n;
  wire rdfint_0n;
  wire [31:0] rdfint_1n;
  wire [3:0] rdfint_2n;
  wire [35:0] rdfint_3n;
  wire rdtint_0n;
  wire [31:0] rdtint_1n;
  wire [3:0] rdtint_2n;
  wire [35:0] rdtint_3n;
  wire [35:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire ig_0n;
  wire [35:0] gif_0n;
  wire [35:0] git_0n;
  wire [35:0] complete1604_0n;
  wire [35:0] gt1603_0n;
  wire [35:0] gf1602_0n;
  assign rgaint_3n = rd_3a;
  assign rd_3r0d[0] = rdfint_3n[0];
  assign rd_3r0d[1] = rdfint_3n[1];
  assign rd_3r0d[2] = rdfint_3n[2];
  assign rd_3r0d[3] = rdfint_3n[3];
  assign rd_3r0d[4] = rdfint_3n[4];
  assign rd_3r0d[5] = rdfint_3n[5];
  assign rd_3r0d[6] = rdfint_3n[6];
  assign rd_3r0d[7] = rdfint_3n[7];
  assign rd_3r0d[8] = rdfint_3n[8];
  assign rd_3r0d[9] = rdfint_3n[9];
  assign rd_3r0d[10] = rdfint_3n[10];
  assign rd_3r0d[11] = rdfint_3n[11];
  assign rd_3r0d[12] = rdfint_3n[12];
  assign rd_3r0d[13] = rdfint_3n[13];
  assign rd_3r0d[14] = rdfint_3n[14];
  assign rd_3r0d[15] = rdfint_3n[15];
  assign rd_3r0d[16] = rdfint_3n[16];
  assign rd_3r0d[17] = rdfint_3n[17];
  assign rd_3r0d[18] = rdfint_3n[18];
  assign rd_3r0d[19] = rdfint_3n[19];
  assign rd_3r0d[20] = rdfint_3n[20];
  assign rd_3r0d[21] = rdfint_3n[21];
  assign rd_3r0d[22] = rdfint_3n[22];
  assign rd_3r0d[23] = rdfint_3n[23];
  assign rd_3r0d[24] = rdfint_3n[24];
  assign rd_3r0d[25] = rdfint_3n[25];
  assign rd_3r0d[26] = rdfint_3n[26];
  assign rd_3r0d[27] = rdfint_3n[27];
  assign rd_3r0d[28] = rdfint_3n[28];
  assign rd_3r0d[29] = rdfint_3n[29];
  assign rd_3r0d[30] = rdfint_3n[30];
  assign rd_3r0d[31] = rdfint_3n[31];
  assign rd_3r0d[32] = rdfint_3n[32];
  assign rd_3r0d[33] = rdfint_3n[33];
  assign rd_3r0d[34] = rdfint_3n[34];
  assign rd_3r0d[35] = rdfint_3n[35];
  assign rd_3r1d[0] = rdtint_3n[0];
  assign rd_3r1d[1] = rdtint_3n[1];
  assign rd_3r1d[2] = rdtint_3n[2];
  assign rd_3r1d[3] = rdtint_3n[3];
  assign rd_3r1d[4] = rdtint_3n[4];
  assign rd_3r1d[5] = rdtint_3n[5];
  assign rd_3r1d[6] = rdtint_3n[6];
  assign rd_3r1d[7] = rdtint_3n[7];
  assign rd_3r1d[8] = rdtint_3n[8];
  assign rd_3r1d[9] = rdtint_3n[9];
  assign rd_3r1d[10] = rdtint_3n[10];
  assign rd_3r1d[11] = rdtint_3n[11];
  assign rd_3r1d[12] = rdtint_3n[12];
  assign rd_3r1d[13] = rdtint_3n[13];
  assign rd_3r1d[14] = rdtint_3n[14];
  assign rd_3r1d[15] = rdtint_3n[15];
  assign rd_3r1d[16] = rdtint_3n[16];
  assign rd_3r1d[17] = rdtint_3n[17];
  assign rd_3r1d[18] = rdtint_3n[18];
  assign rd_3r1d[19] = rdtint_3n[19];
  assign rd_3r1d[20] = rdtint_3n[20];
  assign rd_3r1d[21] = rdtint_3n[21];
  assign rd_3r1d[22] = rdtint_3n[22];
  assign rd_3r1d[23] = rdtint_3n[23];
  assign rd_3r1d[24] = rdtint_3n[24];
  assign rd_3r1d[25] = rdtint_3n[25];
  assign rd_3r1d[26] = rdtint_3n[26];
  assign rd_3r1d[27] = rdtint_3n[27];
  assign rd_3r1d[28] = rdtint_3n[28];
  assign rd_3r1d[29] = rdtint_3n[29];
  assign rd_3r1d[30] = rdtint_3n[30];
  assign rd_3r1d[31] = rdtint_3n[31];
  assign rd_3r1d[32] = rdtint_3n[32];
  assign rd_3r1d[33] = rdtint_3n[33];
  assign rd_3r1d[34] = rdtint_3n[34];
  assign rd_3r1d[35] = rdtint_3n[35];
  assign rgaint_2n = rd_2a;
  assign rd_2r0d[0] = rdfint_2n[0];
  assign rd_2r0d[1] = rdfint_2n[1];
  assign rd_2r0d[2] = rdfint_2n[2];
  assign rd_2r0d[3] = rdfint_2n[3];
  assign rd_2r1d[0] = rdtint_2n[0];
  assign rd_2r1d[1] = rdtint_2n[1];
  assign rd_2r1d[2] = rdtint_2n[2];
  assign rd_2r1d[3] = rdtint_2n[3];
  assign rgaint_1n = rd_1a;
  assign rd_1r0d[0] = rdfint_1n[0];
  assign rd_1r0d[1] = rdfint_1n[1];
  assign rd_1r0d[2] = rdfint_1n[2];
  assign rd_1r0d[3] = rdfint_1n[3];
  assign rd_1r0d[4] = rdfint_1n[4];
  assign rd_1r0d[5] = rdfint_1n[5];
  assign rd_1r0d[6] = rdfint_1n[6];
  assign rd_1r0d[7] = rdfint_1n[7];
  assign rd_1r0d[8] = rdfint_1n[8];
  assign rd_1r0d[9] = rdfint_1n[9];
  assign rd_1r0d[10] = rdfint_1n[10];
  assign rd_1r0d[11] = rdfint_1n[11];
  assign rd_1r0d[12] = rdfint_1n[12];
  assign rd_1r0d[13] = rdfint_1n[13];
  assign rd_1r0d[14] = rdfint_1n[14];
  assign rd_1r0d[15] = rdfint_1n[15];
  assign rd_1r0d[16] = rdfint_1n[16];
  assign rd_1r0d[17] = rdfint_1n[17];
  assign rd_1r0d[18] = rdfint_1n[18];
  assign rd_1r0d[19] = rdfint_1n[19];
  assign rd_1r0d[20] = rdfint_1n[20];
  assign rd_1r0d[21] = rdfint_1n[21];
  assign rd_1r0d[22] = rdfint_1n[22];
  assign rd_1r0d[23] = rdfint_1n[23];
  assign rd_1r0d[24] = rdfint_1n[24];
  assign rd_1r0d[25] = rdfint_1n[25];
  assign rd_1r0d[26] = rdfint_1n[26];
  assign rd_1r0d[27] = rdfint_1n[27];
  assign rd_1r0d[28] = rdfint_1n[28];
  assign rd_1r0d[29] = rdfint_1n[29];
  assign rd_1r0d[30] = rdfint_1n[30];
  assign rd_1r0d[31] = rdfint_1n[31];
  assign rd_1r1d[0] = rdtint_1n[0];
  assign rd_1r1d[1] = rdtint_1n[1];
  assign rd_1r1d[2] = rdtint_1n[2];
  assign rd_1r1d[3] = rdtint_1n[3];
  assign rd_1r1d[4] = rdtint_1n[4];
  assign rd_1r1d[5] = rdtint_1n[5];
  assign rd_1r1d[6] = rdtint_1n[6];
  assign rd_1r1d[7] = rdtint_1n[7];
  assign rd_1r1d[8] = rdtint_1n[8];
  assign rd_1r1d[9] = rdtint_1n[9];
  assign rd_1r1d[10] = rdtint_1n[10];
  assign rd_1r1d[11] = rdtint_1n[11];
  assign rd_1r1d[12] = rdtint_1n[12];
  assign rd_1r1d[13] = rdtint_1n[13];
  assign rd_1r1d[14] = rdtint_1n[14];
  assign rd_1r1d[15] = rdtint_1n[15];
  assign rd_1r1d[16] = rdtint_1n[16];
  assign rd_1r1d[17] = rdtint_1n[17];
  assign rd_1r1d[18] = rdtint_1n[18];
  assign rd_1r1d[19] = rdtint_1n[19];
  assign rd_1r1d[20] = rdtint_1n[20];
  assign rd_1r1d[21] = rdtint_1n[21];
  assign rd_1r1d[22] = rdtint_1n[22];
  assign rd_1r1d[23] = rdtint_1n[23];
  assign rd_1r1d[24] = rdtint_1n[24];
  assign rd_1r1d[25] = rdtint_1n[25];
  assign rd_1r1d[26] = rdtint_1n[26];
  assign rd_1r1d[27] = rdtint_1n[27];
  assign rd_1r1d[28] = rdtint_1n[28];
  assign rd_1r1d[29] = rdtint_1n[29];
  assign rd_1r1d[30] = rdtint_1n[30];
  assign rd_1r1d[31] = rdtint_1n[31];
  assign rgaint_0n = rd_0a;
  assign rd_0r0d = rdfint_0n;
  assign rd_0r1d = rdtint_0n;
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgfint_0n[32] = wg_0r0d[32];
  assign wgfint_0n[33] = wg_0r0d[33];
  assign wgfint_0n[34] = wg_0r0d[34];
  assign wgfint_0n[35] = wg_0r0d[35];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign wgtint_0n[32] = wg_0r1d[32];
  assign wgtint_0n[33] = wg_0r1d[33];
  assign wgtint_0n[34] = wg_0r1d[34];
  assign wgtint_0n[35] = wg_0r1d[35];
  assign rg_3a = rgaint_3n;
  assign rgrint_3n = rg_3r;
  assign rg_2a = rgaint_2n;
  assign rgrint_2n = rg_2r;
  assign rg_1a = rgaint_1n;
  assign rgrint_1n = rg_1r;
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR3 I233 (internal_0n[0], rgrint_0n, rgrint_1n, rgrint_2n);
  NOR3 I234 (internal_0n[1], rgrint_3n, rgaint_0n, rgaint_1n);
  NOR2 I235 (internal_0n[2], rgaint_2n, rgaint_3n);
  AND3 I236 (nanyread_0n, internal_0n[0], internal_0n[1], internal_0n[2]);
  AND2 I237 (rdtint_3n[0], rgrint_3n, dt_0n[0]);
  AND2 I238 (rdtint_3n[1], rgrint_3n, dt_0n[1]);
  AND2 I239 (rdtint_3n[2], rgrint_3n, dt_0n[2]);
  AND2 I240 (rdtint_3n[3], rgrint_3n, dt_0n[3]);
  AND2 I241 (rdtint_3n[4], rgrint_3n, dt_0n[4]);
  AND2 I242 (rdtint_3n[5], rgrint_3n, dt_0n[5]);
  AND2 I243 (rdtint_3n[6], rgrint_3n, dt_0n[6]);
  AND2 I244 (rdtint_3n[7], rgrint_3n, dt_0n[7]);
  AND2 I245 (rdtint_3n[8], rgrint_3n, dt_0n[8]);
  AND2 I246 (rdtint_3n[9], rgrint_3n, dt_0n[9]);
  AND2 I247 (rdtint_3n[10], rgrint_3n, dt_0n[10]);
  AND2 I248 (rdtint_3n[11], rgrint_3n, dt_0n[11]);
  AND2 I249 (rdtint_3n[12], rgrint_3n, dt_0n[12]);
  AND2 I250 (rdtint_3n[13], rgrint_3n, dt_0n[13]);
  AND2 I251 (rdtint_3n[14], rgrint_3n, dt_0n[14]);
  AND2 I252 (rdtint_3n[15], rgrint_3n, dt_0n[15]);
  AND2 I253 (rdtint_3n[16], rgrint_3n, dt_0n[16]);
  AND2 I254 (rdtint_3n[17], rgrint_3n, dt_0n[17]);
  AND2 I255 (rdtint_3n[18], rgrint_3n, dt_0n[18]);
  AND2 I256 (rdtint_3n[19], rgrint_3n, dt_0n[19]);
  AND2 I257 (rdtint_3n[20], rgrint_3n, dt_0n[20]);
  AND2 I258 (rdtint_3n[21], rgrint_3n, dt_0n[21]);
  AND2 I259 (rdtint_3n[22], rgrint_3n, dt_0n[22]);
  AND2 I260 (rdtint_3n[23], rgrint_3n, dt_0n[23]);
  AND2 I261 (rdtint_3n[24], rgrint_3n, dt_0n[24]);
  AND2 I262 (rdtint_3n[25], rgrint_3n, dt_0n[25]);
  AND2 I263 (rdtint_3n[26], rgrint_3n, dt_0n[26]);
  AND2 I264 (rdtint_3n[27], rgrint_3n, dt_0n[27]);
  AND2 I265 (rdtint_3n[28], rgrint_3n, dt_0n[28]);
  AND2 I266 (rdtint_3n[29], rgrint_3n, dt_0n[29]);
  AND2 I267 (rdtint_3n[30], rgrint_3n, dt_0n[30]);
  AND2 I268 (rdtint_3n[31], rgrint_3n, dt_0n[31]);
  AND2 I269 (rdtint_3n[32], rgrint_3n, dt_0n[32]);
  AND2 I270 (rdtint_3n[33], rgrint_3n, dt_0n[33]);
  AND2 I271 (rdtint_3n[34], rgrint_3n, dt_0n[34]);
  AND2 I272 (rdtint_3n[35], rgrint_3n, dt_0n[35]);
  AND2 I273 (rdtint_2n[0], rgrint_2n, dt_0n[0]);
  AND2 I274 (rdtint_2n[1], rgrint_2n, dt_0n[1]);
  AND2 I275 (rdtint_2n[2], rgrint_2n, dt_0n[2]);
  AND2 I276 (rdtint_2n[3], rgrint_2n, dt_0n[3]);
  AND2 I277 (rdtint_1n[0], rgrint_1n, dt_0n[2]);
  AND2 I278 (rdtint_1n[1], rgrint_1n, dt_0n[3]);
  AND2 I279 (rdtint_1n[2], rgrint_1n, dt_0n[4]);
  AND2 I280 (rdtint_1n[3], rgrint_1n, dt_0n[5]);
  AND2 I281 (rdtint_1n[4], rgrint_1n, dt_0n[6]);
  AND2 I282 (rdtint_1n[5], rgrint_1n, dt_0n[7]);
  AND2 I283 (rdtint_1n[6], rgrint_1n, dt_0n[8]);
  AND2 I284 (rdtint_1n[7], rgrint_1n, dt_0n[9]);
  AND2 I285 (rdtint_1n[8], rgrint_1n, dt_0n[10]);
  AND2 I286 (rdtint_1n[9], rgrint_1n, dt_0n[11]);
  AND2 I287 (rdtint_1n[10], rgrint_1n, dt_0n[12]);
  AND2 I288 (rdtint_1n[11], rgrint_1n, dt_0n[13]);
  AND2 I289 (rdtint_1n[12], rgrint_1n, dt_0n[14]);
  AND2 I290 (rdtint_1n[13], rgrint_1n, dt_0n[15]);
  AND2 I291 (rdtint_1n[14], rgrint_1n, dt_0n[16]);
  AND2 I292 (rdtint_1n[15], rgrint_1n, dt_0n[17]);
  AND2 I293 (rdtint_1n[16], rgrint_1n, dt_0n[18]);
  AND2 I294 (rdtint_1n[17], rgrint_1n, dt_0n[19]);
  AND2 I295 (rdtint_1n[18], rgrint_1n, dt_0n[20]);
  AND2 I296 (rdtint_1n[19], rgrint_1n, dt_0n[21]);
  AND2 I297 (rdtint_1n[20], rgrint_1n, dt_0n[22]);
  AND2 I298 (rdtint_1n[21], rgrint_1n, dt_0n[23]);
  AND2 I299 (rdtint_1n[22], rgrint_1n, dt_0n[24]);
  AND2 I300 (rdtint_1n[23], rgrint_1n, dt_0n[25]);
  AND2 I301 (rdtint_1n[24], rgrint_1n, dt_0n[26]);
  AND2 I302 (rdtint_1n[25], rgrint_1n, dt_0n[27]);
  AND2 I303 (rdtint_1n[26], rgrint_1n, dt_0n[28]);
  AND2 I304 (rdtint_1n[27], rgrint_1n, dt_0n[29]);
  AND2 I305 (rdtint_1n[28], rgrint_1n, dt_0n[30]);
  AND2 I306 (rdtint_1n[29], rgrint_1n, dt_0n[31]);
  AND2 I307 (rdtint_1n[30], rgrint_1n, dt_0n[32]);
  AND2 I308 (rdtint_1n[31], rgrint_1n, dt_0n[33]);
  AND2 I309 (rdtint_0n, rgrint_0n, dt_0n[34]);
  AND2 I310 (rdfint_3n[0], rgrint_3n, df_0n[0]);
  AND2 I311 (rdfint_3n[1], rgrint_3n, df_0n[1]);
  AND2 I312 (rdfint_3n[2], rgrint_3n, df_0n[2]);
  AND2 I313 (rdfint_3n[3], rgrint_3n, df_0n[3]);
  AND2 I314 (rdfint_3n[4], rgrint_3n, df_0n[4]);
  AND2 I315 (rdfint_3n[5], rgrint_3n, df_0n[5]);
  AND2 I316 (rdfint_3n[6], rgrint_3n, df_0n[6]);
  AND2 I317 (rdfint_3n[7], rgrint_3n, df_0n[7]);
  AND2 I318 (rdfint_3n[8], rgrint_3n, df_0n[8]);
  AND2 I319 (rdfint_3n[9], rgrint_3n, df_0n[9]);
  AND2 I320 (rdfint_3n[10], rgrint_3n, df_0n[10]);
  AND2 I321 (rdfint_3n[11], rgrint_3n, df_0n[11]);
  AND2 I322 (rdfint_3n[12], rgrint_3n, df_0n[12]);
  AND2 I323 (rdfint_3n[13], rgrint_3n, df_0n[13]);
  AND2 I324 (rdfint_3n[14], rgrint_3n, df_0n[14]);
  AND2 I325 (rdfint_3n[15], rgrint_3n, df_0n[15]);
  AND2 I326 (rdfint_3n[16], rgrint_3n, df_0n[16]);
  AND2 I327 (rdfint_3n[17], rgrint_3n, df_0n[17]);
  AND2 I328 (rdfint_3n[18], rgrint_3n, df_0n[18]);
  AND2 I329 (rdfint_3n[19], rgrint_3n, df_0n[19]);
  AND2 I330 (rdfint_3n[20], rgrint_3n, df_0n[20]);
  AND2 I331 (rdfint_3n[21], rgrint_3n, df_0n[21]);
  AND2 I332 (rdfint_3n[22], rgrint_3n, df_0n[22]);
  AND2 I333 (rdfint_3n[23], rgrint_3n, df_0n[23]);
  AND2 I334 (rdfint_3n[24], rgrint_3n, df_0n[24]);
  AND2 I335 (rdfint_3n[25], rgrint_3n, df_0n[25]);
  AND2 I336 (rdfint_3n[26], rgrint_3n, df_0n[26]);
  AND2 I337 (rdfint_3n[27], rgrint_3n, df_0n[27]);
  AND2 I338 (rdfint_3n[28], rgrint_3n, df_0n[28]);
  AND2 I339 (rdfint_3n[29], rgrint_3n, df_0n[29]);
  AND2 I340 (rdfint_3n[30], rgrint_3n, df_0n[30]);
  AND2 I341 (rdfint_3n[31], rgrint_3n, df_0n[31]);
  AND2 I342 (rdfint_3n[32], rgrint_3n, df_0n[32]);
  AND2 I343 (rdfint_3n[33], rgrint_3n, df_0n[33]);
  AND2 I344 (rdfint_3n[34], rgrint_3n, df_0n[34]);
  AND2 I345 (rdfint_3n[35], rgrint_3n, df_0n[35]);
  AND2 I346 (rdfint_2n[0], rgrint_2n, df_0n[0]);
  AND2 I347 (rdfint_2n[1], rgrint_2n, df_0n[1]);
  AND2 I348 (rdfint_2n[2], rgrint_2n, df_0n[2]);
  AND2 I349 (rdfint_2n[3], rgrint_2n, df_0n[3]);
  AND2 I350 (rdfint_1n[0], rgrint_1n, df_0n[2]);
  AND2 I351 (rdfint_1n[1], rgrint_1n, df_0n[3]);
  AND2 I352 (rdfint_1n[2], rgrint_1n, df_0n[4]);
  AND2 I353 (rdfint_1n[3], rgrint_1n, df_0n[5]);
  AND2 I354 (rdfint_1n[4], rgrint_1n, df_0n[6]);
  AND2 I355 (rdfint_1n[5], rgrint_1n, df_0n[7]);
  AND2 I356 (rdfint_1n[6], rgrint_1n, df_0n[8]);
  AND2 I357 (rdfint_1n[7], rgrint_1n, df_0n[9]);
  AND2 I358 (rdfint_1n[8], rgrint_1n, df_0n[10]);
  AND2 I359 (rdfint_1n[9], rgrint_1n, df_0n[11]);
  AND2 I360 (rdfint_1n[10], rgrint_1n, df_0n[12]);
  AND2 I361 (rdfint_1n[11], rgrint_1n, df_0n[13]);
  AND2 I362 (rdfint_1n[12], rgrint_1n, df_0n[14]);
  AND2 I363 (rdfint_1n[13], rgrint_1n, df_0n[15]);
  AND2 I364 (rdfint_1n[14], rgrint_1n, df_0n[16]);
  AND2 I365 (rdfint_1n[15], rgrint_1n, df_0n[17]);
  AND2 I366 (rdfint_1n[16], rgrint_1n, df_0n[18]);
  AND2 I367 (rdfint_1n[17], rgrint_1n, df_0n[19]);
  AND2 I368 (rdfint_1n[18], rgrint_1n, df_0n[20]);
  AND2 I369 (rdfint_1n[19], rgrint_1n, df_0n[21]);
  AND2 I370 (rdfint_1n[20], rgrint_1n, df_0n[22]);
  AND2 I371 (rdfint_1n[21], rgrint_1n, df_0n[23]);
  AND2 I372 (rdfint_1n[22], rgrint_1n, df_0n[24]);
  AND2 I373 (rdfint_1n[23], rgrint_1n, df_0n[25]);
  AND2 I374 (rdfint_1n[24], rgrint_1n, df_0n[26]);
  AND2 I375 (rdfint_1n[25], rgrint_1n, df_0n[27]);
  AND2 I376 (rdfint_1n[26], rgrint_1n, df_0n[28]);
  AND2 I377 (rdfint_1n[27], rgrint_1n, df_0n[29]);
  AND2 I378 (rdfint_1n[28], rgrint_1n, df_0n[30]);
  AND2 I379 (rdfint_1n[29], rgrint_1n, df_0n[31]);
  AND2 I380 (rdfint_1n[30], rgrint_1n, df_0n[32]);
  AND2 I381 (rdfint_1n[31], rgrint_1n, df_0n[33]);
  AND2 I382 (rdfint_0n, rgrint_0n, df_0n[34]);
  C3 I383 (internal_0n[3], wc_0n, wacks_0n[35], wacks_0n[34]);
  C3 I384 (internal_0n[4], wacks_0n[33], wacks_0n[32], wacks_0n[31]);
  C3 I385 (internal_0n[5], wacks_0n[30], wacks_0n[29], wacks_0n[28]);
  C3 I386 (internal_0n[6], wacks_0n[27], wacks_0n[26], wacks_0n[25]);
  C3 I387 (internal_0n[7], wacks_0n[24], wacks_0n[23], wacks_0n[22]);
  C3 I388 (internal_0n[8], wacks_0n[21], wacks_0n[20], wacks_0n[19]);
  C3 I389 (internal_0n[9], wacks_0n[18], wacks_0n[17], wacks_0n[16]);
  C3 I390 (internal_0n[10], wacks_0n[15], wacks_0n[14], wacks_0n[13]);
  C3 I391 (internal_0n[11], wacks_0n[12], wacks_0n[11], wacks_0n[10]);
  C3 I392 (internal_0n[12], wacks_0n[9], wacks_0n[8], wacks_0n[7]);
  C3 I393 (internal_0n[13], wacks_0n[6], wacks_0n[5], wacks_0n[4]);
  C2 I394 (internal_0n[14], wacks_0n[3], wacks_0n[2]);
  C2 I395 (internal_0n[15], wacks_0n[1], wacks_0n[0]);
  C3 I396 (internal_0n[16], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I397 (internal_0n[17], internal_0n[6], internal_0n[7], internal_0n[8]);
  C3 I398 (internal_0n[18], internal_0n[9], internal_0n[10], internal_0n[11]);
  C2 I399 (internal_0n[19], internal_0n[12], internal_0n[13]);
  C2 I400 (internal_0n[20], internal_0n[14], internal_0n[15]);
  C3 I401 (internal_0n[21], internal_0n[16], internal_0n[17], internal_0n[18]);
  C2 I402 (internal_0n[22], internal_0n[19], internal_0n[20]);
  C2 I403 (wdrint_0n, internal_0n[21], internal_0n[22]);
  assign wen_0n[35] = wc_0n;
  assign wen_0n[34] = wc_0n;
  assign wen_0n[33] = wc_0n;
  assign wen_0n[32] = wc_0n;
  assign wen_0n[31] = wc_0n;
  assign wen_0n[30] = wc_0n;
  assign wen_0n[29] = wc_0n;
  assign wen_0n[28] = wc_0n;
  assign wen_0n[27] = wc_0n;
  assign wen_0n[26] = wc_0n;
  assign wen_0n[25] = wc_0n;
  assign wen_0n[24] = wc_0n;
  assign wen_0n[23] = wc_0n;
  assign wen_0n[22] = wc_0n;
  assign wen_0n[21] = wc_0n;
  assign wen_0n[20] = wc_0n;
  assign wen_0n[19] = wc_0n;
  assign wen_0n[18] = wc_0n;
  assign wen_0n[17] = wc_0n;
  assign wen_0n[16] = wc_0n;
  assign wen_0n[15] = wc_0n;
  assign wen_0n[14] = wc_0n;
  assign wen_0n[13] = wc_0n;
  assign wen_0n[12] = wc_0n;
  assign wen_0n[11] = wc_0n;
  assign wen_0n[10] = wc_0n;
  assign wen_0n[9] = wc_0n;
  assign wen_0n[8] = wc_0n;
  assign wen_0n[7] = wc_0n;
  assign wen_0n[6] = wc_0n;
  assign wen_0n[5] = wc_0n;
  assign wen_0n[4] = wc_0n;
  assign wen_0n[3] = wc_0n;
  assign wen_0n[2] = wc_0n;
  assign wen_0n[1] = wc_0n;
  assign wen_0n[0] = wc_0n;
  assign wt_0n[35] = git_0n[35];
  assign wt_0n[34] = git_0n[34];
  assign wt_0n[33] = git_0n[33];
  assign wt_0n[32] = git_0n[32];
  assign wt_0n[31] = git_0n[31];
  assign wt_0n[30] = git_0n[30];
  assign wt_0n[29] = git_0n[29];
  assign wt_0n[28] = git_0n[28];
  assign wt_0n[27] = git_0n[27];
  assign wt_0n[26] = git_0n[26];
  assign wt_0n[25] = git_0n[25];
  assign wt_0n[24] = git_0n[24];
  assign wt_0n[23] = git_0n[23];
  assign wt_0n[22] = git_0n[22];
  assign wt_0n[21] = git_0n[21];
  assign wt_0n[20] = git_0n[20];
  assign wt_0n[19] = git_0n[19];
  assign wt_0n[18] = git_0n[18];
  assign wt_0n[17] = git_0n[17];
  assign wt_0n[16] = git_0n[16];
  assign wt_0n[15] = git_0n[15];
  assign wt_0n[14] = git_0n[14];
  assign wt_0n[13] = git_0n[13];
  assign wt_0n[12] = git_0n[12];
  assign wt_0n[11] = git_0n[11];
  assign wt_0n[10] = git_0n[10];
  assign wt_0n[9] = git_0n[9];
  assign wt_0n[8] = git_0n[8];
  assign wt_0n[7] = git_0n[7];
  assign wt_0n[6] = git_0n[6];
  assign wt_0n[5] = git_0n[5];
  assign wt_0n[4] = git_0n[4];
  assign wt_0n[3] = git_0n[3];
  assign wt_0n[2] = git_0n[2];
  assign wt_0n[1] = git_0n[1];
  assign wt_0n[0] = git_0n[0];
  assign wf_0n[35] = gif_0n[35];
  assign wf_0n[34] = gif_0n[34];
  assign wf_0n[33] = gif_0n[33];
  assign wf_0n[32] = gif_0n[32];
  assign wf_0n[31] = gif_0n[31];
  assign wf_0n[30] = gif_0n[30];
  assign wf_0n[29] = gif_0n[29];
  assign wf_0n[28] = gif_0n[28];
  assign wf_0n[27] = gif_0n[27];
  assign wf_0n[26] = gif_0n[26];
  assign wf_0n[25] = gif_0n[25];
  assign wf_0n[24] = gif_0n[24];
  assign wf_0n[23] = gif_0n[23];
  assign wf_0n[22] = gif_0n[22];
  assign wf_0n[21] = gif_0n[21];
  assign wf_0n[20] = gif_0n[20];
  assign wf_0n[19] = gif_0n[19];
  assign wf_0n[18] = gif_0n[18];
  assign wf_0n[17] = gif_0n[17];
  assign wf_0n[16] = gif_0n[16];
  assign wf_0n[15] = gif_0n[15];
  assign wf_0n[14] = gif_0n[14];
  assign wf_0n[13] = gif_0n[13];
  assign wf_0n[12] = gif_0n[12];
  assign wf_0n[11] = gif_0n[11];
  assign wf_0n[10] = gif_0n[10];
  assign wf_0n[9] = gif_0n[9];
  assign wf_0n[8] = gif_0n[8];
  assign wf_0n[7] = gif_0n[7];
  assign wf_0n[6] = gif_0n[6];
  assign wf_0n[5] = gif_0n[5];
  assign wf_0n[4] = gif_0n[4];
  assign wf_0n[3] = gif_0n[3];
  assign wf_0n[2] = gif_0n[2];
  assign wf_0n[1] = gif_0n[1];
  assign wf_0n[0] = gif_0n[0];
  AC2 I512 (ig_0n, igc_0n, nanyread_0n);
  assign igc_0n = wc_0n;
  AND2 I514 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I515 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I516 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I517 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I518 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I519 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I520 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I521 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I522 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I523 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I524 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I525 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I526 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I527 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I528 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I529 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I530 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I531 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I532 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I533 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I534 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I535 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I536 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I537 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I538 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I539 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I540 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I541 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I542 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I543 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I544 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I545 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I546 (git_0n[32], wgtint_0n[32], ig_0n);
  AND2 I547 (git_0n[33], wgtint_0n[33], ig_0n);
  AND2 I548 (git_0n[34], wgtint_0n[34], ig_0n);
  AND2 I549 (git_0n[35], wgtint_0n[35], ig_0n);
  AND2 I550 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I551 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I552 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I553 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I554 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I555 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I556 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I557 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I558 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I559 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I560 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I561 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I562 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I563 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I564 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I565 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I566 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I567 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I568 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I569 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I570 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I571 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I572 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I573 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I574 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I575 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I576 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I577 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I578 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I579 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I580 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I581 (gif_0n[31], wgfint_0n[31], ig_0n);
  AND2 I582 (gif_0n[32], wgfint_0n[32], ig_0n);
  AND2 I583 (gif_0n[33], wgfint_0n[33], ig_0n);
  AND2 I584 (gif_0n[34], wgfint_0n[34], ig_0n);
  AND2 I585 (gif_0n[35], wgfint_0n[35], ig_0n);
  C3 I586 (internal_0n[23], complete1604_0n[0], complete1604_0n[1], complete1604_0n[2]);
  C3 I587 (internal_0n[24], complete1604_0n[3], complete1604_0n[4], complete1604_0n[5]);
  C3 I588 (internal_0n[25], complete1604_0n[6], complete1604_0n[7], complete1604_0n[8]);
  C3 I589 (internal_0n[26], complete1604_0n[9], complete1604_0n[10], complete1604_0n[11]);
  C3 I590 (internal_0n[27], complete1604_0n[12], complete1604_0n[13], complete1604_0n[14]);
  C3 I591 (internal_0n[28], complete1604_0n[15], complete1604_0n[16], complete1604_0n[17]);
  C3 I592 (internal_0n[29], complete1604_0n[18], complete1604_0n[19], complete1604_0n[20]);
  C3 I593 (internal_0n[30], complete1604_0n[21], complete1604_0n[22], complete1604_0n[23]);
  C3 I594 (internal_0n[31], complete1604_0n[24], complete1604_0n[25], complete1604_0n[26]);
  C3 I595 (internal_0n[32], complete1604_0n[27], complete1604_0n[28], complete1604_0n[29]);
  C3 I596 (internal_0n[33], complete1604_0n[30], complete1604_0n[31], complete1604_0n[32]);
  C3 I597 (internal_0n[34], complete1604_0n[33], complete1604_0n[34], complete1604_0n[35]);
  C3 I598 (internal_0n[35], internal_0n[23], internal_0n[24], internal_0n[25]);
  C3 I599 (internal_0n[36], internal_0n[26], internal_0n[27], internal_0n[28]);
  C3 I600 (internal_0n[37], internal_0n[29], internal_0n[30], internal_0n[31]);
  C3 I601 (internal_0n[38], internal_0n[32], internal_0n[33], internal_0n[34]);
  C2 I602 (internal_0n[39], internal_0n[35], internal_0n[36]);
  C2 I603 (internal_0n[40], internal_0n[37], internal_0n[38]);
  C2 I604 (wc_0n, internal_0n[39], internal_0n[40]);
  OR2 I605 (complete1604_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I606 (complete1604_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I607 (complete1604_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I608 (complete1604_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I609 (complete1604_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I610 (complete1604_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I611 (complete1604_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I612 (complete1604_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I613 (complete1604_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I614 (complete1604_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I615 (complete1604_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I616 (complete1604_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I617 (complete1604_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I618 (complete1604_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I619 (complete1604_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I620 (complete1604_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I621 (complete1604_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I622 (complete1604_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I623 (complete1604_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I624 (complete1604_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I625 (complete1604_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I626 (complete1604_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I627 (complete1604_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I628 (complete1604_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I629 (complete1604_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I630 (complete1604_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I631 (complete1604_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I632 (complete1604_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I633 (complete1604_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I634 (complete1604_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I635 (complete1604_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I636 (complete1604_0n[31], wgfint_0n[31], wgtint_0n[31]);
  OR2 I637 (complete1604_0n[32], wgfint_0n[32], wgtint_0n[32]);
  OR2 I638 (complete1604_0n[33], wgfint_0n[33], wgtint_0n[33]);
  OR2 I639 (complete1604_0n[34], wgfint_0n[34], wgtint_0n[34]);
  OR2 I640 (complete1604_0n[35], wgfint_0n[35], wgtint_0n[35]);
  AO22 I641 (wacks_0n[35], gf1602_0n[35], df_0n[35], gt1603_0n[35], dt_0n[35]);
  NOR2 I642 (dt_0n[35], df_0n[35], gf1602_0n[35]);
  NOR3 I643 (df_0n[35], dt_0n[35], gt1603_0n[35], init_0n);
  AND2 I644 (gt1603_0n[35], wt_0n[35], wen_0n[35]);
  AND2 I645 (gf1602_0n[35], wf_0n[35], wen_0n[35]);
  AO22 I646 (wacks_0n[34], gf1602_0n[34], df_0n[34], gt1603_0n[34], dt_0n[34]);
  NOR2 I647 (dt_0n[34], df_0n[34], gf1602_0n[34]);
  NOR3 I648 (df_0n[34], dt_0n[34], gt1603_0n[34], init_0n);
  AND2 I649 (gt1603_0n[34], wt_0n[34], wen_0n[34]);
  AND2 I650 (gf1602_0n[34], wf_0n[34], wen_0n[34]);
  AO22 I651 (wacks_0n[33], gf1602_0n[33], df_0n[33], gt1603_0n[33], dt_0n[33]);
  NOR2 I652 (dt_0n[33], df_0n[33], gf1602_0n[33]);
  NOR3 I653 (df_0n[33], dt_0n[33], gt1603_0n[33], init_0n);
  AND2 I654 (gt1603_0n[33], wt_0n[33], wen_0n[33]);
  AND2 I655 (gf1602_0n[33], wf_0n[33], wen_0n[33]);
  AO22 I656 (wacks_0n[32], gf1602_0n[32], df_0n[32], gt1603_0n[32], dt_0n[32]);
  NOR2 I657 (dt_0n[32], df_0n[32], gf1602_0n[32]);
  NOR3 I658 (df_0n[32], dt_0n[32], gt1603_0n[32], init_0n);
  AND2 I659 (gt1603_0n[32], wt_0n[32], wen_0n[32]);
  AND2 I660 (gf1602_0n[32], wf_0n[32], wen_0n[32]);
  AO22 I661 (wacks_0n[31], gf1602_0n[31], df_0n[31], gt1603_0n[31], dt_0n[31]);
  NOR2 I662 (dt_0n[31], df_0n[31], gf1602_0n[31]);
  NOR3 I663 (df_0n[31], dt_0n[31], gt1603_0n[31], init_0n);
  AND2 I664 (gt1603_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I665 (gf1602_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I666 (wacks_0n[30], gf1602_0n[30], df_0n[30], gt1603_0n[30], dt_0n[30]);
  NOR2 I667 (dt_0n[30], df_0n[30], gf1602_0n[30]);
  NOR3 I668 (df_0n[30], dt_0n[30], gt1603_0n[30], init_0n);
  AND2 I669 (gt1603_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I670 (gf1602_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I671 (wacks_0n[29], gf1602_0n[29], df_0n[29], gt1603_0n[29], dt_0n[29]);
  NOR2 I672 (dt_0n[29], df_0n[29], gf1602_0n[29]);
  NOR3 I673 (df_0n[29], dt_0n[29], gt1603_0n[29], init_0n);
  AND2 I674 (gt1603_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I675 (gf1602_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I676 (wacks_0n[28], gf1602_0n[28], df_0n[28], gt1603_0n[28], dt_0n[28]);
  NOR2 I677 (dt_0n[28], df_0n[28], gf1602_0n[28]);
  NOR3 I678 (df_0n[28], dt_0n[28], gt1603_0n[28], init_0n);
  AND2 I679 (gt1603_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I680 (gf1602_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I681 (wacks_0n[27], gf1602_0n[27], df_0n[27], gt1603_0n[27], dt_0n[27]);
  NOR2 I682 (dt_0n[27], df_0n[27], gf1602_0n[27]);
  NOR3 I683 (df_0n[27], dt_0n[27], gt1603_0n[27], init_0n);
  AND2 I684 (gt1603_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I685 (gf1602_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I686 (wacks_0n[26], gf1602_0n[26], df_0n[26], gt1603_0n[26], dt_0n[26]);
  NOR2 I687 (dt_0n[26], df_0n[26], gf1602_0n[26]);
  NOR3 I688 (df_0n[26], dt_0n[26], gt1603_0n[26], init_0n);
  AND2 I689 (gt1603_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I690 (gf1602_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I691 (wacks_0n[25], gf1602_0n[25], df_0n[25], gt1603_0n[25], dt_0n[25]);
  NOR2 I692 (dt_0n[25], df_0n[25], gf1602_0n[25]);
  NOR3 I693 (df_0n[25], dt_0n[25], gt1603_0n[25], init_0n);
  AND2 I694 (gt1603_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I695 (gf1602_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I696 (wacks_0n[24], gf1602_0n[24], df_0n[24], gt1603_0n[24], dt_0n[24]);
  NOR2 I697 (dt_0n[24], df_0n[24], gf1602_0n[24]);
  NOR3 I698 (df_0n[24], dt_0n[24], gt1603_0n[24], init_0n);
  AND2 I699 (gt1603_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I700 (gf1602_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I701 (wacks_0n[23], gf1602_0n[23], df_0n[23], gt1603_0n[23], dt_0n[23]);
  NOR2 I702 (dt_0n[23], df_0n[23], gf1602_0n[23]);
  NOR3 I703 (df_0n[23], dt_0n[23], gt1603_0n[23], init_0n);
  AND2 I704 (gt1603_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I705 (gf1602_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I706 (wacks_0n[22], gf1602_0n[22], df_0n[22], gt1603_0n[22], dt_0n[22]);
  NOR2 I707 (dt_0n[22], df_0n[22], gf1602_0n[22]);
  NOR3 I708 (df_0n[22], dt_0n[22], gt1603_0n[22], init_0n);
  AND2 I709 (gt1603_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I710 (gf1602_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I711 (wacks_0n[21], gf1602_0n[21], df_0n[21], gt1603_0n[21], dt_0n[21]);
  NOR2 I712 (dt_0n[21], df_0n[21], gf1602_0n[21]);
  NOR3 I713 (df_0n[21], dt_0n[21], gt1603_0n[21], init_0n);
  AND2 I714 (gt1603_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I715 (gf1602_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I716 (wacks_0n[20], gf1602_0n[20], df_0n[20], gt1603_0n[20], dt_0n[20]);
  NOR2 I717 (dt_0n[20], df_0n[20], gf1602_0n[20]);
  NOR3 I718 (df_0n[20], dt_0n[20], gt1603_0n[20], init_0n);
  AND2 I719 (gt1603_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I720 (gf1602_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I721 (wacks_0n[19], gf1602_0n[19], df_0n[19], gt1603_0n[19], dt_0n[19]);
  NOR2 I722 (dt_0n[19], df_0n[19], gf1602_0n[19]);
  NOR3 I723 (df_0n[19], dt_0n[19], gt1603_0n[19], init_0n);
  AND2 I724 (gt1603_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I725 (gf1602_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I726 (wacks_0n[18], gf1602_0n[18], df_0n[18], gt1603_0n[18], dt_0n[18]);
  NOR2 I727 (dt_0n[18], df_0n[18], gf1602_0n[18]);
  NOR3 I728 (df_0n[18], dt_0n[18], gt1603_0n[18], init_0n);
  AND2 I729 (gt1603_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I730 (gf1602_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I731 (wacks_0n[17], gf1602_0n[17], df_0n[17], gt1603_0n[17], dt_0n[17]);
  NOR2 I732 (dt_0n[17], df_0n[17], gf1602_0n[17]);
  NOR3 I733 (df_0n[17], dt_0n[17], gt1603_0n[17], init_0n);
  AND2 I734 (gt1603_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I735 (gf1602_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I736 (wacks_0n[16], gf1602_0n[16], df_0n[16], gt1603_0n[16], dt_0n[16]);
  NOR2 I737 (dt_0n[16], df_0n[16], gf1602_0n[16]);
  NOR3 I738 (df_0n[16], dt_0n[16], gt1603_0n[16], init_0n);
  AND2 I739 (gt1603_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I740 (gf1602_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I741 (wacks_0n[15], gf1602_0n[15], df_0n[15], gt1603_0n[15], dt_0n[15]);
  NOR2 I742 (dt_0n[15], df_0n[15], gf1602_0n[15]);
  NOR3 I743 (df_0n[15], dt_0n[15], gt1603_0n[15], init_0n);
  AND2 I744 (gt1603_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I745 (gf1602_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I746 (wacks_0n[14], gf1602_0n[14], df_0n[14], gt1603_0n[14], dt_0n[14]);
  NOR2 I747 (dt_0n[14], df_0n[14], gf1602_0n[14]);
  NOR3 I748 (df_0n[14], dt_0n[14], gt1603_0n[14], init_0n);
  AND2 I749 (gt1603_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I750 (gf1602_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I751 (wacks_0n[13], gf1602_0n[13], df_0n[13], gt1603_0n[13], dt_0n[13]);
  NOR2 I752 (dt_0n[13], df_0n[13], gf1602_0n[13]);
  NOR3 I753 (df_0n[13], dt_0n[13], gt1603_0n[13], init_0n);
  AND2 I754 (gt1603_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I755 (gf1602_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I756 (wacks_0n[12], gf1602_0n[12], df_0n[12], gt1603_0n[12], dt_0n[12]);
  NOR2 I757 (dt_0n[12], df_0n[12], gf1602_0n[12]);
  NOR3 I758 (df_0n[12], dt_0n[12], gt1603_0n[12], init_0n);
  AND2 I759 (gt1603_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I760 (gf1602_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I761 (wacks_0n[11], gf1602_0n[11], df_0n[11], gt1603_0n[11], dt_0n[11]);
  NOR2 I762 (dt_0n[11], df_0n[11], gf1602_0n[11]);
  NOR3 I763 (df_0n[11], dt_0n[11], gt1603_0n[11], init_0n);
  AND2 I764 (gt1603_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I765 (gf1602_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I766 (wacks_0n[10], gf1602_0n[10], df_0n[10], gt1603_0n[10], dt_0n[10]);
  NOR2 I767 (dt_0n[10], df_0n[10], gf1602_0n[10]);
  NOR3 I768 (df_0n[10], dt_0n[10], gt1603_0n[10], init_0n);
  AND2 I769 (gt1603_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I770 (gf1602_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I771 (wacks_0n[9], gf1602_0n[9], df_0n[9], gt1603_0n[9], dt_0n[9]);
  NOR2 I772 (dt_0n[9], df_0n[9], gf1602_0n[9]);
  NOR3 I773 (df_0n[9], dt_0n[9], gt1603_0n[9], init_0n);
  AND2 I774 (gt1603_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I775 (gf1602_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I776 (wacks_0n[8], gf1602_0n[8], df_0n[8], gt1603_0n[8], dt_0n[8]);
  NOR2 I777 (dt_0n[8], df_0n[8], gf1602_0n[8]);
  NOR3 I778 (df_0n[8], dt_0n[8], gt1603_0n[8], init_0n);
  AND2 I779 (gt1603_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I780 (gf1602_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I781 (wacks_0n[7], gf1602_0n[7], df_0n[7], gt1603_0n[7], dt_0n[7]);
  NOR2 I782 (dt_0n[7], df_0n[7], gf1602_0n[7]);
  NOR3 I783 (df_0n[7], dt_0n[7], gt1603_0n[7], init_0n);
  AND2 I784 (gt1603_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I785 (gf1602_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I786 (wacks_0n[6], gf1602_0n[6], df_0n[6], gt1603_0n[6], dt_0n[6]);
  NOR2 I787 (dt_0n[6], df_0n[6], gf1602_0n[6]);
  NOR3 I788 (df_0n[6], dt_0n[6], gt1603_0n[6], init_0n);
  AND2 I789 (gt1603_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I790 (gf1602_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I791 (wacks_0n[5], gf1602_0n[5], df_0n[5], gt1603_0n[5], dt_0n[5]);
  NOR2 I792 (dt_0n[5], df_0n[5], gf1602_0n[5]);
  NOR3 I793 (df_0n[5], dt_0n[5], gt1603_0n[5], init_0n);
  AND2 I794 (gt1603_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I795 (gf1602_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I796 (wacks_0n[4], gf1602_0n[4], df_0n[4], gt1603_0n[4], dt_0n[4]);
  NOR2 I797 (dt_0n[4], df_0n[4], gf1602_0n[4]);
  NOR3 I798 (df_0n[4], dt_0n[4], gt1603_0n[4], init_0n);
  AND2 I799 (gt1603_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I800 (gf1602_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I801 (wacks_0n[3], gf1602_0n[3], df_0n[3], gt1603_0n[3], dt_0n[3]);
  NOR2 I802 (dt_0n[3], df_0n[3], gf1602_0n[3]);
  NOR3 I803 (df_0n[3], dt_0n[3], gt1603_0n[3], init_0n);
  AND2 I804 (gt1603_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I805 (gf1602_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I806 (wacks_0n[2], gf1602_0n[2], df_0n[2], gt1603_0n[2], dt_0n[2]);
  NOR2 I807 (dt_0n[2], df_0n[2], gf1602_0n[2]);
  NOR3 I808 (df_0n[2], dt_0n[2], gt1603_0n[2], init_0n);
  AND2 I809 (gt1603_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I810 (gf1602_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I811 (wacks_0n[1], gf1602_0n[1], df_0n[1], gt1603_0n[1], dt_0n[1]);
  NOR2 I812 (dt_0n[1], df_0n[1], gf1602_0n[1]);
  NOR3 I813 (df_0n[1], dt_0n[1], gt1603_0n[1], init_0n);
  AND2 I814 (gt1603_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I815 (gf1602_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I816 (wacks_0n[0], gf1602_0n[0], df_0n[0], gt1603_0n[0], dt_0n[0]);
  NOR2 I817 (dt_0n[0], df_0n[0], gf1602_0n[0]);
  NOR3 I818 (df_0n[0], dt_0n[0], gt1603_0n[0], init_0n);
  AND2 I819 (gt1603_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I820 (gf1602_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I821 (init_0n, initialise);
endmodule

module BrzV_36_l6__28_29_l45__28_28_280_2036_29_2_m98m (
  wg_0r0d, wg_0r1d, wg_0a,
  wg_1r0d, wg_1r1d, wg_1a,
  wd_0r, wd_0a,
  wd_1r, wd_1a,
  rg_0r, rg_0a,
  rd_0r0d, rd_0r1d, rd_0a,
  initialise
);
  input [35:0] wg_0r0d;
  input [35:0] wg_0r1d;
  output wg_0a;
  input [35:0] wg_1r0d;
  input [35:0] wg_1r1d;
  output wg_1a;
  output wd_0r;
  input wd_0a;
  output wd_1r;
  input wd_1a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0d;
  output [31:0] rd_0r1d;
  input rd_0a;
  input initialise;
  wire [75:0] internal_0n;
  wire [35:0] wf_0n;
  wire [35:0] wt_0n;
  wire [35:0] df_0n;
  wire [35:0] dt_0n;
  wire rgrint_0n;
  wire wc_0n;
  wire wc_1n;
  wire [35:0] wacks_0n;
  wire wdrint_0n;
  wire wdrint_1n;
  wire wgaint_0n;
  wire wgaint_1n;
  wire [35:0] wgfint_0n;
  wire [35:0] wgfint_1n;
  wire [35:0] wgtint_0n;
  wire [35:0] wgtint_1n;
  wire rgaint_0n;
  wire [31:0] rdfint_0n;
  wire [31:0] rdtint_0n;
  wire [35:0] wen_0n;
  wire init_0n;
  wire nanyread_0n;
  wire igc_0n;
  wire igc_1n;
  wire ig_0n;
  wire ig_1n;
  wire [35:0] gif_0n;
  wire [35:0] gif_1n;
  wire [35:0] git_0n;
  wire [35:0] git_1n;
  wire [35:0] complete1628_0n;
  wire [35:0] complete1627_0n;
  wire [35:0] gt1626_0n;
  wire [35:0] gf1625_0n;
  assign rgaint_0n = rd_0a;
  assign rd_0r0d[0] = rdfint_0n[0];
  assign rd_0r0d[1] = rdfint_0n[1];
  assign rd_0r0d[2] = rdfint_0n[2];
  assign rd_0r0d[3] = rdfint_0n[3];
  assign rd_0r0d[4] = rdfint_0n[4];
  assign rd_0r0d[5] = rdfint_0n[5];
  assign rd_0r0d[6] = rdfint_0n[6];
  assign rd_0r0d[7] = rdfint_0n[7];
  assign rd_0r0d[8] = rdfint_0n[8];
  assign rd_0r0d[9] = rdfint_0n[9];
  assign rd_0r0d[10] = rdfint_0n[10];
  assign rd_0r0d[11] = rdfint_0n[11];
  assign rd_0r0d[12] = rdfint_0n[12];
  assign rd_0r0d[13] = rdfint_0n[13];
  assign rd_0r0d[14] = rdfint_0n[14];
  assign rd_0r0d[15] = rdfint_0n[15];
  assign rd_0r0d[16] = rdfint_0n[16];
  assign rd_0r0d[17] = rdfint_0n[17];
  assign rd_0r0d[18] = rdfint_0n[18];
  assign rd_0r0d[19] = rdfint_0n[19];
  assign rd_0r0d[20] = rdfint_0n[20];
  assign rd_0r0d[21] = rdfint_0n[21];
  assign rd_0r0d[22] = rdfint_0n[22];
  assign rd_0r0d[23] = rdfint_0n[23];
  assign rd_0r0d[24] = rdfint_0n[24];
  assign rd_0r0d[25] = rdfint_0n[25];
  assign rd_0r0d[26] = rdfint_0n[26];
  assign rd_0r0d[27] = rdfint_0n[27];
  assign rd_0r0d[28] = rdfint_0n[28];
  assign rd_0r0d[29] = rdfint_0n[29];
  assign rd_0r0d[30] = rdfint_0n[30];
  assign rd_0r0d[31] = rdfint_0n[31];
  assign rd_0r1d[0] = rdtint_0n[0];
  assign rd_0r1d[1] = rdtint_0n[1];
  assign rd_0r1d[2] = rdtint_0n[2];
  assign rd_0r1d[3] = rdtint_0n[3];
  assign rd_0r1d[4] = rdtint_0n[4];
  assign rd_0r1d[5] = rdtint_0n[5];
  assign rd_0r1d[6] = rdtint_0n[6];
  assign rd_0r1d[7] = rdtint_0n[7];
  assign rd_0r1d[8] = rdtint_0n[8];
  assign rd_0r1d[9] = rdtint_0n[9];
  assign rd_0r1d[10] = rdtint_0n[10];
  assign rd_0r1d[11] = rdtint_0n[11];
  assign rd_0r1d[12] = rdtint_0n[12];
  assign rd_0r1d[13] = rdtint_0n[13];
  assign rd_0r1d[14] = rdtint_0n[14];
  assign rd_0r1d[15] = rdtint_0n[15];
  assign rd_0r1d[16] = rdtint_0n[16];
  assign rd_0r1d[17] = rdtint_0n[17];
  assign rd_0r1d[18] = rdtint_0n[18];
  assign rd_0r1d[19] = rdtint_0n[19];
  assign rd_0r1d[20] = rdtint_0n[20];
  assign rd_0r1d[21] = rdtint_0n[21];
  assign rd_0r1d[22] = rdtint_0n[22];
  assign rd_0r1d[23] = rdtint_0n[23];
  assign rd_0r1d[24] = rdtint_0n[24];
  assign rd_0r1d[25] = rdtint_0n[25];
  assign rd_0r1d[26] = rdtint_0n[26];
  assign rd_0r1d[27] = rdtint_0n[27];
  assign rd_0r1d[28] = rdtint_0n[28];
  assign rd_0r1d[29] = rdtint_0n[29];
  assign rd_0r1d[30] = rdtint_0n[30];
  assign rd_0r1d[31] = rdtint_0n[31];
  assign wg_1a = wgaint_1n;
  assign wgfint_1n[0] = wg_1r0d[0];
  assign wgfint_1n[1] = wg_1r0d[1];
  assign wgfint_1n[2] = wg_1r0d[2];
  assign wgfint_1n[3] = wg_1r0d[3];
  assign wgfint_1n[4] = wg_1r0d[4];
  assign wgfint_1n[5] = wg_1r0d[5];
  assign wgfint_1n[6] = wg_1r0d[6];
  assign wgfint_1n[7] = wg_1r0d[7];
  assign wgfint_1n[8] = wg_1r0d[8];
  assign wgfint_1n[9] = wg_1r0d[9];
  assign wgfint_1n[10] = wg_1r0d[10];
  assign wgfint_1n[11] = wg_1r0d[11];
  assign wgfint_1n[12] = wg_1r0d[12];
  assign wgfint_1n[13] = wg_1r0d[13];
  assign wgfint_1n[14] = wg_1r0d[14];
  assign wgfint_1n[15] = wg_1r0d[15];
  assign wgfint_1n[16] = wg_1r0d[16];
  assign wgfint_1n[17] = wg_1r0d[17];
  assign wgfint_1n[18] = wg_1r0d[18];
  assign wgfint_1n[19] = wg_1r0d[19];
  assign wgfint_1n[20] = wg_1r0d[20];
  assign wgfint_1n[21] = wg_1r0d[21];
  assign wgfint_1n[22] = wg_1r0d[22];
  assign wgfint_1n[23] = wg_1r0d[23];
  assign wgfint_1n[24] = wg_1r0d[24];
  assign wgfint_1n[25] = wg_1r0d[25];
  assign wgfint_1n[26] = wg_1r0d[26];
  assign wgfint_1n[27] = wg_1r0d[27];
  assign wgfint_1n[28] = wg_1r0d[28];
  assign wgfint_1n[29] = wg_1r0d[29];
  assign wgfint_1n[30] = wg_1r0d[30];
  assign wgfint_1n[31] = wg_1r0d[31];
  assign wgfint_1n[32] = wg_1r0d[32];
  assign wgfint_1n[33] = wg_1r0d[33];
  assign wgfint_1n[34] = wg_1r0d[34];
  assign wgfint_1n[35] = wg_1r0d[35];
  assign wgtint_1n[0] = wg_1r1d[0];
  assign wgtint_1n[1] = wg_1r1d[1];
  assign wgtint_1n[2] = wg_1r1d[2];
  assign wgtint_1n[3] = wg_1r1d[3];
  assign wgtint_1n[4] = wg_1r1d[4];
  assign wgtint_1n[5] = wg_1r1d[5];
  assign wgtint_1n[6] = wg_1r1d[6];
  assign wgtint_1n[7] = wg_1r1d[7];
  assign wgtint_1n[8] = wg_1r1d[8];
  assign wgtint_1n[9] = wg_1r1d[9];
  assign wgtint_1n[10] = wg_1r1d[10];
  assign wgtint_1n[11] = wg_1r1d[11];
  assign wgtint_1n[12] = wg_1r1d[12];
  assign wgtint_1n[13] = wg_1r1d[13];
  assign wgtint_1n[14] = wg_1r1d[14];
  assign wgtint_1n[15] = wg_1r1d[15];
  assign wgtint_1n[16] = wg_1r1d[16];
  assign wgtint_1n[17] = wg_1r1d[17];
  assign wgtint_1n[18] = wg_1r1d[18];
  assign wgtint_1n[19] = wg_1r1d[19];
  assign wgtint_1n[20] = wg_1r1d[20];
  assign wgtint_1n[21] = wg_1r1d[21];
  assign wgtint_1n[22] = wg_1r1d[22];
  assign wgtint_1n[23] = wg_1r1d[23];
  assign wgtint_1n[24] = wg_1r1d[24];
  assign wgtint_1n[25] = wg_1r1d[25];
  assign wgtint_1n[26] = wg_1r1d[26];
  assign wgtint_1n[27] = wg_1r1d[27];
  assign wgtint_1n[28] = wg_1r1d[28];
  assign wgtint_1n[29] = wg_1r1d[29];
  assign wgtint_1n[30] = wg_1r1d[30];
  assign wgtint_1n[31] = wg_1r1d[31];
  assign wgtint_1n[32] = wg_1r1d[32];
  assign wgtint_1n[33] = wg_1r1d[33];
  assign wgtint_1n[34] = wg_1r1d[34];
  assign wgtint_1n[35] = wg_1r1d[35];
  assign wg_0a = wgaint_0n;
  assign wgfint_0n[0] = wg_0r0d[0];
  assign wgfint_0n[1] = wg_0r0d[1];
  assign wgfint_0n[2] = wg_0r0d[2];
  assign wgfint_0n[3] = wg_0r0d[3];
  assign wgfint_0n[4] = wg_0r0d[4];
  assign wgfint_0n[5] = wg_0r0d[5];
  assign wgfint_0n[6] = wg_0r0d[6];
  assign wgfint_0n[7] = wg_0r0d[7];
  assign wgfint_0n[8] = wg_0r0d[8];
  assign wgfint_0n[9] = wg_0r0d[9];
  assign wgfint_0n[10] = wg_0r0d[10];
  assign wgfint_0n[11] = wg_0r0d[11];
  assign wgfint_0n[12] = wg_0r0d[12];
  assign wgfint_0n[13] = wg_0r0d[13];
  assign wgfint_0n[14] = wg_0r0d[14];
  assign wgfint_0n[15] = wg_0r0d[15];
  assign wgfint_0n[16] = wg_0r0d[16];
  assign wgfint_0n[17] = wg_0r0d[17];
  assign wgfint_0n[18] = wg_0r0d[18];
  assign wgfint_0n[19] = wg_0r0d[19];
  assign wgfint_0n[20] = wg_0r0d[20];
  assign wgfint_0n[21] = wg_0r0d[21];
  assign wgfint_0n[22] = wg_0r0d[22];
  assign wgfint_0n[23] = wg_0r0d[23];
  assign wgfint_0n[24] = wg_0r0d[24];
  assign wgfint_0n[25] = wg_0r0d[25];
  assign wgfint_0n[26] = wg_0r0d[26];
  assign wgfint_0n[27] = wg_0r0d[27];
  assign wgfint_0n[28] = wg_0r0d[28];
  assign wgfint_0n[29] = wg_0r0d[29];
  assign wgfint_0n[30] = wg_0r0d[30];
  assign wgfint_0n[31] = wg_0r0d[31];
  assign wgfint_0n[32] = wg_0r0d[32];
  assign wgfint_0n[33] = wg_0r0d[33];
  assign wgfint_0n[34] = wg_0r0d[34];
  assign wgfint_0n[35] = wg_0r0d[35];
  assign wgtint_0n[0] = wg_0r1d[0];
  assign wgtint_0n[1] = wg_0r1d[1];
  assign wgtint_0n[2] = wg_0r1d[2];
  assign wgtint_0n[3] = wg_0r1d[3];
  assign wgtint_0n[4] = wg_0r1d[4];
  assign wgtint_0n[5] = wg_0r1d[5];
  assign wgtint_0n[6] = wg_0r1d[6];
  assign wgtint_0n[7] = wg_0r1d[7];
  assign wgtint_0n[8] = wg_0r1d[8];
  assign wgtint_0n[9] = wg_0r1d[9];
  assign wgtint_0n[10] = wg_0r1d[10];
  assign wgtint_0n[11] = wg_0r1d[11];
  assign wgtint_0n[12] = wg_0r1d[12];
  assign wgtint_0n[13] = wg_0r1d[13];
  assign wgtint_0n[14] = wg_0r1d[14];
  assign wgtint_0n[15] = wg_0r1d[15];
  assign wgtint_0n[16] = wg_0r1d[16];
  assign wgtint_0n[17] = wg_0r1d[17];
  assign wgtint_0n[18] = wg_0r1d[18];
  assign wgtint_0n[19] = wg_0r1d[19];
  assign wgtint_0n[20] = wg_0r1d[20];
  assign wgtint_0n[21] = wg_0r1d[21];
  assign wgtint_0n[22] = wg_0r1d[22];
  assign wgtint_0n[23] = wg_0r1d[23];
  assign wgtint_0n[24] = wg_0r1d[24];
  assign wgtint_0n[25] = wg_0r1d[25];
  assign wgtint_0n[26] = wg_0r1d[26];
  assign wgtint_0n[27] = wg_0r1d[27];
  assign wgtint_0n[28] = wg_0r1d[28];
  assign wgtint_0n[29] = wg_0r1d[29];
  assign wgtint_0n[30] = wg_0r1d[30];
  assign wgtint_0n[31] = wg_0r1d[31];
  assign wgtint_0n[32] = wg_0r1d[32];
  assign wgtint_0n[33] = wg_0r1d[33];
  assign wgtint_0n[34] = wg_0r1d[34];
  assign wgtint_0n[35] = wg_0r1d[35];
  assign rg_0a = rgaint_0n;
  assign rgrint_0n = rg_0r;
  assign wgaint_1n = wd_1a;
  assign wd_1r = wdrint_1n;
  assign wgaint_0n = wd_0a;
  assign wd_0r = wdrint_0n;
  NOR2 I217 (nanyread_0n, rgrint_0n, rgaint_0n);
  AND2 I218 (rdtint_0n[0], rgrint_0n, dt_0n[3]);
  AND2 I219 (rdtint_0n[1], rgrint_0n, dt_0n[4]);
  AND2 I220 (rdtint_0n[2], rgrint_0n, dt_0n[5]);
  AND2 I221 (rdtint_0n[3], rgrint_0n, dt_0n[6]);
  AND2 I222 (rdtint_0n[4], rgrint_0n, dt_0n[7]);
  AND2 I223 (rdtint_0n[5], rgrint_0n, dt_0n[8]);
  AND2 I224 (rdtint_0n[6], rgrint_0n, dt_0n[9]);
  AND2 I225 (rdtint_0n[7], rgrint_0n, dt_0n[10]);
  AND2 I226 (rdtint_0n[8], rgrint_0n, dt_0n[11]);
  AND2 I227 (rdtint_0n[9], rgrint_0n, dt_0n[12]);
  AND2 I228 (rdtint_0n[10], rgrint_0n, dt_0n[13]);
  AND2 I229 (rdtint_0n[11], rgrint_0n, dt_0n[14]);
  AND2 I230 (rdtint_0n[12], rgrint_0n, dt_0n[15]);
  AND2 I231 (rdtint_0n[13], rgrint_0n, dt_0n[16]);
  AND2 I232 (rdtint_0n[14], rgrint_0n, dt_0n[17]);
  AND2 I233 (rdtint_0n[15], rgrint_0n, dt_0n[18]);
  AND2 I234 (rdtint_0n[16], rgrint_0n, dt_0n[19]);
  AND2 I235 (rdtint_0n[17], rgrint_0n, dt_0n[20]);
  AND2 I236 (rdtint_0n[18], rgrint_0n, dt_0n[21]);
  AND2 I237 (rdtint_0n[19], rgrint_0n, dt_0n[22]);
  AND2 I238 (rdtint_0n[20], rgrint_0n, dt_0n[23]);
  AND2 I239 (rdtint_0n[21], rgrint_0n, dt_0n[24]);
  AND2 I240 (rdtint_0n[22], rgrint_0n, dt_0n[25]);
  AND2 I241 (rdtint_0n[23], rgrint_0n, dt_0n[26]);
  AND2 I242 (rdtint_0n[24], rgrint_0n, dt_0n[27]);
  AND2 I243 (rdtint_0n[25], rgrint_0n, dt_0n[28]);
  AND2 I244 (rdtint_0n[26], rgrint_0n, dt_0n[29]);
  AND2 I245 (rdtint_0n[27], rgrint_0n, dt_0n[30]);
  AND2 I246 (rdtint_0n[28], rgrint_0n, dt_0n[31]);
  AND2 I247 (rdtint_0n[29], rgrint_0n, dt_0n[32]);
  AND2 I248 (rdtint_0n[30], rgrint_0n, dt_0n[33]);
  AND2 I249 (rdtint_0n[31], rgrint_0n, dt_0n[34]);
  AND2 I250 (rdfint_0n[0], rgrint_0n, df_0n[3]);
  AND2 I251 (rdfint_0n[1], rgrint_0n, df_0n[4]);
  AND2 I252 (rdfint_0n[2], rgrint_0n, df_0n[5]);
  AND2 I253 (rdfint_0n[3], rgrint_0n, df_0n[6]);
  AND2 I254 (rdfint_0n[4], rgrint_0n, df_0n[7]);
  AND2 I255 (rdfint_0n[5], rgrint_0n, df_0n[8]);
  AND2 I256 (rdfint_0n[6], rgrint_0n, df_0n[9]);
  AND2 I257 (rdfint_0n[7], rgrint_0n, df_0n[10]);
  AND2 I258 (rdfint_0n[8], rgrint_0n, df_0n[11]);
  AND2 I259 (rdfint_0n[9], rgrint_0n, df_0n[12]);
  AND2 I260 (rdfint_0n[10], rgrint_0n, df_0n[13]);
  AND2 I261 (rdfint_0n[11], rgrint_0n, df_0n[14]);
  AND2 I262 (rdfint_0n[12], rgrint_0n, df_0n[15]);
  AND2 I263 (rdfint_0n[13], rgrint_0n, df_0n[16]);
  AND2 I264 (rdfint_0n[14], rgrint_0n, df_0n[17]);
  AND2 I265 (rdfint_0n[15], rgrint_0n, df_0n[18]);
  AND2 I266 (rdfint_0n[16], rgrint_0n, df_0n[19]);
  AND2 I267 (rdfint_0n[17], rgrint_0n, df_0n[20]);
  AND2 I268 (rdfint_0n[18], rgrint_0n, df_0n[21]);
  AND2 I269 (rdfint_0n[19], rgrint_0n, df_0n[22]);
  AND2 I270 (rdfint_0n[20], rgrint_0n, df_0n[23]);
  AND2 I271 (rdfint_0n[21], rgrint_0n, df_0n[24]);
  AND2 I272 (rdfint_0n[22], rgrint_0n, df_0n[25]);
  AND2 I273 (rdfint_0n[23], rgrint_0n, df_0n[26]);
  AND2 I274 (rdfint_0n[24], rgrint_0n, df_0n[27]);
  AND2 I275 (rdfint_0n[25], rgrint_0n, df_0n[28]);
  AND2 I276 (rdfint_0n[26], rgrint_0n, df_0n[29]);
  AND2 I277 (rdfint_0n[27], rgrint_0n, df_0n[30]);
  AND2 I278 (rdfint_0n[28], rgrint_0n, df_0n[31]);
  AND2 I279 (rdfint_0n[29], rgrint_0n, df_0n[32]);
  AND2 I280 (rdfint_0n[30], rgrint_0n, df_0n[33]);
  AND2 I281 (rdfint_0n[31], rgrint_0n, df_0n[34]);
  C3 I282 (internal_0n[0], wc_1n, wacks_0n[35], wacks_0n[34]);
  C3 I283 (internal_0n[1], wacks_0n[33], wacks_0n[32], wacks_0n[31]);
  C3 I284 (internal_0n[2], wacks_0n[30], wacks_0n[29], wacks_0n[28]);
  C3 I285 (internal_0n[3], wacks_0n[27], wacks_0n[26], wacks_0n[25]);
  C3 I286 (internal_0n[4], wacks_0n[24], wacks_0n[23], wacks_0n[22]);
  C3 I287 (internal_0n[5], wacks_0n[21], wacks_0n[20], wacks_0n[19]);
  C3 I288 (internal_0n[6], wacks_0n[18], wacks_0n[17], wacks_0n[16]);
  C3 I289 (internal_0n[7], wacks_0n[15], wacks_0n[14], wacks_0n[13]);
  C3 I290 (internal_0n[8], wacks_0n[12], wacks_0n[11], wacks_0n[10]);
  C3 I291 (internal_0n[9], wacks_0n[9], wacks_0n[8], wacks_0n[7]);
  C3 I292 (internal_0n[10], wacks_0n[6], wacks_0n[5], wacks_0n[4]);
  C2 I293 (internal_0n[11], wacks_0n[3], wacks_0n[2]);
  C2 I294 (internal_0n[12], wacks_0n[1], wacks_0n[0]);
  C3 I295 (internal_0n[13], internal_0n[0], internal_0n[1], internal_0n[2]);
  C3 I296 (internal_0n[14], internal_0n[3], internal_0n[4], internal_0n[5]);
  C3 I297 (internal_0n[15], internal_0n[6], internal_0n[7], internal_0n[8]);
  C2 I298 (internal_0n[16], internal_0n[9], internal_0n[10]);
  C2 I299 (internal_0n[17], internal_0n[11], internal_0n[12]);
  C3 I300 (internal_0n[18], internal_0n[13], internal_0n[14], internal_0n[15]);
  C2 I301 (internal_0n[19], internal_0n[16], internal_0n[17]);
  C2 I302 (wdrint_1n, internal_0n[18], internal_0n[19]);
  C3 I303 (internal_0n[20], wc_0n, wacks_0n[35], wacks_0n[34]);
  C3 I304 (internal_0n[21], wacks_0n[33], wacks_0n[32], wacks_0n[31]);
  C3 I305 (internal_0n[22], wacks_0n[30], wacks_0n[29], wacks_0n[28]);
  C3 I306 (internal_0n[23], wacks_0n[27], wacks_0n[26], wacks_0n[25]);
  C3 I307 (internal_0n[24], wacks_0n[24], wacks_0n[23], wacks_0n[22]);
  C3 I308 (internal_0n[25], wacks_0n[21], wacks_0n[20], wacks_0n[19]);
  C3 I309 (internal_0n[26], wacks_0n[18], wacks_0n[17], wacks_0n[16]);
  C3 I310 (internal_0n[27], wacks_0n[15], wacks_0n[14], wacks_0n[13]);
  C3 I311 (internal_0n[28], wacks_0n[12], wacks_0n[11], wacks_0n[10]);
  C3 I312 (internal_0n[29], wacks_0n[9], wacks_0n[8], wacks_0n[7]);
  C3 I313 (internal_0n[30], wacks_0n[6], wacks_0n[5], wacks_0n[4]);
  C2 I314 (internal_0n[31], wacks_0n[3], wacks_0n[2]);
  C2 I315 (internal_0n[32], wacks_0n[1], wacks_0n[0]);
  C3 I316 (internal_0n[33], internal_0n[20], internal_0n[21], internal_0n[22]);
  C3 I317 (internal_0n[34], internal_0n[23], internal_0n[24], internal_0n[25]);
  C3 I318 (internal_0n[35], internal_0n[26], internal_0n[27], internal_0n[28]);
  C2 I319 (internal_0n[36], internal_0n[29], internal_0n[30]);
  C2 I320 (internal_0n[37], internal_0n[31], internal_0n[32]);
  C3 I321 (internal_0n[38], internal_0n[33], internal_0n[34], internal_0n[35]);
  C2 I322 (internal_0n[39], internal_0n[36], internal_0n[37]);
  C2 I323 (wdrint_0n, internal_0n[38], internal_0n[39]);
  OR2 I324 (wen_0n[35], wc_1n, wc_0n);
  OR2 I325 (wen_0n[34], wc_1n, wc_0n);
  OR2 I326 (wen_0n[33], wc_1n, wc_0n);
  OR2 I327 (wen_0n[32], wc_1n, wc_0n);
  OR2 I328 (wen_0n[31], wc_1n, wc_0n);
  OR2 I329 (wen_0n[30], wc_1n, wc_0n);
  OR2 I330 (wen_0n[29], wc_1n, wc_0n);
  OR2 I331 (wen_0n[28], wc_1n, wc_0n);
  OR2 I332 (wen_0n[27], wc_1n, wc_0n);
  OR2 I333 (wen_0n[26], wc_1n, wc_0n);
  OR2 I334 (wen_0n[25], wc_1n, wc_0n);
  OR2 I335 (wen_0n[24], wc_1n, wc_0n);
  OR2 I336 (wen_0n[23], wc_1n, wc_0n);
  OR2 I337 (wen_0n[22], wc_1n, wc_0n);
  OR2 I338 (wen_0n[21], wc_1n, wc_0n);
  OR2 I339 (wen_0n[20], wc_1n, wc_0n);
  OR2 I340 (wen_0n[19], wc_1n, wc_0n);
  OR2 I341 (wen_0n[18], wc_1n, wc_0n);
  OR2 I342 (wen_0n[17], wc_1n, wc_0n);
  OR2 I343 (wen_0n[16], wc_1n, wc_0n);
  OR2 I344 (wen_0n[15], wc_1n, wc_0n);
  OR2 I345 (wen_0n[14], wc_1n, wc_0n);
  OR2 I346 (wen_0n[13], wc_1n, wc_0n);
  OR2 I347 (wen_0n[12], wc_1n, wc_0n);
  OR2 I348 (wen_0n[11], wc_1n, wc_0n);
  OR2 I349 (wen_0n[10], wc_1n, wc_0n);
  OR2 I350 (wen_0n[9], wc_1n, wc_0n);
  OR2 I351 (wen_0n[8], wc_1n, wc_0n);
  OR2 I352 (wen_0n[7], wc_1n, wc_0n);
  OR2 I353 (wen_0n[6], wc_1n, wc_0n);
  OR2 I354 (wen_0n[5], wc_1n, wc_0n);
  OR2 I355 (wen_0n[4], wc_1n, wc_0n);
  OR2 I356 (wen_0n[3], wc_1n, wc_0n);
  OR2 I357 (wen_0n[2], wc_1n, wc_0n);
  OR2 I358 (wen_0n[1], wc_1n, wc_0n);
  OR2 I359 (wen_0n[0], wc_1n, wc_0n);
  OR2 I360 (wt_0n[35], git_1n[35], git_0n[35]);
  OR2 I361 (wt_0n[34], git_1n[34], git_0n[34]);
  OR2 I362 (wt_0n[33], git_1n[33], git_0n[33]);
  OR2 I363 (wt_0n[32], git_1n[32], git_0n[32]);
  OR2 I364 (wt_0n[31], git_1n[31], git_0n[31]);
  OR2 I365 (wt_0n[30], git_1n[30], git_0n[30]);
  OR2 I366 (wt_0n[29], git_1n[29], git_0n[29]);
  OR2 I367 (wt_0n[28], git_1n[28], git_0n[28]);
  OR2 I368 (wt_0n[27], git_1n[27], git_0n[27]);
  OR2 I369 (wt_0n[26], git_1n[26], git_0n[26]);
  OR2 I370 (wt_0n[25], git_1n[25], git_0n[25]);
  OR2 I371 (wt_0n[24], git_1n[24], git_0n[24]);
  OR2 I372 (wt_0n[23], git_1n[23], git_0n[23]);
  OR2 I373 (wt_0n[22], git_1n[22], git_0n[22]);
  OR2 I374 (wt_0n[21], git_1n[21], git_0n[21]);
  OR2 I375 (wt_0n[20], git_1n[20], git_0n[20]);
  OR2 I376 (wt_0n[19], git_1n[19], git_0n[19]);
  OR2 I377 (wt_0n[18], git_1n[18], git_0n[18]);
  OR2 I378 (wt_0n[17], git_1n[17], git_0n[17]);
  OR2 I379 (wt_0n[16], git_1n[16], git_0n[16]);
  OR2 I380 (wt_0n[15], git_1n[15], git_0n[15]);
  OR2 I381 (wt_0n[14], git_1n[14], git_0n[14]);
  OR2 I382 (wt_0n[13], git_1n[13], git_0n[13]);
  OR2 I383 (wt_0n[12], git_1n[12], git_0n[12]);
  OR2 I384 (wt_0n[11], git_1n[11], git_0n[11]);
  OR2 I385 (wt_0n[10], git_1n[10], git_0n[10]);
  OR2 I386 (wt_0n[9], git_1n[9], git_0n[9]);
  OR2 I387 (wt_0n[8], git_1n[8], git_0n[8]);
  OR2 I388 (wt_0n[7], git_1n[7], git_0n[7]);
  OR2 I389 (wt_0n[6], git_1n[6], git_0n[6]);
  OR2 I390 (wt_0n[5], git_1n[5], git_0n[5]);
  OR2 I391 (wt_0n[4], git_1n[4], git_0n[4]);
  OR2 I392 (wt_0n[3], git_1n[3], git_0n[3]);
  OR2 I393 (wt_0n[2], git_1n[2], git_0n[2]);
  OR2 I394 (wt_0n[1], git_1n[1], git_0n[1]);
  OR2 I395 (wt_0n[0], git_1n[0], git_0n[0]);
  OR2 I396 (wf_0n[35], gif_1n[35], gif_0n[35]);
  OR2 I397 (wf_0n[34], gif_1n[34], gif_0n[34]);
  OR2 I398 (wf_0n[33], gif_1n[33], gif_0n[33]);
  OR2 I399 (wf_0n[32], gif_1n[32], gif_0n[32]);
  OR2 I400 (wf_0n[31], gif_1n[31], gif_0n[31]);
  OR2 I401 (wf_0n[30], gif_1n[30], gif_0n[30]);
  OR2 I402 (wf_0n[29], gif_1n[29], gif_0n[29]);
  OR2 I403 (wf_0n[28], gif_1n[28], gif_0n[28]);
  OR2 I404 (wf_0n[27], gif_1n[27], gif_0n[27]);
  OR2 I405 (wf_0n[26], gif_1n[26], gif_0n[26]);
  OR2 I406 (wf_0n[25], gif_1n[25], gif_0n[25]);
  OR2 I407 (wf_0n[24], gif_1n[24], gif_0n[24]);
  OR2 I408 (wf_0n[23], gif_1n[23], gif_0n[23]);
  OR2 I409 (wf_0n[22], gif_1n[22], gif_0n[22]);
  OR2 I410 (wf_0n[21], gif_1n[21], gif_0n[21]);
  OR2 I411 (wf_0n[20], gif_1n[20], gif_0n[20]);
  OR2 I412 (wf_0n[19], gif_1n[19], gif_0n[19]);
  OR2 I413 (wf_0n[18], gif_1n[18], gif_0n[18]);
  OR2 I414 (wf_0n[17], gif_1n[17], gif_0n[17]);
  OR2 I415 (wf_0n[16], gif_1n[16], gif_0n[16]);
  OR2 I416 (wf_0n[15], gif_1n[15], gif_0n[15]);
  OR2 I417 (wf_0n[14], gif_1n[14], gif_0n[14]);
  OR2 I418 (wf_0n[13], gif_1n[13], gif_0n[13]);
  OR2 I419 (wf_0n[12], gif_1n[12], gif_0n[12]);
  OR2 I420 (wf_0n[11], gif_1n[11], gif_0n[11]);
  OR2 I421 (wf_0n[10], gif_1n[10], gif_0n[10]);
  OR2 I422 (wf_0n[9], gif_1n[9], gif_0n[9]);
  OR2 I423 (wf_0n[8], gif_1n[8], gif_0n[8]);
  OR2 I424 (wf_0n[7], gif_1n[7], gif_0n[7]);
  OR2 I425 (wf_0n[6], gif_1n[6], gif_0n[6]);
  OR2 I426 (wf_0n[5], gif_1n[5], gif_0n[5]);
  OR2 I427 (wf_0n[4], gif_1n[4], gif_0n[4]);
  OR2 I428 (wf_0n[3], gif_1n[3], gif_0n[3]);
  OR2 I429 (wf_0n[2], gif_1n[2], gif_0n[2]);
  OR2 I430 (wf_0n[1], gif_1n[1], gif_0n[1]);
  OR2 I431 (wf_0n[0], gif_1n[0], gif_0n[0]);
  AC2 I432 (ig_0n, igc_0n, nanyread_0n);
  AC2 I433 (ig_1n, igc_1n, nanyread_0n);
  assign igc_0n = wc_0n;
  assign igc_1n = wc_1n;
  AND2 I436 (git_1n[0], wgtint_1n[0], ig_1n);
  AND2 I437 (git_1n[1], wgtint_1n[1], ig_1n);
  AND2 I438 (git_1n[2], wgtint_1n[2], ig_1n);
  AND2 I439 (git_1n[3], wgtint_1n[3], ig_1n);
  AND2 I440 (git_1n[4], wgtint_1n[4], ig_1n);
  AND2 I441 (git_1n[5], wgtint_1n[5], ig_1n);
  AND2 I442 (git_1n[6], wgtint_1n[6], ig_1n);
  AND2 I443 (git_1n[7], wgtint_1n[7], ig_1n);
  AND2 I444 (git_1n[8], wgtint_1n[8], ig_1n);
  AND2 I445 (git_1n[9], wgtint_1n[9], ig_1n);
  AND2 I446 (git_1n[10], wgtint_1n[10], ig_1n);
  AND2 I447 (git_1n[11], wgtint_1n[11], ig_1n);
  AND2 I448 (git_1n[12], wgtint_1n[12], ig_1n);
  AND2 I449 (git_1n[13], wgtint_1n[13], ig_1n);
  AND2 I450 (git_1n[14], wgtint_1n[14], ig_1n);
  AND2 I451 (git_1n[15], wgtint_1n[15], ig_1n);
  AND2 I452 (git_1n[16], wgtint_1n[16], ig_1n);
  AND2 I453 (git_1n[17], wgtint_1n[17], ig_1n);
  AND2 I454 (git_1n[18], wgtint_1n[18], ig_1n);
  AND2 I455 (git_1n[19], wgtint_1n[19], ig_1n);
  AND2 I456 (git_1n[20], wgtint_1n[20], ig_1n);
  AND2 I457 (git_1n[21], wgtint_1n[21], ig_1n);
  AND2 I458 (git_1n[22], wgtint_1n[22], ig_1n);
  AND2 I459 (git_1n[23], wgtint_1n[23], ig_1n);
  AND2 I460 (git_1n[24], wgtint_1n[24], ig_1n);
  AND2 I461 (git_1n[25], wgtint_1n[25], ig_1n);
  AND2 I462 (git_1n[26], wgtint_1n[26], ig_1n);
  AND2 I463 (git_1n[27], wgtint_1n[27], ig_1n);
  AND2 I464 (git_1n[28], wgtint_1n[28], ig_1n);
  AND2 I465 (git_1n[29], wgtint_1n[29], ig_1n);
  AND2 I466 (git_1n[30], wgtint_1n[30], ig_1n);
  AND2 I467 (git_1n[31], wgtint_1n[31], ig_1n);
  AND2 I468 (git_1n[32], wgtint_1n[32], ig_1n);
  AND2 I469 (git_1n[33], wgtint_1n[33], ig_1n);
  AND2 I470 (git_1n[34], wgtint_1n[34], ig_1n);
  AND2 I471 (git_1n[35], wgtint_1n[35], ig_1n);
  AND2 I472 (git_0n[0], wgtint_0n[0], ig_0n);
  AND2 I473 (git_0n[1], wgtint_0n[1], ig_0n);
  AND2 I474 (git_0n[2], wgtint_0n[2], ig_0n);
  AND2 I475 (git_0n[3], wgtint_0n[3], ig_0n);
  AND2 I476 (git_0n[4], wgtint_0n[4], ig_0n);
  AND2 I477 (git_0n[5], wgtint_0n[5], ig_0n);
  AND2 I478 (git_0n[6], wgtint_0n[6], ig_0n);
  AND2 I479 (git_0n[7], wgtint_0n[7], ig_0n);
  AND2 I480 (git_0n[8], wgtint_0n[8], ig_0n);
  AND2 I481 (git_0n[9], wgtint_0n[9], ig_0n);
  AND2 I482 (git_0n[10], wgtint_0n[10], ig_0n);
  AND2 I483 (git_0n[11], wgtint_0n[11], ig_0n);
  AND2 I484 (git_0n[12], wgtint_0n[12], ig_0n);
  AND2 I485 (git_0n[13], wgtint_0n[13], ig_0n);
  AND2 I486 (git_0n[14], wgtint_0n[14], ig_0n);
  AND2 I487 (git_0n[15], wgtint_0n[15], ig_0n);
  AND2 I488 (git_0n[16], wgtint_0n[16], ig_0n);
  AND2 I489 (git_0n[17], wgtint_0n[17], ig_0n);
  AND2 I490 (git_0n[18], wgtint_0n[18], ig_0n);
  AND2 I491 (git_0n[19], wgtint_0n[19], ig_0n);
  AND2 I492 (git_0n[20], wgtint_0n[20], ig_0n);
  AND2 I493 (git_0n[21], wgtint_0n[21], ig_0n);
  AND2 I494 (git_0n[22], wgtint_0n[22], ig_0n);
  AND2 I495 (git_0n[23], wgtint_0n[23], ig_0n);
  AND2 I496 (git_0n[24], wgtint_0n[24], ig_0n);
  AND2 I497 (git_0n[25], wgtint_0n[25], ig_0n);
  AND2 I498 (git_0n[26], wgtint_0n[26], ig_0n);
  AND2 I499 (git_0n[27], wgtint_0n[27], ig_0n);
  AND2 I500 (git_0n[28], wgtint_0n[28], ig_0n);
  AND2 I501 (git_0n[29], wgtint_0n[29], ig_0n);
  AND2 I502 (git_0n[30], wgtint_0n[30], ig_0n);
  AND2 I503 (git_0n[31], wgtint_0n[31], ig_0n);
  AND2 I504 (git_0n[32], wgtint_0n[32], ig_0n);
  AND2 I505 (git_0n[33], wgtint_0n[33], ig_0n);
  AND2 I506 (git_0n[34], wgtint_0n[34], ig_0n);
  AND2 I507 (git_0n[35], wgtint_0n[35], ig_0n);
  AND2 I508 (gif_1n[0], wgfint_1n[0], ig_1n);
  AND2 I509 (gif_1n[1], wgfint_1n[1], ig_1n);
  AND2 I510 (gif_1n[2], wgfint_1n[2], ig_1n);
  AND2 I511 (gif_1n[3], wgfint_1n[3], ig_1n);
  AND2 I512 (gif_1n[4], wgfint_1n[4], ig_1n);
  AND2 I513 (gif_1n[5], wgfint_1n[5], ig_1n);
  AND2 I514 (gif_1n[6], wgfint_1n[6], ig_1n);
  AND2 I515 (gif_1n[7], wgfint_1n[7], ig_1n);
  AND2 I516 (gif_1n[8], wgfint_1n[8], ig_1n);
  AND2 I517 (gif_1n[9], wgfint_1n[9], ig_1n);
  AND2 I518 (gif_1n[10], wgfint_1n[10], ig_1n);
  AND2 I519 (gif_1n[11], wgfint_1n[11], ig_1n);
  AND2 I520 (gif_1n[12], wgfint_1n[12], ig_1n);
  AND2 I521 (gif_1n[13], wgfint_1n[13], ig_1n);
  AND2 I522 (gif_1n[14], wgfint_1n[14], ig_1n);
  AND2 I523 (gif_1n[15], wgfint_1n[15], ig_1n);
  AND2 I524 (gif_1n[16], wgfint_1n[16], ig_1n);
  AND2 I525 (gif_1n[17], wgfint_1n[17], ig_1n);
  AND2 I526 (gif_1n[18], wgfint_1n[18], ig_1n);
  AND2 I527 (gif_1n[19], wgfint_1n[19], ig_1n);
  AND2 I528 (gif_1n[20], wgfint_1n[20], ig_1n);
  AND2 I529 (gif_1n[21], wgfint_1n[21], ig_1n);
  AND2 I530 (gif_1n[22], wgfint_1n[22], ig_1n);
  AND2 I531 (gif_1n[23], wgfint_1n[23], ig_1n);
  AND2 I532 (gif_1n[24], wgfint_1n[24], ig_1n);
  AND2 I533 (gif_1n[25], wgfint_1n[25], ig_1n);
  AND2 I534 (gif_1n[26], wgfint_1n[26], ig_1n);
  AND2 I535 (gif_1n[27], wgfint_1n[27], ig_1n);
  AND2 I536 (gif_1n[28], wgfint_1n[28], ig_1n);
  AND2 I537 (gif_1n[29], wgfint_1n[29], ig_1n);
  AND2 I538 (gif_1n[30], wgfint_1n[30], ig_1n);
  AND2 I539 (gif_1n[31], wgfint_1n[31], ig_1n);
  AND2 I540 (gif_1n[32], wgfint_1n[32], ig_1n);
  AND2 I541 (gif_1n[33], wgfint_1n[33], ig_1n);
  AND2 I542 (gif_1n[34], wgfint_1n[34], ig_1n);
  AND2 I543 (gif_1n[35], wgfint_1n[35], ig_1n);
  AND2 I544 (gif_0n[0], wgfint_0n[0], ig_0n);
  AND2 I545 (gif_0n[1], wgfint_0n[1], ig_0n);
  AND2 I546 (gif_0n[2], wgfint_0n[2], ig_0n);
  AND2 I547 (gif_0n[3], wgfint_0n[3], ig_0n);
  AND2 I548 (gif_0n[4], wgfint_0n[4], ig_0n);
  AND2 I549 (gif_0n[5], wgfint_0n[5], ig_0n);
  AND2 I550 (gif_0n[6], wgfint_0n[6], ig_0n);
  AND2 I551 (gif_0n[7], wgfint_0n[7], ig_0n);
  AND2 I552 (gif_0n[8], wgfint_0n[8], ig_0n);
  AND2 I553 (gif_0n[9], wgfint_0n[9], ig_0n);
  AND2 I554 (gif_0n[10], wgfint_0n[10], ig_0n);
  AND2 I555 (gif_0n[11], wgfint_0n[11], ig_0n);
  AND2 I556 (gif_0n[12], wgfint_0n[12], ig_0n);
  AND2 I557 (gif_0n[13], wgfint_0n[13], ig_0n);
  AND2 I558 (gif_0n[14], wgfint_0n[14], ig_0n);
  AND2 I559 (gif_0n[15], wgfint_0n[15], ig_0n);
  AND2 I560 (gif_0n[16], wgfint_0n[16], ig_0n);
  AND2 I561 (gif_0n[17], wgfint_0n[17], ig_0n);
  AND2 I562 (gif_0n[18], wgfint_0n[18], ig_0n);
  AND2 I563 (gif_0n[19], wgfint_0n[19], ig_0n);
  AND2 I564 (gif_0n[20], wgfint_0n[20], ig_0n);
  AND2 I565 (gif_0n[21], wgfint_0n[21], ig_0n);
  AND2 I566 (gif_0n[22], wgfint_0n[22], ig_0n);
  AND2 I567 (gif_0n[23], wgfint_0n[23], ig_0n);
  AND2 I568 (gif_0n[24], wgfint_0n[24], ig_0n);
  AND2 I569 (gif_0n[25], wgfint_0n[25], ig_0n);
  AND2 I570 (gif_0n[26], wgfint_0n[26], ig_0n);
  AND2 I571 (gif_0n[27], wgfint_0n[27], ig_0n);
  AND2 I572 (gif_0n[28], wgfint_0n[28], ig_0n);
  AND2 I573 (gif_0n[29], wgfint_0n[29], ig_0n);
  AND2 I574 (gif_0n[30], wgfint_0n[30], ig_0n);
  AND2 I575 (gif_0n[31], wgfint_0n[31], ig_0n);
  AND2 I576 (gif_0n[32], wgfint_0n[32], ig_0n);
  AND2 I577 (gif_0n[33], wgfint_0n[33], ig_0n);
  AND2 I578 (gif_0n[34], wgfint_0n[34], ig_0n);
  AND2 I579 (gif_0n[35], wgfint_0n[35], ig_0n);
  C3 I580 (internal_0n[40], complete1628_0n[0], complete1628_0n[1], complete1628_0n[2]);
  C3 I581 (internal_0n[41], complete1628_0n[3], complete1628_0n[4], complete1628_0n[5]);
  C3 I582 (internal_0n[42], complete1628_0n[6], complete1628_0n[7], complete1628_0n[8]);
  C3 I583 (internal_0n[43], complete1628_0n[9], complete1628_0n[10], complete1628_0n[11]);
  C3 I584 (internal_0n[44], complete1628_0n[12], complete1628_0n[13], complete1628_0n[14]);
  C3 I585 (internal_0n[45], complete1628_0n[15], complete1628_0n[16], complete1628_0n[17]);
  C3 I586 (internal_0n[46], complete1628_0n[18], complete1628_0n[19], complete1628_0n[20]);
  C3 I587 (internal_0n[47], complete1628_0n[21], complete1628_0n[22], complete1628_0n[23]);
  C3 I588 (internal_0n[48], complete1628_0n[24], complete1628_0n[25], complete1628_0n[26]);
  C3 I589 (internal_0n[49], complete1628_0n[27], complete1628_0n[28], complete1628_0n[29]);
  C3 I590 (internal_0n[50], complete1628_0n[30], complete1628_0n[31], complete1628_0n[32]);
  C3 I591 (internal_0n[51], complete1628_0n[33], complete1628_0n[34], complete1628_0n[35]);
  C3 I592 (internal_0n[52], internal_0n[40], internal_0n[41], internal_0n[42]);
  C3 I593 (internal_0n[53], internal_0n[43], internal_0n[44], internal_0n[45]);
  C3 I594 (internal_0n[54], internal_0n[46], internal_0n[47], internal_0n[48]);
  C3 I595 (internal_0n[55], internal_0n[49], internal_0n[50], internal_0n[51]);
  C2 I596 (internal_0n[56], internal_0n[52], internal_0n[53]);
  C2 I597 (internal_0n[57], internal_0n[54], internal_0n[55]);
  C2 I598 (wc_1n, internal_0n[56], internal_0n[57]);
  OR2 I599 (complete1628_0n[0], wgfint_1n[0], wgtint_1n[0]);
  OR2 I600 (complete1628_0n[1], wgfint_1n[1], wgtint_1n[1]);
  OR2 I601 (complete1628_0n[2], wgfint_1n[2], wgtint_1n[2]);
  OR2 I602 (complete1628_0n[3], wgfint_1n[3], wgtint_1n[3]);
  OR2 I603 (complete1628_0n[4], wgfint_1n[4], wgtint_1n[4]);
  OR2 I604 (complete1628_0n[5], wgfint_1n[5], wgtint_1n[5]);
  OR2 I605 (complete1628_0n[6], wgfint_1n[6], wgtint_1n[6]);
  OR2 I606 (complete1628_0n[7], wgfint_1n[7], wgtint_1n[7]);
  OR2 I607 (complete1628_0n[8], wgfint_1n[8], wgtint_1n[8]);
  OR2 I608 (complete1628_0n[9], wgfint_1n[9], wgtint_1n[9]);
  OR2 I609 (complete1628_0n[10], wgfint_1n[10], wgtint_1n[10]);
  OR2 I610 (complete1628_0n[11], wgfint_1n[11], wgtint_1n[11]);
  OR2 I611 (complete1628_0n[12], wgfint_1n[12], wgtint_1n[12]);
  OR2 I612 (complete1628_0n[13], wgfint_1n[13], wgtint_1n[13]);
  OR2 I613 (complete1628_0n[14], wgfint_1n[14], wgtint_1n[14]);
  OR2 I614 (complete1628_0n[15], wgfint_1n[15], wgtint_1n[15]);
  OR2 I615 (complete1628_0n[16], wgfint_1n[16], wgtint_1n[16]);
  OR2 I616 (complete1628_0n[17], wgfint_1n[17], wgtint_1n[17]);
  OR2 I617 (complete1628_0n[18], wgfint_1n[18], wgtint_1n[18]);
  OR2 I618 (complete1628_0n[19], wgfint_1n[19], wgtint_1n[19]);
  OR2 I619 (complete1628_0n[20], wgfint_1n[20], wgtint_1n[20]);
  OR2 I620 (complete1628_0n[21], wgfint_1n[21], wgtint_1n[21]);
  OR2 I621 (complete1628_0n[22], wgfint_1n[22], wgtint_1n[22]);
  OR2 I622 (complete1628_0n[23], wgfint_1n[23], wgtint_1n[23]);
  OR2 I623 (complete1628_0n[24], wgfint_1n[24], wgtint_1n[24]);
  OR2 I624 (complete1628_0n[25], wgfint_1n[25], wgtint_1n[25]);
  OR2 I625 (complete1628_0n[26], wgfint_1n[26], wgtint_1n[26]);
  OR2 I626 (complete1628_0n[27], wgfint_1n[27], wgtint_1n[27]);
  OR2 I627 (complete1628_0n[28], wgfint_1n[28], wgtint_1n[28]);
  OR2 I628 (complete1628_0n[29], wgfint_1n[29], wgtint_1n[29]);
  OR2 I629 (complete1628_0n[30], wgfint_1n[30], wgtint_1n[30]);
  OR2 I630 (complete1628_0n[31], wgfint_1n[31], wgtint_1n[31]);
  OR2 I631 (complete1628_0n[32], wgfint_1n[32], wgtint_1n[32]);
  OR2 I632 (complete1628_0n[33], wgfint_1n[33], wgtint_1n[33]);
  OR2 I633 (complete1628_0n[34], wgfint_1n[34], wgtint_1n[34]);
  OR2 I634 (complete1628_0n[35], wgfint_1n[35], wgtint_1n[35]);
  C3 I635 (internal_0n[58], complete1627_0n[0], complete1627_0n[1], complete1627_0n[2]);
  C3 I636 (internal_0n[59], complete1627_0n[3], complete1627_0n[4], complete1627_0n[5]);
  C3 I637 (internal_0n[60], complete1627_0n[6], complete1627_0n[7], complete1627_0n[8]);
  C3 I638 (internal_0n[61], complete1627_0n[9], complete1627_0n[10], complete1627_0n[11]);
  C3 I639 (internal_0n[62], complete1627_0n[12], complete1627_0n[13], complete1627_0n[14]);
  C3 I640 (internal_0n[63], complete1627_0n[15], complete1627_0n[16], complete1627_0n[17]);
  C3 I641 (internal_0n[64], complete1627_0n[18], complete1627_0n[19], complete1627_0n[20]);
  C3 I642 (internal_0n[65], complete1627_0n[21], complete1627_0n[22], complete1627_0n[23]);
  C3 I643 (internal_0n[66], complete1627_0n[24], complete1627_0n[25], complete1627_0n[26]);
  C3 I644 (internal_0n[67], complete1627_0n[27], complete1627_0n[28], complete1627_0n[29]);
  C3 I645 (internal_0n[68], complete1627_0n[30], complete1627_0n[31], complete1627_0n[32]);
  C3 I646 (internal_0n[69], complete1627_0n[33], complete1627_0n[34], complete1627_0n[35]);
  C3 I647 (internal_0n[70], internal_0n[58], internal_0n[59], internal_0n[60]);
  C3 I648 (internal_0n[71], internal_0n[61], internal_0n[62], internal_0n[63]);
  C3 I649 (internal_0n[72], internal_0n[64], internal_0n[65], internal_0n[66]);
  C3 I650 (internal_0n[73], internal_0n[67], internal_0n[68], internal_0n[69]);
  C2 I651 (internal_0n[74], internal_0n[70], internal_0n[71]);
  C2 I652 (internal_0n[75], internal_0n[72], internal_0n[73]);
  C2 I653 (wc_0n, internal_0n[74], internal_0n[75]);
  OR2 I654 (complete1627_0n[0], wgfint_0n[0], wgtint_0n[0]);
  OR2 I655 (complete1627_0n[1], wgfint_0n[1], wgtint_0n[1]);
  OR2 I656 (complete1627_0n[2], wgfint_0n[2], wgtint_0n[2]);
  OR2 I657 (complete1627_0n[3], wgfint_0n[3], wgtint_0n[3]);
  OR2 I658 (complete1627_0n[4], wgfint_0n[4], wgtint_0n[4]);
  OR2 I659 (complete1627_0n[5], wgfint_0n[5], wgtint_0n[5]);
  OR2 I660 (complete1627_0n[6], wgfint_0n[6], wgtint_0n[6]);
  OR2 I661 (complete1627_0n[7], wgfint_0n[7], wgtint_0n[7]);
  OR2 I662 (complete1627_0n[8], wgfint_0n[8], wgtint_0n[8]);
  OR2 I663 (complete1627_0n[9], wgfint_0n[9], wgtint_0n[9]);
  OR2 I664 (complete1627_0n[10], wgfint_0n[10], wgtint_0n[10]);
  OR2 I665 (complete1627_0n[11], wgfint_0n[11], wgtint_0n[11]);
  OR2 I666 (complete1627_0n[12], wgfint_0n[12], wgtint_0n[12]);
  OR2 I667 (complete1627_0n[13], wgfint_0n[13], wgtint_0n[13]);
  OR2 I668 (complete1627_0n[14], wgfint_0n[14], wgtint_0n[14]);
  OR2 I669 (complete1627_0n[15], wgfint_0n[15], wgtint_0n[15]);
  OR2 I670 (complete1627_0n[16], wgfint_0n[16], wgtint_0n[16]);
  OR2 I671 (complete1627_0n[17], wgfint_0n[17], wgtint_0n[17]);
  OR2 I672 (complete1627_0n[18], wgfint_0n[18], wgtint_0n[18]);
  OR2 I673 (complete1627_0n[19], wgfint_0n[19], wgtint_0n[19]);
  OR2 I674 (complete1627_0n[20], wgfint_0n[20], wgtint_0n[20]);
  OR2 I675 (complete1627_0n[21], wgfint_0n[21], wgtint_0n[21]);
  OR2 I676 (complete1627_0n[22], wgfint_0n[22], wgtint_0n[22]);
  OR2 I677 (complete1627_0n[23], wgfint_0n[23], wgtint_0n[23]);
  OR2 I678 (complete1627_0n[24], wgfint_0n[24], wgtint_0n[24]);
  OR2 I679 (complete1627_0n[25], wgfint_0n[25], wgtint_0n[25]);
  OR2 I680 (complete1627_0n[26], wgfint_0n[26], wgtint_0n[26]);
  OR2 I681 (complete1627_0n[27], wgfint_0n[27], wgtint_0n[27]);
  OR2 I682 (complete1627_0n[28], wgfint_0n[28], wgtint_0n[28]);
  OR2 I683 (complete1627_0n[29], wgfint_0n[29], wgtint_0n[29]);
  OR2 I684 (complete1627_0n[30], wgfint_0n[30], wgtint_0n[30]);
  OR2 I685 (complete1627_0n[31], wgfint_0n[31], wgtint_0n[31]);
  OR2 I686 (complete1627_0n[32], wgfint_0n[32], wgtint_0n[32]);
  OR2 I687 (complete1627_0n[33], wgfint_0n[33], wgtint_0n[33]);
  OR2 I688 (complete1627_0n[34], wgfint_0n[34], wgtint_0n[34]);
  OR2 I689 (complete1627_0n[35], wgfint_0n[35], wgtint_0n[35]);
  AO22 I690 (wacks_0n[35], gf1625_0n[35], df_0n[35], gt1626_0n[35], dt_0n[35]);
  NOR2 I691 (dt_0n[35], df_0n[35], gf1625_0n[35]);
  NOR3 I692 (df_0n[35], dt_0n[35], gt1626_0n[35], init_0n);
  AND2 I693 (gt1626_0n[35], wt_0n[35], wen_0n[35]);
  AND2 I694 (gf1625_0n[35], wf_0n[35], wen_0n[35]);
  AO22 I695 (wacks_0n[34], gf1625_0n[34], df_0n[34], gt1626_0n[34], dt_0n[34]);
  NOR2 I696 (dt_0n[34], df_0n[34], gf1625_0n[34]);
  NOR3 I697 (df_0n[34], dt_0n[34], gt1626_0n[34], init_0n);
  AND2 I698 (gt1626_0n[34], wt_0n[34], wen_0n[34]);
  AND2 I699 (gf1625_0n[34], wf_0n[34], wen_0n[34]);
  AO22 I700 (wacks_0n[33], gf1625_0n[33], df_0n[33], gt1626_0n[33], dt_0n[33]);
  NOR2 I701 (dt_0n[33], df_0n[33], gf1625_0n[33]);
  NOR3 I702 (df_0n[33], dt_0n[33], gt1626_0n[33], init_0n);
  AND2 I703 (gt1626_0n[33], wt_0n[33], wen_0n[33]);
  AND2 I704 (gf1625_0n[33], wf_0n[33], wen_0n[33]);
  AO22 I705 (wacks_0n[32], gf1625_0n[32], df_0n[32], gt1626_0n[32], dt_0n[32]);
  NOR2 I706 (dt_0n[32], df_0n[32], gf1625_0n[32]);
  NOR3 I707 (df_0n[32], dt_0n[32], gt1626_0n[32], init_0n);
  AND2 I708 (gt1626_0n[32], wt_0n[32], wen_0n[32]);
  AND2 I709 (gf1625_0n[32], wf_0n[32], wen_0n[32]);
  AO22 I710 (wacks_0n[31], gf1625_0n[31], df_0n[31], gt1626_0n[31], dt_0n[31]);
  NOR2 I711 (dt_0n[31], df_0n[31], gf1625_0n[31]);
  NOR3 I712 (df_0n[31], dt_0n[31], gt1626_0n[31], init_0n);
  AND2 I713 (gt1626_0n[31], wt_0n[31], wen_0n[31]);
  AND2 I714 (gf1625_0n[31], wf_0n[31], wen_0n[31]);
  AO22 I715 (wacks_0n[30], gf1625_0n[30], df_0n[30], gt1626_0n[30], dt_0n[30]);
  NOR2 I716 (dt_0n[30], df_0n[30], gf1625_0n[30]);
  NOR3 I717 (df_0n[30], dt_0n[30], gt1626_0n[30], init_0n);
  AND2 I718 (gt1626_0n[30], wt_0n[30], wen_0n[30]);
  AND2 I719 (gf1625_0n[30], wf_0n[30], wen_0n[30]);
  AO22 I720 (wacks_0n[29], gf1625_0n[29], df_0n[29], gt1626_0n[29], dt_0n[29]);
  NOR2 I721 (dt_0n[29], df_0n[29], gf1625_0n[29]);
  NOR3 I722 (df_0n[29], dt_0n[29], gt1626_0n[29], init_0n);
  AND2 I723 (gt1626_0n[29], wt_0n[29], wen_0n[29]);
  AND2 I724 (gf1625_0n[29], wf_0n[29], wen_0n[29]);
  AO22 I725 (wacks_0n[28], gf1625_0n[28], df_0n[28], gt1626_0n[28], dt_0n[28]);
  NOR2 I726 (dt_0n[28], df_0n[28], gf1625_0n[28]);
  NOR3 I727 (df_0n[28], dt_0n[28], gt1626_0n[28], init_0n);
  AND2 I728 (gt1626_0n[28], wt_0n[28], wen_0n[28]);
  AND2 I729 (gf1625_0n[28], wf_0n[28], wen_0n[28]);
  AO22 I730 (wacks_0n[27], gf1625_0n[27], df_0n[27], gt1626_0n[27], dt_0n[27]);
  NOR2 I731 (dt_0n[27], df_0n[27], gf1625_0n[27]);
  NOR3 I732 (df_0n[27], dt_0n[27], gt1626_0n[27], init_0n);
  AND2 I733 (gt1626_0n[27], wt_0n[27], wen_0n[27]);
  AND2 I734 (gf1625_0n[27], wf_0n[27], wen_0n[27]);
  AO22 I735 (wacks_0n[26], gf1625_0n[26], df_0n[26], gt1626_0n[26], dt_0n[26]);
  NOR2 I736 (dt_0n[26], df_0n[26], gf1625_0n[26]);
  NOR3 I737 (df_0n[26], dt_0n[26], gt1626_0n[26], init_0n);
  AND2 I738 (gt1626_0n[26], wt_0n[26], wen_0n[26]);
  AND2 I739 (gf1625_0n[26], wf_0n[26], wen_0n[26]);
  AO22 I740 (wacks_0n[25], gf1625_0n[25], df_0n[25], gt1626_0n[25], dt_0n[25]);
  NOR2 I741 (dt_0n[25], df_0n[25], gf1625_0n[25]);
  NOR3 I742 (df_0n[25], dt_0n[25], gt1626_0n[25], init_0n);
  AND2 I743 (gt1626_0n[25], wt_0n[25], wen_0n[25]);
  AND2 I744 (gf1625_0n[25], wf_0n[25], wen_0n[25]);
  AO22 I745 (wacks_0n[24], gf1625_0n[24], df_0n[24], gt1626_0n[24], dt_0n[24]);
  NOR2 I746 (dt_0n[24], df_0n[24], gf1625_0n[24]);
  NOR3 I747 (df_0n[24], dt_0n[24], gt1626_0n[24], init_0n);
  AND2 I748 (gt1626_0n[24], wt_0n[24], wen_0n[24]);
  AND2 I749 (gf1625_0n[24], wf_0n[24], wen_0n[24]);
  AO22 I750 (wacks_0n[23], gf1625_0n[23], df_0n[23], gt1626_0n[23], dt_0n[23]);
  NOR2 I751 (dt_0n[23], df_0n[23], gf1625_0n[23]);
  NOR3 I752 (df_0n[23], dt_0n[23], gt1626_0n[23], init_0n);
  AND2 I753 (gt1626_0n[23], wt_0n[23], wen_0n[23]);
  AND2 I754 (gf1625_0n[23], wf_0n[23], wen_0n[23]);
  AO22 I755 (wacks_0n[22], gf1625_0n[22], df_0n[22], gt1626_0n[22], dt_0n[22]);
  NOR2 I756 (dt_0n[22], df_0n[22], gf1625_0n[22]);
  NOR3 I757 (df_0n[22], dt_0n[22], gt1626_0n[22], init_0n);
  AND2 I758 (gt1626_0n[22], wt_0n[22], wen_0n[22]);
  AND2 I759 (gf1625_0n[22], wf_0n[22], wen_0n[22]);
  AO22 I760 (wacks_0n[21], gf1625_0n[21], df_0n[21], gt1626_0n[21], dt_0n[21]);
  NOR2 I761 (dt_0n[21], df_0n[21], gf1625_0n[21]);
  NOR3 I762 (df_0n[21], dt_0n[21], gt1626_0n[21], init_0n);
  AND2 I763 (gt1626_0n[21], wt_0n[21], wen_0n[21]);
  AND2 I764 (gf1625_0n[21], wf_0n[21], wen_0n[21]);
  AO22 I765 (wacks_0n[20], gf1625_0n[20], df_0n[20], gt1626_0n[20], dt_0n[20]);
  NOR2 I766 (dt_0n[20], df_0n[20], gf1625_0n[20]);
  NOR3 I767 (df_0n[20], dt_0n[20], gt1626_0n[20], init_0n);
  AND2 I768 (gt1626_0n[20], wt_0n[20], wen_0n[20]);
  AND2 I769 (gf1625_0n[20], wf_0n[20], wen_0n[20]);
  AO22 I770 (wacks_0n[19], gf1625_0n[19], df_0n[19], gt1626_0n[19], dt_0n[19]);
  NOR2 I771 (dt_0n[19], df_0n[19], gf1625_0n[19]);
  NOR3 I772 (df_0n[19], dt_0n[19], gt1626_0n[19], init_0n);
  AND2 I773 (gt1626_0n[19], wt_0n[19], wen_0n[19]);
  AND2 I774 (gf1625_0n[19], wf_0n[19], wen_0n[19]);
  AO22 I775 (wacks_0n[18], gf1625_0n[18], df_0n[18], gt1626_0n[18], dt_0n[18]);
  NOR2 I776 (dt_0n[18], df_0n[18], gf1625_0n[18]);
  NOR3 I777 (df_0n[18], dt_0n[18], gt1626_0n[18], init_0n);
  AND2 I778 (gt1626_0n[18], wt_0n[18], wen_0n[18]);
  AND2 I779 (gf1625_0n[18], wf_0n[18], wen_0n[18]);
  AO22 I780 (wacks_0n[17], gf1625_0n[17], df_0n[17], gt1626_0n[17], dt_0n[17]);
  NOR2 I781 (dt_0n[17], df_0n[17], gf1625_0n[17]);
  NOR3 I782 (df_0n[17], dt_0n[17], gt1626_0n[17], init_0n);
  AND2 I783 (gt1626_0n[17], wt_0n[17], wen_0n[17]);
  AND2 I784 (gf1625_0n[17], wf_0n[17], wen_0n[17]);
  AO22 I785 (wacks_0n[16], gf1625_0n[16], df_0n[16], gt1626_0n[16], dt_0n[16]);
  NOR2 I786 (dt_0n[16], df_0n[16], gf1625_0n[16]);
  NOR3 I787 (df_0n[16], dt_0n[16], gt1626_0n[16], init_0n);
  AND2 I788 (gt1626_0n[16], wt_0n[16], wen_0n[16]);
  AND2 I789 (gf1625_0n[16], wf_0n[16], wen_0n[16]);
  AO22 I790 (wacks_0n[15], gf1625_0n[15], df_0n[15], gt1626_0n[15], dt_0n[15]);
  NOR2 I791 (dt_0n[15], df_0n[15], gf1625_0n[15]);
  NOR3 I792 (df_0n[15], dt_0n[15], gt1626_0n[15], init_0n);
  AND2 I793 (gt1626_0n[15], wt_0n[15], wen_0n[15]);
  AND2 I794 (gf1625_0n[15], wf_0n[15], wen_0n[15]);
  AO22 I795 (wacks_0n[14], gf1625_0n[14], df_0n[14], gt1626_0n[14], dt_0n[14]);
  NOR2 I796 (dt_0n[14], df_0n[14], gf1625_0n[14]);
  NOR3 I797 (df_0n[14], dt_0n[14], gt1626_0n[14], init_0n);
  AND2 I798 (gt1626_0n[14], wt_0n[14], wen_0n[14]);
  AND2 I799 (gf1625_0n[14], wf_0n[14], wen_0n[14]);
  AO22 I800 (wacks_0n[13], gf1625_0n[13], df_0n[13], gt1626_0n[13], dt_0n[13]);
  NOR2 I801 (dt_0n[13], df_0n[13], gf1625_0n[13]);
  NOR3 I802 (df_0n[13], dt_0n[13], gt1626_0n[13], init_0n);
  AND2 I803 (gt1626_0n[13], wt_0n[13], wen_0n[13]);
  AND2 I804 (gf1625_0n[13], wf_0n[13], wen_0n[13]);
  AO22 I805 (wacks_0n[12], gf1625_0n[12], df_0n[12], gt1626_0n[12], dt_0n[12]);
  NOR2 I806 (dt_0n[12], df_0n[12], gf1625_0n[12]);
  NOR3 I807 (df_0n[12], dt_0n[12], gt1626_0n[12], init_0n);
  AND2 I808 (gt1626_0n[12], wt_0n[12], wen_0n[12]);
  AND2 I809 (gf1625_0n[12], wf_0n[12], wen_0n[12]);
  AO22 I810 (wacks_0n[11], gf1625_0n[11], df_0n[11], gt1626_0n[11], dt_0n[11]);
  NOR2 I811 (dt_0n[11], df_0n[11], gf1625_0n[11]);
  NOR3 I812 (df_0n[11], dt_0n[11], gt1626_0n[11], init_0n);
  AND2 I813 (gt1626_0n[11], wt_0n[11], wen_0n[11]);
  AND2 I814 (gf1625_0n[11], wf_0n[11], wen_0n[11]);
  AO22 I815 (wacks_0n[10], gf1625_0n[10], df_0n[10], gt1626_0n[10], dt_0n[10]);
  NOR2 I816 (dt_0n[10], df_0n[10], gf1625_0n[10]);
  NOR3 I817 (df_0n[10], dt_0n[10], gt1626_0n[10], init_0n);
  AND2 I818 (gt1626_0n[10], wt_0n[10], wen_0n[10]);
  AND2 I819 (gf1625_0n[10], wf_0n[10], wen_0n[10]);
  AO22 I820 (wacks_0n[9], gf1625_0n[9], df_0n[9], gt1626_0n[9], dt_0n[9]);
  NOR2 I821 (dt_0n[9], df_0n[9], gf1625_0n[9]);
  NOR3 I822 (df_0n[9], dt_0n[9], gt1626_0n[9], init_0n);
  AND2 I823 (gt1626_0n[9], wt_0n[9], wen_0n[9]);
  AND2 I824 (gf1625_0n[9], wf_0n[9], wen_0n[9]);
  AO22 I825 (wacks_0n[8], gf1625_0n[8], df_0n[8], gt1626_0n[8], dt_0n[8]);
  NOR2 I826 (dt_0n[8], df_0n[8], gf1625_0n[8]);
  NOR3 I827 (df_0n[8], dt_0n[8], gt1626_0n[8], init_0n);
  AND2 I828 (gt1626_0n[8], wt_0n[8], wen_0n[8]);
  AND2 I829 (gf1625_0n[8], wf_0n[8], wen_0n[8]);
  AO22 I830 (wacks_0n[7], gf1625_0n[7], df_0n[7], gt1626_0n[7], dt_0n[7]);
  NOR2 I831 (dt_0n[7], df_0n[7], gf1625_0n[7]);
  NOR3 I832 (df_0n[7], dt_0n[7], gt1626_0n[7], init_0n);
  AND2 I833 (gt1626_0n[7], wt_0n[7], wen_0n[7]);
  AND2 I834 (gf1625_0n[7], wf_0n[7], wen_0n[7]);
  AO22 I835 (wacks_0n[6], gf1625_0n[6], df_0n[6], gt1626_0n[6], dt_0n[6]);
  NOR2 I836 (dt_0n[6], df_0n[6], gf1625_0n[6]);
  NOR3 I837 (df_0n[6], dt_0n[6], gt1626_0n[6], init_0n);
  AND2 I838 (gt1626_0n[6], wt_0n[6], wen_0n[6]);
  AND2 I839 (gf1625_0n[6], wf_0n[6], wen_0n[6]);
  AO22 I840 (wacks_0n[5], gf1625_0n[5], df_0n[5], gt1626_0n[5], dt_0n[5]);
  NOR2 I841 (dt_0n[5], df_0n[5], gf1625_0n[5]);
  NOR3 I842 (df_0n[5], dt_0n[5], gt1626_0n[5], init_0n);
  AND2 I843 (gt1626_0n[5], wt_0n[5], wen_0n[5]);
  AND2 I844 (gf1625_0n[5], wf_0n[5], wen_0n[5]);
  AO22 I845 (wacks_0n[4], gf1625_0n[4], df_0n[4], gt1626_0n[4], dt_0n[4]);
  NOR2 I846 (dt_0n[4], df_0n[4], gf1625_0n[4]);
  NOR3 I847 (df_0n[4], dt_0n[4], gt1626_0n[4], init_0n);
  AND2 I848 (gt1626_0n[4], wt_0n[4], wen_0n[4]);
  AND2 I849 (gf1625_0n[4], wf_0n[4], wen_0n[4]);
  AO22 I850 (wacks_0n[3], gf1625_0n[3], df_0n[3], gt1626_0n[3], dt_0n[3]);
  NOR2 I851 (dt_0n[3], df_0n[3], gf1625_0n[3]);
  NOR3 I852 (df_0n[3], dt_0n[3], gt1626_0n[3], init_0n);
  AND2 I853 (gt1626_0n[3], wt_0n[3], wen_0n[3]);
  AND2 I854 (gf1625_0n[3], wf_0n[3], wen_0n[3]);
  AO22 I855 (wacks_0n[2], gf1625_0n[2], df_0n[2], gt1626_0n[2], dt_0n[2]);
  NOR2 I856 (dt_0n[2], df_0n[2], gf1625_0n[2]);
  NOR3 I857 (df_0n[2], dt_0n[2], gt1626_0n[2], init_0n);
  AND2 I858 (gt1626_0n[2], wt_0n[2], wen_0n[2]);
  AND2 I859 (gf1625_0n[2], wf_0n[2], wen_0n[2]);
  AO22 I860 (wacks_0n[1], gf1625_0n[1], df_0n[1], gt1626_0n[1], dt_0n[1]);
  NOR2 I861 (dt_0n[1], df_0n[1], gf1625_0n[1]);
  NOR3 I862 (df_0n[1], dt_0n[1], gt1626_0n[1], init_0n);
  AND2 I863 (gt1626_0n[1], wt_0n[1], wen_0n[1]);
  AND2 I864 (gf1625_0n[1], wf_0n[1], wen_0n[1]);
  AO22 I865 (wacks_0n[0], gf1625_0n[0], df_0n[0], gt1626_0n[0], dt_0n[0]);
  NOR2 I866 (dt_0n[0], df_0n[0], gf1625_0n[0]);
  NOR3 I867 (df_0n[0], dt_0n[0], gt1626_0n[0], init_0n);
  AND2 I868 (gt1626_0n[0], wt_0n[0], wen_0n[0]);
  AND2 I869 (gf1625_0n[0], wf_0n[0], wen_0n[0]);
  GIVE_INIT I870 (init_0n, initialise);
endmodule

module Balsa_signAdj (
  go_0r, go_0a,
  mType_0r0d, mType_0r1d, mType_0a,
  a_0r0d, a_0r1d, a_0a,
  b_0r0d, b_0r1d, b_0a,
  c_0r0d, c_0r1d, c_0a,
  aa_0r0d, aa_0r1d, aa_0a,
  ba_0r0d, ba_0r1d, ba_0a,
  ca_0r0d, ca_0r1d, ca_0a,
  mlength_0r0d, mlength_0r1d, mlength_0a,
  macc_0r0d, macc_0r1d, macc_0a,
  initialise
);
  input go_0r;
  output go_0a;
  input [2:0] mType_0r0d;
  input [2:0] mType_0r1d;
  output mType_0a;
  input [31:0] a_0r0d;
  input [31:0] a_0r1d;
  output a_0a;
  input [31:0] b_0r0d;
  input [31:0] b_0r1d;
  output b_0a;
  input [31:0] c_0r0d;
  input [31:0] c_0r1d;
  output c_0a;
  output [34:0] aa_0r0d;
  output [34:0] aa_0r1d;
  input aa_0a;
  output [35:0] ba_0r0d;
  output [35:0] ba_0r1d;
  input ba_0a;
  output [34:0] ca_0r0d;
  output [34:0] ca_0r1d;
  input ca_0a;
  output mlength_0r0d;
  output mlength_0r1d;
  input mlength_0a;
  output macc_0r0d;
  output macc_0r1d;
  input macc_0a;
  input initialise;
  wire [1:0] c86_r0d;
  wire [1:0] c86_r1d;
  wire c86_a;
  wire [1:0] c85_r0d;
  wire [1:0] c85_r1d;
  wire c85_a;
  wire [1:0] c84_r0d;
  wire [1:0] c84_r1d;
  wire c84_a;
  wire [1:0] c83_r0d;
  wire [1:0] c83_r1d;
  wire c83_a;
  wire c82_r;
  wire c82_a;
  wire [35:0] c81_r0d;
  wire [35:0] c81_r1d;
  wire c81_a;
  wire [35:0] c80_r0d;
  wire [35:0] c80_r1d;
  wire c80_a;
  wire c79_r;
  wire c79_a;
  wire [35:0] c78_r0d;
  wire [35:0] c78_r1d;
  wire c78_a;
  wire c77_r;
  wire c77_a;
  wire [1:0] c76_r0d;
  wire [1:0] c76_r1d;
  wire c76_a;
  wire [1:0] c75_r0d;
  wire [1:0] c75_r1d;
  wire c75_a;
  wire [1:0] c74_r0d;
  wire [1:0] c74_r1d;
  wire c74_a;
  wire [1:0] c73_r0d;
  wire [1:0] c73_r1d;
  wire c73_a;
  wire c72_r;
  wire c72_a;
  wire [34:0] c71_r0d;
  wire [34:0] c71_r1d;
  wire c71_a;
  wire [34:0] c70_r0d;
  wire [34:0] c70_r1d;
  wire c70_a;
  wire c69_r;
  wire c69_a;
  wire [34:0] c68_r0d;
  wire [34:0] c68_r1d;
  wire c68_a;
  wire c67_r;
  wire c67_a;
  wire c66_r;
  wire c66_a;
  wire c65_r;
  wire c65_a;
  wire c64_r;
  wire c64_a;
  wire c63_r;
  wire c63_a;
  wire c62_r;
  wire c62_a;
  wire c61_r;
  wire c61_a;
  wire c60_r;
  wire c60_a;
  wire [31:0] c59_r0d;
  wire [31:0] c59_r1d;
  wire c59_a;
  wire c58_r;
  wire c58_a;
  wire [31:0] c57_r0d;
  wire [31:0] c57_r1d;
  wire c57_a;
  wire c56_r;
  wire c56_a;
  wire [31:0] c55_r0d;
  wire [31:0] c55_r1d;
  wire c55_a;
  wire c54_r;
  wire c54_a;
  wire [2:0] c53_r0d;
  wire [2:0] c53_r1d;
  wire c53_a;
  wire c52_r;
  wire c52_a;
  wire c51_r;
  wire c51_a;
  wire c50_r;
  wire c50_a;
  wire c49_r0d;
  wire c49_r1d;
  wire c49_a;
  wire c48_r;
  wire c48_a;
  wire c47_r;
  wire c47_a;
  wire c46_r0d;
  wire c46_r1d;
  wire c46_a;
  wire c45_r;
  wire c45_a;
  wire c44_r;
  wire c44_a;
  wire [31:0] c43_r0d;
  wire [31:0] c43_r1d;
  wire c43_a;
  wire [34:0] c42_r0d;
  wire [34:0] c42_r1d;
  wire c42_a;
  wire c41_r;
  wire c41_a;
  wire c40_r;
  wire c40_a;
  wire c39_r;
  wire c39_a;
  wire c38_r;
  wire c38_a;
  wire c37_r;
  wire c37_a;
  wire [32:0] c36_r0d;
  wire [32:0] c36_r1d;
  wire c36_a;
  wire c35_r;
  wire c35_a;
  wire [31:0] c34_r0d;
  wire [31:0] c34_r1d;
  wire c34_a;
  wire c33_r0d;
  wire c33_r1d;
  wire c33_a;
  wire c32_r;
  wire c32_a;
  wire [35:0] c31_r0d;
  wire [35:0] c31_r1d;
  wire c31_a;
  wire c30_r;
  wire c30_a;
  wire c29_r;
  wire c29_a;
  wire [31:0] c28_r0d;
  wire [31:0] c28_r1d;
  wire c28_a;
  wire [34:0] c27_r0d;
  wire [34:0] c27_r1d;
  wire c27_a;
  wire c26_r;
  wire c26_a;
  wire c25_r;
  wire c25_a;
  wire c24_r;
  wire c24_a;
  wire c23_r;
  wire c23_a;
  wire [32:0] c22_r0d;
  wire [32:0] c22_r1d;
  wire c22_a;
  wire c21_r;
  wire c21_a;
  wire [31:0] c20_r0d;
  wire [31:0] c20_r1d;
  wire c20_a;
  wire c19_r0d;
  wire c19_r1d;
  wire c19_a;
  wire c18_r;
  wire c18_a;
  wire [35:0] c17_r0d;
  wire [35:0] c17_r1d;
  wire c17_a;
  wire c16_r;
  wire c16_a;
  wire c15_r;
  wire c15_a;
  wire [31:0] c14_r0d;
  wire [31:0] c14_r1d;
  wire c14_a;
  wire [34:0] c13_r0d;
  wire [34:0] c13_r1d;
  wire c13_a;
  wire c12_r;
  wire c12_a;
  wire [2:0] c11_r0d;
  wire [2:0] c11_r1d;
  wire c11_a;
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I0 (c49_r0d, c49_r1d, c49_a, c51_r, c51_a, macc_0r0d, macc_0r1d, macc_0a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I1 (c46_r0d, c46_r1d, c46_a, c48_r, c48_a, mlength_0r0d, mlength_0r1d, mlength_0a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I2 (c42_r0d, c42_r1d, c42_a, c45_r, c45_a, ca_0r0d, ca_0r1d, ca_0a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I3 (c86_r0d, c86_r1d, c86_a, c24_r, c24_a, c38_r, c38_a, initialise);
  BrzJ_l11__280_202_29 I4 (c82_r, c82_a, c85_r0d, c85_r1d, c85_a, c86_r0d, c86_r1d, c86_a, initialise);
  BrzM_2_2 I5 (c83_r0d, c83_r1d, c83_a, c84_r0d, c84_r1d, c84_a, c85_r0d, c85_r1d, c85_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I6 (c79_r, c79_a, c84_r0d, c84_r1d, c84_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I7 (c77_r, c77_a, c83_r0d, c83_r1d, c83_a);
  BrzF_36_l32__28_280_200_29_20_280_2036_29__m44m I8 (c81_r0d, c81_r1d, c81_a, c82_r, c82_a, ba_0r0d, ba_0r1d, ba_0a, initialise);
  BrzM_36_2 I9 (c78_r0d, c78_r1d, c78_a, c80_r0d, c80_r1d, c80_a, c81_r0d, c81_r1d, c81_a, initialise);
  BrzF_36_l32__28_280_200_29_20_280_2036_29__m44m I10 (c31_r0d, c31_r1d, c31_a, c79_r, c79_a, c80_r0d, c80_r1d, c80_a, initialise);
  BrzF_36_l32__28_280_200_29_20_280_2036_29__m44m I11 (c17_r0d, c17_r1d, c17_a, c77_r, c77_a, c78_r0d, c78_r1d, c78_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I12 (c76_r0d, c76_r1d, c76_a, c16_r, c16_a, c30_r, c30_a, initialise);
  BrzJ_l11__280_202_29 I13 (c72_r, c72_a, c75_r0d, c75_r1d, c75_a, c76_r0d, c76_r1d, c76_a, initialise);
  BrzM_2_2 I14 (c73_r0d, c73_r1d, c73_a, c74_r0d, c74_r1d, c74_a, c75_r0d, c75_r1d, c75_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I15 (c69_r, c69_a, c74_r0d, c74_r1d, c74_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I16 (c67_r, c67_a, c73_r0d, c73_r1d, c73_a);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I17 (c71_r0d, c71_r1d, c71_a, c72_r, c72_a, aa_0r0d, aa_0r1d, aa_0a, initialise);
  BrzM_35_2 I18 (c68_r0d, c68_r1d, c68_a, c70_r0d, c70_r1d, c70_a, c71_r0d, c71_r1d, c71_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I19 (c27_r0d, c27_r1d, c27_a, c69_r, c69_a, c70_r0d, c70_r1d, c70_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I20 (c13_r0d, c13_r1d, c13_a, c67_r, c67_a, c68_r0d, c68_r1d, c68_a, initialise);
  BrzJ_l12__2832_200_29 I21 (c_0r0d, c_0r1d, c_0a, c65_r, c65_a, c59_r0d, c59_r1d, c59_a, initialise);
  BrzJ_l12__2832_200_29 I22 (b_0r0d, b_0r1d, b_0a, c64_r, c64_a, c57_r0d, c57_r1d, c57_a, initialise);
  BrzJ_l12__2832_200_29 I23 (a_0r0d, a_0r1d, a_0a, c63_r, c63_a, c55_r0d, c55_r1d, c55_a, initialise);
  BrzJ_l11__283_200_29 I24 (mType_0r0d, mType_0r1d, mType_0a, c62_r, c62_a, c53_r0d, c53_r1d, c53_a, initialise);
  BrzM_0_2 I25 (go_0r, go_0a, c52_r, c52_a, c66_r, c66_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I26 (c66_r, c66_a, c62_r, c62_a, c63_r, c63_a, c64_r, c64_a, c65_r, c65_a, initialise);
  BrzJ_l19__280_200_200_200_29 I27 (c54_r, c54_a, c56_r, c56_a, c58_r, c58_a, c60_r, c60_a, c61_r, c61_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I28 (c59_r0d, c59_r1d, c59_a, c60_r, c60_a, c44_r, c44_a, c43_r0d, c43_r1d, c43_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m81m I29 (c57_r0d, c57_r1d, c57_a, c58_r, c58_a, c21_r, c21_a, c35_r, c35_a, c20_r0d, c20_r1d, c20_a, c34_r0d, c34_r1d, c34_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m81m I30 (c55_r0d, c55_r1d, c55_a, c56_r, c56_a, c15_r, c15_a, c29_r, c29_a, c14_r0d, c14_r1d, c14_a, c28_r0d, c28_r1d, c28_a, initialise);
  BrzV_3_l6__28_29_l23__28_28_280_203_29_29__m76m I31 (c53_r0d, c53_r1d, c53_a, c54_r, c54_a, c12_r, c12_a, c47_r, c47_a, c50_r, c50_a, c11_r0d, c11_r1d, c11_a, c46_r0d, c46_r1d, c46_a, c49_r0d, c49_r1d, c49_a, initialise);
  BrzJ_l19__280_200_200_200_29 I32 (c41_r, c41_a, c45_r, c45_a, c48_r, c48_a, c51_r, c51_a, c52_r, c52_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I33 (c61_r, c61_a, c12_r, c12_a, c44_r, c44_a, c47_r, c47_a, c50_r, c50_a, initialise);
  BrzO_32_35_l76__28_28num_203_200_29_20_28a_m51m I34 (c43_r0d, c43_r1d, c43_a, c42_r0d, c42_r1d, c42_a);
  BrzM_0_2 I35 (c26_r, c26_a, c40_r, c40_a, c41_r, c41_a, initialise);
  BrzS_3_l11__280_203_29_l151__28_28_28_281__m65m I36 (c11_r0d, c11_r1d, c11_a, c25_r, c25_a, c39_r, c39_a, initialise);
  BrzJ_l11__280_200_29 I37 (c30_r, c30_a, c38_r, c38_a, c40_r, c40_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I38 (c39_r, c39_a, c29_r, c29_a, c37_r, c37_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I39 (c37_r, c37_a, c32_r, c32_a, c35_r, c35_a, initialise);
  BrzO_33_36_l76__28_28num_203_200_29_20_28a_m54m I40 (c36_r0d, c36_r1d, c36_a, c31_r0d, c31_r1d, c31_a);
  BrzJ_l12__281_2032_29 I41 (c33_r0d, c33_r1d, c33_a, c34_r0d, c34_r1d, c34_a, c36_r0d, c36_r1d, c36_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I42 (c32_r, c32_a, c33_r0d, c33_r1d, c33_a);
  BrzO_32_35_l76__28_28num_203_200_29_20_28a_m51m I43 (c28_r0d, c28_r1d, c28_a, c27_r0d, c27_r1d, c27_a);
  BrzJ_l11__280_200_29 I44 (c16_r, c16_a, c24_r, c24_a, c26_r, c26_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I45 (c25_r, c25_a, c15_r, c15_a, c23_r, c23_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I46 (c23_r, c23_a, c18_r, c18_a, c21_r, c21_a, initialise);
  BrzO_33_36_l91__28_28app_203_20_280_2032_2_m53m I47 (c22_r0d, c22_r1d, c22_a, c17_r0d, c17_r1d, c17_a);
  BrzJ_l12__281_2032_29 I48 (c19_r0d, c19_r1d, c19_a, c20_r0d, c20_r1d, c20_a, c22_r0d, c22_r1d, c22_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I49 (c18_r, c18_a, c19_r0d, c19_r1d, c19_a);
  BrzO_32_35_l91__28_28app_203_20_280_2031_2_m50m I50 (c14_r0d, c14_r1d, c14_a, c13_r0d, c13_r1d, c13_a);
endmodule

module Balsa_doByPass (
  go_0r, go_0a,
  bH_0r0d, bH_0r1d, bH_0a,
  bL_0r0d, bL_0r1d, bL_0a,
  bpH_0r0d, bpH_0r1d, bpH_0a,
  bpL_0r0d, bpL_0r1d, bpL_0a,
  bmZ_0r0d, bmZ_0r1d, bmZ_0a,
  bmN_0r0d, bmN_0r1d, bmN_0a,
  mpH_0r0d, mpH_0r1d, mpH_0a,
  mpL_0r0d, mpL_0r1d, mpL_0a,
  mZ_0r0d, mZ_0r1d, mZ_0a,
  mN_0r0d, mN_0r1d, mN_0a,
  initialise
);
  input go_0r;
  output go_0a;
  input bH_0r0d;
  input bH_0r1d;
  output bH_0a;
  input bL_0r0d;
  input bL_0r1d;
  output bL_0a;
  input [31:0] bpH_0r0d;
  input [31:0] bpH_0r1d;
  output bpH_0a;
  input [31:0] bpL_0r0d;
  input [31:0] bpL_0r1d;
  output bpL_0a;
  input bmZ_0r0d;
  input bmZ_0r1d;
  output bmZ_0a;
  input bmN_0r0d;
  input bmN_0r1d;
  output bmN_0a;
  output [31:0] mpH_0r0d;
  output [31:0] mpH_0r1d;
  input mpH_0a;
  output [31:0] mpL_0r0d;
  output [31:0] mpL_0r1d;
  input mpL_0a;
  output mZ_0r0d;
  output mZ_0r1d;
  input mZ_0a;
  output mN_0r0d;
  output mN_0r1d;
  input mN_0a;
  input initialise;
  wire [1:0] c105_r0d;
  wire [1:0] c105_r1d;
  wire c105_a;
  wire [1:0] c104_r0d;
  wire [1:0] c104_r1d;
  wire c104_a;
  wire [1:0] c103_r0d;
  wire [1:0] c103_r1d;
  wire c103_a;
  wire [1:0] c102_r0d;
  wire [1:0] c102_r1d;
  wire c102_a;
  wire c101_r;
  wire c101_a;
  wire c100_r0d;
  wire c100_r1d;
  wire c100_a;
  wire c99_r0d;
  wire c99_r1d;
  wire c99_a;
  wire c98_r;
  wire c98_a;
  wire c97_r0d;
  wire c97_r1d;
  wire c97_a;
  wire c96_r;
  wire c96_a;
  wire [1:0] c95_r0d;
  wire [1:0] c95_r1d;
  wire c95_a;
  wire [1:0] c94_r0d;
  wire [1:0] c94_r1d;
  wire c94_a;
  wire [1:0] c93_r0d;
  wire [1:0] c93_r1d;
  wire c93_a;
  wire [1:0] c92_r0d;
  wire [1:0] c92_r1d;
  wire c92_a;
  wire c91_r;
  wire c91_a;
  wire c90_r0d;
  wire c90_r1d;
  wire c90_a;
  wire c89_r0d;
  wire c89_r1d;
  wire c89_a;
  wire c88_r;
  wire c88_a;
  wire c87_r0d;
  wire c87_r1d;
  wire c87_a;
  wire c86_r;
  wire c86_a;
  wire [1:0] c85_r0d;
  wire [1:0] c85_r1d;
  wire c85_a;
  wire [1:0] c84_r0d;
  wire [1:0] c84_r1d;
  wire c84_a;
  wire [1:0] c83_r0d;
  wire [1:0] c83_r1d;
  wire c83_a;
  wire [1:0] c82_r0d;
  wire [1:0] c82_r1d;
  wire c82_a;
  wire c81_r;
  wire c81_a;
  wire [31:0] c80_r0d;
  wire [31:0] c80_r1d;
  wire c80_a;
  wire [31:0] c79_r0d;
  wire [31:0] c79_r1d;
  wire c79_a;
  wire c78_r;
  wire c78_a;
  wire [31:0] c77_r0d;
  wire [31:0] c77_r1d;
  wire c77_a;
  wire c76_r;
  wire c76_a;
  wire [1:0] c75_r0d;
  wire [1:0] c75_r1d;
  wire c75_a;
  wire [1:0] c74_r0d;
  wire [1:0] c74_r1d;
  wire c74_a;
  wire [1:0] c73_r0d;
  wire [1:0] c73_r1d;
  wire c73_a;
  wire [1:0] c72_r0d;
  wire [1:0] c72_r1d;
  wire c72_a;
  wire c71_r;
  wire c71_a;
  wire [31:0] c70_r0d;
  wire [31:0] c70_r1d;
  wire c70_a;
  wire [31:0] c69_r0d;
  wire [31:0] c69_r1d;
  wire c69_a;
  wire c68_r;
  wire c68_a;
  wire [31:0] c67_r0d;
  wire [31:0] c67_r1d;
  wire c67_a;
  wire c66_r;
  wire c66_a;
  wire c65_r;
  wire c65_a;
  wire c64_r;
  wire c64_a;
  wire c63_r;
  wire c63_a;
  wire c62_r;
  wire c62_a;
  wire c61_r;
  wire c61_a;
  wire c60_r0d;
  wire c60_r1d;
  wire c60_a;
  wire c59_r;
  wire c59_a;
  wire c58_r0d;
  wire c58_r1d;
  wire c58_a;
  wire c57_r;
  wire c57_a;
  wire c56_r;
  wire c56_a;
  wire c55_r;
  wire c55_a;
  wire c54_r;
  wire c54_a;
  wire c53_r;
  wire c53_a;
  wire [31:0] c52_r0d;
  wire [31:0] c52_r1d;
  wire c52_a;
  wire c51_r;
  wire c51_a;
  wire c50_r;
  wire c50_a;
  wire c49_r;
  wire c49_a;
  wire c48_r0d;
  wire c48_r1d;
  wire c48_a;
  wire c47_r;
  wire c47_a;
  wire c46_r0d;
  wire c46_r1d;
  wire c46_a;
  wire c45_r;
  wire c45_a;
  wire c44_r;
  wire c44_a;
  wire c43_r0d;
  wire c43_r1d;
  wire c43_a;
  wire c42_r;
  wire c42_a;
  wire c41_r;
  wire c41_a;
  wire [31:0] c40_r0d;
  wire [31:0] c40_r1d;
  wire c40_a;
  wire c39_r;
  wire c39_a;
  wire c38_r;
  wire c38_a;
  wire c37_r;
  wire c37_a;
  wire c36_r;
  wire c36_a;
  wire c35_r;
  wire c35_a;
  wire c34_r;
  wire c34_a;
  wire [31:0] c33_r0d;
  wire [31:0] c33_r1d;
  wire c33_a;
  wire c32_r;
  wire c32_a;
  wire [31:0] c31_r0d;
  wire [31:0] c31_r1d;
  wire c31_a;
  wire c30_r;
  wire c30_a;
  wire c29_r;
  wire c29_a;
  wire c28_r0d;
  wire c28_r1d;
  wire c28_a;
  wire c27_r;
  wire c27_a;
  wire c26_r;
  wire c26_a;
  wire c25_r0d;
  wire c25_r1d;
  wire c25_a;
  wire c24_r;
  wire c24_a;
  wire c23_r0d;
  wire c23_r1d;
  wire c23_a;
  wire c22_r;
  wire c22_a;
  wire c21_r;
  wire c21_a;
  wire c20_r0d;
  wire c20_r1d;
  wire c20_a;
  wire c19_r;
  wire c19_a;
  wire c18_r0d;
  wire c18_r1d;
  wire c18_a;
  wire c17_r;
  wire c17_a;
  wire c16_r;
  wire c16_a;
  wire [31:0] c15_r0d;
  wire [31:0] c15_r1d;
  wire c15_a;
  wire c14_r;
  wire c14_a;
  wire [31:0] c13_r0d;
  wire [31:0] c13_r1d;
  wire c13_a;
  wire c12_r0d;
  wire c12_r1d;
  wire c12_a;
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I0 (c105_r0d, c105_r1d, c105_a, c24_r, c24_a, c47_r, c47_a, initialise);
  BrzJ_l11__280_202_29 I1 (c101_r, c101_a, c104_r0d, c104_r1d, c104_a, c105_r0d, c105_r1d, c105_a, initialise);
  BrzM_2_2 I2 (c102_r0d, c102_r1d, c102_a, c103_r0d, c103_r1d, c103_a, c104_r0d, c104_r1d, c104_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I3 (c98_r, c98_a, c103_r0d, c103_r1d, c103_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I4 (c96_r, c96_a, c102_r0d, c102_r1d, c102_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I5 (c100_r0d, c100_r1d, c100_a, c101_r, c101_a, mN_0r0d, mN_0r1d, mN_0a, initialise);
  BrzM_1_2 I6 (c97_r0d, c97_r1d, c97_a, c99_r0d, c99_r1d, c99_a, c100_r0d, c100_r1d, c100_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I7 (c46_r0d, c46_r1d, c46_a, c98_r, c98_a, c99_r0d, c99_r1d, c99_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I8 (c23_r0d, c23_r1d, c23_a, c96_r, c96_a, c97_r0d, c97_r1d, c97_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I9 (c95_r0d, c95_r1d, c95_a, c19_r, c19_a, c44_r, c44_a, initialise);
  BrzJ_l11__280_202_29 I10 (c91_r, c91_a, c94_r0d, c94_r1d, c94_a, c95_r0d, c95_r1d, c95_a, initialise);
  BrzM_2_2 I11 (c92_r0d, c92_r1d, c92_a, c93_r0d, c93_r1d, c93_a, c94_r0d, c94_r1d, c94_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I12 (c88_r, c88_a, c93_r0d, c93_r1d, c93_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I13 (c86_r, c86_a, c92_r0d, c92_r1d, c92_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I14 (c90_r0d, c90_r1d, c90_a, c91_r, c91_a, mZ_0r0d, mZ_0r1d, mZ_0a, initialise);
  BrzM_1_2 I15 (c87_r0d, c87_r1d, c87_a, c89_r0d, c89_r1d, c89_a, c90_r0d, c90_r1d, c90_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I16 (c43_r0d, c43_r1d, c43_a, c88_r, c88_a, c89_r0d, c89_r1d, c89_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I17 (c18_r0d, c18_r1d, c18_a, c86_r, c86_a, c87_r0d, c87_r1d, c87_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I18 (c85_r0d, c85_r1d, c85_a, c14_r, c14_a, c41_r, c41_a, initialise);
  BrzJ_l11__280_202_29 I19 (c81_r, c81_a, c84_r0d, c84_r1d, c84_a, c85_r0d, c85_r1d, c85_a, initialise);
  BrzM_2_2 I20 (c82_r0d, c82_r1d, c82_a, c83_r0d, c83_r1d, c83_a, c84_r0d, c84_r1d, c84_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I21 (c78_r, c78_a, c83_r0d, c83_r1d, c83_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I22 (c76_r, c76_a, c82_r0d, c82_r1d, c82_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I23 (c80_r0d, c80_r1d, c80_a, c81_r, c81_a, mpL_0r0d, mpL_0r1d, mpL_0a, initialise);
  BrzM_32_2 I24 (c77_r0d, c77_r1d, c77_a, c79_r0d, c79_r1d, c79_a, c80_r0d, c80_r1d, c80_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I25 (c40_r0d, c40_r1d, c40_a, c78_r, c78_a, c79_r0d, c79_r1d, c79_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I26 (c13_r0d, c13_r1d, c13_a, c76_r, c76_a, c77_r0d, c77_r1d, c77_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I27 (c75_r0d, c75_r1d, c75_a, c32_r, c32_a, c53_r, c53_a, initialise);
  BrzJ_l11__280_202_29 I28 (c71_r, c71_a, c74_r0d, c74_r1d, c74_a, c75_r0d, c75_r1d, c75_a, initialise);
  BrzM_2_2 I29 (c72_r0d, c72_r1d, c72_a, c73_r0d, c73_r1d, c73_a, c74_r0d, c74_r1d, c74_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I30 (c68_r, c68_a, c73_r0d, c73_r1d, c73_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I31 (c66_r, c66_a, c72_r0d, c72_r1d, c72_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I32 (c70_r0d, c70_r1d, c70_a, c71_r, c71_a, mpH_0r0d, mpH_0r1d, mpH_0a, initialise);
  BrzM_32_2 I33 (c67_r0d, c67_r1d, c67_a, c69_r0d, c69_r1d, c69_a, c70_r0d, c70_r1d, c70_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I34 (c52_r0d, c52_r1d, c52_a, c68_r, c68_a, c69_r0d, c69_r1d, c69_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I35 (c31_r0d, c31_r1d, c31_a, c66_r, c66_a, c67_r0d, c67_r1d, c67_a, initialise);
  BrzJ_l11__281_200_29 I36 (bmN_0r0d, bmN_0r1d, bmN_0a, c27_r, c27_a, c25_r0d, c25_r1d, c25_a, initialise);
  BrzJ_l11__281_200_29 I37 (bmZ_0r0d, bmZ_0r1d, bmZ_0a, c22_r, c22_a, c20_r0d, c20_r1d, c20_a, initialise);
  BrzJ_l12__2832_200_29 I38 (bpL_0r0d, bpL_0r1d, bpL_0a, c17_r, c17_a, c15_r0d, c15_r1d, c15_a, initialise);
  BrzJ_l12__2832_200_29 I39 (bpH_0r0d, bpH_0r1d, bpH_0a, c35_r, c35_a, c33_r0d, c33_r1d, c33_a, initialise);
  BrzJ_l11__281_200_29 I40 (bL_0r0d, bL_0r1d, bL_0a, c64_r, c64_a, c60_r0d, c60_r1d, c60_a, initialise);
  BrzJ_l11__281_200_29 I41 (bH_0r0d, bH_0r1d, bH_0a, c63_r, c63_a, c58_r0d, c58_r1d, c58_a, initialise);
  BrzM_0_2 I42 (go_0r, go_0a, c57_r, c57_a, c65_r, c65_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I43 (c65_r, c65_a, c63_r, c63_a, c64_r, c64_a, initialise);
  BrzJ_l11__280_200_29 I44 (c59_r, c59_a, c61_r, c61_a, c62_r, c62_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I45 (c60_r0d, c60_r1d, c60_a, c61_r, c61_a, c62_r, c62_a, c12_r0d, c12_r1d, c12_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m72m I46 (c58_r0d, c58_r1d, c58_a, c59_r, c59_a, c29_r, c29_a, c49_r, c49_a, c28_r0d, c28_r1d, c28_a, c48_r0d, c48_r1d, c48_a, initialise);
  BrzM_0_2 I47 (c38_r, c38_a, c56_r, c56_a, c57_r, c57_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I48 (c12_r0d, c12_r1d, c12_a, c37_r, c37_a, c55_r, c55_a, initialise);
  BrzJ_l19__280_200_200_200_29 I49 (c41_r, c41_a, c44_r, c44_a, c47_r, c47_a, c54_r, c54_a, c56_r, c56_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I50 (c55_r, c55_a, c39_r, c39_a, c42_r, c42_a, c45_r, c45_a, c49_r, c49_a, initialise);
  BrzM_0_2 I51 (c50_r, c50_a, c53_r, c53_a, c54_r, c54_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I52 (c48_r0d, c48_r1d, c48_a, c50_r, c50_a, c51_r, c51_a, initialise);
  BrzO_0_32_l24__28_28num_2032_200_29_29 I53 (c51_r, c51_a, c52_r0d, c52_r1d, c52_a);
  BrzO_0_1_l23__28_28num_201_200_29_29 I54 (c45_r, c45_a, c46_r0d, c46_r1d, c46_a);
  BrzO_0_1_l23__28_28num_201_200_29_29 I55 (c42_r, c42_a, c43_r0d, c43_r1d, c43_a);
  BrzO_0_32_l24__28_28num_2032_200_29_29 I56 (c39_r, c39_a, c40_r0d, c40_r1d, c40_a);
  BrzJ_l19__280_200_200_200_29 I57 (c14_r, c14_a, c19_r, c19_a, c24_r, c24_a, c36_r, c36_a, c38_r, c38_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I58 (c37_r, c37_a, c17_r, c17_a, c22_r, c22_a, c27_r, c27_a, c29_r, c29_a, initialise);
  BrzM_0_2 I59 (c30_r, c30_a, c32_r, c32_a, c36_r, c36_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I60 (c28_r0d, c28_r1d, c28_a, c30_r, c30_a, c35_r, c35_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I61 (c33_r0d, c33_r1d, c33_a, c34_r, c34_a, c34_r, c34_a, c31_r0d, c31_r1d, c31_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I62 (c25_r0d, c25_r1d, c25_a, c26_r, c26_a, c26_r, c26_a, c23_r0d, c23_r1d, c23_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I63 (c20_r0d, c20_r1d, c20_a, c21_r, c21_a, c21_r, c21_a, c18_r0d, c18_r1d, c18_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I64 (c15_r0d, c15_r1d, c15_a, c16_r, c16_a, c16_r, c16_a, c13_r0d, c13_r1d, c13_a, initialise);
endmodule

module Balsa_bypassMul (
  go_0r, go_0a,
  bypass_0r0d, bypass_0r1d, bypass_0a,
  bypassH_0r0d, bypassH_0r1d, bypassH_0a,
  mulOpA_0r0d, mulOpA_0r1d, mulOpA_0a,
  mulOpB_0r0d, mulOpB_0r1d, mulOpB_0a,
  mulOpC_0r0d, mulOpC_0r1d, mulOpC_0a,
  mulType_0r0d, mulType_0r1d, mulType_0a,
  mulOpAo_0r0d, mulOpAo_0r1d, mulOpAo_0a,
  mulOpBo_0r0d, mulOpBo_0r1d, mulOpBo_0a,
  mulOpCo_0r0d, mulOpCo_0r1d, mulOpCo_0a,
  mulTypeo_0r0d, mulTypeo_0r1d, mulTypeo_0a,
  bH_0r0d, bH_0r1d, bH_0a,
  bL_0r0d, bL_0r1d, bL_0a,
  initialise
);
  input go_0r;
  output go_0a;
  input bypass_0r0d;
  input bypass_0r1d;
  output bypass_0a;
  input bypassH_0r0d;
  input bypassH_0r1d;
  output bypassH_0a;
  input [31:0] mulOpA_0r0d;
  input [31:0] mulOpA_0r1d;
  output mulOpA_0a;
  input [31:0] mulOpB_0r0d;
  input [31:0] mulOpB_0r1d;
  output mulOpB_0a;
  input [31:0] mulOpC_0r0d;
  input [31:0] mulOpC_0r1d;
  output mulOpC_0a;
  input [2:0] mulType_0r0d;
  input [2:0] mulType_0r1d;
  output mulType_0a;
  output [31:0] mulOpAo_0r0d;
  output [31:0] mulOpAo_0r1d;
  input mulOpAo_0a;
  output [31:0] mulOpBo_0r0d;
  output [31:0] mulOpBo_0r1d;
  input mulOpBo_0a;
  output [31:0] mulOpCo_0r0d;
  output [31:0] mulOpCo_0r1d;
  input mulOpCo_0a;
  output [2:0] mulTypeo_0r0d;
  output [2:0] mulTypeo_0r1d;
  input mulTypeo_0a;
  output bH_0r0d;
  output bH_0r1d;
  input bH_0a;
  output bL_0r0d;
  output bL_0r1d;
  input bL_0a;
  input initialise;
  wire [1:0] c84_r0d;
  wire [1:0] c84_r1d;
  wire c84_a;
  wire [1:0] c83_r0d;
  wire [1:0] c83_r1d;
  wire c83_a;
  wire [1:0] c82_r0d;
  wire [1:0] c82_r1d;
  wire c82_a;
  wire [1:0] c81_r0d;
  wire [1:0] c81_r1d;
  wire c81_a;
  wire c80_r;
  wire c80_a;
  wire [31:0] c79_r0d;
  wire [31:0] c79_r1d;
  wire c79_a;
  wire [31:0] c78_r0d;
  wire [31:0] c78_r1d;
  wire c78_a;
  wire c77_r;
  wire c77_a;
  wire [31:0] c76_r0d;
  wire [31:0] c76_r1d;
  wire c76_a;
  wire c75_r;
  wire c75_a;
  wire [33:0] c74_r0d;
  wire [33:0] c74_r1d;
  wire c74_a;
  wire [1:0] c73_r0d;
  wire [1:0] c73_r1d;
  wire c73_a;
  wire [1:0] c72_r0d;
  wire [1:0] c72_r1d;
  wire c72_a;
  wire [1:0] c71_r0d;
  wire [1:0] c71_r1d;
  wire c71_a;
  wire c70_r;
  wire c70_a;
  wire c69_r;
  wire c69_a;
  wire c68_r;
  wire c68_a;
  wire c67_r;
  wire c67_a;
  wire c66_r;
  wire c66_a;
  wire c65_r;
  wire c65_a;
  wire [2:0] c64_r0d;
  wire [2:0] c64_r1d;
  wire c64_a;
  wire c63_r;
  wire c63_a;
  wire c62_r0d;
  wire c62_r1d;
  wire c62_a;
  wire c61_r;
  wire c61_a;
  wire c60_r0d;
  wire c60_r1d;
  wire c60_a;
  wire c59_r;
  wire c59_a;
  wire c58_r;
  wire c58_a;
  wire c57_r;
  wire c57_a;
  wire c56_r0d;
  wire c56_r1d;
  wire c56_a;
  wire c55_r;
  wire c55_a;
  wire c54_r;
  wire c54_a;
  wire c53_r0d;
  wire c53_r1d;
  wire c53_a;
  wire c52_r;
  wire c52_a;
  wire c51_r;
  wire c51_a;
  wire c50_r;
  wire c50_a;
  wire c49_r;
  wire c49_a;
  wire c48_r;
  wire c48_a;
  wire [31:0] c47_r0d;
  wire [31:0] c47_r1d;
  wire c47_a;
  wire c46_r;
  wire c46_a;
  wire [31:0] c45_r0d;
  wire [31:0] c45_r1d;
  wire c45_a;
  wire c44_r;
  wire c44_a;
  wire c43_r;
  wire c43_a;
  wire c42_r;
  wire c42_a;
  wire c41_r;
  wire c41_a;
  wire [31:0] c40_r0d;
  wire [31:0] c40_r1d;
  wire c40_a;
  wire c39_r;
  wire c39_a;
  wire c38_r;
  wire c38_a;
  wire [2:0] c37_r0d;
  wire [2:0] c37_r1d;
  wire c37_a;
  wire c36_r;
  wire c36_a;
  wire c35_r;
  wire c35_a;
  wire c34_r;
  wire c34_a;
  wire c33_r;
  wire c33_a;
  wire c32_r;
  wire c32_a;
  wire [31:0] c31_r0d;
  wire [31:0] c31_r1d;
  wire c31_a;
  wire c30_r;
  wire c30_a;
  wire [31:0] c29_r0d;
  wire [31:0] c29_r1d;
  wire c29_a;
  wire c28_r;
  wire c28_a;
  wire [31:0] c27_r0d;
  wire [31:0] c27_r1d;
  wire c27_a;
  wire c26_r;
  wire c26_a;
  wire c25_r;
  wire c25_a;
  wire [2:0] c24_r0d;
  wire [2:0] c24_r1d;
  wire c24_a;
  wire c23_r;
  wire c23_a;
  wire c22_r;
  wire c22_a;
  wire [2:0] c21_r0d;
  wire [2:0] c21_r1d;
  wire c21_a;
  wire c20_r;
  wire c20_a;
  wire c19_r;
  wire c19_a;
  wire [31:0] c18_r0d;
  wire [31:0] c18_r1d;
  wire c18_a;
  wire c17_r;
  wire c17_a;
  wire c16_r;
  wire c16_a;
  wire [31:0] c15_r0d;
  wire [31:0] c15_r1d;
  wire c15_a;
  wire c14_r0d;
  wire c14_r1d;
  wire c14_a;
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I0 (c53_r0d, c53_r1d, c53_a, c55_r, c55_a, bL_0r0d, bL_0r1d, bL_0a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I1 (c56_r0d, c56_r1d, c56_a, c58_r, c58_a, bH_0r0d, bH_0r1d, bH_0a, initialise);
  BrzF_3_l31__28_280_200_29_20_280_203_29_29 I2 (c21_r0d, c21_r1d, c21_a, c23_r, c23_a, mulTypeo_0r0d, mulTypeo_0r1d, mulTypeo_0a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I3 (c84_r0d, c84_r1d, c84_a, c28_r, c28_a, c30_r, c30_a, initialise);
  BrzJ_l11__280_202_29 I4 (c80_r, c80_a, c83_r0d, c83_r1d, c83_a, c84_r0d, c84_r1d, c84_a, initialise);
  BrzM_2_2 I5 (c81_r0d, c81_r1d, c81_a, c82_r0d, c82_r1d, c82_a, c83_r0d, c83_r1d, c83_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I6 (c77_r, c77_a, c82_r0d, c82_r1d, c82_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I7 (c75_r, c75_a, c81_r0d, c81_r1d, c81_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I8 (c79_r0d, c79_r1d, c79_a, c80_r, c80_a, mulOpCo_0r0d, mulOpCo_0r1d, mulOpCo_0a, initialise);
  BrzM_32_2 I9 (c76_r0d, c76_r1d, c76_a, c78_r0d, c78_r1d, c78_a, c79_r0d, c79_r1d, c79_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I10 (c29_r0d, c29_r1d, c29_a, c77_r, c77_a, c78_r0d, c78_r1d, c78_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I11 (c27_r0d, c27_r1d, c27_a, c75_r, c75_a, c76_r0d, c76_r1d, c76_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I12 (c18_r0d, c18_r1d, c18_a, c20_r, c20_a, mulOpBo_0r0d, mulOpBo_0r1d, mulOpBo_0a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I13 (c15_r0d, c15_r1d, c15_a, c17_r, c17_a, mulOpAo_0r0d, mulOpAo_0r1d, mulOpAo_0a, initialise);
  BrzJ_l11__283_200_29 I14 (mulType_0r0d, mulType_0r1d, mulType_0a, c69_r, c69_a, c64_r0d, c64_r1d, c64_a, initialise);
  BrzS_34_l12__2832_202_29_l97__28_28_28_281_m69m I15 (c74_r0d, c74_r1d, c74_a, c31_r0d, c31_r1d, c31_a, c40_r0d, c40_r1d, c40_a, initialise);
  BrzJ_l12__2832_202_29 I16 (mulOpC_0r0d, mulOpC_0r1d, mulOpC_0a, c73_r0d, c73_r1d, c73_a, c74_r0d, c74_r1d, c74_a, initialise);
  BrzM_2_2 I17 (c71_r0d, c71_r1d, c71_a, c72_r0d, c72_r1d, c72_a, c73_r0d, c73_r1d, c73_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I18 (c42_r, c42_a, c72_r0d, c72_r1d, c72_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I19 (c33_r, c33_a, c71_r0d, c71_r1d, c71_a);
  BrzJ_l12__2832_200_29 I20 (mulOpB_0r0d, mulOpB_0r1d, mulOpB_0a, c51_r, c51_a, c47_r0d, c47_r1d, c47_a, initialise);
  BrzJ_l12__2832_200_29 I21 (mulOpA_0r0d, mulOpA_0r1d, mulOpA_0a, c50_r, c50_a, c45_r0d, c45_r1d, c45_a, initialise);
  BrzJ_l11__281_200_29 I22 (bypassH_0r0d, bypassH_0r1d, bypassH_0a, c68_r, c68_a, c62_r0d, c62_r1d, c62_a, initialise);
  BrzJ_l11__281_200_29 I23 (bypass_0r0d, bypass_0r1d, bypass_0a, c67_r, c67_a, c60_r0d, c60_r1d, c60_a, initialise);
  BrzM_0_2 I24 (go_0r, go_0a, c59_r, c59_a, c70_r, c70_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I25 (c70_r, c70_a, c67_r, c67_a, c68_r, c68_a, c69_r, c69_a, initialise);
  BrzJ_l15__280_200_200_29 I26 (c61_r, c61_a, c63_r, c63_a, c65_r, c65_a, c66_r, c66_a, initialise);
  BrzV_3_l6__28_29_l23__28_28_280_203_29_29__m75m I27 (c64_r0d, c64_r1d, c64_a, c65_r, c65_a, c22_r, c22_a, c25_r, c25_a, c38_r, c38_a, c21_r0d, c21_r1d, c21_a, c24_r0d, c24_r1d, c24_a, c37_r0d, c37_r1d, c37_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I28 (c62_r0d, c62_r1d, c62_a, c63_r, c63_a, c57_r, c57_a, c56_r0d, c56_r1d, c56_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m72m I29 (c60_r0d, c60_r1d, c60_a, c61_r, c61_a, c49_r, c49_a, c54_r, c54_a, c14_r0d, c14_r1d, c14_a, c53_r0d, c53_r1d, c53_a, initialise);
  BrzJ_l15__280_200_200_29 I30 (c44_r, c44_a, c55_r, c55_a, c58_r, c58_a, c59_r, c59_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I31 (c66_r, c66_a, c52_r, c52_a, c54_r, c54_a, c57_r, c57_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I32 (c52_r, c52_a, c50_r, c50_a, c51_r, c51_a, initialise);
  BrzJ_l11__280_200_29 I33 (c46_r, c46_a, c48_r, c48_a, c49_r, c49_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I34 (c47_r0d, c47_r1d, c47_a, c48_r, c48_a, c19_r, c19_a, c18_r0d, c18_r1d, c18_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I35 (c45_r0d, c45_r1d, c45_a, c46_r, c46_a, c16_r, c16_a, c15_r0d, c15_r1d, c15_a, initialise);
  BrzM_0_2 I36 (c36_r, c36_a, c43_r, c43_a, c44_r, c44_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I37 (c14_r0d, c14_r1d, c14_a, c35_r, c35_a, c38_r, c38_a, initialise);
  BrzM_0_2 I38 (c39_r, c39_a, c41_r, c41_a, c43_r, c43_a, initialise);
  BrzS_3_l11__280_203_29_l137__28_28_28_280__m63m I39 (c37_r0d, c37_r1d, c37_a, c39_r, c39_a, c42_r, c42_a, initialise);
  BrzF_32_l17__28_280_200_29_29 I40 (c40_r0d, c40_r1d, c40_a, c41_r, c41_a, initialise);
  BrzJ_l19__280_200_200_200_29 I41 (c17_r, c17_a, c20_r, c20_a, c23_r, c23_a, c34_r, c34_a, c36_r, c36_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I42 (c35_r, c35_a, c16_r, c16_a, c19_r, c19_a, c22_r, c22_a, c25_r, c25_a, initialise);
  BrzM_0_2 I43 (c28_r, c28_a, c30_r, c30_a, c34_r, c34_a, initialise);
  BrzS_3_l11__280_203_29_l137__28_28_28_280__m63m I44 (c24_r0d, c24_r1d, c24_a, c26_r, c26_a, c33_r, c33_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I45 (c31_r0d, c31_r1d, c31_a, c32_r, c32_a, c32_r, c32_a, c29_r0d, c29_r1d, c29_a, initialise);
  BrzO_0_32_l24__28_28num_2032_200_29_29 I46 (c26_r, c26_a, c27_r0d, c27_r1d, c27_a);
endmodule

module Balsa_mControl10 (
  go_0r, go_0a,
  load_0r0d, load_0r1d, load_0a,
  done_0r0d, done_0r1d, done_0a,
  initialise
);
  input go_0r;
  output go_0a;
  input load_0r0d;
  input load_0r1d;
  output load_0a;
  output done_0r0d;
  output done_0r1d;
  input done_0a;
  input initialise;
  wire [1:0] c39_r0d;
  wire [1:0] c39_r1d;
  wire c39_a;
  wire [1:0] c38_r0d;
  wire [1:0] c38_r1d;
  wire c38_a;
  wire [1:0] c37_r0d;
  wire [1:0] c37_r1d;
  wire c37_a;
  wire [1:0] c36_r0d;
  wire [1:0] c36_r1d;
  wire c36_a;
  wire c35_r;
  wire c35_a;
  wire c34_r0d;
  wire c34_r1d;
  wire c34_a;
  wire c33_r0d;
  wire c33_r1d;
  wire c33_a;
  wire c32_r;
  wire c32_a;
  wire c31_r0d;
  wire c31_r1d;
  wire c31_a;
  wire c30_r;
  wire c30_a;
  wire c29_r;
  wire c29_a;
  wire c28_r;
  wire c28_a;
  wire c27_r;
  wire c27_a;
  wire c26_r;
  wire c26_a;
  wire c25_r0d;
  wire c25_r1d;
  wire c25_a;
  wire c24_r;
  wire c24_a;
  wire c23_r;
  wire c23_a;
  wire [9:0] c22_r0d;
  wire [9:0] c22_r1d;
  wire c22_a;
  wire c21_r;
  wire c21_a;
  wire c20_r;
  wire c20_a;
  wire [9:0] c19_r0d;
  wire [9:0] c19_r1d;
  wire c19_a;
  wire c18_r;
  wire c18_a;
  wire c17_r;
  wire c17_a;
  wire c16_r;
  wire c16_a;
  wire [8:0] c15_r0d;
  wire [8:0] c15_r1d;
  wire c15_a;
  wire [9:0] c14_r0d;
  wire [9:0] c14_r1d;
  wire c14_a;
  wire c13_r;
  wire c13_a;
  wire c12_r;
  wire c12_a;
  wire c11_r0d;
  wire c11_r1d;
  wire c11_a;
  wire c10_r;
  wire c10_a;
  wire c9_r0d;
  wire c9_r1d;
  wire c9_a;
  wire c8_r;
  wire c8_a;
  wire c7_r0d;
  wire c7_r1d;
  wire c7_a;
  wire c6_r;
  wire c6_a;
  wire c5_r0d;
  wire c5_r1d;
  wire c5_a;
  wire c4_r;
  wire c4_a;
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I0 (c39_r0d, c39_r1d, c39_a, c13_r, c13_a, c26_r, c26_a, initialise);
  BrzJ_l11__280_202_29 I1 (c35_r, c35_a, c38_r0d, c38_r1d, c38_a, c39_r0d, c39_r1d, c39_a, initialise);
  BrzM_2_2 I2 (c36_r0d, c36_r1d, c36_a, c37_r0d, c37_r1d, c37_a, c38_r0d, c38_r1d, c38_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I3 (c32_r, c32_a, c37_r0d, c37_r1d, c37_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I4 (c30_r, c30_a, c36_r0d, c36_r1d, c36_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I5 (c34_r0d, c34_r1d, c34_a, c35_r, c35_a, done_0r0d, done_0r1d, done_0a, initialise);
  BrzM_1_2 I6 (c31_r0d, c31_r1d, c31_a, c33_r0d, c33_r1d, c33_a, c34_r0d, c34_r1d, c34_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I7 (c25_r0d, c25_r1d, c25_a, c32_r, c32_a, c33_r0d, c33_r1d, c33_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I8 (c11_r0d, c11_r1d, c11_a, c30_r, c30_a, c31_r0d, c31_r1d, c31_a, initialise);
  BrzJ_l11__281_200_29 I9 (load_0r0d, load_0r1d, load_0a, c4_r, c4_a, c7_r0d, c7_r1d, c7_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I10 (c5_r0d, c5_r1d, c5_a, c6_r, c6_a, c6_r, c6_a, c9_r0d, c9_r1d, c9_a, initialise);
  BrzV_10_l6__28_29_l45__28_28_280_2010_29_2_m79m I11 (c22_r0d, c22_r1d, c22_a, c19_r0d, c19_r1d, c19_a, c23_r, c23_a, c20_r, c20_a, c16_r, c16_a, c12_r, c12_a, c15_r0d, c15_r1d, c15_a, c11_r0d, c11_r1d, c11_a, initialise);
  BrzV_10_l6__28_29_l24__28_28_280_2010_29_2_m78m I12 (c14_r0d, c14_r1d, c14_a, c17_r, c17_a, c18_r, c18_a, c19_r0d, c19_r1d, c19_a, initialise);
  BrzM_0_2 I13 (go_0r, go_0a, c29_r, c29_a, c4_r, c4_a, initialise);
  BrzM_0_2 I14 (c20_r, c20_a, c28_r, c28_a, c29_r, c29_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I15 (c9_r0d, c9_r1d, c9_a, c10_r, c10_a, c27_r, c27_a, initialise);
  BrzJ_l11__280_200_29 I16 (c23_r, c23_a, c26_r, c26_a, c28_r, c28_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I17 (c27_r, c27_a, c21_r, c21_a, c24_r, c24_a, initialise);
  BrzO_0_1_l23__28_28num_201_201_29_29 I18 (c24_r, c24_a, c25_r0d, c25_r1d, c25_a);
  BrzO_0_10_l26__28_28num_2010_20256_29_29 I19 (c21_r, c21_a, c22_r0d, c22_r1d, c22_a);
  BrzJ_l11__280_200_29 I20 (c13_r, c13_a, c17_r, c17_a, c18_r, c18_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I21 (c10_r, c10_a, c12_r, c12_a, c16_r, c16_a, initialise);
  BrzO_9_10_l75__28_28num_201_200_29_20_28ap_m49m I22 (c15_r0d, c15_r1d, c15_a, c14_r0d, c14_r1d, c14_a);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I23 (c7_r0d, c7_r1d, c7_a, c8_r, c8_a, c8_r, c8_a, c5_r0d, c5_r1d, c5_a, initialise);
endmodule

module Balsa_nanoMBoothR3rolled (
  go_0r, go_0a,
  cin_0r0d, cin_0r1d, cin_0a,
  res_0r0d, res_0r1d, res_0a,
  a_0r0d, a_0r1d, a_0a,
  b_0r0d, b_0r1d, b_0a,
  c_0r0d, c_0r1d, c_0a,
  mlength_0r0d, mlength_0r1d, mlength_0a,
  macc_0r0d, macc_0r1d, macc_0a,
  load_0r0d, load_0r1d, load_0a,
  done_0r0d, done_0r1d, done_0a,
  opA_0r0d, opA_0r1d, opA_0a,
  opB_0r0d, opB_0r1d, opB_0a,
  cs_0r0d, cs_0r1d, cs_0a,
  raA_0r0d, raA_0r1d, raA_0a,
  raB_0r0d, raB_0r1d, raB_0a,
  rac0_0r0d, rac0_0r1d, rac0_0a,
  raS_0r0d, raS_0r1d, raS_0a,
  racN_0r0d, racN_0r1d, racN_0a,
  pH_0r0d, pH_0r1d, pH_0a,
  pL_0r0d, pL_0r1d, pL_0a,
  z_0r0d, z_0r1d, z_0a,
  n_0r0d, n_0r1d, n_0a,
  initialise
);
  input go_0r;
  output go_0a;
  input [34:0] cin_0r0d;
  input [34:0] cin_0r1d;
  output cin_0a;
  input [34:0] res_0r0d;
  input [34:0] res_0r1d;
  output res_0a;
  input [34:0] a_0r0d;
  input [34:0] a_0r1d;
  output a_0a;
  input [35:0] b_0r0d;
  input [35:0] b_0r1d;
  output b_0a;
  input [34:0] c_0r0d;
  input [34:0] c_0r1d;
  output c_0a;
  input mlength_0r0d;
  input mlength_0r1d;
  output mlength_0a;
  input macc_0r0d;
  input macc_0r1d;
  output macc_0a;
  output load_0r0d;
  output load_0r1d;
  input load_0a;
  input done_0r0d;
  input done_0r1d;
  output done_0a;
  output [34:0] opA_0r0d;
  output [34:0] opA_0r1d;
  input opA_0a;
  output [34:0] opB_0r0d;
  output [34:0] opB_0r1d;
  input opB_0a;
  output [34:0] cs_0r0d;
  output [34:0] cs_0r1d;
  input cs_0a;
  output [31:0] raA_0r0d;
  output [31:0] raA_0r1d;
  input raA_0a;
  output [31:0] raB_0r0d;
  output [31:0] raB_0r1d;
  input raB_0a;
  output rac0_0r0d;
  output rac0_0r1d;
  input rac0_0a;
  input [31:0] raS_0r0d;
  input [31:0] raS_0r1d;
  output raS_0a;
  input racN_0r0d;
  input racN_0r1d;
  output racN_0a;
  output [31:0] pH_0r0d;
  output [31:0] pH_0r1d;
  input pH_0a;
  output [31:0] pL_0r0d;
  output [31:0] pL_0r1d;
  input pL_0a;
  output z_0r0d;
  output z_0r1d;
  input z_0a;
  output n_0r0d;
  output n_0r1d;
  input n_0a;
  input initialise;
  wire [1:0] c479_r0d;
  wire [1:0] c479_r1d;
  wire c479_a;
  wire [1:0] c478_r0d;
  wire [1:0] c478_r1d;
  wire c478_a;
  wire [1:0] c477_r0d;
  wire [1:0] c477_r1d;
  wire c477_a;
  wire [1:0] c476_r0d;
  wire [1:0] c476_r1d;
  wire c476_a;
  wire c475_r;
  wire c475_a;
  wire c474_r0d;
  wire c474_r1d;
  wire c474_a;
  wire c473_r0d;
  wire c473_r1d;
  wire c473_a;
  wire c472_r;
  wire c472_a;
  wire c471_r0d;
  wire c471_r1d;
  wire c471_a;
  wire c470_r;
  wire c470_a;
  wire [2:0] c469_r0d;
  wire [2:0] c469_r1d;
  wire c469_a;
  wire [2:0] c468_r0d;
  wire [2:0] c468_r1d;
  wire c468_a;
  wire [2:0] c467_r0d;
  wire [2:0] c467_r1d;
  wire c467_a;
  wire [2:0] c466_r0d;
  wire [2:0] c466_r1d;
  wire c466_a;
  wire [2:0] c465_r0d;
  wire [2:0] c465_r1d;
  wire c465_a;
  wire c464_r;
  wire c464_a;
  wire c463_r0d;
  wire c463_r1d;
  wire c463_a;
  wire c462_r0d;
  wire c462_r1d;
  wire c462_a;
  wire c461_r;
  wire c461_a;
  wire c460_r0d;
  wire c460_r1d;
  wire c460_a;
  wire c459_r;
  wire c459_a;
  wire c458_r0d;
  wire c458_r1d;
  wire c458_a;
  wire c457_r;
  wire c457_a;
  wire [1:0] c456_r0d;
  wire [1:0] c456_r1d;
  wire c456_a;
  wire [1:0] c455_r0d;
  wire [1:0] c455_r1d;
  wire c455_a;
  wire [1:0] c454_r0d;
  wire [1:0] c454_r1d;
  wire c454_a;
  wire [1:0] c453_r0d;
  wire [1:0] c453_r1d;
  wire c453_a;
  wire c452_r;
  wire c452_a;
  wire [31:0] c451_r0d;
  wire [31:0] c451_r1d;
  wire c451_a;
  wire [31:0] c450_r0d;
  wire [31:0] c450_r1d;
  wire c450_a;
  wire c449_r;
  wire c449_a;
  wire [31:0] c448_r0d;
  wire [31:0] c448_r1d;
  wire c448_a;
  wire c447_r;
  wire c447_a;
  wire [3:0] c446_r0d;
  wire [3:0] c446_r1d;
  wire c446_a;
  wire [2:0] c445_r0d;
  wire [2:0] c445_r1d;
  wire c445_a;
  wire [2:0] c444_r0d;
  wire [2:0] c444_r1d;
  wire c444_a;
  wire [2:0] c443_r0d;
  wire [2:0] c443_r1d;
  wire c443_a;
  wire [2:0] c442_r0d;
  wire [2:0] c442_r1d;
  wire c442_a;
  wire [34:0] c441_r0d;
  wire [34:0] c441_r1d;
  wire c441_a;
  wire [2:0] c440_r0d;
  wire [2:0] c440_r1d;
  wire c440_a;
  wire [2:0] c439_r0d;
  wire [2:0] c439_r1d;
  wire c439_a;
  wire [2:0] c438_r0d;
  wire [2:0] c438_r1d;
  wire c438_a;
  wire [2:0] c437_r0d;
  wire [2:0] c437_r1d;
  wire c437_a;
  wire [2:0] c436_r0d;
  wire [2:0] c436_r1d;
  wire c436_a;
  wire [2:0] c435_r0d;
  wire [2:0] c435_r1d;
  wire c435_a;
  wire [2:0] c434_r0d;
  wire [2:0] c434_r1d;
  wire c434_a;
  wire [2:0] c433_r0d;
  wire [2:0] c433_r1d;
  wire c433_a;
  wire [2:0] c432_r0d;
  wire [2:0] c432_r1d;
  wire c432_a;
  wire c431_r;
  wire c431_a;
  wire c430_r0d;
  wire c430_r1d;
  wire c430_a;
  wire c429_r0d;
  wire c429_r1d;
  wire c429_a;
  wire c428_r;
  wire c428_a;
  wire c427_r0d;
  wire c427_r1d;
  wire c427_a;
  wire c426_r;
  wire c426_a;
  wire c425_r0d;
  wire c425_r1d;
  wire c425_a;
  wire c424_r;
  wire c424_a;
  wire [2:0] c423_r0d;
  wire [2:0] c423_r1d;
  wire c423_a;
  wire [2:0] c422_r0d;
  wire [2:0] c422_r1d;
  wire c422_a;
  wire [2:0] c421_r0d;
  wire [2:0] c421_r1d;
  wire c421_a;
  wire [2:0] c420_r0d;
  wire [2:0] c420_r1d;
  wire c420_a;
  wire [2:0] c419_r0d;
  wire [2:0] c419_r1d;
  wire c419_a;
  wire c418_r;
  wire c418_a;
  wire [31:0] c417_r0d;
  wire [31:0] c417_r1d;
  wire c417_a;
  wire [31:0] c416_r0d;
  wire [31:0] c416_r1d;
  wire c416_a;
  wire c415_r;
  wire c415_a;
  wire [31:0] c414_r0d;
  wire [31:0] c414_r1d;
  wire c414_a;
  wire c413_r;
  wire c413_a;
  wire [31:0] c412_r0d;
  wire [31:0] c412_r1d;
  wire c412_a;
  wire c411_r;
  wire c411_a;
  wire [2:0] c410_r0d;
  wire [2:0] c410_r1d;
  wire c410_a;
  wire [2:0] c409_r0d;
  wire [2:0] c409_r1d;
  wire c409_a;
  wire [2:0] c408_r0d;
  wire [2:0] c408_r1d;
  wire c408_a;
  wire [2:0] c407_r0d;
  wire [2:0] c407_r1d;
  wire c407_a;
  wire [2:0] c406_r0d;
  wire [2:0] c406_r1d;
  wire c406_a;
  wire c405_r;
  wire c405_a;
  wire [31:0] c404_r0d;
  wire [31:0] c404_r1d;
  wire c404_a;
  wire [31:0] c403_r0d;
  wire [31:0] c403_r1d;
  wire c403_a;
  wire c402_r;
  wire c402_a;
  wire [31:0] c401_r0d;
  wire [31:0] c401_r1d;
  wire c401_a;
  wire c400_r;
  wire c400_a;
  wire [31:0] c399_r0d;
  wire [31:0] c399_r1d;
  wire c399_a;
  wire c398_r;
  wire c398_a;
  wire [8:0] c397_r0d;
  wire [8:0] c397_r1d;
  wire c397_a;
  wire [8:0] c396_r0d;
  wire [8:0] c396_r1d;
  wire c396_a;
  wire [8:0] c395_r0d;
  wire [8:0] c395_r1d;
  wire c395_a;
  wire [8:0] c394_r0d;
  wire [8:0] c394_r1d;
  wire c394_a;
  wire [8:0] c393_r0d;
  wire [8:0] c393_r1d;
  wire c393_a;
  wire [8:0] c392_r0d;
  wire [8:0] c392_r1d;
  wire c392_a;
  wire [8:0] c391_r0d;
  wire [8:0] c391_r1d;
  wire c391_a;
  wire [8:0] c390_r0d;
  wire [8:0] c390_r1d;
  wire c390_a;
  wire [8:0] c389_r0d;
  wire [8:0] c389_r1d;
  wire c389_a;
  wire [8:0] c388_r0d;
  wire [8:0] c388_r1d;
  wire c388_a;
  wire [8:0] c387_r0d;
  wire [8:0] c387_r1d;
  wire c387_a;
  wire c386_r;
  wire c386_a;
  wire [34:0] c385_r0d;
  wire [34:0] c385_r1d;
  wire c385_a;
  wire [34:0] c384_r0d;
  wire [34:0] c384_r1d;
  wire c384_a;
  wire c383_r;
  wire c383_a;
  wire [34:0] c382_r0d;
  wire [34:0] c382_r1d;
  wire c382_a;
  wire c381_r;
  wire c381_a;
  wire [34:0] c380_r0d;
  wire [34:0] c380_r1d;
  wire c380_a;
  wire c379_r;
  wire c379_a;
  wire [34:0] c378_r0d;
  wire [34:0] c378_r1d;
  wire c378_a;
  wire c377_r;
  wire c377_a;
  wire [34:0] c376_r0d;
  wire [34:0] c376_r1d;
  wire c376_a;
  wire c375_r;
  wire c375_a;
  wire [34:0] c374_r0d;
  wire [34:0] c374_r1d;
  wire c374_a;
  wire c373_r;
  wire c373_a;
  wire [34:0] c372_r0d;
  wire [34:0] c372_r1d;
  wire c372_a;
  wire c371_r;
  wire c371_a;
  wire [34:0] c370_r0d;
  wire [34:0] c370_r1d;
  wire c370_a;
  wire c369_r;
  wire c369_a;
  wire [34:0] c368_r0d;
  wire [34:0] c368_r1d;
  wire c368_a;
  wire c367_r;
  wire c367_a;
  wire [1:0] c366_r0d;
  wire [1:0] c366_r1d;
  wire c366_a;
  wire [1:0] c365_r0d;
  wire [1:0] c365_r1d;
  wire c365_a;
  wire [1:0] c364_r0d;
  wire [1:0] c364_r1d;
  wire c364_a;
  wire [1:0] c363_r0d;
  wire [1:0] c363_r1d;
  wire c363_a;
  wire c362_r;
  wire c362_a;
  wire c361_r0d;
  wire c361_r1d;
  wire c361_a;
  wire c360_r0d;
  wire c360_r1d;
  wire c360_a;
  wire c359_r;
  wire c359_a;
  wire c358_r0d;
  wire c358_r1d;
  wire c358_a;
  wire c357_r;
  wire c357_a;
  wire [34:0] c356_r0d;
  wire [34:0] c356_r1d;
  wire c356_a;
  wire [34:0] c355_r0d;
  wire [34:0] c355_r1d;
  wire c355_a;
  wire c354_r0d;
  wire c354_r1d;
  wire c354_a;
  wire c353_r;
  wire c353_a;
  wire c352_r;
  wire c352_a;
  wire c351_r;
  wire c351_a;
  wire c350_r;
  wire c350_a;
  wire c349_r0d;
  wire c349_r1d;
  wire c349_a;
  wire c348_r;
  wire c348_a;
  wire c347_r;
  wire c347_a;
  wire c346_r;
  wire c346_a;
  wire c345_r0d;
  wire c345_r1d;
  wire c345_a;
  wire c344_r;
  wire c344_a;
  wire c343_r;
  wire c343_a;
  wire c342_r0d;
  wire c342_r1d;
  wire c342_a;
  wire [1:0] c341_r0d;
  wire [1:0] c341_r1d;
  wire c341_a;
  wire c340_r;
  wire c340_a;
  wire c339_r0d;
  wire c339_r1d;
  wire c339_a;
  wire c338_r0d;
  wire c338_r1d;
  wire c338_a;
  wire [32:0] c337_r0d;
  wire [32:0] c337_r1d;
  wire c337_a;
  wire c336_r0d;
  wire c336_r1d;
  wire c336_a;
  wire c335_r;
  wire c335_a;
  wire c334_r;
  wire c334_a;
  wire [31:0] c333_r0d;
  wire [31:0] c333_r1d;
  wire c333_a;
  wire c332_r;
  wire c332_a;
  wire c331_r0d;
  wire c331_r1d;
  wire c331_a;
  wire c330_r;
  wire c330_a;
  wire c329_r;
  wire c329_a;
  wire [31:0] c328_r0d;
  wire [31:0] c328_r1d;
  wire c328_a;
  wire c327_r;
  wire c327_a;
  wire c326_r;
  wire c326_a;
  wire [31:0] c325_r0d;
  wire [31:0] c325_r1d;
  wire c325_a;
  wire c324_r;
  wire c324_a;
  wire c323_r;
  wire c323_a;
  wire c322_r;
  wire c322_a;
  wire c321_r;
  wire c321_a;
  wire c320_r;
  wire c320_a;
  wire c319_r;
  wire c319_a;
  wire c318_r0d;
  wire c318_r1d;
  wire c318_a;
  wire c317_r;
  wire c317_a;
  wire [31:0] c316_r0d;
  wire [31:0] c316_r1d;
  wire c316_a;
  wire c315_r;
  wire c315_a;
  wire [31:0] c314_r0d;
  wire [31:0] c314_r1d;
  wire c314_a;
  wire c313_r;
  wire c313_a;
  wire c312_r;
  wire c312_a;
  wire c311_r0d;
  wire c311_r1d;
  wire c311_a;
  wire c310_r;
  wire c310_a;
  wire c309_r;
  wire c309_a;
  wire [31:0] c308_r0d;
  wire [31:0] c308_r1d;
  wire c308_a;
  wire c307_r;
  wire c307_a;
  wire c306_r;
  wire c306_a;
  wire [31:0] c305_r0d;
  wire [31:0] c305_r1d;
  wire c305_a;
  wire c304_r;
  wire c304_a;
  wire [30:0] c303_r0d;
  wire [30:0] c303_r1d;
  wire c303_a;
  wire c302_r;
  wire c302_a;
  wire c301_r0d;
  wire c301_r1d;
  wire c301_a;
  wire c300_r;
  wire c300_a;
  wire c299_r;
  wire c299_a;
  wire c298_r;
  wire c298_a;
  wire c297_r;
  wire c297_a;
  wire c296_r;
  wire c296_a;
  wire c295_r0d;
  wire c295_r1d;
  wire c295_a;
  wire c294_r;
  wire c294_a;
  wire c293_r;
  wire c293_a;
  wire c292_r0d;
  wire c292_r1d;
  wire c292_a;
  wire c291_r;
  wire c291_a;
  wire c290_r;
  wire c290_a;
  wire [31:0] c289_r0d;
  wire [31:0] c289_r1d;
  wire c289_a;
  wire c288_r0d;
  wire c288_r1d;
  wire c288_a;
  wire c287_r;
  wire c287_a;
  wire c286_r;
  wire c286_a;
  wire c285_r;
  wire c285_a;
  wire c284_r;
  wire c284_a;
  wire c283_r;
  wire c283_a;
  wire c282_r;
  wire c282_a;
  wire c281_r0d;
  wire c281_r1d;
  wire c281_a;
  wire c280_r;
  wire c280_a;
  wire [31:0] c279_r0d;
  wire [31:0] c279_r1d;
  wire c279_a;
  wire c278_r;
  wire c278_a;
  wire c277_r;
  wire c277_a;
  wire c276_r;
  wire c276_a;
  wire c275_r0d;
  wire c275_r1d;
  wire c275_a;
  wire [32:0] c274_r0d;
  wire [32:0] c274_r1d;
  wire c274_a;
  wire c273_r0d;
  wire c273_r1d;
  wire c273_a;
  wire c272_r;
  wire c272_a;
  wire c271_r;
  wire c271_a;
  wire [31:0] c270_r0d;
  wire [31:0] c270_r1d;
  wire c270_a;
  wire c269_r;
  wire c269_a;
  wire c268_r;
  wire c268_a;
  wire c267_r0d;
  wire c267_r1d;
  wire c267_a;
  wire c266_r;
  wire c266_a;
  wire c265_r;
  wire c265_a;
  wire c264_r0d;
  wire c264_r1d;
  wire c264_a;
  wire c263_r;
  wire c263_a;
  wire c262_r;
  wire c262_a;
  wire [31:0] c261_r0d;
  wire [31:0] c261_r1d;
  wire c261_a;
  wire c260_r;
  wire c260_a;
  wire c259_r0d;
  wire c259_r1d;
  wire c259_a;
  wire c258_r;
  wire c258_a;
  wire c257_r;
  wire c257_a;
  wire c256_r;
  wire c256_a;
  wire [31:0] c255_r0d;
  wire [31:0] c255_r1d;
  wire c255_a;
  wire c254_r;
  wire c254_a;
  wire c253_r;
  wire c253_a;
  wire [31:0] c252_r0d;
  wire [31:0] c252_r1d;
  wire c252_a;
  wire c251_r;
  wire c251_a;
  wire c250_r;
  wire c250_a;
  wire c249_r;
  wire c249_a;
  wire c248_r;
  wire c248_a;
  wire c247_r0d;
  wire c247_r1d;
  wire c247_a;
  wire c246_r;
  wire c246_a;
  wire c245_r;
  wire c245_a;
  wire c244_r;
  wire c244_a;
  wire [3:0] c243_r0d;
  wire [3:0] c243_r1d;
  wire c243_a;
  wire c242_r;
  wire c242_a;
  wire c241_r;
  wire c241_a;
  wire [35:0] c240_r0d;
  wire [35:0] c240_r1d;
  wire c240_a;
  wire c239_r;
  wire c239_a;
  wire c238_r;
  wire c238_a;
  wire [34:0] c237_r0d;
  wire [34:0] c237_r1d;
  wire c237_a;
  wire c236_r;
  wire c236_a;
  wire c235_r;
  wire c235_a;
  wire [35:0] c234_r0d;
  wire [35:0] c234_r1d;
  wire c234_a;
  wire c233_r;
  wire c233_a;
  wire c232_r;
  wire c232_a;
  wire [34:0] c231_r0d;
  wire [34:0] c231_r1d;
  wire c231_a;
  wire c230_r;
  wire c230_a;
  wire c229_r0d;
  wire c229_r1d;
  wire c229_a;
  wire [33:0] c228_r0d;
  wire [33:0] c228_r1d;
  wire c228_a;
  wire c227_r;
  wire c227_a;
  wire c226_r0d;
  wire c226_r1d;
  wire c226_a;
  wire c225_r;
  wire c225_a;
  wire [32:0] c224_r0d;
  wire [32:0] c224_r1d;
  wire c224_a;
  wire c223_r;
  wire c223_a;
  wire c222_r;
  wire c222_a;
  wire c221_r;
  wire c221_a;
  wire c220_r;
  wire c220_a;
  wire c219_r0d;
  wire c219_r1d;
  wire c219_a;
  wire c218_r;
  wire c218_a;
  wire c217_r0d;
  wire c217_r1d;
  wire c217_a;
  wire c216_r;
  wire c216_a;
  wire c215_r;
  wire c215_a;
  wire c214_r;
  wire c214_a;
  wire c213_r;
  wire c213_a;
  wire c212_r;
  wire c212_a;
  wire c211_r;
  wire c211_a;
  wire c210_r0d;
  wire c210_r1d;
  wire c210_a;
  wire c209_r;
  wire c209_a;
  wire [34:0] c208_r0d;
  wire [34:0] c208_r1d;
  wire c208_a;
  wire c207_r;
  wire c207_a;
  wire [34:0] c206_r0d;
  wire [34:0] c206_r1d;
  wire c206_a;
  wire c205_r;
  wire c205_a;
  wire c204_r;
  wire c204_a;
  wire c203_r;
  wire c203_a;
  wire [34:0] c202_r0d;
  wire [34:0] c202_r1d;
  wire c202_a;
  wire c201_r;
  wire c201_a;
  wire [2:0] c200_r0d;
  wire [2:0] c200_r1d;
  wire c200_a;
  wire c199_r;
  wire c199_a;
  wire [31:0] c198_r0d;
  wire [31:0] c198_r1d;
  wire c198_a;
  wire [35:0] c197_r0d;
  wire [35:0] c197_r1d;
  wire c197_a;
  wire c196_r;
  wire c196_a;
  wire c195_r;
  wire c195_a;
  wire [31:0] c194_r0d;
  wire [31:0] c194_r1d;
  wire c194_a;
  wire [34:0] c193_r0d;
  wire [34:0] c193_r1d;
  wire c193_a;
  wire c192_r;
  wire c192_a;
  wire c191_r;
  wire c191_a;
  wire [34:0] c190_r0d;
  wire [34:0] c190_r1d;
  wire c190_a;
  wire c189_r;
  wire c189_a;
  wire [1:0] c188_r0d;
  wire [1:0] c188_r1d;
  wire c188_a;
  wire [32:0] c187_r0d;
  wire [32:0] c187_r1d;
  wire c187_a;
  wire c186_r;
  wire c186_a;
  wire c185_r0d;
  wire c185_r1d;
  wire c185_a;
  wire c184_r;
  wire c184_a;
  wire [31:0] c183_r0d;
  wire [31:0] c183_r1d;
  wire c183_a;
  wire [35:0] c182_r0d;
  wire [35:0] c182_r1d;
  wire c182_a;
  wire c181_r;
  wire c181_a;
  wire c180_r;
  wire c180_a;
  wire [34:0] c179_r0d;
  wire [34:0] c179_r1d;
  wire c179_a;
  wire c178_r;
  wire c178_a;
  wire c177_r;
  wire c177_a;
  wire c176_r;
  wire c176_a;
  wire [34:0] c175_r0d;
  wire [34:0] c175_r1d;
  wire c175_a;
  wire c174_r;
  wire c174_a;
  wire c173_r;
  wire c173_a;
  wire [34:0] c172_r0d;
  wire [34:0] c172_r1d;
  wire c172_a;
  wire c171_r;
  wire c171_a;
  wire c170_r;
  wire c170_a;
  wire [34:0] c169_r0d;
  wire [34:0] c169_r1d;
  wire c169_a;
  wire c168_r;
  wire c168_a;
  wire c167_r;
  wire c167_a;
  wire [34:0] c166_r0d;
  wire [34:0] c166_r1d;
  wire c166_a;
  wire c165_r;
  wire c165_a;
  wire c164_r;
  wire c164_a;
  wire [34:0] c163_r0d;
  wire [34:0] c163_r1d;
  wire c163_a;
  wire c162_r;
  wire c162_a;
  wire c161_r;
  wire c161_a;
  wire [34:0] c160_r0d;
  wire [34:0] c160_r1d;
  wire c160_a;
  wire c159_r;
  wire c159_a;
  wire c158_r;
  wire c158_a;
  wire [34:0] c157_r0d;
  wire [34:0] c157_r1d;
  wire c157_a;
  wire c156_r;
  wire c156_a;
  wire c155_r;
  wire c155_a;
  wire [34:0] c154_r0d;
  wire [34:0] c154_r1d;
  wire c154_a;
  wire c153_r;
  wire c153_a;
  wire c152_r;
  wire c152_a;
  wire [3:0] c151_r0d;
  wire [3:0] c151_r1d;
  wire c151_a;
  wire [34:0] c150_r0d;
  wire [34:0] c150_r1d;
  wire c150_a;
  wire c149_r;
  wire c149_a;
  wire [3:0] c148_r0d;
  wire [3:0] c148_r1d;
  wire c148_a;
  wire c147_r;
  wire c147_a;
  wire c146_r;
  wire c146_a;
  wire c145_r0d;
  wire c145_r1d;
  wire c145_a;
  wire c144_r;
  wire c144_a;
  wire c143_r;
  wire c143_a;
  wire [34:0] c142_r0d;
  wire [34:0] c142_r1d;
  wire c142_a;
  wire c141_r;
  wire c141_a;
  wire [34:0] c140_r0d;
  wire [34:0] c140_r1d;
  wire c140_a;
  wire c139_r;
  wire c139_a;
  wire c138_r;
  wire c138_a;
  wire [34:0] c137_r0d;
  wire [34:0] c137_r1d;
  wire c137_a;
  wire c136_r;
  wire c136_a;
  wire [34:0] c135_r0d;
  wire [34:0] c135_r1d;
  wire c135_a;
  wire c134_r;
  wire c134_a;
  wire c133_r;
  wire c133_a;
  wire [34:0] c132_r0d;
  wire [34:0] c132_r1d;
  wire c132_a;
  wire c131_r;
  wire c131_a;
  wire c130_r;
  wire c130_a;
  wire [34:0] c129_r0d;
  wire [34:0] c129_r1d;
  wire c129_a;
  wire c128_r0d;
  wire c128_r1d;
  wire c128_a;
  wire c127_r;
  wire c127_a;
  wire c126_r;
  wire c126_a;
  wire c125_r0d;
  wire c125_r1d;
  wire c125_a;
  wire c124_r;
  wire c124_a;
  wire c123_r;
  wire c123_a;
  wire c122_r;
  wire c122_a;
  wire [34:0] c121_r0d;
  wire [34:0] c121_r1d;
  wire c121_a;
  wire [34:0] c120_r0d;
  wire [34:0] c120_r1d;
  wire c120_a;
  wire c119_r;
  wire c119_a;
  wire c118_r;
  wire c118_a;
  wire [34:0] c117_r0d;
  wire [34:0] c117_r1d;
  wire c117_a;
  wire [34:0] c116_r0d;
  wire [34:0] c116_r1d;
  wire c116_a;
  wire c115_r;
  wire c115_a;
  wire c114_r;
  wire c114_a;
  wire [34:0] c113_r0d;
  wire [34:0] c113_r1d;
  wire c113_a;
  wire [34:0] c112_r0d;
  wire [34:0] c112_r1d;
  wire c112_a;
  wire c111_r;
  wire c111_a;
  wire c110_r;
  wire c110_a;
  wire [34:0] c109_r0d;
  wire [34:0] c109_r1d;
  wire c109_a;
  wire [34:0] c108_r0d;
  wire [34:0] c108_r1d;
  wire c108_a;
  wire c107_r;
  wire c107_a;
  wire c106_r;
  wire c106_a;
  wire c105_r;
  wire c105_a;
  wire c104_r;
  wire c104_a;
  wire c103_r;
  wire c103_a;
  wire c102_r;
  wire c102_a;
  wire c101_r;
  wire c101_a;
  wire c100_r0d;
  wire c100_r1d;
  wire c100_a;
  wire c99_r;
  wire c99_a;
  wire c98_r0d;
  wire c98_r1d;
  wire c98_a;
  wire c97_r;
  wire c97_a;
  wire [34:0] c96_r0d;
  wire [34:0] c96_r1d;
  wire c96_a;
  wire c95_r;
  wire c95_a;
  wire [35:0] c94_r0d;
  wire [35:0] c94_r1d;
  wire c94_a;
  wire c93_r;
  wire c93_a;
  wire [34:0] c92_r0d;
  wire [34:0] c92_r1d;
  wire c92_a;
  wire c91_r;
  wire c91_a;
  wire c90_r;
  wire c90_a;
  wire [35:0] c89_r0d;
  wire [35:0] c89_r1d;
  wire c89_a;
  wire c88_r;
  wire c88_a;
  wire c87_r;
  wire c87_a;
  wire [34:0] c86_r0d;
  wire [34:0] c86_r1d;
  wire c86_a;
  wire c85_r;
  wire c85_a;
  wire c84_r;
  wire c84_a;
  wire c83_r;
  wire c83_a;
  wire [3:0] c82_r0d;
  wire [3:0] c82_r1d;
  wire c82_a;
  wire c81_r;
  wire c81_a;
  wire c80_r;
  wire c80_a;
  wire [34:0] c79_r0d;
  wire [34:0] c79_r1d;
  wire c79_a;
  wire c78_r;
  wire c78_a;
  wire c77_r;
  wire c77_a;
  wire [35:0] c76_r0d;
  wire [35:0] c76_r1d;
  wire c76_a;
  wire c75_r;
  wire c75_a;
  wire c74_r;
  wire c74_a;
  wire c73_r;
  wire c73_a;
  wire c72_r;
  wire c72_a;
  wire c71_r;
  wire c71_a;
  wire c70_r0d;
  wire c70_r1d;
  wire c70_a;
  wire c69_r;
  wire c69_a;
  wire [31:0] c68_r0d;
  wire [31:0] c68_r1d;
  wire c68_a;
  wire c67_r;
  wire c67_a;
  wire [34:0] c66_r0d;
  wire [34:0] c66_r1d;
  wire c66_a;
  wire c65_r;
  wire c65_a;
  wire c64_r0d;
  wire c64_r1d;
  wire c64_a;
  wire [33:0] c63_r0d;
  wire [33:0] c63_r1d;
  wire c63_a;
  wire c62_r;
  wire c62_a;
  wire c61_r0d;
  wire c61_r1d;
  wire c61_a;
  wire [32:0] c60_r0d;
  wire [32:0] c60_r1d;
  wire c60_a;
  wire c59_r;
  wire c59_a;
  wire [31:0] c58_r0d;
  wire [31:0] c58_r1d;
  wire c58_a;
  wire c57_r;
  wire c57_a;
  wire c56_r0d;
  wire c56_r1d;
  wire c56_a;
  wire c55_r;
  wire c55_a;
  wire c54_r0d;
  wire c54_r1d;
  wire c54_a;
  wire c53_r;
  wire c53_a;
  wire c52_r;
  wire c52_a;
  wire c51_r;
  wire c51_a;
  wire [31:0] c50_r0d;
  wire [31:0] c50_r1d;
  wire c50_a;
  wire c49_r;
  wire c49_a;
  wire c48_r;
  wire c48_a;
  wire [31:0] c47_r0d;
  wire [31:0] c47_r1d;
  wire c47_a;
  wire c46_r;
  wire c46_a;
  wire c45_r;
  wire c45_a;
  wire [34:0] c44_r0d;
  wire [34:0] c44_r1d;
  wire c44_a;
  wire c43_r;
  wire c43_a;
  wire [32:0] c42_r0d;
  wire [32:0] c42_r1d;
  wire c42_a;
  wire [1:0] c41_r0d;
  wire [1:0] c41_r1d;
  wire c41_a;
  wire c40_r;
  wire c40_a;
  wire c39_r;
  wire c39_a;
  wire c38_r;
  wire c38_a;
  wire [34:0] c37_r0d;
  wire [34:0] c37_r1d;
  wire c37_a;
  wire c36_r;
  wire c36_a;
  wire [33:0] c35_r0d;
  wire [33:0] c35_r1d;
  wire c35_a;
  wire c34_r0d;
  wire c34_r1d;
  wire c34_a;
  wire c33_r;
  wire c33_a;
  wire c32_r;
  wire c32_a;
  wire c31_r;
  wire c31_a;
  wire [34:0] c30_r0d;
  wire [34:0] c30_r1d;
  wire c30_a;
  wire c29_r;
  wire c29_a;
  wire c28_r;
  wire c28_a;
  wire c27_r0d;
  wire c27_r1d;
  wire c27_a;
  wire c26_r;
  wire c26_a;
  wire c25_r;
  wire c25_a;
  wire c24_r0d;
  wire c24_r1d;
  wire c24_a;
  wire c23_r;
  wire c23_a;
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I0 (c479_r0d, c479_r1d, c479_a, c297_r, c297_a, c351_r, c351_a, initialise);
  BrzJ_l11__280_202_29 I1 (c475_r, c475_a, c478_r0d, c478_r1d, c478_a, c479_r0d, c479_r1d, c479_a, initialise);
  BrzM_2_2 I2 (c476_r0d, c476_r1d, c476_a, c477_r0d, c477_r1d, c477_a, c478_r0d, c478_r1d, c478_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I3 (c472_r, c472_a, c477_r0d, c477_r1d, c477_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I4 (c470_r, c470_a, c476_r0d, c476_r1d, c476_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I5 (c474_r0d, c474_r1d, c474_a, c475_r, c475_a, n_0r0d, n_0r1d, n_0a, initialise);
  BrzM_1_2 I6 (c471_r0d, c471_r1d, c471_a, c473_r0d, c473_r1d, c473_a, c474_r0d, c474_r1d, c474_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I7 (c349_r0d, c349_r1d, c349_a, c472_r, c472_a, c473_r0d, c473_r1d, c473_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I8 (c295_r0d, c295_r1d, c295_a, c470_r, c470_a, c471_r0d, c471_r1d, c471_a, initialise);
  BrzS_3_l11__280_203_29_l141__28_28_28_281__m64m I9 (c469_r0d, c469_r1d, c469_a, c294_r, c294_a, c344_r, c344_a, c347_r, c347_a, initialise);
  BrzJ_l11__280_203_29 I10 (c464_r, c464_a, c468_r0d, c468_r1d, c468_a, c469_r0d, c469_r1d, c469_a, initialise);
  BrzM_3_3 I11 (c465_r0d, c465_r1d, c465_a, c466_r0d, c466_r1d, c466_a, c467_r0d, c467_r1d, c467_a, c468_r0d, c468_r1d, c468_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I12 (c461_r, c461_a, c467_r0d, c467_r1d, c467_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I13 (c459_r, c459_a, c466_r0d, c466_r1d, c466_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I14 (c457_r, c457_a, c465_r0d, c465_r1d, c465_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I15 (c463_r0d, c463_r1d, c463_a, c464_r, c464_a, z_0r0d, z_0r1d, z_0a, initialise);
  BrzM_1_3 I16 (c458_r0d, c458_r1d, c458_a, c460_r0d, c460_r1d, c460_a, c462_r0d, c462_r1d, c462_a, c463_r0d, c463_r1d, c463_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I17 (c345_r0d, c345_r1d, c345_a, c461_r, c461_a, c462_r0d, c462_r1d, c462_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I18 (c342_r0d, c342_r1d, c342_a, c459_r, c459_a, c460_r0d, c460_r1d, c460_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I19 (c292_r0d, c292_r1d, c292_a, c457_r, c457_a, c458_r0d, c458_r1d, c458_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I20 (c456_r0d, c456_r1d, c456_a, c291_r, c291_a, c330_r, c330_a, initialise);
  BrzJ_l11__280_202_29 I21 (c452_r, c452_a, c455_r0d, c455_r1d, c455_a, c456_r0d, c456_r1d, c456_a, initialise);
  BrzM_2_2 I22 (c453_r0d, c453_r1d, c453_a, c454_r0d, c454_r1d, c454_a, c455_r0d, c455_r1d, c455_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I23 (c449_r, c449_a, c454_r0d, c454_r1d, c454_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I24 (c447_r, c447_a, c453_r0d, c453_r1d, c453_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I25 (c451_r0d, c451_r1d, c451_a, c452_r, c452_a, pL_0r0d, pL_0r1d, pL_0a, initialise);
  BrzM_32_2 I26 (c448_r0d, c448_r1d, c448_a, c450_r0d, c450_r1d, c450_a, c451_r0d, c451_r1d, c451_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I27 (c328_r0d, c328_r1d, c328_a, c449_r, c449_a, c450_r0d, c450_r1d, c450_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I28 (c289_r0d, c289_r1d, c289_a, c447_r, c447_a, c448_r0d, c448_r1d, c448_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I29 (c325_r0d, c325_r1d, c325_a, c327_r, c327_a, pH_0r0d, pH_0r1d, pH_0a, initialise);
  BrzS_4_l11__281_203_29_l141__28_28_28_281__m67m I30 (c446_r0d, c446_r1d, c446_a, c70_r0d, c70_r1d, c70_a, c281_r0d, c281_r1d, c281_a, c318_r0d, c318_r1d, c318_a, initialise);
  BrzJ_l11__281_203_29 I31 (racN_0r0d, racN_0r1d, racN_0a, c445_r0d, c445_r1d, c445_a, c446_r0d, c446_r1d, c446_a, initialise);
  BrzM_3_3 I32 (c442_r0d, c442_r1d, c442_a, c443_r0d, c443_r1d, c443_a, c444_r0d, c444_r1d, c444_a, c445_r0d, c445_r1d, c445_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I33 (c322_r, c322_a, c444_r0d, c444_r1d, c444_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I34 (c285_r, c285_a, c443_r0d, c443_r1d, c443_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I35 (c74_r, c74_a, c442_r0d, c442_r1d, c442_a);
  BrzS_35_l12__2832_203_29_l144__28_28_28_28_m70m I36 (c441_r0d, c441_r1d, c441_a, c68_r0d, c68_r1d, c68_a, c279_r0d, c279_r1d, c279_a, c316_r0d, c316_r1d, c316_a, initialise);
  BrzJ_l12__2832_203_29 I37 (raS_0r0d, raS_0r1d, raS_0a, c440_r0d, c440_r1d, c440_a, c441_r0d, c441_r1d, c441_a, initialise);
  BrzM_3_3 I38 (c437_r0d, c437_r1d, c437_a, c438_r0d, c438_r1d, c438_a, c439_r0d, c439_r1d, c439_a, c440_r0d, c440_r1d, c440_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I39 (c321_r, c321_a, c439_r0d, c439_r1d, c439_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I40 (c284_r, c284_a, c438_r0d, c438_r1d, c438_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I41 (c73_r, c73_a, c437_r0d, c437_r1d, c437_a);
  BrzS_3_l11__280_203_29_l141__28_28_28_281__m64m I42 (c436_r0d, c436_r1d, c436_a, c55_r, c55_a, c260_r, c260_a, c313_r, c313_a, initialise);
  BrzJ_l11__280_203_29 I43 (c431_r, c431_a, c435_r0d, c435_r1d, c435_a, c436_r0d, c436_r1d, c436_a, initialise);
  BrzM_3_3 I44 (c432_r0d, c432_r1d, c432_a, c433_r0d, c433_r1d, c433_a, c434_r0d, c434_r1d, c434_a, c435_r0d, c435_r1d, c435_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I45 (c428_r, c428_a, c434_r0d, c434_r1d, c434_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I46 (c426_r, c426_a, c433_r0d, c433_r1d, c433_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I47 (c424_r, c424_a, c432_r0d, c432_r1d, c432_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I48 (c430_r0d, c430_r1d, c430_a, c431_r, c431_a, rac0_0r0d, rac0_0r1d, rac0_0a, initialise);
  BrzM_1_3 I49 (c425_r0d, c425_r1d, c425_a, c427_r0d, c427_r1d, c427_a, c429_r0d, c429_r1d, c429_a, c430_r0d, c430_r1d, c430_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I50 (c311_r0d, c311_r1d, c311_a, c428_r, c428_a, c429_r0d, c429_r1d, c429_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I51 (c259_r0d, c259_r1d, c259_a, c426_r, c426_a, c427_r0d, c427_r1d, c427_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I52 (c54_r0d, c54_r1d, c54_a, c424_r, c424_a, c425_r0d, c425_r1d, c425_a, initialise);
  BrzS_3_l11__280_203_29_l141__28_28_28_281__m64m I53 (c423_r0d, c423_r1d, c423_a, c52_r, c52_a, c257_r, c257_a, c310_r, c310_a, initialise);
  BrzJ_l11__280_203_29 I54 (c418_r, c418_a, c422_r0d, c422_r1d, c422_a, c423_r0d, c423_r1d, c423_a, initialise);
  BrzM_3_3 I55 (c419_r0d, c419_r1d, c419_a, c420_r0d, c420_r1d, c420_a, c421_r0d, c421_r1d, c421_a, c422_r0d, c422_r1d, c422_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I56 (c415_r, c415_a, c421_r0d, c421_r1d, c421_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I57 (c413_r, c413_a, c420_r0d, c420_r1d, c420_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I58 (c411_r, c411_a, c419_r0d, c419_r1d, c419_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I59 (c417_r0d, c417_r1d, c417_a, c418_r, c418_a, raB_0r0d, raB_0r1d, raB_0a, initialise);
  BrzM_32_3 I60 (c412_r0d, c412_r1d, c412_a, c414_r0d, c414_r1d, c414_a, c416_r0d, c416_r1d, c416_a, c417_r0d, c417_r1d, c417_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I61 (c308_r0d, c308_r1d, c308_a, c415_r, c415_a, c416_r0d, c416_r1d, c416_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I62 (c255_r0d, c255_r1d, c255_a, c413_r, c413_a, c414_r0d, c414_r1d, c414_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I63 (c50_r0d, c50_r1d, c50_a, c411_r, c411_a, c412_r0d, c412_r1d, c412_a, initialise);
  BrzS_3_l11__280_203_29_l141__28_28_28_281__m64m I64 (c410_r0d, c410_r1d, c410_a, c49_r, c49_a, c254_r, c254_a, c307_r, c307_a, initialise);
  BrzJ_l11__280_203_29 I65 (c405_r, c405_a, c409_r0d, c409_r1d, c409_a, c410_r0d, c410_r1d, c410_a, initialise);
  BrzM_3_3 I66 (c406_r0d, c406_r1d, c406_a, c407_r0d, c407_r1d, c407_a, c408_r0d, c408_r1d, c408_a, c409_r0d, c409_r1d, c409_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I67 (c402_r, c402_a, c408_r0d, c408_r1d, c408_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I68 (c400_r, c400_a, c407_r0d, c407_r1d, c407_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I69 (c398_r, c398_a, c406_r0d, c406_r1d, c406_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I70 (c404_r0d, c404_r1d, c404_a, c405_r, c405_a, raA_0r0d, raA_0r1d, raA_0a, initialise);
  BrzM_32_3 I71 (c399_r0d, c399_r1d, c399_a, c401_r0d, c401_r1d, c401_a, c403_r0d, c403_r1d, c403_a, c404_r0d, c404_r1d, c404_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I72 (c305_r0d, c305_r1d, c305_a, c402_r, c402_a, c403_r0d, c403_r1d, c403_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I73 (c252_r0d, c252_r1d, c252_a, c400_r, c400_a, c401_r0d, c401_r1d, c401_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I74 (c47_r0d, c47_r1d, c47_a, c398_r, c398_a, c399_r0d, c399_r1d, c399_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I75 (c132_r0d, c132_r1d, c132_a, c134_r, c134_a, cs_0r0d, cs_0r1d, cs_0a, initialise);
  BrzS_9_l11__280_209_29_l424__28_28_28_281__m68m I76 (c397_r0d, c397_r1d, c397_a, c153_r, c153_a, c156_r, c156_a, c159_r, c159_a, c162_r, c162_a, c165_r, c165_a, c168_r, c168_a, c171_r, c171_a, c174_r, c174_a, c177_r, c177_a, initialise);
  BrzJ_l11__280_209_29 I77 (c386_r, c386_a, c396_r0d, c396_r1d, c396_a, c397_r0d, c397_r1d, c397_a, initialise);
  BrzM_9_9 I78 (c387_r0d, c387_r1d, c387_a, c388_r0d, c388_r1d, c388_a, c389_r0d, c389_r1d, c389_a, c390_r0d, c390_r1d, c390_a, c391_r0d, c391_r1d, c391_a, c392_r0d, c392_r1d, c392_a, c393_r0d, c393_r1d, c393_a, c394_r0d, c394_r1d, c394_a, c395_r0d, c395_r1d, c395_a, c396_r0d, c396_r1d, c396_a, initialise);
  BrzO_0_9_l25__28_28num_209_20256_29_29 I79 (c383_r, c383_a, c395_r0d, c395_r1d, c395_a);
  BrzO_0_9_l25__28_28num_209_20128_29_29 I80 (c381_r, c381_a, c394_r0d, c394_r1d, c394_a);
  BrzO_0_9_l24__28_28num_209_2064_29_29 I81 (c379_r, c379_a, c393_r0d, c393_r1d, c393_a);
  BrzO_0_9_l24__28_28num_209_2032_29_29 I82 (c377_r, c377_a, c392_r0d, c392_r1d, c392_a);
  BrzO_0_9_l24__28_28num_209_2016_29_29 I83 (c375_r, c375_a, c391_r0d, c391_r1d, c391_a);
  BrzO_0_9_l23__28_28num_209_208_29_29 I84 (c373_r, c373_a, c390_r0d, c390_r1d, c390_a);
  BrzO_0_9_l23__28_28num_209_204_29_29 I85 (c371_r, c371_a, c389_r0d, c389_r1d, c389_a);
  BrzO_0_9_l23__28_28num_209_202_29_29 I86 (c369_r, c369_a, c388_r0d, c388_r1d, c388_a);
  BrzO_0_9_l23__28_28num_209_201_29_29 I87 (c367_r, c367_a, c387_r0d, c387_r1d, c387_a);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I88 (c385_r0d, c385_r1d, c385_a, c386_r, c386_a, opB_0r0d, opB_0r1d, opB_0a, initialise);
  BrzM_35_9 I89 (c368_r0d, c368_r1d, c368_a, c370_r0d, c370_r1d, c370_a, c372_r0d, c372_r1d, c372_a, c374_r0d, c374_r1d, c374_a, c376_r0d, c376_r1d, c376_a, c378_r0d, c378_r1d, c378_a, c380_r0d, c380_r1d, c380_a, c382_r0d, c382_r1d, c382_a, c384_r0d, c384_r1d, c384_a, c385_r0d, c385_r1d, c385_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I90 (c175_r0d, c175_r1d, c175_a, c383_r, c383_a, c384_r0d, c384_r1d, c384_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I91 (c172_r0d, c172_r1d, c172_a, c381_r, c381_a, c382_r0d, c382_r1d, c382_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I92 (c169_r0d, c169_r1d, c169_a, c379_r, c379_a, c380_r0d, c380_r1d, c380_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I93 (c166_r0d, c166_r1d, c166_a, c377_r, c377_a, c378_r0d, c378_r1d, c378_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I94 (c163_r0d, c163_r1d, c163_a, c375_r, c375_a, c376_r0d, c376_r1d, c376_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I95 (c160_r0d, c160_r1d, c160_a, c373_r, c373_a, c374_r0d, c374_r1d, c374_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I96 (c157_r0d, c157_r1d, c157_a, c371_r, c371_a, c372_r0d, c372_r1d, c372_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I97 (c154_r0d, c154_r1d, c154_a, c369_r, c369_a, c370_r0d, c370_r1d, c370_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I98 (c150_r0d, c150_r1d, c150_a, c367_r, c367_a, c368_r0d, c368_r1d, c368_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I99 (c129_r0d, c129_r1d, c129_a, c131_r, c131_a, opA_0r0d, opA_0r1d, opA_0a, initialise);
  BrzJ_l11__281_200_29 I100 (done_0r0d, done_0r1d, done_0a, c221_r, c221_a, c219_r0d, c219_r1d, c219_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I101 (c366_r0d, c366_r1d, c366_a, c126_r, c126_a, c248_r, c248_a, initialise);
  BrzJ_l11__280_202_29 I102 (c362_r, c362_a, c365_r0d, c365_r1d, c365_a, c366_r0d, c366_r1d, c366_a, initialise);
  BrzM_2_2 I103 (c363_r0d, c363_r1d, c363_a, c364_r0d, c364_r1d, c364_a, c365_r0d, c365_r1d, c365_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I104 (c359_r, c359_a, c364_r0d, c364_r1d, c364_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I105 (c357_r, c357_a, c363_r0d, c363_r1d, c363_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I106 (c361_r0d, c361_r1d, c361_a, c362_r, c362_a, load_0r0d, load_0r1d, load_0a, initialise);
  BrzM_1_2 I107 (c358_r0d, c358_r1d, c358_a, c360_r0d, c360_r1d, c360_a, c361_r0d, c361_r1d, c361_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I108 (c247_r0d, c247_r1d, c247_a, c359_r, c359_a, c360_r0d, c360_r1d, c360_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I109 (c125_r0d, c125_r1d, c125_a, c357_r, c357_a, c358_r0d, c358_r1d, c358_a, initialise);
  BrzJ_l11__281_200_29 I110 (macc_0r0d, macc_0r1d, macc_0a, c107_r, c107_a, c100_r0d, c100_r1d, c100_a, initialise);
  BrzJ_l11__281_200_29 I111 (mlength_0r0d, mlength_0r1d, mlength_0a, c106_r, c106_a, c98_r0d, c98_r1d, c98_a, initialise);
  BrzJ_l12__2835_200_29 I112 (c_0r0d, c_0r1d, c_0a, c105_r, c105_a, c96_r0d, c96_r1d, c96_a, initialise);
  BrzJ_l12__2836_200_29 I113 (b_0r0d, b_0r1d, b_0a, c104_r, c104_a, c94_r0d, c94_r1d, c94_a, initialise);
  BrzJ_l12__2835_200_29 I114 (a_0r0d, a_0r1d, a_0a, c103_r, c103_a, c92_r0d, c92_r1d, c92_a, initialise);
  BrzJ_l12__2835_200_29 I115 (res_0r0d, res_0r1d, res_0a, c139_r, c139_a, c137_r0d, c137_r1d, c137_a, initialise);
  BrzJ_l12__2835_200_29 I116 (cin_0r0d, cin_0r1d, cin_0a, c144_r, c144_a, c142_r0d, c142_r1d, c142_a, initialise);
  BrzJ_l12__2835_200_29 I117 (c356_r0d, c356_r1d, c356_a, c213_r, c213_a, c206_r0d, c206_r1d, c206_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I118 (c135_r0d, c135_r1d, c135_a, c136_r, c136_a, c356_r0d, c356_r1d, c356_a, initialise);
  BrzJ_l12__2835_200_29 I119 (c355_r0d, c355_r1d, c355_a, c214_r, c214_a, c208_r0d, c208_r1d, c208_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I120 (c140_r0d, c140_r1d, c140_a, c141_r, c141_a, c355_r0d, c355_r1d, c355_a, initialise);
  BrzJ_l11__281_200_29 I121 (c354_r0d, c354_r1d, c354_a, c215_r, c215_a, c210_r0d, c210_r1d, c210_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I122 (c145_r0d, c145_r1d, c145_a, c147_r, c147_a, c354_r0d, c354_r1d, c354_a, initialise);
  BrzV_4_l6__28_29_l43__28_28_280_204_29_29__m77m I123 (c243_r0d, c243_r1d, c243_a, c82_r0d, c82_r1d, c82_a, c245_r, c245_a, c84_r, c84_a, c152_r, c152_a, c149_r, c149_a, c146_r, c146_a, c151_r0d, c151_r1d, c151_a, c148_r0d, c148_r1d, c148_a, c145_r0d, c145_r1d, c145_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m83m I124 (c314_r0d, c314_r1d, c314_a, c315_r, c315_a, c350_r, c350_a, c334_r, c334_a, c326_r, c326_a, c349_r0d, c349_r1d, c349_a, c333_r0d, c333_r1d, c333_a, c325_r0d, c325_r1d, c325_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m81m I125 (c261_r0d, c261_r1d, c261_a, c263_r, c263_a, c329_r, c329_a, c290_r, c290_a, c328_r0d, c328_r1d, c328_a, c289_r0d, c289_r1d, c289_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m90m I126 (c30_r0d, c30_r1d, c30_a, c32_r, c32_a, c155_r, c155_a, c110_r, c110_a, c154_r0d, c154_r1d, c154_a, c109_r0d, c109_r1d, c109_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m90m I127 (c37_r0d, c37_r1d, c37_a, c39_r, c39_a, c158_r, c158_a, c114_r, c114_a, c157_r0d, c157_r1d, c157_a, c113_r0d, c113_r1d, c113_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m90m I128 (c66_r0d, c66_r1d, c66_a, c67_r, c67_a, c161_r, c161_a, c118_r, c118_a, c160_r0d, c160_r1d, c160_a, c117_r0d, c117_r1d, c117_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m90m I129 (c44_r0d, c44_r1d, c44_a, c46_r, c46_a, c164_r, c164_a, c122_r, c122_a, c163_r0d, c163_r1d, c163_a, c121_r0d, c121_r1d, c121_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I130 (c108_r0d, c108_r1d, c108_a, c111_r, c111_a, c176_r, c176_a, c175_r0d, c175_r1d, c175_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I131 (c112_r0d, c112_r1d, c112_a, c115_r, c115_a, c173_r, c173_a, c172_r0d, c172_r1d, c172_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I132 (c116_r0d, c116_r1d, c116_a, c119_r, c119_a, c170_r, c170_a, c169_r0d, c169_r1d, c169_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I133 (c120_r0d, c120_r1d, c120_a, c123_r, c123_a, c167_r, c167_a, c166_r0d, c166_r1d, c166_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m92m I134 (c179_r0d, c179_r1d, c179_a, c181_r, c181_a, c309_r, c309_a, c230_r, c230_a, c227_r, c227_a, c225_r, c225_a, c308_r0d, c308_r1d, c308_a, c229_r0d, c229_r1d, c229_a, c226_r0d, c226_r1d, c226_a, c224_r0d, c224_r1d, c224_a, initialise);
  BrzV_36_l6__28_29_l24__28_28_280_2036_29_2_m96m I135 (c182_r0d, c182_r1d, c182_a, c192_r, c192_a, c256_r, c256_a, c235_r, c235_a, c255_r0d, c255_r1d, c255_a, c234_r0d, c234_r1d, c234_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m86m I136 (c193_r0d, c193_r1d, c193_a, c196_r, c196_a, c304_r, c304_a, c238_r, c238_a, c303_r0d, c303_r1d, c303_a, c237_r0d, c237_r1d, c237_a, initialise);
  BrzV_36_l6__28_29_l24__28_28_280_2036_29_2_m97m I137 (c197_r0d, c197_r1d, c197_a, c204_r, c204_a, c302_r, c302_a, c253_r, c253_a, c244_r, c244_a, c241_r, c241_a, c301_r0d, c301_r1d, c301_a, c252_r0d, c252_r1d, c252_a, c243_r0d, c243_r1d, c243_a, c240_r0d, c240_r1d, c240_a, initialise);
  BrzV_35_l6__28_29_l45__28_28_280_2035_29_2_m94m I138 (c237_r0d, c237_r1d, c237_a, c79_r0d, c79_r1d, c79_a, c239_r, c239_a, c81_r, c81_a, c130_r, c130_a, c129_r0d, c129_r1d, c129_a, initialise);
  BrzV_35_l6__28_29_l45__28_28_280_2035_29_2_m94m I139 (c231_r0d, c231_r1d, c231_a, c86_r0d, c86_r1d, c86_a, c233_r, c233_a, c87_r, c87_a, c133_r, c133_a, c132_r0d, c132_r1d, c132_a, initialise);
  BrzV_36_l6__28_29_l45__28_28_280_2036_29_2_m98m I140 (c234_r0d, c234_r1d, c234_a, c89_r0d, c89_r1d, c89_a, c236_r, c236_a, c90_r, c90_a, c184_r, c184_a, c183_r0d, c183_r1d, c183_a, initialise);
  BrzV_36_l6__28_29_l45__28_28_280_2036_29_2_m98m I141 (c240_r0d, c240_r1d, c240_a, c76_r0d, c76_r1d, c76_a, c242_r, c242_a, c78_r, c78_a, c199_r, c199_a, c198_r0d, c198_r1d, c198_a, initialise);
  BrzV_1_l6__28_29_l43__28_28_280_201_29_29__m74m I142 (c264_r0d, c264_r1d, c264_a, c217_r0d, c217_r1d, c217_a, c266_r, c266_a, c218_r, c218_a, c312_r, c312_a, c223_r, c223_a, c311_r0d, c311_r1d, c311_a, c128_r0d, c128_r1d, c128_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I143 (c24_r0d, c24_r1d, c24_a, c26_r, c26_a, c287_r, c287_a, c288_r0d, c288_r1d, c288_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I144 (c27_r0d, c27_r1d, c27_a, c29_r, c29_a, c332_r, c332_a, c331_r0d, c331_r1d, c331_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m73m I145 (c275_r0d, c275_r1d, c275_a, c277_r, c277_a, c346_r, c346_a, c340_r, c340_a, c293_r, c293_a, c345_r0d, c345_r1d, c345_a, c339_r0d, c339_r1d, c339_a, c292_r0d, c292_r1d, c292_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I146 (c267_r0d, c267_r1d, c267_a, c269_r, c269_a, c296_r, c296_a, c295_r0d, c295_r1d, c295_a, initialise);
  BrzM_0_2 I147 (go_0r, go_0a, c353_r, c353_a, c23_r, c23_a, initialise);
  BrzM_0_2 I148 (c299_r, c299_a, c352_r, c352_a, c353_r, c353_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I149 (c288_r0d, c288_r1d, c288_a, c298_r, c298_a, c300_r, c300_a, initialise);
  BrzJ_l19__280_200_200_200_29 I150 (c327_r, c327_a, c330_r, c330_a, c348_r, c348_a, c351_r, c351_a, c352_r, c352_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I151 (c324_r, c324_a, c326_r, c326_a, c329_r, c329_a, c332_r, c332_a, c350_r, c350_a, initialise);
  BrzM_0_2 I152 (c344_r, c344_a, c347_r, c347_a, c348_r, c348_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I153 (c331_r0d, c331_r1d, c331_a, c343_r, c343_a, c346_r, c346_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I154 (c343_r, c343_a, c334_r, c334_a, c335_r, c335_a, c340_r, c340_a, initialise);
  BrzO_2_1_l119__28_28app_201_20_280_200_201_m47m I155 (c341_r0d, c341_r1d, c341_a, c342_r0d, c342_r1d, c342_a);
  BrzJ_l11__281_201_29 I156 (c338_r0d, c338_r1d, c338_a, c339_r0d, c339_r1d, c339_a, c341_r0d, c341_r1d, c341_a, initialise);
  BrzO_33_1_l196__28_28app_201_20_280_200_20_m52m I157 (c337_r0d, c337_r1d, c337_a, c338_r0d, c338_r1d, c338_a);
  BrzJ_l12__2832_201_29 I158 (c333_r0d, c333_r1d, c333_a, c336_r0d, c336_r1d, c336_a, c337_r0d, c337_r1d, c337_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I159 (c335_r, c335_a, c336_r0d, c336_r1d, c336_a);
  BrzJ_l19__280_200_200_200_29 I160 (c307_r, c307_a, c310_r, c310_a, c313_r, c313_a, c315_r, c315_a, c324_r, c324_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I161 (c300_r, c300_a, c306_r, c306_a, c309_r, c309_a, c312_r, c312_a, c323_r, c323_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I162 (c323_r, c323_a, c321_r, c321_a, c322_r, c322_a, initialise);
  BrzJ_l11__280_200_29 I163 (c317_r, c317_a, c319_r, c319_a, c320_r, c320_a, initialise);
  BrzF_1_l17__28_280_200_29_29 I164 (c318_r0d, c318_r1d, c318_a, c319_r, c319_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I165 (c316_r0d, c316_r1d, c316_a, c317_r, c317_a, c320_r, c320_a, c314_r0d, c314_r1d, c314_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I166 (c306_r, c306_a, c302_r, c302_a, c304_r, c304_a, initialise);
  BrzJ_l12__281_2031_29 I167 (c301_r0d, c301_r1d, c301_a, c303_r0d, c303_r1d, c303_a, c305_r0d, c305_r1d, c305_a, initialise);
  BrzJ_l15__280_200_200_29 I168 (c291_r, c291_a, c294_r, c294_a, c297_r, c297_a, c299_r, c299_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I169 (c298_r, c298_a, c290_r, c290_a, c293_r, c293_a, c296_r, c296_a, initialise);
  BrzJ_l19__280_200_200_200_29 I170 (c254_r, c254_a, c257_r, c257_a, c260_r, c260_a, c278_r, c278_a, c287_r, c287_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I171 (c251_r, c251_a, c253_r, c253_a, c256_r, c256_a, c258_r, c258_a, c286_r, c286_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I172 (c286_r, c286_a, c284_r, c284_a, c285_r, c285_a, initialise);
  BrzJ_l11__280_200_29 I173 (c280_r, c280_a, c282_r, c282_a, c283_r, c283_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I174 (c281_r0d, c281_r1d, c281_a, c282_r, c282_a, c265_r, c265_a, c264_r0d, c264_r1d, c264_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m82m I175 (c279_r0d, c279_r1d, c279_a, c280_r, c280_a, c262_r, c262_a, c268_r, c268_a, c271_r, c271_a, c261_r0d, c261_r1d, c261_a, c267_r0d, c267_r1d, c267_a, c270_r0d, c270_r1d, c270_a, initialise);
  BrzJ_l19__280_200_200_200_29 I176 (c263_r, c263_a, c266_r, c266_a, c269_r, c269_a, c277_r, c277_a, c278_r, c278_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I177 (c283_r, c283_a, c262_r, c262_a, c265_r, c265_a, c268_r, c268_a, c276_r, c276_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I178 (c276_r, c276_a, c271_r, c271_a, c272_r, c272_a, initialise);
  BrzO_33_1_l196__28_28app_201_20_280_200_20_m52m I179 (c274_r0d, c274_r1d, c274_a, c275_r0d, c275_r1d, c275_a);
  BrzJ_l12__2832_201_29 I180 (c270_r0d, c270_r1d, c270_a, c273_r0d, c273_r1d, c273_a, c274_r0d, c274_r1d, c274_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I181 (c272_r, c272_a, c273_r0d, c273_r1d, c273_a);
  BrzO_0_1_l23__28_28num_201_200_29_29 I182 (c258_r, c258_a, c259_r0d, c259_r1d, c259_a);
  BrzM_0_2 I183 (c127_r, c127_a, c250_r, c250_a, c222_r, c222_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I184 (c128_r0d, c128_r1d, c128_a, c251_r, c251_a, c249_r, c249_a, initialise);
  BrzJ_l27__280_200_200_200_200_200_29 I185 (c233_r, c233_a, c236_r, c236_a, c239_r, c239_a, c242_r, c242_a, c245_r, c245_a, c248_r, c248_a, c250_r, c250_a, initialise);
  BrzF_0_l87__28_280_200_29_20_280_200_29_20_m36m I186 (c249_r, c249_a, c232_r, c232_a, c235_r, c235_a, c238_r, c238_a, c241_r, c241_a, c244_r, c244_a, c246_r, c246_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I187 (c246_r, c246_a, c247_r0d, c247_r1d, c247_a);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I188 (c232_r, c232_a, c225_r, c225_a, c227_r, c227_a, c230_r, c230_a, initialise);
  BrzJ_l12__2834_201_29 I189 (c228_r0d, c228_r1d, c228_a, c229_r0d, c229_r1d, c229_a, c231_r0d, c231_r1d, c231_a, initialise);
  BrzJ_l12__2833_201_29 I190 (c224_r0d, c224_r1d, c224_a, c226_r0d, c226_r1d, c226_a, c228_r0d, c228_r1d, c228_a, initialise);
  BrzJ_l35__280_200_200_200_200_200_200_200__m45m I191 (c131_r, c131_a, c134_r, c134_a, c136_r, c136_a, c141_r, c141_a, c147_r, c147_a, c178_r, c178_a, c205_r, c205_a, c218_r, c218_a, c223_r, c223_a, initialise);
  BrzF_0_l115__28_280_200_29_20_280_200_29_2_m38m I192 (c222_r, c222_a, c130_r, c130_a, c133_r, c133_a, c139_r, c139_a, c144_r, c144_a, c146_r, c146_a, c149_r, c149_a, c216_r, c216_a, c221_r, c221_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I193 (c219_r0d, c219_r1d, c219_a, c220_r, c220_a, c220_r, c220_a, c217_r0d, c217_r1d, c217_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I194 (c216_r, c216_a, c213_r, c213_a, c214_r, c214_a, c215_r, c215_a, initialise);
  BrzJ_l15__280_200_200_29 I195 (c207_r, c207_a, c209_r, c209_a, c211_r, c211_a, c212_r, c212_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I196 (c210_r0d, c210_r1d, c210_a, c211_r, c211_a, c186_r, c186_a, c185_r0d, c185_r1d, c185_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m88m I197 (c208_r0d, c208_r1d, c208_a, c209_r, c209_a, c180_r, c180_a, c189_r, c189_a, c179_r0d, c179_r1d, c179_a, c188_r0d, c188_r1d, c188_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m93m I198 (c206_r0d, c206_r1d, c206_a, c207_r, c207_a, c195_r, c195_a, c201_r, c201_a, c194_r0d, c194_r1d, c194_a, c200_r0d, c200_r1d, c200_a, initialise);
  BrzJ_l19__280_200_200_200_29 I199 (c181_r, c181_a, c192_r, c192_a, c196_r, c196_a, c204_r, c204_a, c205_r, c205_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I200 (c212_r, c212_a, c180_r, c180_a, c191_r, c191_a, c195_r, c195_a, c203_r, c203_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I201 (c203_r, c203_a, c199_r, c199_a, c201_r, c201_a, initialise);
  BrzO_35_36_l76__28_28num_201_200_29_20_28a_m56m I202 (c202_r0d, c202_r1d, c202_a, c197_r0d, c197_r1d, c197_a);
  BrzJ_l12__2832_203_29 I203 (c198_r0d, c198_r1d, c198_a, c200_r0d, c200_r1d, c200_a, c202_r0d, c202_r1d, c202_a, initialise);
  BrzO_32_35_l91__28_28app_203_20_280_2031_2_m50m I204 (c194_r0d, c194_r1d, c194_a, c193_r0d, c193_r1d, c193_a);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I205 (c191_r, c191_a, c184_r, c184_a, c186_r, c186_a, c189_r, c189_a, initialise);
  BrzO_35_36_l76__28_28num_201_200_29_20_28a_m56m I206 (c190_r0d, c190_r1d, c190_a, c182_r0d, c182_r1d, c182_a);
  BrzJ_l12__2833_202_29 I207 (c187_r0d, c187_r1d, c187_a, c188_r0d, c188_r1d, c188_a, c190_r0d, c190_r1d, c190_a, initialise);
  BrzJ_l12__2832_201_29 I208 (c183_r0d, c183_r1d, c183_a, c185_r0d, c185_r1d, c185_a, c187_r0d, c187_r1d, c187_a, initialise);
  BrzM_0_9 I209 (c153_r, c153_a, c156_r, c156_a, c159_r, c159_a, c162_r, c162_a, c165_r, c165_a, c168_r, c168_a, c171_r, c171_a, c174_r, c174_a, c177_r, c177_a, c178_r, c178_a, initialise);
  BrzS_4_l11__280_204_29_l521__28_28_28_280__m66m I210 (c148_r0d, c148_r1d, c148_a, c152_r, c152_a, c155_r, c155_a, c158_r, c158_a, c161_r, c161_a, c164_r, c164_a, c167_r, c167_a, c170_r, c170_a, c173_r, c173_a, c176_r, c176_a, initialise);
  BrzO_4_35_l91__28_28app_2031_20_280_203_20_m48m I211 (c151_r0d, c151_r1d, c151_a, c150_r0d, c150_r1d, c150_a);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I212 (c142_r0d, c142_r1d, c142_a, c143_r, c143_a, c143_r, c143_a, c140_r0d, c140_r1d, c140_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I213 (c137_r0d, c137_r1d, c137_a, c138_r, c138_a, c138_r, c138_a, c135_r0d, c135_r1d, c135_a, initialise);
  BrzJ_l23__280_200_200_200_200_29 I214 (c111_r, c111_a, c115_r, c115_a, c119_r, c119_a, c123_r, c123_a, c126_r, c126_a, c127_r, c127_a, initialise);
  BrzF_0_l73__28_280_200_29_20_280_200_29_20_m35m I215 (c91_r, c91_a, c110_r, c110_a, c114_r, c114_a, c118_r, c118_a, c122_r, c122_a, c124_r, c124_a, initialise);
  BrzO_0_1_l23__28_28num_201_201_29_29 I216 (c124_r, c124_a, c125_r0d, c125_r1d, c125_a);
  BrzO_35_35_l34__28_28not_20_280_200_2035_2_m55m I217 (c121_r0d, c121_r1d, c121_a, c120_r0d, c120_r1d, c120_a);
  BrzO_35_35_l34__28_28not_20_280_200_2035_2_m55m I218 (c117_r0d, c117_r1d, c117_a, c116_r0d, c116_r1d, c116_a);
  BrzO_35_35_l34__28_28not_20_280_200_2035_2_m55m I219 (c113_r0d, c113_r1d, c113_a, c112_r0d, c112_r1d, c112_a);
  BrzO_35_35_l34__28_28not_20_280_200_2035_2_m55m I220 (c109_r0d, c109_r1d, c109_a, c108_r0d, c108_r1d, c108_a);
  BrzF_0_l73__28_280_200_29_20_280_200_29_20_m35m I221 (c23_r, c23_a, c103_r, c103_a, c104_r, c104_a, c105_r, c105_a, c106_r, c106_a, c107_r, c107_a, initialise);
  BrzJ_l23__280_200_200_200_200_29 I222 (c93_r, c93_a, c95_r, c95_a, c97_r, c97_a, c99_r, c99_a, c101_r, c101_a, c102_r, c102_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I223 (c100_r0d, c100_r1d, c100_a, c101_r, c101_a, c28_r, c28_a, c27_r0d, c27_r1d, c27_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I224 (c98_r0d, c98_r1d, c98_a, c99_r, c99_a, c25_r, c25_a, c24_r0d, c24_r1d, c24_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I225 (c96_r0d, c96_r1d, c96_a, c97_r, c97_a, c80_r, c80_a, c79_r0d, c79_r1d, c79_a, initialise);
  BrzV_36_l6__28_29_l24__28_28_280_2036_29_2_m95m I226 (c94_r0d, c94_r1d, c94_a, c95_r, c95_a, c77_r, c77_a, c83_r, c83_a, c76_r0d, c76_r1d, c76_a, c82_r0d, c82_r1d, c82_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m89m I227 (c92_r0d, c92_r1d, c92_a, c93_r, c93_a, c31_r, c31_a, c36_r, c36_a, c43_r, c43_a, c48_r, c48_a, c51_r, c51_a, c57_r, c57_a, c65_r, c65_a, c30_r0d, c30_r1d, c30_a, c35_r0d, c35_r1d, c35_a, c42_r0d, c42_r1d, c42_a, c47_r0d, c47_r1d, c47_a, c50_r0d, c50_r1d, c50_a, c56_r0d, c56_r1d, c56_a, c64_r0d, c64_r1d, c64_a, initialise);
  BrzJ_l59__280_200_200_200_200_200_200_200__m46m I228 (c26_r, c26_a, c29_r, c29_a, c32_r, c32_a, c39_r, c39_a, c46_r, c46_a, c49_r, c49_a, c52_r, c52_a, c55_r, c55_a, c67_r, c67_a, c78_r, c78_a, c81_r, c81_a, c84_r, c84_a, c87_r, c87_a, c90_r, c90_a, c91_r, c91_a, initialise);
  BrzF_0_l199__28_280_200_29_20_280_200_29_2_m39m I229 (c102_r, c102_a, c25_r, c25_a, c28_r, c28_a, c31_r, c31_a, c38_r, c38_a, c45_r, c45_a, c48_r, c48_a, c51_r, c51_a, c53_r, c53_a, c75_r, c75_a, c77_r, c77_a, c80_r, c80_a, c83_r, c83_a, c85_r, c85_a, c88_r, c88_a, initialise);
  BrzO_0_36_l24__28_28num_2036_200_29_29 I230 (c88_r, c88_a, c89_r0d, c89_r1d, c89_a);
  BrzO_0_35_l24__28_28num_2035_200_29_29 I231 (c85_r, c85_a, c86_r0d, c86_r1d, c86_a);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I232 (c75_r, c75_a, c73_r, c73_a, c74_r, c74_a, initialise);
  BrzJ_l11__280_200_29 I233 (c69_r, c69_a, c71_r, c71_a, c72_r, c72_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I234 (c70_r0d, c70_r1d, c70_a, c71_r, c71_a, c62_r, c62_a, c61_r0d, c61_r1d, c61_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I235 (c68_r0d, c68_r1d, c68_a, c69_r, c69_a, c59_r, c59_a, c58_r0d, c58_r1d, c58_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I236 (c72_r, c72_a, c57_r, c57_a, c59_r, c59_a, c62_r, c62_a, c65_r, c65_a, initialise);
  BrzJ_l12__2834_201_29 I237 (c63_r0d, c63_r1d, c63_a, c64_r0d, c64_r1d, c64_a, c66_r0d, c66_r1d, c66_a, initialise);
  BrzJ_l12__2833_201_29 I238 (c60_r0d, c60_r1d, c60_a, c61_r0d, c61_r1d, c61_a, c63_r0d, c63_r1d, c63_a, initialise);
  BrzJ_l12__281_2032_29 I239 (c56_r0d, c56_r1d, c56_a, c58_r0d, c58_r1d, c58_a, c60_r0d, c60_r1d, c60_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I240 (c53_r, c53_a, c54_r0d, c54_r1d, c54_a);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I241 (c45_r, c45_a, c40_r, c40_a, c43_r, c43_a, initialise);
  BrzJ_l12__282_2033_29 I242 (c41_r0d, c41_r1d, c41_a, c42_r0d, c42_r1d, c42_a, c44_r0d, c44_r1d, c44_a, initialise);
  BrzO_0_2_l23__28_28num_202_200_29_29 I243 (c40_r, c40_a, c41_r0d, c41_r1d, c41_a);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I244 (c38_r, c38_a, c33_r, c33_a, c36_r, c36_a, initialise);
  BrzJ_l12__281_2034_29 I245 (c34_r0d, c34_r1d, c34_a, c35_r0d, c35_r1d, c35_a, c37_r0d, c37_r1d, c37_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I246 (c33_r, c33_a, c34_r0d, c34_r1d, c34_a);
endmodule

module Balsa_CSAdder__DP2 (
  go_0r, go_0a,
  a_0r0d, a_0r1d, a_0a,
  b_0r0d, b_0r1d, b_0a,
  cs_0r0d, cs_0r1d, cs_0a,
  cout_0r0d, cout_0r1d, cout_0a,
  s_0r0d, s_0r1d, s_0a,
  initialise
);
  input go_0r;
  output go_0a;
  input [34:0] a_0r0d;
  input [34:0] a_0r1d;
  output a_0a;
  input [34:0] b_0r0d;
  input [34:0] b_0r1d;
  output b_0a;
  input [34:0] cs_0r0d;
  input [34:0] cs_0r1d;
  output cs_0a;
  output [34:0] cout_0r0d;
  output [34:0] cout_0r1d;
  input cout_0a;
  output [34:0] s_0r0d;
  output [34:0] s_0r1d;
  input s_0a;
  input initialise;
  wire c54_r;
  wire c54_a;
  wire c53_r;
  wire c53_a;
  wire c52_r;
  wire c52_a;
  wire c51_r;
  wire c51_a;
  wire c50_r;
  wire c50_a;
  wire c49_r;
  wire c49_a;
  wire [34:0] c48_r0d;
  wire [34:0] c48_r1d;
  wire c48_a;
  wire c47_r;
  wire c47_a;
  wire [34:0] c46_r0d;
  wire [34:0] c46_r1d;
  wire c46_a;
  wire c45_r;
  wire c45_a;
  wire [34:0] c44_r0d;
  wire [34:0] c44_r1d;
  wire c44_a;
  wire c43_r;
  wire c43_a;
  wire c42_r;
  wire c42_a;
  wire c41_r;
  wire c41_a;
  wire [34:0] c40_r0d;
  wire [34:0] c40_r1d;
  wire c40_a;
  wire [69:0] c39_r0d;
  wire [69:0] c39_r1d;
  wire c39_a;
  wire [34:0] c38_r0d;
  wire [34:0] c38_r1d;
  wire c38_a;
  wire [69:0] c37_r0d;
  wire [69:0] c37_r1d;
  wire c37_a;
  wire c36_r;
  wire c36_a;
  wire [34:0] c35_r0d;
  wire [34:0] c35_r1d;
  wire c35_a;
  wire c34_r;
  wire c34_a;
  wire [34:0] c33_r0d;
  wire [34:0] c33_r1d;
  wire c33_a;
  wire [34:0] c32_r0d;
  wire [34:0] c32_r1d;
  wire c32_a;
  wire [69:0] c31_r0d;
  wire [69:0] c31_r1d;
  wire c31_a;
  wire [34:0] c30_r0d;
  wire [34:0] c30_r1d;
  wire c30_a;
  wire [69:0] c29_r0d;
  wire [69:0] c29_r1d;
  wire c29_a;
  wire c28_r;
  wire c28_a;
  wire [34:0] c27_r0d;
  wire [34:0] c27_r1d;
  wire c27_a;
  wire c26_r;
  wire c26_a;
  wire [34:0] c25_r0d;
  wire [34:0] c25_r1d;
  wire c25_a;
  wire [34:0] c24_r0d;
  wire [34:0] c24_r1d;
  wire c24_a;
  wire [69:0] c23_r0d;
  wire [69:0] c23_r1d;
  wire c23_a;
  wire c22_r;
  wire c22_a;
  wire [34:0] c21_r0d;
  wire [34:0] c21_r1d;
  wire c21_a;
  wire c20_r;
  wire c20_a;
  wire [34:0] c19_r0d;
  wire [34:0] c19_r1d;
  wire c19_a;
  wire c18_r;
  wire c18_a;
  wire c17_r;
  wire c17_a;
  wire [34:0] c16_r0d;
  wire [34:0] c16_r1d;
  wire c16_a;
  wire [69:0] c15_r0d;
  wire [69:0] c15_r1d;
  wire c15_a;
  wire c14_r;
  wire c14_a;
  wire [34:0] c13_r0d;
  wire [34:0] c13_r1d;
  wire c13_a;
  wire [34:0] c12_r0d;
  wire [34:0] c12_r1d;
  wire c12_a;
  wire [69:0] c11_r0d;
  wire [69:0] c11_r1d;
  wire c11_a;
  wire c10_r;
  wire c10_a;
  wire [34:0] c9_r0d;
  wire [34:0] c9_r1d;
  wire c9_a;
  wire c8_r;
  wire c8_a;
  wire [34:0] c7_r0d;
  wire [34:0] c7_r1d;
  wire c7_a;
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I0 (c16_r0d, c16_r1d, c16_a, c18_r, c18_a, s_0r0d, s_0r1d, s_0a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I1 (c40_r0d, c40_r1d, c40_a, c42_r, c42_a, cout_0r0d, cout_0r1d, cout_0a, initialise);
  BrzJ_l12__2835_200_29 I2 (cs_0r0d, cs_0r1d, cs_0a, c53_r, c53_a, c48_r0d, c48_r1d, c48_a, initialise);
  BrzJ_l12__2835_200_29 I3 (b_0r0d, b_0r1d, b_0a, c52_r, c52_a, c46_r0d, c46_r1d, c46_a, initialise);
  BrzJ_l12__2835_200_29 I4 (a_0r0d, a_0r1d, a_0a, c51_r, c51_a, c44_r0d, c44_r1d, c44_a, initialise);
  BrzM_0_2 I5 (go_0r, go_0a, c43_r, c43_a, c54_r, c54_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I6 (c54_r, c54_a, c51_r, c51_a, c52_r, c52_a, c53_r, c53_a, initialise);
  BrzJ_l15__280_200_200_29 I7 (c45_r, c45_a, c47_r, c47_a, c49_r, c49_a, c50_r, c50_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m91m I8 (c48_r0d, c48_r1d, c48_a, c49_r, c49_a, c14_r, c14_a, c26_r, c26_a, c34_r, c34_a, c13_r0d, c13_r1d, c13_a, c25_r0d, c25_r1d, c25_a, c33_r0d, c33_r1d, c33_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m91m I9 (c46_r0d, c46_r1d, c46_a, c47_r, c47_a, c10_r, c10_a, c22_r, c22_a, c36_r, c36_a, c9_r0d, c9_r1d, c9_a, c21_r0d, c21_r1d, c21_a, c35_r0d, c35_r1d, c35_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m91m I10 (c44_r0d, c44_r1d, c44_a, c45_r, c45_a, c8_r, c8_a, c20_r, c20_a, c28_r, c28_a, c7_r0d, c7_r1d, c7_a, c19_r0d, c19_r1d, c19_a, c27_r0d, c27_r1d, c27_a, initialise);
  BrzJ_l11__280_200_29 I11 (c18_r, c18_a, c42_r, c42_a, c43_r, c43_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I12 (c50_r, c50_a, c17_r, c17_a, c41_r, c41_a, initialise);
  BrzF_0_l87__28_280_200_29_20_280_200_29_20_m36m I13 (c41_r, c41_a, c20_r, c20_a, c22_r, c22_a, c26_r, c26_a, c28_r, c28_a, c34_r, c34_a, c36_r, c36_a, initialise);
  BrzO_70_35_l123__28_28app_201_20_280_200_2_m59m I14 (c39_r0d, c39_r1d, c39_a, c40_r0d, c40_r1d, c40_a);
  BrzJ_l13__2835_2035_29 I15 (c32_r0d, c32_r1d, c32_a, c38_r0d, c38_r1d, c38_a, c39_r0d, c39_r1d, c39_a, initialise);
  BrzO_70_35_l124__28_28app_201_20_280_200_2_m58m I16 (c37_r0d, c37_r1d, c37_a, c38_r0d, c38_r1d, c38_a);
  BrzJ_l13__2835_2035_29 I17 (c33_r0d, c33_r1d, c33_a, c35_r0d, c35_r1d, c35_a, c37_r0d, c37_r1d, c37_a, initialise);
  BrzO_70_35_l123__28_28app_201_20_280_200_2_m59m I18 (c31_r0d, c31_r1d, c31_a, c32_r0d, c32_r1d, c32_a);
  BrzJ_l13__2835_2035_29 I19 (c24_r0d, c24_r1d, c24_a, c30_r0d, c30_r1d, c30_a, c31_r0d, c31_r1d, c31_a, initialise);
  BrzO_70_35_l124__28_28app_201_20_280_200_2_m58m I20 (c29_r0d, c29_r1d, c29_a, c30_r0d, c30_r1d, c30_a);
  BrzJ_l13__2835_2035_29 I21 (c25_r0d, c25_r1d, c25_a, c27_r0d, c27_r1d, c27_a, c29_r0d, c29_r1d, c29_a, initialise);
  BrzO_70_35_l124__28_28app_201_20_280_200_2_m58m I22 (c23_r0d, c23_r1d, c23_a, c24_r0d, c24_r1d, c24_a);
  BrzJ_l13__2835_2035_29 I23 (c19_r0d, c19_r1d, c19_a, c21_r0d, c21_r1d, c21_a, c23_r0d, c23_r1d, c23_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I24 (c17_r, c17_a, c8_r, c8_a, c10_r, c10_a, c14_r, c14_a, initialise);
  BrzO_70_35_l124__28_28app_201_20_280_200_2_m60m I25 (c15_r0d, c15_r1d, c15_a, c16_r0d, c16_r1d, c16_a);
  BrzJ_l13__2835_2035_29 I26 (c12_r0d, c12_r1d, c12_a, c13_r0d, c13_r1d, c13_a, c15_r0d, c15_r1d, c15_a, initialise);
  BrzO_70_35_l124__28_28app_201_20_280_200_2_m60m I27 (c11_r0d, c11_r1d, c11_a, c12_r0d, c12_r1d, c12_a);
  BrzJ_l13__2835_2035_29 I28 (c7_r0d, c7_r1d, c7_a, c9_r0d, c9_r1d, c9_a, c11_r0d, c11_r1d, c11_a, initialise);
endmodule

module Balsa_CPadder (
  go_0r, go_0a,
  a_0r0d, a_0r1d, a_0a,
  b_0r0d, b_0r1d, b_0a,
  c0_0r0d, c0_0r1d, c0_0a,
  s_0r0d, s_0r1d, s_0a,
  cN_0r0d, cN_0r1d, cN_0a,
  initialise
);
  input go_0r;
  output go_0a;
  input [31:0] a_0r0d;
  input [31:0] a_0r1d;
  output a_0a;
  input [31:0] b_0r0d;
  input [31:0] b_0r1d;
  output b_0a;
  input c0_0r0d;
  input c0_0r1d;
  output c0_0a;
  output [31:0] s_0r0d;
  output [31:0] s_0r1d;
  input s_0a;
  output cN_0r0d;
  output cN_0r1d;
  input cN_0a;
  input initialise;
  wire [32:0] c62_r0d;
  wire [32:0] c62_r1d;
  wire c62_a;
  wire [32:0] c61_r0d;
  wire [32:0] c61_r1d;
  wire c61_a;
  wire [33:0] c60_r0d;
  wire [33:0] c60_r1d;
  wire c60_a;
  wire c59_r;
  wire c59_a;
  wire c58_r;
  wire c58_a;
  wire c57_r;
  wire c57_a;
  wire c56_r;
  wire c56_a;
  wire [33:0] c55_r0d;
  wire [33:0] c55_r1d;
  wire c55_a;
  wire c54_r;
  wire c54_a;
  wire c53_r;
  wire c53_a;
  wire c52_r;
  wire c52_a;
  wire c51_r0d;
  wire c51_r1d;
  wire c51_a;
  wire c50_r;
  wire c50_a;
  wire c49_r;
  wire c49_a;
  wire [31:0] c48_r0d;
  wire [31:0] c48_r1d;
  wire c48_a;
  wire c47_r;
  wire c47_a;
  wire c46_r;
  wire c46_a;
  wire c45_r;
  wire c45_a;
  wire c44_r;
  wire c44_a;
  wire c43_r;
  wire c43_a;
  wire [32:0] c42_r0d;
  wire [32:0] c42_r1d;
  wire c42_a;
  wire c41_r;
  wire c41_a;
  wire [32:0] c40_r0d;
  wire [32:0] c40_r1d;
  wire c40_a;
  wire c39_r;
  wire c39_a;
  wire [33:0] c38_r0d;
  wire [33:0] c38_r1d;
  wire c38_a;
  wire [65:0] c37_r0d;
  wire [65:0] c37_r1d;
  wire c37_a;
  wire c36_r;
  wire c36_a;
  wire [32:0] c35_r0d;
  wire [32:0] c35_r1d;
  wire c35_a;
  wire c34_r;
  wire c34_a;
  wire [32:0] c33_r0d;
  wire [32:0] c33_r1d;
  wire c33_a;
  wire c32_r;
  wire c32_a;
  wire c31_r;
  wire c31_a;
  wire c30_r;
  wire c30_a;
  wire c29_r;
  wire c29_a;
  wire c28_r;
  wire c28_a;
  wire c27_r;
  wire c27_a;
  wire c26_r0d;
  wire c26_r1d;
  wire c26_a;
  wire c25_r;
  wire c25_a;
  wire [31:0] c24_r0d;
  wire [31:0] c24_r1d;
  wire c24_a;
  wire c23_r;
  wire c23_a;
  wire [31:0] c22_r0d;
  wire [31:0] c22_r1d;
  wire c22_a;
  wire c21_r;
  wire c21_a;
  wire c20_r;
  wire c20_a;
  wire c19_r;
  wire c19_a;
  wire [32:0] c18_r0d;
  wire [32:0] c18_r1d;
  wire c18_a;
  wire c17_r;
  wire c17_a;
  wire [31:0] c16_r0d;
  wire [31:0] c16_r1d;
  wire c16_a;
  wire c15_r;
  wire c15_a;
  wire c14_r0d;
  wire c14_r1d;
  wire c14_a;
  wire c13_r;
  wire c13_a;
  wire c12_r;
  wire c12_a;
  wire [32:0] c11_r0d;
  wire [32:0] c11_r1d;
  wire c11_a;
  wire c10_r;
  wire c10_a;
  wire [31:0] c9_r0d;
  wire [31:0] c9_r1d;
  wire c9_a;
  wire c8_r;
  wire c8_a;
  wire c7_r0d;
  wire c7_r1d;
  wire c7_a;
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I0 (c51_r0d, c51_r1d, c51_a, c53_r, c53_a, cN_0r0d, cN_0r1d, cN_0a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I1 (c48_r0d, c48_r1d, c48_a, c50_r, c50_a, s_0r0d, s_0r1d, s_0a, initialise);
  BrzJ_l11__281_200_29 I2 (c0_0r0d, c0_0r1d, c0_0a, c31_r, c31_a, c26_r0d, c26_r1d, c26_a, initialise);
  BrzJ_l12__2832_200_29 I3 (b_0r0d, b_0r1d, b_0a, c30_r, c30_a, c24_r0d, c24_r1d, c24_a, initialise);
  BrzJ_l12__2832_200_29 I4 (a_0r0d, a_0r1d, a_0a, c29_r, c29_a, c22_r0d, c22_r1d, c22_a, initialise);
  BrzJ_l12__2833_200_29 I5 (c62_r0d, c62_r1d, c62_a, c45_r, c45_a, c40_r0d, c40_r1d, c40_a, initialise);
  BrzF_33_l32__28_280_200_29_20_280_2033_29__m41m I6 (c11_r0d, c11_r1d, c11_a, c13_r, c13_a, c62_r0d, c62_r1d, c62_a, initialise);
  BrzJ_l12__2833_200_29 I7 (c61_r0d, c61_r1d, c61_a, c46_r, c46_a, c42_r0d, c42_r1d, c42_a, initialise);
  BrzF_33_l32__28_280_200_29_20_280_2033_29__m41m I8 (c18_r0d, c18_r1d, c18_a, c20_r, c20_a, c61_r0d, c61_r1d, c61_a, initialise);
  BrzJ_l12__2834_200_29 I9 (c60_r0d, c60_r1d, c60_a, c57_r, c57_a, c55_r0d, c55_r1d, c55_a, initialise);
  BrzF_34_l32__28_280_200_29_20_280_2034_29__m42m I10 (c38_r0d, c38_r1d, c38_a, c39_r, c39_a, c60_r0d, c60_r1d, c60_a, initialise);
  BrzM_0_2 I11 (go_0r, go_0a, c59_r, c59_a, c58_r, c58_a, initialise);
  BrzJ_l15__280_200_200_29 I12 (c21_r, c21_a, c39_r, c39_a, c54_r, c54_a, c59_r, c59_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I13 (c58_r, c58_a, c32_r, c32_a, c47_r, c47_a, c57_r, c57_a, initialise);
  BrzV_34_l6__28_29_l24__28_28_280_2034_29_2_m85m I14 (c55_r0d, c55_r1d, c55_a, c56_r, c56_a, c49_r, c49_a, c52_r, c52_a, c48_r0d, c48_r1d, c48_a, c51_r0d, c51_r1d, c51_a, initialise);
  BrzJ_l11__280_200_29 I15 (c50_r, c50_a, c53_r, c53_a, c54_r, c54_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I16 (c56_r, c56_a, c49_r, c49_a, c52_r, c52_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I17 (c47_r, c47_a, c45_r, c45_a, c46_r, c46_a, initialise);
  BrzJ_l11__280_200_29 I18 (c41_r, c41_a, c43_r, c43_a, c44_r, c44_a, initialise);
  BrzV_33_l6__28_29_l24__28_28_280_2033_29_2_m84m I19 (c42_r0d, c42_r1d, c42_a, c43_r, c43_a, c36_r, c36_a, c35_r0d, c35_r1d, c35_a, initialise);
  BrzV_33_l6__28_29_l24__28_28_280_2033_29_2_m84m I20 (c40_r0d, c40_r1d, c40_a, c41_r, c41_a, c34_r, c34_a, c33_r0d, c33_r1d, c33_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I21 (c44_r, c44_a, c34_r, c34_a, c36_r, c36_a, initialise);
  BrzO_66_34_l270__28_28app_201_20_280_200_2_m57m I22 (c37_r0d, c37_r1d, c37_a, c38_r0d, c38_r1d, c38_a);
  BrzJ_l13__2833_2033_29 I23 (c33_r0d, c33_r1d, c33_a, c35_r0d, c35_r1d, c35_a, c37_r0d, c37_r1d, c37_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I24 (c32_r, c32_a, c29_r, c29_a, c30_r, c30_a, c31_r, c31_a, initialise);
  BrzJ_l15__280_200_200_29 I25 (c23_r, c23_a, c25_r, c25_a, c27_r, c27_a, c28_r, c28_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m72m I26 (c26_r0d, c26_r1d, c26_a, c27_r, c27_a, c8_r, c8_a, c15_r, c15_a, c7_r0d, c7_r1d, c7_a, c14_r0d, c14_r1d, c14_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I27 (c24_r0d, c24_r1d, c24_a, c25_r, c25_a, c17_r, c17_a, c16_r0d, c16_r1d, c16_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I28 (c22_r0d, c22_r1d, c22_a, c23_r, c23_a, c10_r, c10_a, c9_r0d, c9_r1d, c9_a, initialise);
  BrzJ_l11__280_200_29 I29 (c13_r, c13_a, c20_r, c20_a, c21_r, c21_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I30 (c28_r, c28_a, c12_r, c12_a, c19_r, c19_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I31 (c19_r, c19_a, c15_r, c15_a, c17_r, c17_a, initialise);
  BrzJ_l12__281_2032_29 I32 (c14_r0d, c14_r1d, c14_a, c16_r0d, c16_r1d, c16_a, c18_r0d, c18_r1d, c18_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I33 (c12_r, c12_a, c8_r, c8_a, c10_r, c10_a, initialise);
  BrzJ_l12__281_2032_29 I34 (c7_r0d, c7_r1d, c7_a, c9_r0d, c9_r1d, c9_a, c11_r0d, c11_r1d, c11_a, initialise);
endmodule

module Balsa_nanoSpaMultiplier (
  go_0r, go_0a,
  bypass_0r0d, bypass_0r1d, bypass_0a,
  bypassH_0r0d, bypassH_0r1d, bypassH_0a,
  mType_0r0d, mType_0r1d, mType_0a,
  a_0r0d, a_0r1d, a_0a,
  b_0r0d, b_0r1d, b_0a,
  c_0r0d, c_0r1d, c_0a,
  mpH_0r0d, mpH_0r1d, mpH_0a,
  mpL_0r0d, mpL_0r1d, mpL_0a,
  mZ_0r0d, mZ_0r1d, mZ_0a,
  mN_0r0d, mN_0r1d, mN_0a,
  initialise
);
  input go_0r;
  output go_0a;
  input bypass_0r0d;
  input bypass_0r1d;
  output bypass_0a;
  input bypassH_0r0d;
  input bypassH_0r1d;
  output bypassH_0a;
  input [2:0] mType_0r0d;
  input [2:0] mType_0r1d;
  output mType_0a;
  input [31:0] a_0r0d;
  input [31:0] a_0r1d;
  output a_0a;
  input [31:0] b_0r0d;
  input [31:0] b_0r1d;
  output b_0a;
  input [31:0] c_0r0d;
  input [31:0] c_0r1d;
  output c_0a;
  output [31:0] mpH_0r0d;
  output [31:0] mpH_0r1d;
  input mpH_0a;
  output [31:0] mpL_0r0d;
  output [31:0] mpL_0r1d;
  input mpL_0a;
  output mZ_0r0d;
  output mZ_0r1d;
  input mZ_0a;
  output mN_0r0d;
  output mN_0r1d;
  input mN_0a;
  input initialise;
  wire [1:0] c883_r0d;
  wire [1:0] c883_r1d;
  wire c883_a;
  wire [1:0] c882_r0d;
  wire [1:0] c882_r1d;
  wire c882_a;
  wire [1:0] c881_r0d;
  wire [1:0] c881_r1d;
  wire c881_a;
  wire [1:0] c880_r0d;
  wire [1:0] c880_r1d;
  wire c880_a;
  wire c879_r;
  wire c879_a;
  wire c878_r0d;
  wire c878_r1d;
  wire c878_a;
  wire c877_r0d;
  wire c877_r1d;
  wire c877_a;
  wire c876_r;
  wire c876_a;
  wire c875_r0d;
  wire c875_r1d;
  wire c875_a;
  wire c874_r;
  wire c874_a;
  wire [1:0] c873_r0d;
  wire [1:0] c873_r1d;
  wire c873_a;
  wire [1:0] c872_r0d;
  wire [1:0] c872_r1d;
  wire c872_a;
  wire [1:0] c871_r0d;
  wire [1:0] c871_r1d;
  wire c871_a;
  wire [1:0] c870_r0d;
  wire [1:0] c870_r1d;
  wire c870_a;
  wire c869_r;
  wire c869_a;
  wire c868_r0d;
  wire c868_r1d;
  wire c868_a;
  wire c867_r0d;
  wire c867_r1d;
  wire c867_a;
  wire c866_r;
  wire c866_a;
  wire c865_r0d;
  wire c865_r1d;
  wire c865_a;
  wire c864_r;
  wire c864_a;
  wire [1:0] c863_r0d;
  wire [1:0] c863_r1d;
  wire c863_a;
  wire [1:0] c862_r0d;
  wire [1:0] c862_r1d;
  wire c862_a;
  wire [1:0] c861_r0d;
  wire [1:0] c861_r1d;
  wire c861_a;
  wire [1:0] c860_r0d;
  wire [1:0] c860_r1d;
  wire c860_a;
  wire c859_r;
  wire c859_a;
  wire [31:0] c858_r0d;
  wire [31:0] c858_r1d;
  wire c858_a;
  wire [31:0] c857_r0d;
  wire [31:0] c857_r1d;
  wire c857_a;
  wire c856_r;
  wire c856_a;
  wire [31:0] c855_r0d;
  wire [31:0] c855_r1d;
  wire c855_a;
  wire c854_r;
  wire c854_a;
  wire [1:0] c853_r0d;
  wire [1:0] c853_r1d;
  wire c853_a;
  wire [1:0] c852_r0d;
  wire [1:0] c852_r1d;
  wire c852_a;
  wire [1:0] c851_r0d;
  wire [1:0] c851_r1d;
  wire c851_a;
  wire [1:0] c850_r0d;
  wire [1:0] c850_r1d;
  wire c850_a;
  wire c849_r;
  wire c849_a;
  wire [31:0] c848_r0d;
  wire [31:0] c848_r1d;
  wire c848_a;
  wire [31:0] c847_r0d;
  wire [31:0] c847_r1d;
  wire c847_a;
  wire c846_r;
  wire c846_a;
  wire [31:0] c845_r0d;
  wire [31:0] c845_r1d;
  wire c845_a;
  wire c844_r;
  wire c844_a;
  wire [33:0] c843_r0d;
  wire [33:0] c843_r1d;
  wire c843_a;
  wire [1:0] c842_r0d;
  wire [1:0] c842_r1d;
  wire c842_a;
  wire [1:0] c841_r0d;
  wire [1:0] c841_r1d;
  wire c841_a;
  wire [1:0] c840_r0d;
  wire [1:0] c840_r1d;
  wire c840_a;
  wire [1:0] c839_r0d;
  wire [1:0] c839_r1d;
  wire c839_a;
  wire [1:0] c838_r0d;
  wire [1:0] c838_r1d;
  wire c838_a;
  wire [1:0] c837_r0d;
  wire [1:0] c837_r1d;
  wire c837_a;
  wire [1:0] c836_r0d;
  wire [1:0] c836_r1d;
  wire c836_a;
  wire [34:0] c835_r0d;
  wire [34:0] c835_r1d;
  wire c835_a;
  wire c834_r;
  wire c834_a;
  wire [34:0] c833_r0d;
  wire [34:0] c833_r1d;
  wire c833_a;
  wire [34:0] c832_r0d;
  wire [34:0] c832_r1d;
  wire c832_a;
  wire c831_r;
  wire c831_a;
  wire [34:0] c830_r0d;
  wire [34:0] c830_r1d;
  wire c830_a;
  wire c829_r;
  wire c829_a;
  wire [1:0] c828_r0d;
  wire [1:0] c828_r1d;
  wire c828_a;
  wire [1:0] c827_r0d;
  wire [1:0] c827_r1d;
  wire c827_a;
  wire [1:0] c826_r0d;
  wire [1:0] c826_r1d;
  wire c826_a;
  wire [1:0] c825_r0d;
  wire [1:0] c825_r1d;
  wire c825_a;
  wire [35:0] c824_r0d;
  wire [35:0] c824_r1d;
  wire c824_a;
  wire c823_r;
  wire c823_a;
  wire [35:0] c822_r0d;
  wire [35:0] c822_r1d;
  wire c822_a;
  wire [35:0] c821_r0d;
  wire [35:0] c821_r1d;
  wire c821_a;
  wire c820_r;
  wire c820_a;
  wire [35:0] c819_r0d;
  wire [35:0] c819_r1d;
  wire c819_a;
  wire c818_r;
  wire c818_a;
  wire [34:0] c817_r0d;
  wire [34:0] c817_r1d;
  wire c817_a;
  wire c816_r0d;
  wire c816_r1d;
  wire c816_a;
  wire c815_r0d;
  wire c815_r1d;
  wire c815_a;
  wire [31:0] c814_r0d;
  wire [31:0] c814_r1d;
  wire c814_a;
  wire [31:0] c813_r0d;
  wire [31:0] c813_r1d;
  wire c813_a;
  wire [1:0] c812_r0d;
  wire [1:0] c812_r1d;
  wire c812_a;
  wire [1:0] c811_r0d;
  wire [1:0] c811_r1d;
  wire c811_a;
  wire [1:0] c810_r0d;
  wire [1:0] c810_r1d;
  wire c810_a;
  wire [1:0] c809_r0d;
  wire [1:0] c809_r1d;
  wire c809_a;
  wire [31:0] c808_r0d;
  wire [31:0] c808_r1d;
  wire c808_a;
  wire c807_r;
  wire c807_a;
  wire [31:0] c806_r0d;
  wire [31:0] c806_r1d;
  wire c806_a;
  wire [31:0] c805_r0d;
  wire [31:0] c805_r1d;
  wire c805_a;
  wire c804_r;
  wire c804_a;
  wire [31:0] c803_r0d;
  wire [31:0] c803_r1d;
  wire c803_a;
  wire c802_r;
  wire c802_a;
  wire [2:0] c801_r0d;
  wire [2:0] c801_r1d;
  wire c801_a;
  wire [34:0] c800_r0d;
  wire [34:0] c800_r1d;
  wire c800_a;
  wire [8:0] c799_r0d;
  wire [8:0] c799_r1d;
  wire c799_a;
  wire [8:0] c798_r0d;
  wire [8:0] c798_r1d;
  wire c798_a;
  wire [8:0] c797_r0d;
  wire [8:0] c797_r1d;
  wire c797_a;
  wire [8:0] c796_r0d;
  wire [8:0] c796_r1d;
  wire c796_a;
  wire [8:0] c795_r0d;
  wire [8:0] c795_r1d;
  wire c795_a;
  wire [8:0] c794_r0d;
  wire [8:0] c794_r1d;
  wire c794_a;
  wire [8:0] c793_r0d;
  wire [8:0] c793_r1d;
  wire c793_a;
  wire [8:0] c792_r0d;
  wire [8:0] c792_r1d;
  wire c792_a;
  wire [8:0] c791_r0d;
  wire [8:0] c791_r1d;
  wire c791_a;
  wire [8:0] c790_r0d;
  wire [8:0] c790_r1d;
  wire c790_a;
  wire [8:0] c789_r0d;
  wire [8:0] c789_r1d;
  wire c789_a;
  wire [34:0] c788_r0d;
  wire [34:0] c788_r1d;
  wire c788_a;
  wire c787_r;
  wire c787_a;
  wire [34:0] c786_r0d;
  wire [34:0] c786_r1d;
  wire c786_a;
  wire [34:0] c785_r0d;
  wire [34:0] c785_r1d;
  wire c785_a;
  wire c784_r;
  wire c784_a;
  wire [34:0] c783_r0d;
  wire [34:0] c783_r1d;
  wire c783_a;
  wire c782_r;
  wire c782_a;
  wire [34:0] c781_r0d;
  wire [34:0] c781_r1d;
  wire c781_a;
  wire c780_r;
  wire c780_a;
  wire [34:0] c779_r0d;
  wire [34:0] c779_r1d;
  wire c779_a;
  wire c778_r;
  wire c778_a;
  wire [34:0] c777_r0d;
  wire [34:0] c777_r1d;
  wire c777_a;
  wire c776_r;
  wire c776_a;
  wire [34:0] c775_r0d;
  wire [34:0] c775_r1d;
  wire c775_a;
  wire c774_r;
  wire c774_a;
  wire [34:0] c773_r0d;
  wire [34:0] c773_r1d;
  wire c773_a;
  wire c772_r;
  wire c772_a;
  wire [34:0] c771_r0d;
  wire [34:0] c771_r1d;
  wire c771_a;
  wire c770_r;
  wire c770_a;
  wire [34:0] c769_r0d;
  wire [34:0] c769_r1d;
  wire c769_a;
  wire c768_r;
  wire c768_a;
  wire [34:0] c767_r0d;
  wire [34:0] c767_r1d;
  wire c767_a;
  wire [34:0] c766_r0d;
  wire [34:0] c766_r1d;
  wire c766_a;
  wire [34:0] c765_r0d;
  wire [34:0] c765_r1d;
  wire c765_a;
  wire [2:0] c764_r0d;
  wire [2:0] c764_r1d;
  wire c764_a;
  wire [2:0] c763_r0d;
  wire [2:0] c763_r1d;
  wire c763_a;
  wire [2:0] c762_r0d;
  wire [2:0] c762_r1d;
  wire c762_a;
  wire [2:0] c761_r0d;
  wire [2:0] c761_r1d;
  wire c761_a;
  wire [2:0] c760_r0d;
  wire [2:0] c760_r1d;
  wire c760_a;
  wire [31:0] c759_r0d;
  wire [31:0] c759_r1d;
  wire c759_a;
  wire c758_r;
  wire c758_a;
  wire [31:0] c757_r0d;
  wire [31:0] c757_r1d;
  wire c757_a;
  wire [31:0] c756_r0d;
  wire [31:0] c756_r1d;
  wire c756_a;
  wire c755_r;
  wire c755_a;
  wire [31:0] c754_r0d;
  wire [31:0] c754_r1d;
  wire c754_a;
  wire c753_r;
  wire c753_a;
  wire [31:0] c752_r0d;
  wire [31:0] c752_r1d;
  wire c752_a;
  wire c751_r;
  wire c751_a;
  wire [2:0] c750_r0d;
  wire [2:0] c750_r1d;
  wire c750_a;
  wire [2:0] c749_r0d;
  wire [2:0] c749_r1d;
  wire c749_a;
  wire [2:0] c748_r0d;
  wire [2:0] c748_r1d;
  wire c748_a;
  wire [2:0] c747_r0d;
  wire [2:0] c747_r1d;
  wire c747_a;
  wire [2:0] c746_r0d;
  wire [2:0] c746_r1d;
  wire c746_a;
  wire [31:0] c745_r0d;
  wire [31:0] c745_r1d;
  wire c745_a;
  wire c744_r;
  wire c744_a;
  wire [31:0] c743_r0d;
  wire [31:0] c743_r1d;
  wire c743_a;
  wire [31:0] c742_r0d;
  wire [31:0] c742_r1d;
  wire c742_a;
  wire c741_r;
  wire c741_a;
  wire [31:0] c740_r0d;
  wire [31:0] c740_r1d;
  wire c740_a;
  wire c739_r;
  wire c739_a;
  wire [31:0] c738_r0d;
  wire [31:0] c738_r1d;
  wire c738_a;
  wire c737_r;
  wire c737_a;
  wire [2:0] c736_r0d;
  wire [2:0] c736_r1d;
  wire c736_a;
  wire [2:0] c735_r0d;
  wire [2:0] c735_r1d;
  wire c735_a;
  wire [2:0] c734_r0d;
  wire [2:0] c734_r1d;
  wire c734_a;
  wire [2:0] c733_r0d;
  wire [2:0] c733_r1d;
  wire c733_a;
  wire [2:0] c732_r0d;
  wire [2:0] c732_r1d;
  wire c732_a;
  wire c731_r0d;
  wire c731_r1d;
  wire c731_a;
  wire c730_r;
  wire c730_a;
  wire c729_r0d;
  wire c729_r1d;
  wire c729_a;
  wire c728_r0d;
  wire c728_r1d;
  wire c728_a;
  wire c727_r;
  wire c727_a;
  wire c726_r0d;
  wire c726_r1d;
  wire c726_a;
  wire c725_r;
  wire c725_a;
  wire c724_r0d;
  wire c724_r1d;
  wire c724_a;
  wire c723_r;
  wire c723_a;
  wire [34:0] c722_r0d;
  wire [34:0] c722_r1d;
  wire c722_a;
  wire [2:0] c721_r0d;
  wire [2:0] c721_r1d;
  wire c721_a;
  wire [2:0] c720_r0d;
  wire [2:0] c720_r1d;
  wire c720_a;
  wire [2:0] c719_r0d;
  wire [2:0] c719_r1d;
  wire c719_a;
  wire [2:0] c718_r0d;
  wire [2:0] c718_r1d;
  wire c718_a;
  wire [31:0] c717_r0d;
  wire [31:0] c717_r1d;
  wire c717_a;
  wire [3:0] c716_r0d;
  wire [3:0] c716_r1d;
  wire c716_a;
  wire [2:0] c715_r0d;
  wire [2:0] c715_r1d;
  wire c715_a;
  wire [2:0] c714_r0d;
  wire [2:0] c714_r1d;
  wire c714_a;
  wire [2:0] c713_r0d;
  wire [2:0] c713_r1d;
  wire c713_a;
  wire [2:0] c712_r0d;
  wire [2:0] c712_r1d;
  wire c712_a;
  wire c711_r0d;
  wire c711_r1d;
  wire c711_a;
  wire [1:0] c710_r0d;
  wire [1:0] c710_r1d;
  wire c710_a;
  wire [1:0] c709_r0d;
  wire [1:0] c709_r1d;
  wire c709_a;
  wire [1:0] c708_r0d;
  wire [1:0] c708_r1d;
  wire c708_a;
  wire [1:0] c707_r0d;
  wire [1:0] c707_r1d;
  wire c707_a;
  wire c706_r0d;
  wire c706_r1d;
  wire c706_a;
  wire c705_r;
  wire c705_a;
  wire c704_r0d;
  wire c704_r1d;
  wire c704_a;
  wire c703_r0d;
  wire c703_r1d;
  wire c703_a;
  wire c702_r;
  wire c702_a;
  wire c701_r0d;
  wire c701_r1d;
  wire c701_a;
  wire c700_r;
  wire c700_a;
  wire [1:0] c699_r0d;
  wire [1:0] c699_r1d;
  wire c699_a;
  wire [1:0] c698_r0d;
  wire [1:0] c698_r1d;
  wire c698_a;
  wire [1:0] c697_r0d;
  wire [1:0] c697_r1d;
  wire c697_a;
  wire [1:0] c696_r0d;
  wire [1:0] c696_r1d;
  wire c696_a;
  wire c695_r0d;
  wire c695_r1d;
  wire c695_a;
  wire c694_r;
  wire c694_a;
  wire c693_r0d;
  wire c693_r1d;
  wire c693_a;
  wire c692_r0d;
  wire c692_r1d;
  wire c692_a;
  wire c691_r;
  wire c691_a;
  wire c690_r0d;
  wire c690_r1d;
  wire c690_a;
  wire c689_r;
  wire c689_a;
  wire [31:0] c688_r0d;
  wire [31:0] c688_r1d;
  wire c688_a;
  wire [1:0] c687_r0d;
  wire [1:0] c687_r1d;
  wire c687_a;
  wire [1:0] c686_r0d;
  wire [1:0] c686_r1d;
  wire c686_a;
  wire [1:0] c685_r0d;
  wire [1:0] c685_r1d;
  wire c685_a;
  wire [1:0] c684_r0d;
  wire [1:0] c684_r1d;
  wire c684_a;
  wire [31:0] c683_r0d;
  wire [31:0] c683_r1d;
  wire c683_a;
  wire c682_r;
  wire c682_a;
  wire [31:0] c681_r0d;
  wire [31:0] c681_r1d;
  wire c681_a;
  wire [31:0] c680_r0d;
  wire [31:0] c680_r1d;
  wire c680_a;
  wire c679_r;
  wire c679_a;
  wire [31:0] c678_r0d;
  wire [31:0] c678_r1d;
  wire c678_a;
  wire c677_r;
  wire c677_a;
  wire [2:0] c676_r0d;
  wire [2:0] c676_r1d;
  wire c676_a;
  wire [2:0] c675_r0d;
  wire [2:0] c675_r1d;
  wire c675_a;
  wire [2:0] c674_r0d;
  wire [2:0] c674_r1d;
  wire c674_a;
  wire [2:0] c673_r0d;
  wire [2:0] c673_r1d;
  wire c673_a;
  wire [2:0] c672_r0d;
  wire [2:0] c672_r1d;
  wire c672_a;
  wire c671_r0d;
  wire c671_r1d;
  wire c671_a;
  wire c670_r;
  wire c670_a;
  wire c669_r0d;
  wire c669_r1d;
  wire c669_a;
  wire c668_r0d;
  wire c668_r1d;
  wire c668_a;
  wire c667_r;
  wire c667_a;
  wire c666_r0d;
  wire c666_r1d;
  wire c666_a;
  wire c665_r;
  wire c665_a;
  wire c664_r0d;
  wire c664_r1d;
  wire c664_a;
  wire c663_r;
  wire c663_a;
  wire [1:0] c662_r0d;
  wire [1:0] c662_r1d;
  wire c662_a;
  wire [1:0] c661_r0d;
  wire [1:0] c661_r1d;
  wire c661_a;
  wire [1:0] c660_r0d;
  wire [1:0] c660_r1d;
  wire c660_a;
  wire [1:0] c659_r0d;
  wire [1:0] c659_r1d;
  wire c659_a;
  wire c658_r0d;
  wire c658_r1d;
  wire c658_a;
  wire c657_r;
  wire c657_a;
  wire c656_r0d;
  wire c656_r1d;
  wire c656_a;
  wire c655_r0d;
  wire c655_r1d;
  wire c655_a;
  wire c654_r;
  wire c654_a;
  wire c653_r0d;
  wire c653_r1d;
  wire c653_a;
  wire c652_r;
  wire c652_a;
  wire c651_r0d;
  wire c651_r1d;
  wire c651_a;
  wire c650_r0d;
  wire c650_r1d;
  wire c650_a;
  wire c649_r;
  wire c649_a;
  wire c648_r;
  wire c648_a;
  wire c647_r;
  wire c647_a;
  wire c646_r;
  wire c646_a;
  wire c645_r;
  wire c645_a;
  wire c644_r;
  wire c644_a;
  wire c643_r0d;
  wire c643_r1d;
  wire c643_a;
  wire c642_r;
  wire c642_a;
  wire c641_r0d;
  wire c641_r1d;
  wire c641_a;
  wire c640_r;
  wire c640_a;
  wire c639_r;
  wire c639_a;
  wire c638_r;
  wire c638_a;
  wire c637_r;
  wire c637_a;
  wire c636_r;
  wire c636_a;
  wire [31:0] c635_r0d;
  wire [31:0] c635_r1d;
  wire c635_a;
  wire c634_r;
  wire c634_a;
  wire c633_r;
  wire c633_a;
  wire c632_r;
  wire c632_a;
  wire c631_r0d;
  wire c631_r1d;
  wire c631_a;
  wire c630_r;
  wire c630_a;
  wire c629_r0d;
  wire c629_r1d;
  wire c629_a;
  wire c628_r;
  wire c628_a;
  wire c627_r;
  wire c627_a;
  wire c626_r0d;
  wire c626_r1d;
  wire c626_a;
  wire c625_r;
  wire c625_a;
  wire c624_r;
  wire c624_a;
  wire [31:0] c623_r0d;
  wire [31:0] c623_r1d;
  wire c623_a;
  wire c622_r;
  wire c622_a;
  wire c621_r;
  wire c621_a;
  wire c620_r;
  wire c620_a;
  wire c619_r;
  wire c619_a;
  wire c618_r;
  wire c618_a;
  wire c617_r;
  wire c617_a;
  wire [31:0] c616_r0d;
  wire [31:0] c616_r1d;
  wire c616_a;
  wire c615_r;
  wire c615_a;
  wire [31:0] c614_r0d;
  wire [31:0] c614_r1d;
  wire c614_a;
  wire c613_r;
  wire c613_a;
  wire c612_r;
  wire c612_a;
  wire c611_r0d;
  wire c611_r1d;
  wire c611_a;
  wire c610_r;
  wire c610_a;
  wire c609_r;
  wire c609_a;
  wire c608_r0d;
  wire c608_r1d;
  wire c608_a;
  wire c607_r;
  wire c607_a;
  wire c606_r0d;
  wire c606_r1d;
  wire c606_a;
  wire c605_r;
  wire c605_a;
  wire c604_r;
  wire c604_a;
  wire c603_r0d;
  wire c603_r1d;
  wire c603_a;
  wire c602_r;
  wire c602_a;
  wire c601_r0d;
  wire c601_r1d;
  wire c601_a;
  wire c600_r;
  wire c600_a;
  wire c599_r;
  wire c599_a;
  wire [31:0] c598_r0d;
  wire [31:0] c598_r1d;
  wire c598_a;
  wire c597_r;
  wire c597_a;
  wire [31:0] c596_r0d;
  wire [31:0] c596_r1d;
  wire c596_a;
  wire c595_r0d;
  wire c595_r1d;
  wire c595_a;
  wire c594_r;
  wire c594_a;
  wire c593_r;
  wire c593_a;
  wire c592_r;
  wire c592_a;
  wire c591_r;
  wire c591_a;
  wire c590_r;
  wire c590_a;
  wire c589_r;
  wire c589_a;
  wire c588_r;
  wire c588_a;
  wire [2:0] c587_r0d;
  wire [2:0] c587_r1d;
  wire c587_a;
  wire c586_r;
  wire c586_a;
  wire c585_r0d;
  wire c585_r1d;
  wire c585_a;
  wire c584_r;
  wire c584_a;
  wire c583_r0d;
  wire c583_r1d;
  wire c583_a;
  wire c582_r;
  wire c582_a;
  wire c581_r;
  wire c581_a;
  wire c580_r;
  wire c580_a;
  wire c579_r0d;
  wire c579_r1d;
  wire c579_a;
  wire c578_r;
  wire c578_a;
  wire c577_r;
  wire c577_a;
  wire c576_r0d;
  wire c576_r1d;
  wire c576_a;
  wire c575_r;
  wire c575_a;
  wire c574_r;
  wire c574_a;
  wire c573_r;
  wire c573_a;
  wire c572_r;
  wire c572_a;
  wire c571_r;
  wire c571_a;
  wire [31:0] c570_r0d;
  wire [31:0] c570_r1d;
  wire c570_a;
  wire c569_r;
  wire c569_a;
  wire [31:0] c568_r0d;
  wire [31:0] c568_r1d;
  wire c568_a;
  wire c567_r;
  wire c567_a;
  wire c566_r;
  wire c566_a;
  wire c565_r;
  wire c565_a;
  wire c564_r;
  wire c564_a;
  wire [31:0] c563_r0d;
  wire [31:0] c563_r1d;
  wire c563_a;
  wire c562_r;
  wire c562_a;
  wire c561_r;
  wire c561_a;
  wire [2:0] c560_r0d;
  wire [2:0] c560_r1d;
  wire c560_a;
  wire c559_r;
  wire c559_a;
  wire c558_r;
  wire c558_a;
  wire c557_r;
  wire c557_a;
  wire c556_r;
  wire c556_a;
  wire c555_r;
  wire c555_a;
  wire [31:0] c554_r0d;
  wire [31:0] c554_r1d;
  wire c554_a;
  wire c553_r;
  wire c553_a;
  wire [31:0] c552_r0d;
  wire [31:0] c552_r1d;
  wire c552_a;
  wire c551_r;
  wire c551_a;
  wire [31:0] c550_r0d;
  wire [31:0] c550_r1d;
  wire c550_a;
  wire c549_r;
  wire c549_a;
  wire c548_r;
  wire c548_a;
  wire [2:0] c547_r0d;
  wire [2:0] c547_r1d;
  wire c547_a;
  wire c546_r;
  wire c546_a;
  wire c545_r;
  wire c545_a;
  wire [2:0] c544_r0d;
  wire [2:0] c544_r1d;
  wire c544_a;
  wire c543_r;
  wire c543_a;
  wire c542_r;
  wire c542_a;
  wire [31:0] c541_r0d;
  wire [31:0] c541_r1d;
  wire c541_a;
  wire c540_r;
  wire c540_a;
  wire c539_r;
  wire c539_a;
  wire [31:0] c538_r0d;
  wire [31:0] c538_r1d;
  wire c538_a;
  wire c537_r0d;
  wire c537_r1d;
  wire c537_a;
  wire c536_r;
  wire c536_a;
  wire c535_r;
  wire c535_a;
  wire c534_r;
  wire c534_a;
  wire c533_r;
  wire c533_a;
  wire c532_r;
  wire c532_a;
  wire c531_r;
  wire c531_a;
  wire c530_r;
  wire c530_a;
  wire c529_r;
  wire c529_a;
  wire [31:0] c528_r0d;
  wire [31:0] c528_r1d;
  wire c528_a;
  wire c527_r;
  wire c527_a;
  wire [31:0] c526_r0d;
  wire [31:0] c526_r1d;
  wire c526_a;
  wire c525_r;
  wire c525_a;
  wire [31:0] c524_r0d;
  wire [31:0] c524_r1d;
  wire c524_a;
  wire c523_r;
  wire c523_a;
  wire [2:0] c522_r0d;
  wire [2:0] c522_r1d;
  wire c522_a;
  wire c521_r;
  wire c521_a;
  wire c520_r;
  wire c520_a;
  wire c519_r;
  wire c519_a;
  wire c518_r0d;
  wire c518_r1d;
  wire c518_a;
  wire c517_r;
  wire c517_a;
  wire c516_r;
  wire c516_a;
  wire c515_r0d;
  wire c515_r1d;
  wire c515_a;
  wire c514_r;
  wire c514_a;
  wire c513_r;
  wire c513_a;
  wire [31:0] c512_r0d;
  wire [31:0] c512_r1d;
  wire c512_a;
  wire [34:0] c511_r0d;
  wire [34:0] c511_r1d;
  wire c511_a;
  wire c510_r;
  wire c510_a;
  wire c509_r;
  wire c509_a;
  wire c508_r;
  wire c508_a;
  wire c507_r;
  wire c507_a;
  wire c506_r;
  wire c506_a;
  wire [32:0] c505_r0d;
  wire [32:0] c505_r1d;
  wire c505_a;
  wire c504_r;
  wire c504_a;
  wire [31:0] c503_r0d;
  wire [31:0] c503_r1d;
  wire c503_a;
  wire c502_r0d;
  wire c502_r1d;
  wire c502_a;
  wire c501_r;
  wire c501_a;
  wire [35:0] c500_r0d;
  wire [35:0] c500_r1d;
  wire c500_a;
  wire c499_r;
  wire c499_a;
  wire c498_r;
  wire c498_a;
  wire [31:0] c497_r0d;
  wire [31:0] c497_r1d;
  wire c497_a;
  wire [34:0] c496_r0d;
  wire [34:0] c496_r1d;
  wire c496_a;
  wire c495_r;
  wire c495_a;
  wire c494_r;
  wire c494_a;
  wire c493_r;
  wire c493_a;
  wire c492_r;
  wire c492_a;
  wire [32:0] c491_r0d;
  wire [32:0] c491_r1d;
  wire c491_a;
  wire c490_r;
  wire c490_a;
  wire [31:0] c489_r0d;
  wire [31:0] c489_r1d;
  wire c489_a;
  wire c488_r0d;
  wire c488_r1d;
  wire c488_a;
  wire c487_r;
  wire c487_a;
  wire [35:0] c486_r0d;
  wire [35:0] c486_r1d;
  wire c486_a;
  wire c485_r;
  wire c485_a;
  wire c484_r;
  wire c484_a;
  wire [31:0] c483_r0d;
  wire [31:0] c483_r1d;
  wire c483_a;
  wire [34:0] c482_r0d;
  wire [34:0] c482_r1d;
  wire c482_a;
  wire c481_r;
  wire c481_a;
  wire [2:0] c480_r0d;
  wire [2:0] c480_r1d;
  wire c480_a;
  wire c479_r;
  wire c479_a;
  wire c478_r;
  wire c478_a;
  wire c477_r;
  wire c477_a;
  wire c476_r;
  wire c476_a;
  wire c475_r;
  wire c475_a;
  wire c474_r0d;
  wire c474_r1d;
  wire c474_a;
  wire c473_r;
  wire c473_a;
  wire c472_r;
  wire c472_a;
  wire [9:0] c471_r0d;
  wire [9:0] c471_r1d;
  wire c471_a;
  wire c470_r;
  wire c470_a;
  wire c469_r;
  wire c469_a;
  wire [9:0] c468_r0d;
  wire [9:0] c468_r1d;
  wire c468_a;
  wire c467_r;
  wire c467_a;
  wire c466_r;
  wire c466_a;
  wire c465_r;
  wire c465_a;
  wire [8:0] c464_r0d;
  wire [8:0] c464_r1d;
  wire c464_a;
  wire [9:0] c463_r0d;
  wire [9:0] c463_r1d;
  wire c463_a;
  wire c462_r;
  wire c462_a;
  wire c461_r;
  wire c461_a;
  wire c460_r0d;
  wire c460_r1d;
  wire c460_a;
  wire c459_r;
  wire c459_a;
  wire c458_r0d;
  wire c458_r1d;
  wire c458_a;
  wire c457_r;
  wire c457_a;
  wire c456_r0d;
  wire c456_r1d;
  wire c456_a;
  wire c455_r;
  wire c455_a;
  wire c454_r0d;
  wire c454_r1d;
  wire c454_a;
  wire c453_r;
  wire c453_a;
  wire [34:0] c452_r0d;
  wire [34:0] c452_r1d;
  wire c452_a;
  wire [34:0] c451_r0d;
  wire [34:0] c451_r1d;
  wire c451_a;
  wire c450_r0d;
  wire c450_r1d;
  wire c450_a;
  wire c449_r;
  wire c449_a;
  wire c448_r;
  wire c448_a;
  wire c447_r;
  wire c447_a;
  wire c446_r;
  wire c446_a;
  wire c445_r;
  wire c445_a;
  wire c444_r0d;
  wire c444_r1d;
  wire c444_a;
  wire c443_r;
  wire c443_a;
  wire c442_r;
  wire c442_a;
  wire c441_r;
  wire c441_a;
  wire c440_r0d;
  wire c440_r1d;
  wire c440_a;
  wire c439_r;
  wire c439_a;
  wire c438_r;
  wire c438_a;
  wire c437_r0d;
  wire c437_r1d;
  wire c437_a;
  wire [1:0] c436_r0d;
  wire [1:0] c436_r1d;
  wire c436_a;
  wire c435_r;
  wire c435_a;
  wire c434_r0d;
  wire c434_r1d;
  wire c434_a;
  wire c433_r0d;
  wire c433_r1d;
  wire c433_a;
  wire [32:0] c432_r0d;
  wire [32:0] c432_r1d;
  wire c432_a;
  wire c431_r0d;
  wire c431_r1d;
  wire c431_a;
  wire c430_r;
  wire c430_a;
  wire c429_r;
  wire c429_a;
  wire [31:0] c428_r0d;
  wire [31:0] c428_r1d;
  wire c428_a;
  wire c427_r;
  wire c427_a;
  wire c426_r0d;
  wire c426_r1d;
  wire c426_a;
  wire c425_r;
  wire c425_a;
  wire c424_r;
  wire c424_a;
  wire [31:0] c423_r0d;
  wire [31:0] c423_r1d;
  wire c423_a;
  wire c422_r;
  wire c422_a;
  wire c421_r;
  wire c421_a;
  wire [31:0] c420_r0d;
  wire [31:0] c420_r1d;
  wire c420_a;
  wire c419_r;
  wire c419_a;
  wire c418_r;
  wire c418_a;
  wire c417_r;
  wire c417_a;
  wire c416_r;
  wire c416_a;
  wire c415_r;
  wire c415_a;
  wire c414_r;
  wire c414_a;
  wire c413_r0d;
  wire c413_r1d;
  wire c413_a;
  wire c412_r;
  wire c412_a;
  wire [31:0] c411_r0d;
  wire [31:0] c411_r1d;
  wire c411_a;
  wire c410_r;
  wire c410_a;
  wire [31:0] c409_r0d;
  wire [31:0] c409_r1d;
  wire c409_a;
  wire c408_r;
  wire c408_a;
  wire c407_r;
  wire c407_a;
  wire c406_r0d;
  wire c406_r1d;
  wire c406_a;
  wire c405_r;
  wire c405_a;
  wire c404_r;
  wire c404_a;
  wire [31:0] c403_r0d;
  wire [31:0] c403_r1d;
  wire c403_a;
  wire c402_r;
  wire c402_a;
  wire c401_r;
  wire c401_a;
  wire [31:0] c400_r0d;
  wire [31:0] c400_r1d;
  wire c400_a;
  wire c399_r;
  wire c399_a;
  wire [30:0] c398_r0d;
  wire [30:0] c398_r1d;
  wire c398_a;
  wire c397_r;
  wire c397_a;
  wire c396_r0d;
  wire c396_r1d;
  wire c396_a;
  wire c395_r;
  wire c395_a;
  wire c394_r;
  wire c394_a;
  wire c393_r;
  wire c393_a;
  wire c392_r;
  wire c392_a;
  wire c391_r;
  wire c391_a;
  wire c390_r0d;
  wire c390_r1d;
  wire c390_a;
  wire c389_r;
  wire c389_a;
  wire c388_r;
  wire c388_a;
  wire c387_r0d;
  wire c387_r1d;
  wire c387_a;
  wire c386_r;
  wire c386_a;
  wire c385_r;
  wire c385_a;
  wire [31:0] c384_r0d;
  wire [31:0] c384_r1d;
  wire c384_a;
  wire c383_r0d;
  wire c383_r1d;
  wire c383_a;
  wire c382_r;
  wire c382_a;
  wire c381_r;
  wire c381_a;
  wire c380_r;
  wire c380_a;
  wire c379_r;
  wire c379_a;
  wire c378_r;
  wire c378_a;
  wire c377_r;
  wire c377_a;
  wire c376_r0d;
  wire c376_r1d;
  wire c376_a;
  wire c375_r;
  wire c375_a;
  wire [31:0] c374_r0d;
  wire [31:0] c374_r1d;
  wire c374_a;
  wire c373_r;
  wire c373_a;
  wire c372_r;
  wire c372_a;
  wire c371_r;
  wire c371_a;
  wire c370_r0d;
  wire c370_r1d;
  wire c370_a;
  wire [32:0] c369_r0d;
  wire [32:0] c369_r1d;
  wire c369_a;
  wire c368_r0d;
  wire c368_r1d;
  wire c368_a;
  wire c367_r;
  wire c367_a;
  wire c366_r;
  wire c366_a;
  wire [31:0] c365_r0d;
  wire [31:0] c365_r1d;
  wire c365_a;
  wire c364_r;
  wire c364_a;
  wire c363_r;
  wire c363_a;
  wire c362_r0d;
  wire c362_r1d;
  wire c362_a;
  wire c361_r;
  wire c361_a;
  wire c360_r;
  wire c360_a;
  wire c359_r0d;
  wire c359_r1d;
  wire c359_a;
  wire c358_r;
  wire c358_a;
  wire c357_r;
  wire c357_a;
  wire [31:0] c356_r0d;
  wire [31:0] c356_r1d;
  wire c356_a;
  wire c355_r;
  wire c355_a;
  wire c354_r0d;
  wire c354_r1d;
  wire c354_a;
  wire c353_r;
  wire c353_a;
  wire c352_r;
  wire c352_a;
  wire c351_r;
  wire c351_a;
  wire [31:0] c350_r0d;
  wire [31:0] c350_r1d;
  wire c350_a;
  wire c349_r;
  wire c349_a;
  wire c348_r;
  wire c348_a;
  wire [31:0] c347_r0d;
  wire [31:0] c347_r1d;
  wire c347_a;
  wire c346_r;
  wire c346_a;
  wire c345_r;
  wire c345_a;
  wire c344_r;
  wire c344_a;
  wire c343_r;
  wire c343_a;
  wire c342_r0d;
  wire c342_r1d;
  wire c342_a;
  wire c341_r;
  wire c341_a;
  wire c340_r;
  wire c340_a;
  wire c339_r;
  wire c339_a;
  wire [3:0] c338_r0d;
  wire [3:0] c338_r1d;
  wire c338_a;
  wire c337_r;
  wire c337_a;
  wire c336_r;
  wire c336_a;
  wire [35:0] c335_r0d;
  wire [35:0] c335_r1d;
  wire c335_a;
  wire c334_r;
  wire c334_a;
  wire c333_r;
  wire c333_a;
  wire [34:0] c332_r0d;
  wire [34:0] c332_r1d;
  wire c332_a;
  wire c331_r;
  wire c331_a;
  wire c330_r;
  wire c330_a;
  wire [35:0] c329_r0d;
  wire [35:0] c329_r1d;
  wire c329_a;
  wire c328_r;
  wire c328_a;
  wire c327_r;
  wire c327_a;
  wire [34:0] c326_r0d;
  wire [34:0] c326_r1d;
  wire c326_a;
  wire c325_r;
  wire c325_a;
  wire c324_r0d;
  wire c324_r1d;
  wire c324_a;
  wire [33:0] c323_r0d;
  wire [33:0] c323_r1d;
  wire c323_a;
  wire c322_r;
  wire c322_a;
  wire c321_r0d;
  wire c321_r1d;
  wire c321_a;
  wire c320_r;
  wire c320_a;
  wire [32:0] c319_r0d;
  wire [32:0] c319_r1d;
  wire c319_a;
  wire c318_r;
  wire c318_a;
  wire c317_r;
  wire c317_a;
  wire c316_r;
  wire c316_a;
  wire c315_r;
  wire c315_a;
  wire c314_r0d;
  wire c314_r1d;
  wire c314_a;
  wire c313_r;
  wire c313_a;
  wire c312_r0d;
  wire c312_r1d;
  wire c312_a;
  wire c311_r;
  wire c311_a;
  wire c310_r;
  wire c310_a;
  wire c309_r;
  wire c309_a;
  wire c308_r;
  wire c308_a;
  wire c307_r;
  wire c307_a;
  wire c306_r;
  wire c306_a;
  wire c305_r0d;
  wire c305_r1d;
  wire c305_a;
  wire c304_r;
  wire c304_a;
  wire [34:0] c303_r0d;
  wire [34:0] c303_r1d;
  wire c303_a;
  wire c302_r;
  wire c302_a;
  wire [34:0] c301_r0d;
  wire [34:0] c301_r1d;
  wire c301_a;
  wire c300_r;
  wire c300_a;
  wire c299_r;
  wire c299_a;
  wire c298_r;
  wire c298_a;
  wire [34:0] c297_r0d;
  wire [34:0] c297_r1d;
  wire c297_a;
  wire c296_r;
  wire c296_a;
  wire [2:0] c295_r0d;
  wire [2:0] c295_r1d;
  wire c295_a;
  wire c294_r;
  wire c294_a;
  wire [31:0] c293_r0d;
  wire [31:0] c293_r1d;
  wire c293_a;
  wire [35:0] c292_r0d;
  wire [35:0] c292_r1d;
  wire c292_a;
  wire c291_r;
  wire c291_a;
  wire c290_r;
  wire c290_a;
  wire [31:0] c289_r0d;
  wire [31:0] c289_r1d;
  wire c289_a;
  wire [34:0] c288_r0d;
  wire [34:0] c288_r1d;
  wire c288_a;
  wire c287_r;
  wire c287_a;
  wire c286_r;
  wire c286_a;
  wire [34:0] c285_r0d;
  wire [34:0] c285_r1d;
  wire c285_a;
  wire c284_r;
  wire c284_a;
  wire [1:0] c283_r0d;
  wire [1:0] c283_r1d;
  wire c283_a;
  wire [32:0] c282_r0d;
  wire [32:0] c282_r1d;
  wire c282_a;
  wire c281_r;
  wire c281_a;
  wire c280_r0d;
  wire c280_r1d;
  wire c280_a;
  wire c279_r;
  wire c279_a;
  wire [31:0] c278_r0d;
  wire [31:0] c278_r1d;
  wire c278_a;
  wire [35:0] c277_r0d;
  wire [35:0] c277_r1d;
  wire c277_a;
  wire c276_r;
  wire c276_a;
  wire c275_r;
  wire c275_a;
  wire [34:0] c274_r0d;
  wire [34:0] c274_r1d;
  wire c274_a;
  wire c273_r;
  wire c273_a;
  wire c272_r;
  wire c272_a;
  wire c271_r;
  wire c271_a;
  wire [34:0] c270_r0d;
  wire [34:0] c270_r1d;
  wire c270_a;
  wire c269_r;
  wire c269_a;
  wire c268_r;
  wire c268_a;
  wire [34:0] c267_r0d;
  wire [34:0] c267_r1d;
  wire c267_a;
  wire c266_r;
  wire c266_a;
  wire c265_r;
  wire c265_a;
  wire [34:0] c264_r0d;
  wire [34:0] c264_r1d;
  wire c264_a;
  wire c263_r;
  wire c263_a;
  wire c262_r;
  wire c262_a;
  wire [34:0] c261_r0d;
  wire [34:0] c261_r1d;
  wire c261_a;
  wire c260_r;
  wire c260_a;
  wire c259_r;
  wire c259_a;
  wire [34:0] c258_r0d;
  wire [34:0] c258_r1d;
  wire c258_a;
  wire c257_r;
  wire c257_a;
  wire c256_r;
  wire c256_a;
  wire [34:0] c255_r0d;
  wire [34:0] c255_r1d;
  wire c255_a;
  wire c254_r;
  wire c254_a;
  wire c253_r;
  wire c253_a;
  wire [34:0] c252_r0d;
  wire [34:0] c252_r1d;
  wire c252_a;
  wire c251_r;
  wire c251_a;
  wire c250_r;
  wire c250_a;
  wire [34:0] c249_r0d;
  wire [34:0] c249_r1d;
  wire c249_a;
  wire c248_r;
  wire c248_a;
  wire c247_r;
  wire c247_a;
  wire [3:0] c246_r0d;
  wire [3:0] c246_r1d;
  wire c246_a;
  wire [34:0] c245_r0d;
  wire [34:0] c245_r1d;
  wire c245_a;
  wire c244_r;
  wire c244_a;
  wire [3:0] c243_r0d;
  wire [3:0] c243_r1d;
  wire c243_a;
  wire c242_r;
  wire c242_a;
  wire c241_r;
  wire c241_a;
  wire c240_r0d;
  wire c240_r1d;
  wire c240_a;
  wire c239_r;
  wire c239_a;
  wire c238_r;
  wire c238_a;
  wire [34:0] c237_r0d;
  wire [34:0] c237_r1d;
  wire c237_a;
  wire c236_r;
  wire c236_a;
  wire [34:0] c235_r0d;
  wire [34:0] c235_r1d;
  wire c235_a;
  wire c234_r;
  wire c234_a;
  wire c233_r;
  wire c233_a;
  wire [34:0] c232_r0d;
  wire [34:0] c232_r1d;
  wire c232_a;
  wire c231_r;
  wire c231_a;
  wire [34:0] c230_r0d;
  wire [34:0] c230_r1d;
  wire c230_a;
  wire c229_r;
  wire c229_a;
  wire c228_r;
  wire c228_a;
  wire [34:0] c227_r0d;
  wire [34:0] c227_r1d;
  wire c227_a;
  wire c226_r;
  wire c226_a;
  wire c225_r;
  wire c225_a;
  wire [34:0] c224_r0d;
  wire [34:0] c224_r1d;
  wire c224_a;
  wire c223_r0d;
  wire c223_r1d;
  wire c223_a;
  wire c222_r;
  wire c222_a;
  wire c221_r;
  wire c221_a;
  wire c220_r0d;
  wire c220_r1d;
  wire c220_a;
  wire c219_r;
  wire c219_a;
  wire c218_r;
  wire c218_a;
  wire c217_r;
  wire c217_a;
  wire [34:0] c216_r0d;
  wire [34:0] c216_r1d;
  wire c216_a;
  wire [34:0] c215_r0d;
  wire [34:0] c215_r1d;
  wire c215_a;
  wire c214_r;
  wire c214_a;
  wire c213_r;
  wire c213_a;
  wire [34:0] c212_r0d;
  wire [34:0] c212_r1d;
  wire c212_a;
  wire [34:0] c211_r0d;
  wire [34:0] c211_r1d;
  wire c211_a;
  wire c210_r;
  wire c210_a;
  wire c209_r;
  wire c209_a;
  wire [34:0] c208_r0d;
  wire [34:0] c208_r1d;
  wire c208_a;
  wire [34:0] c207_r0d;
  wire [34:0] c207_r1d;
  wire c207_a;
  wire c206_r;
  wire c206_a;
  wire c205_r;
  wire c205_a;
  wire [34:0] c204_r0d;
  wire [34:0] c204_r1d;
  wire c204_a;
  wire [34:0] c203_r0d;
  wire [34:0] c203_r1d;
  wire c203_a;
  wire c202_r;
  wire c202_a;
  wire c201_r;
  wire c201_a;
  wire c200_r;
  wire c200_a;
  wire c199_r;
  wire c199_a;
  wire c198_r;
  wire c198_a;
  wire c197_r;
  wire c197_a;
  wire c196_r;
  wire c196_a;
  wire c195_r0d;
  wire c195_r1d;
  wire c195_a;
  wire c194_r;
  wire c194_a;
  wire c193_r0d;
  wire c193_r1d;
  wire c193_a;
  wire c192_r;
  wire c192_a;
  wire [34:0] c191_r0d;
  wire [34:0] c191_r1d;
  wire c191_a;
  wire c190_r;
  wire c190_a;
  wire [35:0] c189_r0d;
  wire [35:0] c189_r1d;
  wire c189_a;
  wire c188_r;
  wire c188_a;
  wire [34:0] c187_r0d;
  wire [34:0] c187_r1d;
  wire c187_a;
  wire c186_r;
  wire c186_a;
  wire c185_r;
  wire c185_a;
  wire [35:0] c184_r0d;
  wire [35:0] c184_r1d;
  wire c184_a;
  wire c183_r;
  wire c183_a;
  wire c182_r;
  wire c182_a;
  wire [34:0] c181_r0d;
  wire [34:0] c181_r1d;
  wire c181_a;
  wire c180_r;
  wire c180_a;
  wire c179_r;
  wire c179_a;
  wire c178_r;
  wire c178_a;
  wire [3:0] c177_r0d;
  wire [3:0] c177_r1d;
  wire c177_a;
  wire c176_r;
  wire c176_a;
  wire c175_r;
  wire c175_a;
  wire [34:0] c174_r0d;
  wire [34:0] c174_r1d;
  wire c174_a;
  wire c173_r;
  wire c173_a;
  wire c172_r;
  wire c172_a;
  wire [35:0] c171_r0d;
  wire [35:0] c171_r1d;
  wire c171_a;
  wire c170_r;
  wire c170_a;
  wire c169_r;
  wire c169_a;
  wire c168_r;
  wire c168_a;
  wire c167_r;
  wire c167_a;
  wire c166_r;
  wire c166_a;
  wire c165_r0d;
  wire c165_r1d;
  wire c165_a;
  wire c164_r;
  wire c164_a;
  wire [31:0] c163_r0d;
  wire [31:0] c163_r1d;
  wire c163_a;
  wire c162_r;
  wire c162_a;
  wire [34:0] c161_r0d;
  wire [34:0] c161_r1d;
  wire c161_a;
  wire c160_r;
  wire c160_a;
  wire c159_r0d;
  wire c159_r1d;
  wire c159_a;
  wire [33:0] c158_r0d;
  wire [33:0] c158_r1d;
  wire c158_a;
  wire c157_r;
  wire c157_a;
  wire c156_r0d;
  wire c156_r1d;
  wire c156_a;
  wire [32:0] c155_r0d;
  wire [32:0] c155_r1d;
  wire c155_a;
  wire c154_r;
  wire c154_a;
  wire [31:0] c153_r0d;
  wire [31:0] c153_r1d;
  wire c153_a;
  wire c152_r;
  wire c152_a;
  wire c151_r0d;
  wire c151_r1d;
  wire c151_a;
  wire c150_r;
  wire c150_a;
  wire c149_r0d;
  wire c149_r1d;
  wire c149_a;
  wire c148_r;
  wire c148_a;
  wire c147_r;
  wire c147_a;
  wire c146_r;
  wire c146_a;
  wire [31:0] c145_r0d;
  wire [31:0] c145_r1d;
  wire c145_a;
  wire c144_r;
  wire c144_a;
  wire c143_r;
  wire c143_a;
  wire [31:0] c142_r0d;
  wire [31:0] c142_r1d;
  wire c142_a;
  wire c141_r;
  wire c141_a;
  wire c140_r;
  wire c140_a;
  wire [34:0] c139_r0d;
  wire [34:0] c139_r1d;
  wire c139_a;
  wire c138_r;
  wire c138_a;
  wire [32:0] c137_r0d;
  wire [32:0] c137_r1d;
  wire c137_a;
  wire [1:0] c136_r0d;
  wire [1:0] c136_r1d;
  wire c136_a;
  wire c135_r;
  wire c135_a;
  wire c134_r;
  wire c134_a;
  wire c133_r;
  wire c133_a;
  wire [34:0] c132_r0d;
  wire [34:0] c132_r1d;
  wire c132_a;
  wire c131_r;
  wire c131_a;
  wire [33:0] c130_r0d;
  wire [33:0] c130_r1d;
  wire c130_a;
  wire c129_r0d;
  wire c129_r1d;
  wire c129_a;
  wire c128_r;
  wire c128_a;
  wire c127_r;
  wire c127_a;
  wire c126_r;
  wire c126_a;
  wire [34:0] c125_r0d;
  wire [34:0] c125_r1d;
  wire c125_a;
  wire c124_r;
  wire c124_a;
  wire c123_r;
  wire c123_a;
  wire c122_r0d;
  wire c122_r1d;
  wire c122_a;
  wire c121_r;
  wire c121_a;
  wire c120_r;
  wire c120_a;
  wire c119_r0d;
  wire c119_r1d;
  wire c119_a;
  wire c118_r;
  wire c118_a;
  wire [32:0] c117_r0d;
  wire [32:0] c117_r1d;
  wire c117_a;
  wire [32:0] c116_r0d;
  wire [32:0] c116_r1d;
  wire c116_a;
  wire [33:0] c115_r0d;
  wire [33:0] c115_r1d;
  wire c115_a;
  wire c114_r;
  wire c114_a;
  wire c113_r;
  wire c113_a;
  wire c112_r;
  wire c112_a;
  wire c111_r;
  wire c111_a;
  wire c110_r;
  wire c110_a;
  wire [33:0] c109_r0d;
  wire [33:0] c109_r1d;
  wire c109_a;
  wire c108_r;
  wire c108_a;
  wire c107_r;
  wire c107_a;
  wire c106_r;
  wire c106_a;
  wire c105_r0d;
  wire c105_r1d;
  wire c105_a;
  wire c104_r;
  wire c104_a;
  wire c103_r;
  wire c103_a;
  wire [31:0] c102_r0d;
  wire [31:0] c102_r1d;
  wire c102_a;
  wire c101_r;
  wire c101_a;
  wire c100_r;
  wire c100_a;
  wire c99_r;
  wire c99_a;
  wire c98_r;
  wire c98_a;
  wire c97_r;
  wire c97_a;
  wire [32:0] c96_r0d;
  wire [32:0] c96_r1d;
  wire c96_a;
  wire c95_r;
  wire c95_a;
  wire [32:0] c94_r0d;
  wire [32:0] c94_r1d;
  wire c94_a;
  wire c93_r;
  wire c93_a;
  wire [33:0] c92_r0d;
  wire [33:0] c92_r1d;
  wire c92_a;
  wire [65:0] c91_r0d;
  wire [65:0] c91_r1d;
  wire c91_a;
  wire c90_r;
  wire c90_a;
  wire [32:0] c89_r0d;
  wire [32:0] c89_r1d;
  wire c89_a;
  wire c88_r;
  wire c88_a;
  wire [32:0] c87_r0d;
  wire [32:0] c87_r1d;
  wire c87_a;
  wire c86_r;
  wire c86_a;
  wire c85_r;
  wire c85_a;
  wire c84_r;
  wire c84_a;
  wire c83_r;
  wire c83_a;
  wire c82_r;
  wire c82_a;
  wire c81_r;
  wire c81_a;
  wire c80_r0d;
  wire c80_r1d;
  wire c80_a;
  wire c79_r;
  wire c79_a;
  wire [31:0] c78_r0d;
  wire [31:0] c78_r1d;
  wire c78_a;
  wire c77_r;
  wire c77_a;
  wire [31:0] c76_r0d;
  wire [31:0] c76_r1d;
  wire c76_a;
  wire c75_r;
  wire c75_a;
  wire c74_r;
  wire c74_a;
  wire c73_r;
  wire c73_a;
  wire [32:0] c72_r0d;
  wire [32:0] c72_r1d;
  wire c72_a;
  wire c71_r;
  wire c71_a;
  wire [31:0] c70_r0d;
  wire [31:0] c70_r1d;
  wire c70_a;
  wire c69_r;
  wire c69_a;
  wire c68_r0d;
  wire c68_r1d;
  wire c68_a;
  wire c67_r;
  wire c67_a;
  wire c66_r;
  wire c66_a;
  wire [32:0] c65_r0d;
  wire [32:0] c65_r1d;
  wire c65_a;
  wire c64_r;
  wire c64_a;
  wire [31:0] c63_r0d;
  wire [31:0] c63_r1d;
  wire c63_a;
  wire c62_r;
  wire c62_a;
  wire c61_r0d;
  wire c61_r1d;
  wire c61_a;
  wire c60_r;
  wire c60_a;
  wire c59_r;
  wire c59_a;
  wire c58_r;
  wire c58_a;
  wire c57_r;
  wire c57_a;
  wire c56_r;
  wire c56_a;
  wire c55_r;
  wire c55_a;
  wire c54_r;
  wire c54_a;
  wire [34:0] c53_r0d;
  wire [34:0] c53_r1d;
  wire c53_a;
  wire c52_r;
  wire c52_a;
  wire [34:0] c51_r0d;
  wire [34:0] c51_r1d;
  wire c51_a;
  wire c50_r;
  wire c50_a;
  wire [34:0] c49_r0d;
  wire [34:0] c49_r1d;
  wire c49_a;
  wire c48_r;
  wire c48_a;
  wire c47_r;
  wire c47_a;
  wire c46_r;
  wire c46_a;
  wire [34:0] c45_r0d;
  wire [34:0] c45_r1d;
  wire c45_a;
  wire [69:0] c44_r0d;
  wire [69:0] c44_r1d;
  wire c44_a;
  wire [34:0] c43_r0d;
  wire [34:0] c43_r1d;
  wire c43_a;
  wire [69:0] c42_r0d;
  wire [69:0] c42_r1d;
  wire c42_a;
  wire c41_r;
  wire c41_a;
  wire [34:0] c40_r0d;
  wire [34:0] c40_r1d;
  wire c40_a;
  wire c39_r;
  wire c39_a;
  wire [34:0] c38_r0d;
  wire [34:0] c38_r1d;
  wire c38_a;
  wire [34:0] c37_r0d;
  wire [34:0] c37_r1d;
  wire c37_a;
  wire [69:0] c36_r0d;
  wire [69:0] c36_r1d;
  wire c36_a;
  wire [34:0] c35_r0d;
  wire [34:0] c35_r1d;
  wire c35_a;
  wire [69:0] c34_r0d;
  wire [69:0] c34_r1d;
  wire c34_a;
  wire c33_r;
  wire c33_a;
  wire [34:0] c32_r0d;
  wire [34:0] c32_r1d;
  wire c32_a;
  wire c31_r;
  wire c31_a;
  wire [34:0] c30_r0d;
  wire [34:0] c30_r1d;
  wire c30_a;
  wire [34:0] c29_r0d;
  wire [34:0] c29_r1d;
  wire c29_a;
  wire [69:0] c28_r0d;
  wire [69:0] c28_r1d;
  wire c28_a;
  wire c27_r;
  wire c27_a;
  wire [34:0] c26_r0d;
  wire [34:0] c26_r1d;
  wire c26_a;
  wire c25_r;
  wire c25_a;
  wire [34:0] c24_r0d;
  wire [34:0] c24_r1d;
  wire c24_a;
  wire c23_r;
  wire c23_a;
  wire c22_r;
  wire c22_a;
  wire [34:0] c21_r0d;
  wire [34:0] c21_r1d;
  wire c21_a;
  wire [69:0] c20_r0d;
  wire [69:0] c20_r1d;
  wire c20_a;
  wire c19_r;
  wire c19_a;
  wire [34:0] c18_r0d;
  wire [34:0] c18_r1d;
  wire c18_a;
  wire [34:0] c17_r0d;
  wire [34:0] c17_r1d;
  wire c17_a;
  wire [69:0] c16_r0d;
  wire [69:0] c16_r1d;
  wire c16_a;
  wire c15_r;
  wire c15_a;
  wire [34:0] c14_r0d;
  wire [34:0] c14_r1d;
  wire c14_a;
  wire c13_r;
  wire c13_a;
  wire [34:0] c12_r0d;
  wire [34:0] c12_r1d;
  wire c12_a;
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I0 (c883_r0d, c883_r1d, c883_a, c607_r, c607_a, c630_r, c630_a, initialise);
  BrzJ_l11__280_202_29 I1 (c879_r, c879_a, c882_r0d, c882_r1d, c882_a, c883_r0d, c883_r1d, c883_a, initialise);
  BrzM_2_2 I2 (c880_r0d, c880_r1d, c880_a, c881_r0d, c881_r1d, c881_a, c882_r0d, c882_r1d, c882_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I3 (c876_r, c876_a, c881_r0d, c881_r1d, c881_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I4 (c874_r, c874_a, c880_r0d, c880_r1d, c880_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I5 (c878_r0d, c878_r1d, c878_a, c879_r, c879_a, mN_0r0d, mN_0r1d, mN_0a, initialise);
  BrzM_1_2 I6 (c875_r0d, c875_r1d, c875_a, c877_r0d, c877_r1d, c877_a, c878_r0d, c878_r1d, c878_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I7 (c629_r0d, c629_r1d, c629_a, c876_r, c876_a, c877_r0d, c877_r1d, c877_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I8 (c606_r0d, c606_r1d, c606_a, c874_r, c874_a, c875_r0d, c875_r1d, c875_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I9 (c873_r0d, c873_r1d, c873_a, c602_r, c602_a, c627_r, c627_a, initialise);
  BrzJ_l11__280_202_29 I10 (c869_r, c869_a, c872_r0d, c872_r1d, c872_a, c873_r0d, c873_r1d, c873_a, initialise);
  BrzM_2_2 I11 (c870_r0d, c870_r1d, c870_a, c871_r0d, c871_r1d, c871_a, c872_r0d, c872_r1d, c872_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I12 (c866_r, c866_a, c871_r0d, c871_r1d, c871_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I13 (c864_r, c864_a, c870_r0d, c870_r1d, c870_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I14 (c868_r0d, c868_r1d, c868_a, c869_r, c869_a, mZ_0r0d, mZ_0r1d, mZ_0a, initialise);
  BrzM_1_2 I15 (c865_r0d, c865_r1d, c865_a, c867_r0d, c867_r1d, c867_a, c868_r0d, c868_r1d, c868_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I16 (c626_r0d, c626_r1d, c626_a, c866_r, c866_a, c867_r0d, c867_r1d, c867_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I17 (c601_r0d, c601_r1d, c601_a, c864_r, c864_a, c865_r0d, c865_r1d, c865_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I18 (c863_r0d, c863_r1d, c863_a, c597_r, c597_a, c624_r, c624_a, initialise);
  BrzJ_l11__280_202_29 I19 (c859_r, c859_a, c862_r0d, c862_r1d, c862_a, c863_r0d, c863_r1d, c863_a, initialise);
  BrzM_2_2 I20 (c860_r0d, c860_r1d, c860_a, c861_r0d, c861_r1d, c861_a, c862_r0d, c862_r1d, c862_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I21 (c856_r, c856_a, c861_r0d, c861_r1d, c861_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I22 (c854_r, c854_a, c860_r0d, c860_r1d, c860_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I23 (c858_r0d, c858_r1d, c858_a, c859_r, c859_a, mpL_0r0d, mpL_0r1d, mpL_0a, initialise);
  BrzM_32_2 I24 (c855_r0d, c855_r1d, c855_a, c857_r0d, c857_r1d, c857_a, c858_r0d, c858_r1d, c858_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I25 (c623_r0d, c623_r1d, c623_a, c856_r, c856_a, c857_r0d, c857_r1d, c857_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I26 (c596_r0d, c596_r1d, c596_a, c854_r, c854_a, c855_r0d, c855_r1d, c855_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I27 (c853_r0d, c853_r1d, c853_a, c615_r, c615_a, c636_r, c636_a, initialise);
  BrzJ_l11__280_202_29 I28 (c849_r, c849_a, c852_r0d, c852_r1d, c852_a, c853_r0d, c853_r1d, c853_a, initialise);
  BrzM_2_2 I29 (c850_r0d, c850_r1d, c850_a, c851_r0d, c851_r1d, c851_a, c852_r0d, c852_r1d, c852_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I30 (c846_r, c846_a, c851_r0d, c851_r1d, c851_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I31 (c844_r, c844_a, c850_r0d, c850_r1d, c850_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I32 (c848_r0d, c848_r1d, c848_a, c849_r, c849_a, mpH_0r0d, mpH_0r1d, mpH_0a, initialise);
  BrzM_32_2 I33 (c845_r0d, c845_r1d, c845_a, c847_r0d, c847_r1d, c847_a, c848_r0d, c848_r1d, c848_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I34 (c635_r0d, c635_r1d, c635_a, c846_r, c846_a, c847_r0d, c847_r1d, c847_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I35 (c614_r0d, c614_r1d, c614_a, c844_r, c844_a, c845_r0d, c845_r1d, c845_a, initialise);
  BrzS_34_l12__2832_202_29_l97__28_28_28_281_m69m I36 (c843_r0d, c843_r1d, c843_a, c554_r0d, c554_r1d, c554_a, c563_r0d, c563_r1d, c563_a, initialise);
  BrzJ_l12__2832_202_29 I37 (c_0r0d, c_0r1d, c_0a, c842_r0d, c842_r1d, c842_a, c843_r0d, c843_r1d, c843_a, initialise);
  BrzM_2_2 I38 (c840_r0d, c840_r1d, c840_a, c841_r0d, c841_r1d, c841_a, c842_r0d, c842_r1d, c842_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I39 (c565_r, c565_a, c841_r0d, c841_r1d, c841_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I40 (c556_r, c556_a, c840_r0d, c840_r1d, c840_a);
  BrzJ_l12__2832_200_29 I41 (b_0r0d, b_0r1d, b_0a, c574_r, c574_a, c570_r0d, c570_r1d, c570_a, initialise);
  BrzJ_l12__2832_200_29 I42 (a_0r0d, a_0r1d, a_0a, c573_r, c573_a, c568_r0d, c568_r1d, c568_a, initialise);
  BrzJ_l11__283_200_29 I43 (mType_0r0d, mType_0r1d, mType_0a, c592_r, c592_a, c587_r0d, c587_r1d, c587_a, initialise);
  BrzJ_l11__281_200_29 I44 (bypassH_0r0d, bypassH_0r1d, bypassH_0a, c591_r, c591_a, c585_r0d, c585_r1d, c585_a, initialise);
  BrzJ_l11__281_200_29 I45 (bypass_0r0d, bypass_0r1d, bypass_0a, c590_r, c590_a, c583_r0d, c583_r1d, c583_a, initialise);
  BrzJ_l12__2835_200_29 I46 (c835_r0d, c835_r1d, c835_a, c198_r, c198_a, c187_r0d, c187_r1d, c187_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I47 (c839_r0d, c839_r1d, c839_a, c485_r, c485_a, c499_r, c499_a, initialise);
  BrzJ_l11__280_202_29 I48 (c834_r, c834_a, c838_r0d, c838_r1d, c838_a, c839_r0d, c839_r1d, c839_a, initialise);
  BrzM_2_2 I49 (c836_r0d, c836_r1d, c836_a, c837_r0d, c837_r1d, c837_a, c838_r0d, c838_r1d, c838_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I50 (c831_r, c831_a, c837_r0d, c837_r1d, c837_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I51 (c829_r, c829_a, c836_r0d, c836_r1d, c836_a);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I52 (c833_r0d, c833_r1d, c833_a, c834_r, c834_a, c835_r0d, c835_r1d, c835_a, initialise);
  BrzM_35_2 I53 (c830_r0d, c830_r1d, c830_a, c832_r0d, c832_r1d, c832_a, c833_r0d, c833_r1d, c833_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I54 (c496_r0d, c496_r1d, c496_a, c831_r, c831_a, c832_r0d, c832_r1d, c832_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I55 (c482_r0d, c482_r1d, c482_a, c829_r, c829_a, c830_r0d, c830_r1d, c830_a, initialise);
  BrzJ_l12__2836_200_29 I56 (c824_r0d, c824_r1d, c824_a, c199_r, c199_a, c189_r0d, c189_r1d, c189_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I57 (c828_r0d, c828_r1d, c828_a, c493_r, c493_a, c507_r, c507_a, initialise);
  BrzJ_l11__280_202_29 I58 (c823_r, c823_a, c827_r0d, c827_r1d, c827_a, c828_r0d, c828_r1d, c828_a, initialise);
  BrzM_2_2 I59 (c825_r0d, c825_r1d, c825_a, c826_r0d, c826_r1d, c826_a, c827_r0d, c827_r1d, c827_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I60 (c820_r, c820_a, c826_r0d, c826_r1d, c826_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I61 (c818_r, c818_a, c825_r0d, c825_r1d, c825_a);
  BrzF_36_l32__28_280_200_29_20_280_2036_29__m44m I62 (c822_r0d, c822_r1d, c822_a, c823_r, c823_a, c824_r0d, c824_r1d, c824_a, initialise);
  BrzM_36_2 I63 (c819_r0d, c819_r1d, c819_a, c821_r0d, c821_r1d, c821_a, c822_r0d, c822_r1d, c822_a, initialise);
  BrzF_36_l32__28_280_200_29_20_280_2036_29__m44m I64 (c500_r0d, c500_r1d, c500_a, c820_r, c820_a, c821_r0d, c821_r1d, c821_a, initialise);
  BrzF_36_l32__28_280_200_29_20_280_2036_29__m44m I65 (c486_r0d, c486_r1d, c486_a, c818_r, c818_a, c819_r0d, c819_r1d, c819_a, initialise);
  BrzJ_l12__2835_200_29 I66 (c817_r0d, c817_r1d, c817_a, c200_r, c200_a, c191_r0d, c191_r1d, c191_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I67 (c511_r0d, c511_r1d, c511_a, c514_r, c514_a, c817_r0d, c817_r1d, c817_a, initialise);
  BrzJ_l11__281_200_29 I68 (c816_r0d, c816_r1d, c816_a, c201_r, c201_a, c193_r0d, c193_r1d, c193_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I69 (c515_r0d, c515_r1d, c515_a, c517_r, c517_a, c816_r0d, c816_r1d, c816_a, initialise);
  BrzJ_l11__281_200_29 I70 (c815_r0d, c815_r1d, c815_a, c202_r, c202_a, c195_r0d, c195_r1d, c195_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I71 (c518_r0d, c518_r1d, c518_a, c520_r, c520_a, c815_r0d, c815_r1d, c815_a, initialise);
  BrzJ_l12__2832_200_29 I72 (c814_r0d, c814_r1d, c814_a, c532_r, c532_a, c524_r0d, c524_r1d, c524_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I73 (c538_r0d, c538_r1d, c538_a, c540_r, c540_a, c814_r0d, c814_r1d, c814_a, initialise);
  BrzJ_l12__2832_200_29 I74 (c813_r0d, c813_r1d, c813_a, c533_r, c533_a, c526_r0d, c526_r1d, c526_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I75 (c541_r0d, c541_r1d, c541_a, c543_r, c543_a, c813_r0d, c813_r1d, c813_a, initialise);
  BrzJ_l12__2832_200_29 I76 (c808_r0d, c808_r1d, c808_a, c534_r, c534_a, c528_r0d, c528_r1d, c528_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I77 (c812_r0d, c812_r1d, c812_a, c551_r, c551_a, c553_r, c553_a, initialise);
  BrzJ_l11__280_202_29 I78 (c807_r, c807_a, c811_r0d, c811_r1d, c811_a, c812_r0d, c812_r1d, c812_a, initialise);
  BrzM_2_2 I79 (c809_r0d, c809_r1d, c809_a, c810_r0d, c810_r1d, c810_a, c811_r0d, c811_r1d, c811_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I80 (c804_r, c804_a, c810_r0d, c810_r1d, c810_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I81 (c802_r, c802_a, c809_r0d, c809_r1d, c809_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I82 (c806_r0d, c806_r1d, c806_a, c807_r, c807_a, c808_r0d, c808_r1d, c808_a, initialise);
  BrzM_32_2 I83 (c803_r0d, c803_r1d, c803_a, c805_r0d, c805_r1d, c805_a, c806_r0d, c806_r1d, c806_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I84 (c552_r0d, c552_r1d, c552_a, c804_r, c804_a, c805_r0d, c805_r1d, c805_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I85 (c550_r0d, c550_r1d, c550_a, c802_r, c802_a, c803_r0d, c803_r1d, c803_a, initialise);
  BrzJ_l11__283_200_29 I86 (c801_r0d, c801_r1d, c801_a, c531_r, c531_a, c522_r0d, c522_r1d, c522_a, initialise);
  BrzF_3_l31__28_280_200_29_20_280_203_29_29 I87 (c544_r0d, c544_r1d, c544_a, c546_r, c546_a, c801_r0d, c801_r1d, c801_a, initialise);
  BrzJ_l12__2835_200_29 I88 (c800_r0d, c800_r1d, c800_a, c56_r, c56_a, c49_r0d, c49_r1d, c49_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I89 (c224_r0d, c224_r1d, c224_a, c226_r, c226_a, c800_r0d, c800_r1d, c800_a, initialise);
  BrzJ_l12__2835_200_29 I90 (c788_r0d, c788_r1d, c788_a, c57_r, c57_a, c51_r0d, c51_r1d, c51_a, initialise);
  BrzS_9_l11__280_209_29_l424__28_28_28_281__m68m I91 (c799_r0d, c799_r1d, c799_a, c248_r, c248_a, c251_r, c251_a, c254_r, c254_a, c257_r, c257_a, c260_r, c260_a, c263_r, c263_a, c266_r, c266_a, c269_r, c269_a, c272_r, c272_a, initialise);
  BrzJ_l11__280_209_29 I92 (c787_r, c787_a, c798_r0d, c798_r1d, c798_a, c799_r0d, c799_r1d, c799_a, initialise);
  BrzM_9_9 I93 (c789_r0d, c789_r1d, c789_a, c790_r0d, c790_r1d, c790_a, c791_r0d, c791_r1d, c791_a, c792_r0d, c792_r1d, c792_a, c793_r0d, c793_r1d, c793_a, c794_r0d, c794_r1d, c794_a, c795_r0d, c795_r1d, c795_a, c796_r0d, c796_r1d, c796_a, c797_r0d, c797_r1d, c797_a, c798_r0d, c798_r1d, c798_a, initialise);
  BrzO_0_9_l25__28_28num_209_20256_29_29 I94 (c784_r, c784_a, c797_r0d, c797_r1d, c797_a);
  BrzO_0_9_l25__28_28num_209_20128_29_29 I95 (c782_r, c782_a, c796_r0d, c796_r1d, c796_a);
  BrzO_0_9_l24__28_28num_209_2064_29_29 I96 (c780_r, c780_a, c795_r0d, c795_r1d, c795_a);
  BrzO_0_9_l24__28_28num_209_2032_29_29 I97 (c778_r, c778_a, c794_r0d, c794_r1d, c794_a);
  BrzO_0_9_l24__28_28num_209_2016_29_29 I98 (c776_r, c776_a, c793_r0d, c793_r1d, c793_a);
  BrzO_0_9_l23__28_28num_209_208_29_29 I99 (c774_r, c774_a, c792_r0d, c792_r1d, c792_a);
  BrzO_0_9_l23__28_28num_209_204_29_29 I100 (c772_r, c772_a, c791_r0d, c791_r1d, c791_a);
  BrzO_0_9_l23__28_28num_209_202_29_29 I101 (c770_r, c770_a, c790_r0d, c790_r1d, c790_a);
  BrzO_0_9_l23__28_28num_209_201_29_29 I102 (c768_r, c768_a, c789_r0d, c789_r1d, c789_a);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I103 (c786_r0d, c786_r1d, c786_a, c787_r, c787_a, c788_r0d, c788_r1d, c788_a, initialise);
  BrzM_35_9 I104 (c769_r0d, c769_r1d, c769_a, c771_r0d, c771_r1d, c771_a, c773_r0d, c773_r1d, c773_a, c775_r0d, c775_r1d, c775_a, c777_r0d, c777_r1d, c777_a, c779_r0d, c779_r1d, c779_a, c781_r0d, c781_r1d, c781_a, c783_r0d, c783_r1d, c783_a, c785_r0d, c785_r1d, c785_a, c786_r0d, c786_r1d, c786_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I105 (c270_r0d, c270_r1d, c270_a, c784_r, c784_a, c785_r0d, c785_r1d, c785_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I106 (c267_r0d, c267_r1d, c267_a, c782_r, c782_a, c783_r0d, c783_r1d, c783_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I107 (c264_r0d, c264_r1d, c264_a, c780_r, c780_a, c781_r0d, c781_r1d, c781_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I108 (c261_r0d, c261_r1d, c261_a, c778_r, c778_a, c779_r0d, c779_r1d, c779_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I109 (c258_r0d, c258_r1d, c258_a, c776_r, c776_a, c777_r0d, c777_r1d, c777_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I110 (c255_r0d, c255_r1d, c255_a, c774_r, c774_a, c775_r0d, c775_r1d, c775_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I111 (c252_r0d, c252_r1d, c252_a, c772_r, c772_a, c773_r0d, c773_r1d, c773_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I112 (c249_r0d, c249_r1d, c249_a, c770_r, c770_a, c771_r0d, c771_r1d, c771_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I113 (c245_r0d, c245_r1d, c245_a, c768_r, c768_a, c769_r0d, c769_r1d, c769_a, initialise);
  BrzJ_l12__2835_200_29 I114 (c767_r0d, c767_r1d, c767_a, c58_r, c58_a, c53_r0d, c53_r1d, c53_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I115 (c227_r0d, c227_r1d, c227_a, c229_r, c229_a, c767_r0d, c767_r1d, c767_a, initialise);
  BrzJ_l12__2835_200_29 I116 (c766_r0d, c766_r1d, c766_a, c239_r, c239_a, c237_r0d, c237_r1d, c237_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I117 (c45_r0d, c45_r1d, c45_a, c47_r, c47_a, c766_r0d, c766_r1d, c766_a, initialise);
  BrzJ_l12__2835_200_29 I118 (c765_r0d, c765_r1d, c765_a, c234_r, c234_a, c232_r0d, c232_r1d, c232_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I119 (c21_r0d, c21_r1d, c21_a, c23_r, c23_a, c765_r0d, c765_r1d, c765_a, initialise);
  BrzJ_l12__2832_200_29 I120 (c759_r0d, c759_r1d, c759_a, c83_r, c83_a, c76_r0d, c76_r1d, c76_a, initialise);
  BrzS_3_l11__280_203_29_l141__28_28_28_281__m64m I121 (c764_r0d, c764_r1d, c764_a, c144_r, c144_a, c349_r, c349_a, c402_r, c402_a, initialise);
  BrzJ_l11__280_203_29 I122 (c758_r, c758_a, c763_r0d, c763_r1d, c763_a, c764_r0d, c764_r1d, c764_a, initialise);
  BrzM_3_3 I123 (c760_r0d, c760_r1d, c760_a, c761_r0d, c761_r1d, c761_a, c762_r0d, c762_r1d, c762_a, c763_r0d, c763_r1d, c763_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I124 (c755_r, c755_a, c762_r0d, c762_r1d, c762_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I125 (c753_r, c753_a, c761_r0d, c761_r1d, c761_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I126 (c751_r, c751_a, c760_r0d, c760_r1d, c760_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I127 (c757_r0d, c757_r1d, c757_a, c758_r, c758_a, c759_r0d, c759_r1d, c759_a, initialise);
  BrzM_32_3 I128 (c752_r0d, c752_r1d, c752_a, c754_r0d, c754_r1d, c754_a, c756_r0d, c756_r1d, c756_a, c757_r0d, c757_r1d, c757_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I129 (c400_r0d, c400_r1d, c400_a, c755_r, c755_a, c756_r0d, c756_r1d, c756_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I130 (c347_r0d, c347_r1d, c347_a, c753_r, c753_a, c754_r0d, c754_r1d, c754_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I131 (c142_r0d, c142_r1d, c142_a, c751_r, c751_a, c752_r0d, c752_r1d, c752_a, initialise);
  BrzJ_l12__2832_200_29 I132 (c745_r0d, c745_r1d, c745_a, c84_r, c84_a, c78_r0d, c78_r1d, c78_a, initialise);
  BrzS_3_l11__280_203_29_l141__28_28_28_281__m64m I133 (c750_r0d, c750_r1d, c750_a, c147_r, c147_a, c352_r, c352_a, c405_r, c405_a, initialise);
  BrzJ_l11__280_203_29 I134 (c744_r, c744_a, c749_r0d, c749_r1d, c749_a, c750_r0d, c750_r1d, c750_a, initialise);
  BrzM_3_3 I135 (c746_r0d, c746_r1d, c746_a, c747_r0d, c747_r1d, c747_a, c748_r0d, c748_r1d, c748_a, c749_r0d, c749_r1d, c749_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I136 (c741_r, c741_a, c748_r0d, c748_r1d, c748_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I137 (c739_r, c739_a, c747_r0d, c747_r1d, c747_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I138 (c737_r, c737_a, c746_r0d, c746_r1d, c746_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I139 (c743_r0d, c743_r1d, c743_a, c744_r, c744_a, c745_r0d, c745_r1d, c745_a, initialise);
  BrzM_32_3 I140 (c738_r0d, c738_r1d, c738_a, c740_r0d, c740_r1d, c740_a, c742_r0d, c742_r1d, c742_a, c743_r0d, c743_r1d, c743_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I141 (c403_r0d, c403_r1d, c403_a, c741_r, c741_a, c742_r0d, c742_r1d, c742_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I142 (c350_r0d, c350_r1d, c350_a, c739_r, c739_a, c740_r0d, c740_r1d, c740_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I143 (c145_r0d, c145_r1d, c145_a, c737_r, c737_a, c738_r0d, c738_r1d, c738_a, initialise);
  BrzJ_l11__281_200_29 I144 (c731_r0d, c731_r1d, c731_a, c85_r, c85_a, c80_r0d, c80_r1d, c80_a, initialise);
  BrzS_3_l11__280_203_29_l141__28_28_28_281__m64m I145 (c736_r0d, c736_r1d, c736_a, c150_r, c150_a, c355_r, c355_a, c408_r, c408_a, initialise);
  BrzJ_l11__280_203_29 I146 (c730_r, c730_a, c735_r0d, c735_r1d, c735_a, c736_r0d, c736_r1d, c736_a, initialise);
  BrzM_3_3 I147 (c732_r0d, c732_r1d, c732_a, c733_r0d, c733_r1d, c733_a, c734_r0d, c734_r1d, c734_a, c735_r0d, c735_r1d, c735_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I148 (c727_r, c727_a, c734_r0d, c734_r1d, c734_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I149 (c725_r, c725_a, c733_r0d, c733_r1d, c733_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I150 (c723_r, c723_a, c732_r0d, c732_r1d, c732_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I151 (c729_r0d, c729_r1d, c729_a, c730_r, c730_a, c731_r0d, c731_r1d, c731_a, initialise);
  BrzM_1_3 I152 (c724_r0d, c724_r1d, c724_a, c726_r0d, c726_r1d, c726_a, c728_r0d, c728_r1d, c728_a, c729_r0d, c729_r1d, c729_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I153 (c406_r0d, c406_r1d, c406_a, c727_r, c727_a, c728_r0d, c728_r1d, c728_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I154 (c354_r0d, c354_r1d, c354_a, c725_r, c725_a, c726_r0d, c726_r1d, c726_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I155 (c149_r0d, c149_r1d, c149_a, c723_r, c723_a, c724_r0d, c724_r1d, c724_a, initialise);
  BrzS_35_l12__2832_203_29_l144__28_28_28_28_m70m I156 (c722_r0d, c722_r1d, c722_a, c163_r0d, c163_r1d, c163_a, c374_r0d, c374_r1d, c374_a, c411_r0d, c411_r1d, c411_a, initialise);
  BrzJ_l12__2832_203_29 I157 (c717_r0d, c717_r1d, c717_a, c721_r0d, c721_r1d, c721_a, c722_r0d, c722_r1d, c722_a, initialise);
  BrzM_3_3 I158 (c718_r0d, c718_r1d, c718_a, c719_r0d, c719_r1d, c719_a, c720_r0d, c720_r1d, c720_a, c721_r0d, c721_r1d, c721_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I159 (c416_r, c416_a, c720_r0d, c720_r1d, c720_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I160 (c379_r, c379_a, c719_r0d, c719_r1d, c719_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I161 (c168_r, c168_a, c718_r0d, c718_r1d, c718_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I162 (c102_r0d, c102_r1d, c102_a, c104_r, c104_a, c717_r0d, c717_r1d, c717_a, initialise);
  BrzS_4_l11__281_203_29_l141__28_28_28_281__m67m I163 (c716_r0d, c716_r1d, c716_a, c165_r0d, c165_r1d, c165_a, c376_r0d, c376_r1d, c376_a, c413_r0d, c413_r1d, c413_a, initialise);
  BrzJ_l11__281_203_29 I164 (c711_r0d, c711_r1d, c711_a, c715_r0d, c715_r1d, c715_a, c716_r0d, c716_r1d, c716_a, initialise);
  BrzM_3_3 I165 (c712_r0d, c712_r1d, c712_a, c713_r0d, c713_r1d, c713_a, c714_r0d, c714_r1d, c714_a, c715_r0d, c715_r1d, c715_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I166 (c417_r, c417_a, c714_r0d, c714_r1d, c714_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I167 (c380_r, c380_a, c713_r0d, c713_r1d, c713_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I168 (c169_r, c169_a, c712_r0d, c712_r1d, c712_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I169 (c105_r0d, c105_r1d, c105_a, c107_r, c107_a, c711_r0d, c711_r1d, c711_a, initialise);
  BrzJ_l11__281_200_29 I170 (c706_r0d, c706_r1d, c706_a, c453_r, c453_a, c456_r0d, c456_r1d, c456_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I171 (c710_r0d, c710_r1d, c710_a, c221_r, c221_a, c343_r, c343_a, initialise);
  BrzJ_l11__280_202_29 I172 (c705_r, c705_a, c709_r0d, c709_r1d, c709_a, c710_r0d, c710_r1d, c710_a, initialise);
  BrzM_2_2 I173 (c707_r0d, c707_r1d, c707_a, c708_r0d, c708_r1d, c708_a, c709_r0d, c709_r1d, c709_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I174 (c702_r, c702_a, c708_r0d, c708_r1d, c708_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I175 (c700_r, c700_a, c707_r0d, c707_r1d, c707_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I176 (c704_r0d, c704_r1d, c704_a, c705_r, c705_a, c706_r0d, c706_r1d, c706_a, initialise);
  BrzM_1_2 I177 (c701_r0d, c701_r1d, c701_a, c703_r0d, c703_r1d, c703_a, c704_r0d, c704_r1d, c704_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I178 (c342_r0d, c342_r1d, c342_a, c702_r, c702_a, c703_r0d, c703_r1d, c703_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I179 (c220_r0d, c220_r1d, c220_a, c700_r, c700_a, c701_r0d, c701_r1d, c701_a, initialise);
  BrzJ_l11__281_200_29 I180 (c695_r0d, c695_r1d, c695_a, c316_r, c316_a, c314_r0d, c314_r1d, c314_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I181 (c699_r0d, c699_r1d, c699_a, c462_r, c462_a, c475_r, c475_a, initialise);
  BrzJ_l11__280_202_29 I182 (c694_r, c694_a, c698_r0d, c698_r1d, c698_a, c699_r0d, c699_r1d, c699_a, initialise);
  BrzM_2_2 I183 (c696_r0d, c696_r1d, c696_a, c697_r0d, c697_r1d, c697_a, c698_r0d, c698_r1d, c698_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I184 (c691_r, c691_a, c697_r0d, c697_r1d, c697_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I185 (c689_r, c689_a, c696_r0d, c696_r1d, c696_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I186 (c693_r0d, c693_r1d, c693_a, c694_r, c694_a, c695_r0d, c695_r1d, c695_a, initialise);
  BrzM_1_2 I187 (c690_r0d, c690_r1d, c690_a, c692_r0d, c692_r1d, c692_a, c693_r0d, c693_r1d, c693_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I188 (c474_r0d, c474_r1d, c474_a, c691_r, c691_a, c692_r0d, c692_r1d, c692_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I189 (c460_r0d, c460_r1d, c460_a, c689_r, c689_a, c690_r0d, c690_r1d, c690_a, initialise);
  BrzJ_l12__2832_200_29 I190 (c688_r0d, c688_r1d, c688_a, c618_r, c618_a, c616_r0d, c616_r1d, c616_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I191 (c420_r0d, c420_r1d, c420_a, c422_r, c422_a, c688_r0d, c688_r1d, c688_a, initialise);
  BrzJ_l12__2832_200_29 I192 (c683_r0d, c683_r1d, c683_a, c600_r, c600_a, c598_r0d, c598_r1d, c598_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I193 (c687_r0d, c687_r1d, c687_a, c386_r, c386_a, c425_r, c425_a, initialise);
  BrzJ_l11__280_202_29 I194 (c682_r, c682_a, c686_r0d, c686_r1d, c686_a, c687_r0d, c687_r1d, c687_a, initialise);
  BrzM_2_2 I195 (c684_r0d, c684_r1d, c684_a, c685_r0d, c685_r1d, c685_a, c686_r0d, c686_r1d, c686_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I196 (c679_r, c679_a, c685_r0d, c685_r1d, c685_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I197 (c677_r, c677_a, c684_r0d, c684_r1d, c684_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I198 (c681_r0d, c681_r1d, c681_a, c682_r, c682_a, c683_r0d, c683_r1d, c683_a, initialise);
  BrzM_32_2 I199 (c678_r0d, c678_r1d, c678_a, c680_r0d, c680_r1d, c680_a, c681_r0d, c681_r1d, c681_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I200 (c423_r0d, c423_r1d, c423_a, c679_r, c679_a, c680_r0d, c680_r1d, c680_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I201 (c384_r0d, c384_r1d, c384_a, c677_r, c677_a, c678_r0d, c678_r1d, c678_a, initialise);
  BrzJ_l11__281_200_29 I202 (c671_r0d, c671_r1d, c671_a, c605_r, c605_a, c603_r0d, c603_r1d, c603_a, initialise);
  BrzS_3_l11__280_203_29_l141__28_28_28_281__m64m I203 (c676_r0d, c676_r1d, c676_a, c389_r, c389_a, c439_r, c439_a, c442_r, c442_a, initialise);
  BrzJ_l11__280_203_29 I204 (c670_r, c670_a, c675_r0d, c675_r1d, c675_a, c676_r0d, c676_r1d, c676_a, initialise);
  BrzM_3_3 I205 (c672_r0d, c672_r1d, c672_a, c673_r0d, c673_r1d, c673_a, c674_r0d, c674_r1d, c674_a, c675_r0d, c675_r1d, c675_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I206 (c667_r, c667_a, c674_r0d, c674_r1d, c674_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I207 (c665_r, c665_a, c673_r0d, c673_r1d, c673_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I208 (c663_r, c663_a, c672_r0d, c672_r1d, c672_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I209 (c669_r0d, c669_r1d, c669_a, c670_r, c670_a, c671_r0d, c671_r1d, c671_a, initialise);
  BrzM_1_3 I210 (c664_r0d, c664_r1d, c664_a, c666_r0d, c666_r1d, c666_a, c668_r0d, c668_r1d, c668_a, c669_r0d, c669_r1d, c669_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I211 (c440_r0d, c440_r1d, c440_a, c667_r, c667_a, c668_r0d, c668_r1d, c668_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I212 (c437_r0d, c437_r1d, c437_a, c665_r, c665_a, c666_r0d, c666_r1d, c666_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I213 (c387_r0d, c387_r1d, c387_a, c663_r, c663_a, c664_r0d, c664_r1d, c664_a, initialise);
  BrzJ_l11__281_200_29 I214 (c658_r0d, c658_r1d, c658_a, c610_r, c610_a, c608_r0d, c608_r1d, c608_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I215 (c662_r0d, c662_r1d, c662_a, c392_r, c392_a, c446_r, c446_a, initialise);
  BrzJ_l11__280_202_29 I216 (c657_r, c657_a, c661_r0d, c661_r1d, c661_a, c662_r0d, c662_r1d, c662_a, initialise);
  BrzM_2_2 I217 (c659_r0d, c659_r1d, c659_a, c660_r0d, c660_r1d, c660_a, c661_r0d, c661_r1d, c661_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I218 (c654_r, c654_a, c660_r0d, c660_r1d, c660_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I219 (c652_r, c652_a, c659_r0d, c659_r1d, c659_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I220 (c656_r0d, c656_r1d, c656_a, c657_r, c657_a, c658_r0d, c658_r1d, c658_a, initialise);
  BrzM_1_2 I221 (c653_r0d, c653_r1d, c653_a, c655_r0d, c655_r1d, c655_a, c656_r0d, c656_r1d, c656_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I222 (c444_r0d, c444_r1d, c444_a, c654_r, c654_a, c655_r0d, c655_r1d, c655_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I223 (c390_r0d, c390_r1d, c390_a, c652_r, c652_a, c653_r0d, c653_r1d, c653_a, initialise);
  BrzJ_l11__281_200_29 I224 (c651_r0d, c651_r1d, c651_a, c646_r, c646_a, c641_r0d, c641_r1d, c641_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I225 (c579_r0d, c579_r1d, c579_a, c581_r, c581_a, c651_r0d, c651_r1d, c651_a, initialise);
  BrzJ_l11__281_200_29 I226 (c650_r0d, c650_r1d, c650_a, c647_r, c647_a, c643_r0d, c643_r1d, c643_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I227 (c576_r0d, c576_r1d, c576_a, c578_r, c578_a, c650_r0d, c650_r1d, c650_a, initialise);
  BrzF_0_l101__28_280_200_29_20_280_200_29_2_m37m I228 (go_0r, go_0a, c60_r, c60_a, c114_r, c114_a, c449_r, c449_a, c479_r, c479_a, c536_r, c536_a, c594_r, c594_a, c649_r, c649_a, initialise);
  BrzM_0_2 I229 (c649_r, c649_a, c640_r, c640_a, c648_r, c648_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I230 (c648_r, c648_a, c646_r, c646_a, c647_r, c647_a, initialise);
  BrzJ_l11__280_200_29 I231 (c642_r, c642_a, c644_r, c644_a, c645_r, c645_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I232 (c643_r0d, c643_r1d, c643_a, c644_r, c644_a, c645_r, c645_a, c595_r0d, c595_r1d, c595_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m72m I233 (c641_r0d, c641_r1d, c641_a, c642_r, c642_a, c612_r, c612_a, c632_r, c632_a, c611_r0d, c611_r1d, c611_a, c631_r0d, c631_r1d, c631_a, initialise);
  BrzM_0_2 I234 (c621_r, c621_a, c639_r, c639_a, c640_r, c640_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I235 (c595_r0d, c595_r1d, c595_a, c620_r, c620_a, c638_r, c638_a, initialise);
  BrzJ_l19__280_200_200_200_29 I236 (c624_r, c624_a, c627_r, c627_a, c630_r, c630_a, c637_r, c637_a, c639_r, c639_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I237 (c638_r, c638_a, c622_r, c622_a, c625_r, c625_a, c628_r, c628_a, c632_r, c632_a, initialise);
  BrzM_0_2 I238 (c633_r, c633_a, c636_r, c636_a, c637_r, c637_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I239 (c631_r0d, c631_r1d, c631_a, c633_r, c633_a, c634_r, c634_a, initialise);
  BrzO_0_32_l24__28_28num_2032_200_29_29 I240 (c634_r, c634_a, c635_r0d, c635_r1d, c635_a);
  BrzO_0_1_l23__28_28num_201_200_29_29 I241 (c628_r, c628_a, c629_r0d, c629_r1d, c629_a);
  BrzO_0_1_l23__28_28num_201_200_29_29 I242 (c625_r, c625_a, c626_r0d, c626_r1d, c626_a);
  BrzO_0_32_l24__28_28num_2032_200_29_29 I243 (c622_r, c622_a, c623_r0d, c623_r1d, c623_a);
  BrzJ_l19__280_200_200_200_29 I244 (c597_r, c597_a, c602_r, c602_a, c607_r, c607_a, c619_r, c619_a, c621_r, c621_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I245 (c620_r, c620_a, c600_r, c600_a, c605_r, c605_a, c610_r, c610_a, c612_r, c612_a, initialise);
  BrzM_0_2 I246 (c613_r, c613_a, c615_r, c615_a, c619_r, c619_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I247 (c611_r0d, c611_r1d, c611_a, c613_r, c613_a, c618_r, c618_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I248 (c616_r0d, c616_r1d, c616_a, c617_r, c617_a, c617_r, c617_a, c614_r0d, c614_r1d, c614_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I249 (c608_r0d, c608_r1d, c608_a, c609_r, c609_a, c609_r, c609_a, c606_r0d, c606_r1d, c606_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I250 (c603_r0d, c603_r1d, c603_a, c604_r, c604_a, c604_r, c604_a, c601_r0d, c601_r1d, c601_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I251 (c598_r0d, c598_r1d, c598_a, c599_r, c599_a, c599_r, c599_a, c596_r0d, c596_r1d, c596_a, initialise);
  BrzM_0_2 I252 (c594_r, c594_a, c582_r, c582_a, c593_r, c593_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I253 (c593_r, c593_a, c590_r, c590_a, c591_r, c591_a, c592_r, c592_a, initialise);
  BrzJ_l15__280_200_200_29 I254 (c584_r, c584_a, c586_r, c586_a, c588_r, c588_a, c589_r, c589_a, initialise);
  BrzV_3_l6__28_29_l23__28_28_280_203_29_29__m75m I255 (c587_r0d, c587_r1d, c587_a, c588_r, c588_a, c545_r, c545_a, c548_r, c548_a, c561_r, c561_a, c544_r0d, c544_r1d, c544_a, c547_r0d, c547_r1d, c547_a, c560_r0d, c560_r1d, c560_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I256 (c585_r0d, c585_r1d, c585_a, c586_r, c586_a, c580_r, c580_a, c579_r0d, c579_r1d, c579_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m72m I257 (c583_r0d, c583_r1d, c583_a, c584_r, c584_a, c572_r, c572_a, c577_r, c577_a, c537_r0d, c537_r1d, c537_a, c576_r0d, c576_r1d, c576_a, initialise);
  BrzJ_l15__280_200_200_29 I258 (c567_r, c567_a, c578_r, c578_a, c581_r, c581_a, c582_r, c582_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I259 (c589_r, c589_a, c575_r, c575_a, c577_r, c577_a, c580_r, c580_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I260 (c575_r, c575_a, c573_r, c573_a, c574_r, c574_a, initialise);
  BrzJ_l11__280_200_29 I261 (c569_r, c569_a, c571_r, c571_a, c572_r, c572_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I262 (c570_r0d, c570_r1d, c570_a, c571_r, c571_a, c542_r, c542_a, c541_r0d, c541_r1d, c541_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I263 (c568_r0d, c568_r1d, c568_a, c569_r, c569_a, c539_r, c539_a, c538_r0d, c538_r1d, c538_a, initialise);
  BrzM_0_2 I264 (c559_r, c559_a, c566_r, c566_a, c567_r, c567_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I265 (c537_r0d, c537_r1d, c537_a, c558_r, c558_a, c561_r, c561_a, initialise);
  BrzM_0_2 I266 (c562_r, c562_a, c564_r, c564_a, c566_r, c566_a, initialise);
  BrzS_3_l11__280_203_29_l137__28_28_28_280__m63m I267 (c560_r0d, c560_r1d, c560_a, c562_r, c562_a, c565_r, c565_a, initialise);
  BrzF_32_l17__28_280_200_29_29 I268 (c563_r0d, c563_r1d, c563_a, c564_r, c564_a, initialise);
  BrzJ_l19__280_200_200_200_29 I269 (c540_r, c540_a, c543_r, c543_a, c546_r, c546_a, c557_r, c557_a, c559_r, c559_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I270 (c558_r, c558_a, c539_r, c539_a, c542_r, c542_a, c545_r, c545_a, c548_r, c548_a, initialise);
  BrzM_0_2 I271 (c551_r, c551_a, c553_r, c553_a, c557_r, c557_a, initialise);
  BrzS_3_l11__280_203_29_l137__28_28_28_280__m63m I272 (c547_r0d, c547_r1d, c547_a, c549_r, c549_a, c556_r, c556_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I273 (c554_r0d, c554_r1d, c554_a, c555_r, c555_a, c555_r, c555_a, c552_r0d, c552_r1d, c552_a, initialise);
  BrzO_0_32_l24__28_28num_2032_200_29_29 I274 (c549_r, c549_a, c550_r0d, c550_r1d, c550_a);
  BrzM_0_2 I275 (c536_r, c536_a, c521_r, c521_a, c535_r, c535_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I276 (c535_r, c535_a, c531_r, c531_a, c532_r, c532_a, c533_r, c533_a, c534_r, c534_a, initialise);
  BrzJ_l19__280_200_200_200_29 I277 (c523_r, c523_a, c525_r, c525_a, c527_r, c527_a, c529_r, c529_a, c530_r, c530_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I278 (c528_r0d, c528_r1d, c528_a, c529_r, c529_a, c513_r, c513_a, c512_r0d, c512_r1d, c512_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m81m I279 (c526_r0d, c526_r1d, c526_a, c527_r, c527_a, c490_r, c490_a, c504_r, c504_a, c489_r0d, c489_r1d, c489_a, c503_r0d, c503_r1d, c503_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m81m I280 (c524_r0d, c524_r1d, c524_a, c525_r, c525_a, c484_r, c484_a, c498_r, c498_a, c483_r0d, c483_r1d, c483_a, c497_r0d, c497_r1d, c497_a, initialise);
  BrzV_3_l6__28_29_l23__28_28_280_203_29_29__m76m I281 (c522_r0d, c522_r1d, c522_a, c523_r, c523_a, c481_r, c481_a, c516_r, c516_a, c519_r, c519_a, c480_r0d, c480_r1d, c480_a, c515_r0d, c515_r1d, c515_a, c518_r0d, c518_r1d, c518_a, initialise);
  BrzJ_l19__280_200_200_200_29 I282 (c510_r, c510_a, c514_r, c514_a, c517_r, c517_a, c520_r, c520_a, c521_r, c521_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I283 (c530_r, c530_a, c481_r, c481_a, c513_r, c513_a, c516_r, c516_a, c519_r, c519_a, initialise);
  BrzO_32_35_l76__28_28num_203_200_29_20_28a_m51m I284 (c512_r0d, c512_r1d, c512_a, c511_r0d, c511_r1d, c511_a);
  BrzM_0_2 I285 (c495_r, c495_a, c509_r, c509_a, c510_r, c510_a, initialise);
  BrzS_3_l11__280_203_29_l151__28_28_28_281__m65m I286 (c480_r0d, c480_r1d, c480_a, c494_r, c494_a, c508_r, c508_a, initialise);
  BrzJ_l11__280_200_29 I287 (c499_r, c499_a, c507_r, c507_a, c509_r, c509_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I288 (c508_r, c508_a, c498_r, c498_a, c506_r, c506_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I289 (c506_r, c506_a, c501_r, c501_a, c504_r, c504_a, initialise);
  BrzO_33_36_l76__28_28num_203_200_29_20_28a_m54m I290 (c505_r0d, c505_r1d, c505_a, c500_r0d, c500_r1d, c500_a);
  BrzJ_l12__281_2032_29 I291 (c502_r0d, c502_r1d, c502_a, c503_r0d, c503_r1d, c503_a, c505_r0d, c505_r1d, c505_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I292 (c501_r, c501_a, c502_r0d, c502_r1d, c502_a);
  BrzO_32_35_l76__28_28num_203_200_29_20_28a_m51m I293 (c497_r0d, c497_r1d, c497_a, c496_r0d, c496_r1d, c496_a);
  BrzJ_l11__280_200_29 I294 (c485_r, c485_a, c493_r, c493_a, c495_r, c495_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I295 (c494_r, c494_a, c484_r, c484_a, c492_r, c492_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I296 (c492_r, c492_a, c487_r, c487_a, c490_r, c490_a, initialise);
  BrzO_33_36_l91__28_28app_203_20_280_2032_2_m53m I297 (c491_r0d, c491_r1d, c491_a, c486_r0d, c486_r1d, c486_a);
  BrzJ_l12__281_2032_29 I298 (c488_r0d, c488_r1d, c488_a, c489_r0d, c489_r1d, c489_a, c491_r0d, c491_r1d, c491_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I299 (c487_r, c487_a, c488_r0d, c488_r1d, c488_a);
  BrzO_32_35_l91__28_28app_203_20_280_2031_2_m50m I300 (c483_r0d, c483_r1d, c483_a, c482_r0d, c482_r1d, c482_a);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I301 (c454_r0d, c454_r1d, c454_a, c455_r, c455_a, c455_r, c455_a, c458_r0d, c458_r1d, c458_a, initialise);
  BrzV_10_l6__28_29_l45__28_28_280_2010_29_2_m79m I302 (c471_r0d, c471_r1d, c471_a, c468_r0d, c468_r1d, c468_a, c472_r, c472_a, c469_r, c469_a, c465_r, c465_a, c461_r, c461_a, c464_r0d, c464_r1d, c464_a, c460_r0d, c460_r1d, c460_a, initialise);
  BrzV_10_l6__28_29_l24__28_28_280_2010_29_2_m78m I303 (c463_r0d, c463_r1d, c463_a, c466_r, c466_a, c467_r, c467_a, c468_r0d, c468_r1d, c468_a, initialise);
  BrzM_0_2 I304 (c479_r, c479_a, c478_r, c478_a, c453_r, c453_a, initialise);
  BrzM_0_2 I305 (c469_r, c469_a, c477_r, c477_a, c478_r, c478_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I306 (c458_r0d, c458_r1d, c458_a, c459_r, c459_a, c476_r, c476_a, initialise);
  BrzJ_l11__280_200_29 I307 (c472_r, c472_a, c475_r, c475_a, c477_r, c477_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I308 (c476_r, c476_a, c470_r, c470_a, c473_r, c473_a, initialise);
  BrzO_0_1_l23__28_28num_201_201_29_29 I309 (c473_r, c473_a, c474_r0d, c474_r1d, c474_a);
  BrzO_0_10_l26__28_28num_2010_20256_29_29 I310 (c470_r, c470_a, c471_r0d, c471_r1d, c471_a);
  BrzJ_l11__280_200_29 I311 (c462_r, c462_a, c466_r, c466_a, c467_r, c467_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I312 (c459_r, c459_a, c461_r, c461_a, c465_r, c465_a, initialise);
  BrzO_9_10_l75__28_28num_201_200_29_20_28ap_m49m I313 (c464_r0d, c464_r1d, c464_a, c463_r0d, c463_r1d, c463_a);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I314 (c456_r0d, c456_r1d, c456_a, c457_r, c457_a, c457_r, c457_a, c454_r0d, c454_r1d, c454_a, initialise);
  BrzJ_l12__2835_200_29 I315 (c452_r0d, c452_r1d, c452_a, c308_r, c308_a, c301_r0d, c301_r1d, c301_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I316 (c230_r0d, c230_r1d, c230_a, c231_r, c231_a, c452_r0d, c452_r1d, c452_a, initialise);
  BrzJ_l12__2835_200_29 I317 (c451_r0d, c451_r1d, c451_a, c309_r, c309_a, c303_r0d, c303_r1d, c303_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I318 (c235_r0d, c235_r1d, c235_a, c236_r, c236_a, c451_r0d, c451_r1d, c451_a, initialise);
  BrzJ_l11__281_200_29 I319 (c450_r0d, c450_r1d, c450_a, c310_r, c310_a, c305_r0d, c305_r1d, c305_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I320 (c240_r0d, c240_r1d, c240_a, c242_r, c242_a, c450_r0d, c450_r1d, c450_a, initialise);
  BrzV_4_l6__28_29_l43__28_28_280_204_29_29__m77m I321 (c338_r0d, c338_r1d, c338_a, c177_r0d, c177_r1d, c177_a, c340_r, c340_a, c179_r, c179_a, c247_r, c247_a, c244_r, c244_a, c241_r, c241_a, c246_r0d, c246_r1d, c246_a, c243_r0d, c243_r1d, c243_a, c240_r0d, c240_r1d, c240_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m83m I322 (c409_r0d, c409_r1d, c409_a, c410_r, c410_a, c445_r, c445_a, c429_r, c429_a, c421_r, c421_a, c444_r0d, c444_r1d, c444_a, c428_r0d, c428_r1d, c428_a, c420_r0d, c420_r1d, c420_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m81m I323 (c356_r0d, c356_r1d, c356_a, c358_r, c358_a, c424_r, c424_a, c385_r, c385_a, c423_r0d, c423_r1d, c423_a, c384_r0d, c384_r1d, c384_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m90m I324 (c125_r0d, c125_r1d, c125_a, c127_r, c127_a, c250_r, c250_a, c205_r, c205_a, c249_r0d, c249_r1d, c249_a, c204_r0d, c204_r1d, c204_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m90m I325 (c132_r0d, c132_r1d, c132_a, c134_r, c134_a, c253_r, c253_a, c209_r, c209_a, c252_r0d, c252_r1d, c252_a, c208_r0d, c208_r1d, c208_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m90m I326 (c161_r0d, c161_r1d, c161_a, c162_r, c162_a, c256_r, c256_a, c213_r, c213_a, c255_r0d, c255_r1d, c255_a, c212_r0d, c212_r1d, c212_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m90m I327 (c139_r0d, c139_r1d, c139_a, c141_r, c141_a, c259_r, c259_a, c217_r, c217_a, c258_r0d, c258_r1d, c258_a, c216_r0d, c216_r1d, c216_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I328 (c203_r0d, c203_r1d, c203_a, c206_r, c206_a, c271_r, c271_a, c270_r0d, c270_r1d, c270_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I329 (c207_r0d, c207_r1d, c207_a, c210_r, c210_a, c268_r, c268_a, c267_r0d, c267_r1d, c267_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I330 (c211_r0d, c211_r1d, c211_a, c214_r, c214_a, c265_r, c265_a, c264_r0d, c264_r1d, c264_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I331 (c215_r0d, c215_r1d, c215_a, c218_r, c218_a, c262_r, c262_a, c261_r0d, c261_r1d, c261_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m92m I332 (c274_r0d, c274_r1d, c274_a, c276_r, c276_a, c404_r, c404_a, c325_r, c325_a, c322_r, c322_a, c320_r, c320_a, c403_r0d, c403_r1d, c403_a, c324_r0d, c324_r1d, c324_a, c321_r0d, c321_r1d, c321_a, c319_r0d, c319_r1d, c319_a, initialise);
  BrzV_36_l6__28_29_l24__28_28_280_2036_29_2_m96m I333 (c277_r0d, c277_r1d, c277_a, c287_r, c287_a, c351_r, c351_a, c330_r, c330_a, c350_r0d, c350_r1d, c350_a, c329_r0d, c329_r1d, c329_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m86m I334 (c288_r0d, c288_r1d, c288_a, c291_r, c291_a, c399_r, c399_a, c333_r, c333_a, c398_r0d, c398_r1d, c398_a, c332_r0d, c332_r1d, c332_a, initialise);
  BrzV_36_l6__28_29_l24__28_28_280_2036_29_2_m97m I335 (c292_r0d, c292_r1d, c292_a, c299_r, c299_a, c397_r, c397_a, c348_r, c348_a, c339_r, c339_a, c336_r, c336_a, c396_r0d, c396_r1d, c396_a, c347_r0d, c347_r1d, c347_a, c338_r0d, c338_r1d, c338_a, c335_r0d, c335_r1d, c335_a, initialise);
  BrzV_35_l6__28_29_l45__28_28_280_2035_29_2_m94m I336 (c332_r0d, c332_r1d, c332_a, c174_r0d, c174_r1d, c174_a, c334_r, c334_a, c176_r, c176_a, c225_r, c225_a, c224_r0d, c224_r1d, c224_a, initialise);
  BrzV_35_l6__28_29_l45__28_28_280_2035_29_2_m94m I337 (c326_r0d, c326_r1d, c326_a, c181_r0d, c181_r1d, c181_a, c328_r, c328_a, c182_r, c182_a, c228_r, c228_a, c227_r0d, c227_r1d, c227_a, initialise);
  BrzV_36_l6__28_29_l45__28_28_280_2036_29_2_m98m I338 (c329_r0d, c329_r1d, c329_a, c184_r0d, c184_r1d, c184_a, c331_r, c331_a, c185_r, c185_a, c279_r, c279_a, c278_r0d, c278_r1d, c278_a, initialise);
  BrzV_36_l6__28_29_l45__28_28_280_2036_29_2_m98m I339 (c335_r0d, c335_r1d, c335_a, c171_r0d, c171_r1d, c171_a, c337_r, c337_a, c173_r, c173_a, c294_r, c294_a, c293_r0d, c293_r1d, c293_a, initialise);
  BrzV_1_l6__28_29_l43__28_28_280_201_29_29__m74m I340 (c359_r0d, c359_r1d, c359_a, c312_r0d, c312_r1d, c312_a, c361_r, c361_a, c313_r, c313_a, c407_r, c407_a, c318_r, c318_a, c406_r0d, c406_r1d, c406_a, c223_r0d, c223_r1d, c223_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I341 (c119_r0d, c119_r1d, c119_a, c121_r, c121_a, c382_r, c382_a, c383_r0d, c383_r1d, c383_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I342 (c122_r0d, c122_r1d, c122_a, c124_r, c124_a, c427_r, c427_a, c426_r0d, c426_r1d, c426_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m73m I343 (c370_r0d, c370_r1d, c370_a, c372_r, c372_a, c441_r, c441_a, c435_r, c435_a, c388_r, c388_a, c440_r0d, c440_r1d, c440_a, c434_r0d, c434_r1d, c434_a, c387_r0d, c387_r1d, c387_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I344 (c362_r0d, c362_r1d, c362_a, c364_r, c364_a, c391_r, c391_a, c390_r0d, c390_r1d, c390_a, initialise);
  BrzM_0_2 I345 (c449_r, c449_a, c448_r, c448_a, c118_r, c118_a, initialise);
  BrzM_0_2 I346 (c394_r, c394_a, c447_r, c447_a, c448_r, c448_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I347 (c383_r0d, c383_r1d, c383_a, c393_r, c393_a, c395_r, c395_a, initialise);
  BrzJ_l19__280_200_200_200_29 I348 (c422_r, c422_a, c425_r, c425_a, c443_r, c443_a, c446_r, c446_a, c447_r, c447_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I349 (c419_r, c419_a, c421_r, c421_a, c424_r, c424_a, c427_r, c427_a, c445_r, c445_a, initialise);
  BrzM_0_2 I350 (c439_r, c439_a, c442_r, c442_a, c443_r, c443_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I351 (c426_r0d, c426_r1d, c426_a, c438_r, c438_a, c441_r, c441_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I352 (c438_r, c438_a, c429_r, c429_a, c430_r, c430_a, c435_r, c435_a, initialise);
  BrzO_2_1_l119__28_28app_201_20_280_200_201_m47m I353 (c436_r0d, c436_r1d, c436_a, c437_r0d, c437_r1d, c437_a);
  BrzJ_l11__281_201_29 I354 (c433_r0d, c433_r1d, c433_a, c434_r0d, c434_r1d, c434_a, c436_r0d, c436_r1d, c436_a, initialise);
  BrzO_33_1_l196__28_28app_201_20_280_200_20_m52m I355 (c432_r0d, c432_r1d, c432_a, c433_r0d, c433_r1d, c433_a);
  BrzJ_l12__2832_201_29 I356 (c428_r0d, c428_r1d, c428_a, c431_r0d, c431_r1d, c431_a, c432_r0d, c432_r1d, c432_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I357 (c430_r, c430_a, c431_r0d, c431_r1d, c431_a);
  BrzJ_l19__280_200_200_200_29 I358 (c402_r, c402_a, c405_r, c405_a, c408_r, c408_a, c410_r, c410_a, c419_r, c419_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I359 (c395_r, c395_a, c401_r, c401_a, c404_r, c404_a, c407_r, c407_a, c418_r, c418_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I360 (c418_r, c418_a, c416_r, c416_a, c417_r, c417_a, initialise);
  BrzJ_l11__280_200_29 I361 (c412_r, c412_a, c414_r, c414_a, c415_r, c415_a, initialise);
  BrzF_1_l17__28_280_200_29_29 I362 (c413_r0d, c413_r1d, c413_a, c414_r, c414_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I363 (c411_r0d, c411_r1d, c411_a, c412_r, c412_a, c415_r, c415_a, c409_r0d, c409_r1d, c409_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I364 (c401_r, c401_a, c397_r, c397_a, c399_r, c399_a, initialise);
  BrzJ_l12__281_2031_29 I365 (c396_r0d, c396_r1d, c396_a, c398_r0d, c398_r1d, c398_a, c400_r0d, c400_r1d, c400_a, initialise);
  BrzJ_l15__280_200_200_29 I366 (c386_r, c386_a, c389_r, c389_a, c392_r, c392_a, c394_r, c394_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I367 (c393_r, c393_a, c385_r, c385_a, c388_r, c388_a, c391_r, c391_a, initialise);
  BrzJ_l19__280_200_200_200_29 I368 (c349_r, c349_a, c352_r, c352_a, c355_r, c355_a, c373_r, c373_a, c382_r, c382_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I369 (c346_r, c346_a, c348_r, c348_a, c351_r, c351_a, c353_r, c353_a, c381_r, c381_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I370 (c381_r, c381_a, c379_r, c379_a, c380_r, c380_a, initialise);
  BrzJ_l11__280_200_29 I371 (c375_r, c375_a, c377_r, c377_a, c378_r, c378_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I372 (c376_r0d, c376_r1d, c376_a, c377_r, c377_a, c360_r, c360_a, c359_r0d, c359_r1d, c359_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m82m I373 (c374_r0d, c374_r1d, c374_a, c375_r, c375_a, c357_r, c357_a, c363_r, c363_a, c366_r, c366_a, c356_r0d, c356_r1d, c356_a, c362_r0d, c362_r1d, c362_a, c365_r0d, c365_r1d, c365_a, initialise);
  BrzJ_l19__280_200_200_200_29 I374 (c358_r, c358_a, c361_r, c361_a, c364_r, c364_a, c372_r, c372_a, c373_r, c373_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I375 (c378_r, c378_a, c357_r, c357_a, c360_r, c360_a, c363_r, c363_a, c371_r, c371_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I376 (c371_r, c371_a, c366_r, c366_a, c367_r, c367_a, initialise);
  BrzO_33_1_l196__28_28app_201_20_280_200_20_m52m I377 (c369_r0d, c369_r1d, c369_a, c370_r0d, c370_r1d, c370_a);
  BrzJ_l12__2832_201_29 I378 (c365_r0d, c365_r1d, c365_a, c368_r0d, c368_r1d, c368_a, c369_r0d, c369_r1d, c369_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I379 (c367_r, c367_a, c368_r0d, c368_r1d, c368_a);
  BrzO_0_1_l23__28_28num_201_200_29_29 I380 (c353_r, c353_a, c354_r0d, c354_r1d, c354_a);
  BrzM_0_2 I381 (c222_r, c222_a, c345_r, c345_a, c317_r, c317_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I382 (c223_r0d, c223_r1d, c223_a, c346_r, c346_a, c344_r, c344_a, initialise);
  BrzJ_l27__280_200_200_200_200_200_29 I383 (c328_r, c328_a, c331_r, c331_a, c334_r, c334_a, c337_r, c337_a, c340_r, c340_a, c343_r, c343_a, c345_r, c345_a, initialise);
  BrzF_0_l87__28_280_200_29_20_280_200_29_20_m36m I384 (c344_r, c344_a, c327_r, c327_a, c330_r, c330_a, c333_r, c333_a, c336_r, c336_a, c339_r, c339_a, c341_r, c341_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I385 (c341_r, c341_a, c342_r0d, c342_r1d, c342_a);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I386 (c327_r, c327_a, c320_r, c320_a, c322_r, c322_a, c325_r, c325_a, initialise);
  BrzJ_l12__2834_201_29 I387 (c323_r0d, c323_r1d, c323_a, c324_r0d, c324_r1d, c324_a, c326_r0d, c326_r1d, c326_a, initialise);
  BrzJ_l12__2833_201_29 I388 (c319_r0d, c319_r1d, c319_a, c321_r0d, c321_r1d, c321_a, c323_r0d, c323_r1d, c323_a, initialise);
  BrzJ_l35__280_200_200_200_200_200_200_200__m45m I389 (c226_r, c226_a, c229_r, c229_a, c231_r, c231_a, c236_r, c236_a, c242_r, c242_a, c273_r, c273_a, c300_r, c300_a, c313_r, c313_a, c318_r, c318_a, initialise);
  BrzF_0_l115__28_280_200_29_20_280_200_29_2_m38m I390 (c317_r, c317_a, c225_r, c225_a, c228_r, c228_a, c234_r, c234_a, c239_r, c239_a, c241_r, c241_a, c244_r, c244_a, c311_r, c311_a, c316_r, c316_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I391 (c314_r0d, c314_r1d, c314_a, c315_r, c315_a, c315_r, c315_a, c312_r0d, c312_r1d, c312_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I392 (c311_r, c311_a, c308_r, c308_a, c309_r, c309_a, c310_r, c310_a, initialise);
  BrzJ_l15__280_200_200_29 I393 (c302_r, c302_a, c304_r, c304_a, c306_r, c306_a, c307_r, c307_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I394 (c305_r0d, c305_r1d, c305_a, c306_r, c306_a, c281_r, c281_a, c280_r0d, c280_r1d, c280_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m88m I395 (c303_r0d, c303_r1d, c303_a, c304_r, c304_a, c275_r, c275_a, c284_r, c284_a, c274_r0d, c274_r1d, c274_a, c283_r0d, c283_r1d, c283_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m93m I396 (c301_r0d, c301_r1d, c301_a, c302_r, c302_a, c290_r, c290_a, c296_r, c296_a, c289_r0d, c289_r1d, c289_a, c295_r0d, c295_r1d, c295_a, initialise);
  BrzJ_l19__280_200_200_200_29 I397 (c276_r, c276_a, c287_r, c287_a, c291_r, c291_a, c299_r, c299_a, c300_r, c300_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I398 (c307_r, c307_a, c275_r, c275_a, c286_r, c286_a, c290_r, c290_a, c298_r, c298_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I399 (c298_r, c298_a, c294_r, c294_a, c296_r, c296_a, initialise);
  BrzO_35_36_l76__28_28num_201_200_29_20_28a_m56m I400 (c297_r0d, c297_r1d, c297_a, c292_r0d, c292_r1d, c292_a);
  BrzJ_l12__2832_203_29 I401 (c293_r0d, c293_r1d, c293_a, c295_r0d, c295_r1d, c295_a, c297_r0d, c297_r1d, c297_a, initialise);
  BrzO_32_35_l91__28_28app_203_20_280_2031_2_m50m I402 (c289_r0d, c289_r1d, c289_a, c288_r0d, c288_r1d, c288_a);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I403 (c286_r, c286_a, c279_r, c279_a, c281_r, c281_a, c284_r, c284_a, initialise);
  BrzO_35_36_l76__28_28num_201_200_29_20_28a_m56m I404 (c285_r0d, c285_r1d, c285_a, c277_r0d, c277_r1d, c277_a);
  BrzJ_l12__2833_202_29 I405 (c282_r0d, c282_r1d, c282_a, c283_r0d, c283_r1d, c283_a, c285_r0d, c285_r1d, c285_a, initialise);
  BrzJ_l12__2832_201_29 I406 (c278_r0d, c278_r1d, c278_a, c280_r0d, c280_r1d, c280_a, c282_r0d, c282_r1d, c282_a, initialise);
  BrzM_0_9 I407 (c248_r, c248_a, c251_r, c251_a, c254_r, c254_a, c257_r, c257_a, c260_r, c260_a, c263_r, c263_a, c266_r, c266_a, c269_r, c269_a, c272_r, c272_a, c273_r, c273_a, initialise);
  BrzS_4_l11__280_204_29_l521__28_28_28_280__m66m I408 (c243_r0d, c243_r1d, c243_a, c247_r, c247_a, c250_r, c250_a, c253_r, c253_a, c256_r, c256_a, c259_r, c259_a, c262_r, c262_a, c265_r, c265_a, c268_r, c268_a, c271_r, c271_a, initialise);
  BrzO_4_35_l91__28_28app_2031_20_280_203_20_m48m I409 (c246_r0d, c246_r1d, c246_a, c245_r0d, c245_r1d, c245_a);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I410 (c237_r0d, c237_r1d, c237_a, c238_r, c238_a, c238_r, c238_a, c235_r0d, c235_r1d, c235_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I411 (c232_r0d, c232_r1d, c232_a, c233_r, c233_a, c233_r, c233_a, c230_r0d, c230_r1d, c230_a, initialise);
  BrzJ_l23__280_200_200_200_200_29 I412 (c206_r, c206_a, c210_r, c210_a, c214_r, c214_a, c218_r, c218_a, c221_r, c221_a, c222_r, c222_a, initialise);
  BrzF_0_l73__28_280_200_29_20_280_200_29_20_m35m I413 (c186_r, c186_a, c205_r, c205_a, c209_r, c209_a, c213_r, c213_a, c217_r, c217_a, c219_r, c219_a, initialise);
  BrzO_0_1_l23__28_28num_201_201_29_29 I414 (c219_r, c219_a, c220_r0d, c220_r1d, c220_a);
  BrzO_35_35_l34__28_28not_20_280_200_2035_2_m55m I415 (c216_r0d, c216_r1d, c216_a, c215_r0d, c215_r1d, c215_a);
  BrzO_35_35_l34__28_28not_20_280_200_2035_2_m55m I416 (c212_r0d, c212_r1d, c212_a, c211_r0d, c211_r1d, c211_a);
  BrzO_35_35_l34__28_28not_20_280_200_2035_2_m55m I417 (c208_r0d, c208_r1d, c208_a, c207_r0d, c207_r1d, c207_a);
  BrzO_35_35_l34__28_28not_20_280_200_2035_2_m55m I418 (c204_r0d, c204_r1d, c204_a, c203_r0d, c203_r1d, c203_a);
  BrzF_0_l73__28_280_200_29_20_280_200_29_20_m35m I419 (c118_r, c118_a, c198_r, c198_a, c199_r, c199_a, c200_r, c200_a, c201_r, c201_a, c202_r, c202_a, initialise);
  BrzJ_l23__280_200_200_200_200_29 I420 (c188_r, c188_a, c190_r, c190_a, c192_r, c192_a, c194_r, c194_a, c196_r, c196_a, c197_r, c197_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I421 (c195_r0d, c195_r1d, c195_a, c196_r, c196_a, c123_r, c123_a, c122_r0d, c122_r1d, c122_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I422 (c193_r0d, c193_r1d, c193_a, c194_r, c194_a, c120_r, c120_a, c119_r0d, c119_r1d, c119_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I423 (c191_r0d, c191_r1d, c191_a, c192_r, c192_a, c175_r, c175_a, c174_r0d, c174_r1d, c174_a, initialise);
  BrzV_36_l6__28_29_l24__28_28_280_2036_29_2_m95m I424 (c189_r0d, c189_r1d, c189_a, c190_r, c190_a, c172_r, c172_a, c178_r, c178_a, c171_r0d, c171_r1d, c171_a, c177_r0d, c177_r1d, c177_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m89m I425 (c187_r0d, c187_r1d, c187_a, c188_r, c188_a, c126_r, c126_a, c131_r, c131_a, c138_r, c138_a, c143_r, c143_a, c146_r, c146_a, c152_r, c152_a, c160_r, c160_a, c125_r0d, c125_r1d, c125_a, c130_r0d, c130_r1d, c130_a, c137_r0d, c137_r1d, c137_a, c142_r0d, c142_r1d, c142_a, c145_r0d, c145_r1d, c145_a, c151_r0d, c151_r1d, c151_a, c159_r0d, c159_r1d, c159_a, initialise);
  BrzJ_l59__280_200_200_200_200_200_200_200__m46m I426 (c121_r, c121_a, c124_r, c124_a, c127_r, c127_a, c134_r, c134_a, c141_r, c141_a, c144_r, c144_a, c147_r, c147_a, c150_r, c150_a, c162_r, c162_a, c173_r, c173_a, c176_r, c176_a, c179_r, c179_a, c182_r, c182_a, c185_r, c185_a, c186_r, c186_a, initialise);
  BrzF_0_l199__28_280_200_29_20_280_200_29_2_m39m I427 (c197_r, c197_a, c120_r, c120_a, c123_r, c123_a, c126_r, c126_a, c133_r, c133_a, c140_r, c140_a, c143_r, c143_a, c146_r, c146_a, c148_r, c148_a, c170_r, c170_a, c172_r, c172_a, c175_r, c175_a, c178_r, c178_a, c180_r, c180_a, c183_r, c183_a, initialise);
  BrzO_0_36_l24__28_28num_2036_200_29_29 I428 (c183_r, c183_a, c184_r0d, c184_r1d, c184_a);
  BrzO_0_35_l24__28_28num_2035_200_29_29 I429 (c180_r, c180_a, c181_r0d, c181_r1d, c181_a);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I430 (c170_r, c170_a, c168_r, c168_a, c169_r, c169_a, initialise);
  BrzJ_l11__280_200_29 I431 (c164_r, c164_a, c166_r, c166_a, c167_r, c167_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I432 (c165_r0d, c165_r1d, c165_a, c166_r, c166_a, c157_r, c157_a, c156_r0d, c156_r1d, c156_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I433 (c163_r0d, c163_r1d, c163_a, c164_r, c164_a, c154_r, c154_a, c153_r0d, c153_r1d, c153_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I434 (c167_r, c167_a, c152_r, c152_a, c154_r, c154_a, c157_r, c157_a, c160_r, c160_a, initialise);
  BrzJ_l12__2834_201_29 I435 (c158_r0d, c158_r1d, c158_a, c159_r0d, c159_r1d, c159_a, c161_r0d, c161_r1d, c161_a, initialise);
  BrzJ_l12__2833_201_29 I436 (c155_r0d, c155_r1d, c155_a, c156_r0d, c156_r1d, c156_a, c158_r0d, c158_r1d, c158_a, initialise);
  BrzJ_l12__281_2032_29 I437 (c151_r0d, c151_r1d, c151_a, c153_r0d, c153_r1d, c153_a, c155_r0d, c155_r1d, c155_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I438 (c148_r, c148_a, c149_r0d, c149_r1d, c149_a);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I439 (c140_r, c140_a, c135_r, c135_a, c138_r, c138_a, initialise);
  BrzJ_l12__282_2033_29 I440 (c136_r0d, c136_r1d, c136_a, c137_r0d, c137_r1d, c137_a, c139_r0d, c139_r1d, c139_a, initialise);
  BrzO_0_2_l23__28_28num_202_200_29_29 I441 (c135_r, c135_a, c136_r0d, c136_r1d, c136_a);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I442 (c133_r, c133_a, c128_r, c128_a, c131_r, c131_a, initialise);
  BrzJ_l12__281_2034_29 I443 (c129_r0d, c129_r1d, c129_a, c130_r0d, c130_r1d, c130_a, c132_r0d, c132_r1d, c132_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I444 (c128_r, c128_a, c129_r0d, c129_r1d, c129_a);
  BrzJ_l12__2833_200_29 I445 (c117_r0d, c117_r1d, c117_a, c99_r, c99_a, c94_r0d, c94_r1d, c94_a, initialise);
  BrzF_33_l32__28_280_200_29_20_280_2033_29__m41m I446 (c65_r0d, c65_r1d, c65_a, c67_r, c67_a, c117_r0d, c117_r1d, c117_a, initialise);
  BrzJ_l12__2833_200_29 I447 (c116_r0d, c116_r1d, c116_a, c100_r, c100_a, c96_r0d, c96_r1d, c96_a, initialise);
  BrzF_33_l32__28_280_200_29_20_280_2033_29__m41m I448 (c72_r0d, c72_r1d, c72_a, c74_r, c74_a, c116_r0d, c116_r1d, c116_a, initialise);
  BrzJ_l12__2834_200_29 I449 (c115_r0d, c115_r1d, c115_a, c111_r, c111_a, c109_r0d, c109_r1d, c109_a, initialise);
  BrzF_34_l32__28_280_200_29_20_280_2034_29__m42m I450 (c92_r0d, c92_r1d, c92_a, c93_r, c93_a, c115_r0d, c115_r1d, c115_a, initialise);
  BrzM_0_2 I451 (c114_r, c114_a, c113_r, c113_a, c112_r, c112_a, initialise);
  BrzJ_l15__280_200_200_29 I452 (c75_r, c75_a, c93_r, c93_a, c108_r, c108_a, c113_r, c113_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I453 (c112_r, c112_a, c86_r, c86_a, c101_r, c101_a, c111_r, c111_a, initialise);
  BrzV_34_l6__28_29_l24__28_28_280_2034_29_2_m85m I454 (c109_r0d, c109_r1d, c109_a, c110_r, c110_a, c103_r, c103_a, c106_r, c106_a, c102_r0d, c102_r1d, c102_a, c105_r0d, c105_r1d, c105_a, initialise);
  BrzJ_l11__280_200_29 I455 (c104_r, c104_a, c107_r, c107_a, c108_r, c108_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I456 (c110_r, c110_a, c103_r, c103_a, c106_r, c106_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I457 (c101_r, c101_a, c99_r, c99_a, c100_r, c100_a, initialise);
  BrzJ_l11__280_200_29 I458 (c95_r, c95_a, c97_r, c97_a, c98_r, c98_a, initialise);
  BrzV_33_l6__28_29_l24__28_28_280_2033_29_2_m84m I459 (c96_r0d, c96_r1d, c96_a, c97_r, c97_a, c90_r, c90_a, c89_r0d, c89_r1d, c89_a, initialise);
  BrzV_33_l6__28_29_l24__28_28_280_2033_29_2_m84m I460 (c94_r0d, c94_r1d, c94_a, c95_r, c95_a, c88_r, c88_a, c87_r0d, c87_r1d, c87_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I461 (c98_r, c98_a, c88_r, c88_a, c90_r, c90_a, initialise);
  BrzO_66_34_l270__28_28app_201_20_280_200_2_m57m I462 (c91_r0d, c91_r1d, c91_a, c92_r0d, c92_r1d, c92_a);
  BrzJ_l13__2833_2033_29 I463 (c87_r0d, c87_r1d, c87_a, c89_r0d, c89_r1d, c89_a, c91_r0d, c91_r1d, c91_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I464 (c86_r, c86_a, c83_r, c83_a, c84_r, c84_a, c85_r, c85_a, initialise);
  BrzJ_l15__280_200_200_29 I465 (c77_r, c77_a, c79_r, c79_a, c81_r, c81_a, c82_r, c82_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m72m I466 (c80_r0d, c80_r1d, c80_a, c81_r, c81_a, c62_r, c62_a, c69_r, c69_a, c61_r0d, c61_r1d, c61_a, c68_r0d, c68_r1d, c68_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I467 (c78_r0d, c78_r1d, c78_a, c79_r, c79_a, c71_r, c71_a, c70_r0d, c70_r1d, c70_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I468 (c76_r0d, c76_r1d, c76_a, c77_r, c77_a, c64_r, c64_a, c63_r0d, c63_r1d, c63_a, initialise);
  BrzJ_l11__280_200_29 I469 (c67_r, c67_a, c74_r, c74_a, c75_r, c75_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I470 (c82_r, c82_a, c66_r, c66_a, c73_r, c73_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I471 (c73_r, c73_a, c69_r, c69_a, c71_r, c71_a, initialise);
  BrzJ_l12__281_2032_29 I472 (c68_r0d, c68_r1d, c68_a, c70_r0d, c70_r1d, c70_a, c72_r0d, c72_r1d, c72_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I473 (c66_r, c66_a, c62_r, c62_a, c64_r, c64_a, initialise);
  BrzJ_l12__281_2032_29 I474 (c61_r0d, c61_r1d, c61_a, c63_r0d, c63_r1d, c63_a, c65_r0d, c65_r1d, c65_a, initialise);
  BrzM_0_2 I475 (c60_r, c60_a, c48_r, c48_a, c59_r, c59_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I476 (c59_r, c59_a, c56_r, c56_a, c57_r, c57_a, c58_r, c58_a, initialise);
  BrzJ_l15__280_200_200_29 I477 (c50_r, c50_a, c52_r, c52_a, c54_r, c54_a, c55_r, c55_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m91m I478 (c53_r0d, c53_r1d, c53_a, c54_r, c54_a, c19_r, c19_a, c31_r, c31_a, c39_r, c39_a, c18_r0d, c18_r1d, c18_a, c30_r0d, c30_r1d, c30_a, c38_r0d, c38_r1d, c38_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m91m I479 (c51_r0d, c51_r1d, c51_a, c52_r, c52_a, c15_r, c15_a, c27_r, c27_a, c41_r, c41_a, c14_r0d, c14_r1d, c14_a, c26_r0d, c26_r1d, c26_a, c40_r0d, c40_r1d, c40_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m91m I480 (c49_r0d, c49_r1d, c49_a, c50_r, c50_a, c13_r, c13_a, c25_r, c25_a, c33_r, c33_a, c12_r0d, c12_r1d, c12_a, c24_r0d, c24_r1d, c24_a, c32_r0d, c32_r1d, c32_a, initialise);
  BrzJ_l11__280_200_29 I481 (c23_r, c23_a, c47_r, c47_a, c48_r, c48_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I482 (c55_r, c55_a, c22_r, c22_a, c46_r, c46_a, initialise);
  BrzF_0_l87__28_280_200_29_20_280_200_29_20_m36m I483 (c46_r, c46_a, c25_r, c25_a, c27_r, c27_a, c31_r, c31_a, c33_r, c33_a, c39_r, c39_a, c41_r, c41_a, initialise);
  BrzO_70_35_l123__28_28app_201_20_280_200_2_m59m I484 (c44_r0d, c44_r1d, c44_a, c45_r0d, c45_r1d, c45_a);
  BrzJ_l13__2835_2035_29 I485 (c37_r0d, c37_r1d, c37_a, c43_r0d, c43_r1d, c43_a, c44_r0d, c44_r1d, c44_a, initialise);
  BrzO_70_35_l124__28_28app_201_20_280_200_2_m58m I486 (c42_r0d, c42_r1d, c42_a, c43_r0d, c43_r1d, c43_a);
  BrzJ_l13__2835_2035_29 I487 (c38_r0d, c38_r1d, c38_a, c40_r0d, c40_r1d, c40_a, c42_r0d, c42_r1d, c42_a, initialise);
  BrzO_70_35_l123__28_28app_201_20_280_200_2_m59m I488 (c36_r0d, c36_r1d, c36_a, c37_r0d, c37_r1d, c37_a);
  BrzJ_l13__2835_2035_29 I489 (c29_r0d, c29_r1d, c29_a, c35_r0d, c35_r1d, c35_a, c36_r0d, c36_r1d, c36_a, initialise);
  BrzO_70_35_l124__28_28app_201_20_280_200_2_m58m I490 (c34_r0d, c34_r1d, c34_a, c35_r0d, c35_r1d, c35_a);
  BrzJ_l13__2835_2035_29 I491 (c30_r0d, c30_r1d, c30_a, c32_r0d, c32_r1d, c32_a, c34_r0d, c34_r1d, c34_a, initialise);
  BrzO_70_35_l124__28_28app_201_20_280_200_2_m58m I492 (c28_r0d, c28_r1d, c28_a, c29_r0d, c29_r1d, c29_a);
  BrzJ_l13__2835_2035_29 I493 (c24_r0d, c24_r1d, c24_a, c26_r0d, c26_r1d, c26_a, c28_r0d, c28_r1d, c28_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I494 (c22_r, c22_a, c13_r, c13_a, c15_r, c15_a, c19_r, c19_a, initialise);
  BrzO_70_35_l124__28_28app_201_20_280_200_2_m60m I495 (c20_r0d, c20_r1d, c20_a, c21_r0d, c21_r1d, c21_a);
  BrzJ_l13__2835_2035_29 I496 (c17_r0d, c17_r1d, c17_a, c18_r0d, c18_r1d, c18_a, c20_r0d, c20_r1d, c20_a, initialise);
  BrzO_70_35_l124__28_28app_201_20_280_200_2_m60m I497 (c16_r0d, c16_r1d, c16_a, c17_r0d, c17_r1d, c17_a);
  BrzJ_l13__2835_2035_29 I498 (c12_r0d, c12_r1d, c12_a, c14_r0d, c14_r1d, c14_a, c16_r0d, c16_r1d, c16_a, initialise);
endmodule

module Balsa_nmult (
  go_0r, go_0a,
  bypass_0r0d, bypass_0r1d, bypass_0a,
  bypassH_0r0d, bypassH_0r1d, bypassH_0a,
  mType_0r0d, mType_0r1d, mType_0a,
  a_0r0d, a_0r1d, a_0a,
  b_0r0d, b_0r1d, b_0a,
  c_0r0d, c_0r1d, c_0a,
  mpH_0r0d, mpH_0r1d, mpH_0a,
  mpL_0r0d, mpL_0r1d, mpL_0a,
  mZ_0r0d, mZ_0r1d, mZ_0a,
  mN_0r0d, mN_0r1d, mN_0a,
  initialise
);
  input go_0r;
  output go_0a;
  input bypass_0r0d;
  input bypass_0r1d;
  output bypass_0a;
  input bypassH_0r0d;
  input bypassH_0r1d;
  output bypassH_0a;
  input [2:0] mType_0r0d;
  input [2:0] mType_0r1d;
  output mType_0a;
  input [31:0] a_0r0d;
  input [31:0] a_0r1d;
  output a_0a;
  input [31:0] b_0r0d;
  input [31:0] b_0r1d;
  output b_0a;
  input [31:0] c_0r0d;
  input [31:0] c_0r1d;
  output c_0a;
  output [31:0] mpH_0r0d;
  output [31:0] mpH_0r1d;
  input mpH_0a;
  output [31:0] mpL_0r0d;
  output [31:0] mpL_0r1d;
  input mpL_0a;
  output mZ_0r0d;
  output mZ_0r1d;
  input mZ_0a;
  output mN_0r0d;
  output mN_0r1d;
  input mN_0a;
  input initialise;
  wire [1:0] c883_r0d;
  wire [1:0] c883_r1d;
  wire c883_a;
  wire [1:0] c882_r0d;
  wire [1:0] c882_r1d;
  wire c882_a;
  wire [1:0] c881_r0d;
  wire [1:0] c881_r1d;
  wire c881_a;
  wire [1:0] c880_r0d;
  wire [1:0] c880_r1d;
  wire c880_a;
  wire c879_r;
  wire c879_a;
  wire c878_r0d;
  wire c878_r1d;
  wire c878_a;
  wire c877_r0d;
  wire c877_r1d;
  wire c877_a;
  wire c876_r;
  wire c876_a;
  wire c875_r0d;
  wire c875_r1d;
  wire c875_a;
  wire c874_r;
  wire c874_a;
  wire [1:0] c873_r0d;
  wire [1:0] c873_r1d;
  wire c873_a;
  wire [1:0] c872_r0d;
  wire [1:0] c872_r1d;
  wire c872_a;
  wire [1:0] c871_r0d;
  wire [1:0] c871_r1d;
  wire c871_a;
  wire [1:0] c870_r0d;
  wire [1:0] c870_r1d;
  wire c870_a;
  wire c869_r;
  wire c869_a;
  wire c868_r0d;
  wire c868_r1d;
  wire c868_a;
  wire c867_r0d;
  wire c867_r1d;
  wire c867_a;
  wire c866_r;
  wire c866_a;
  wire c865_r0d;
  wire c865_r1d;
  wire c865_a;
  wire c864_r;
  wire c864_a;
  wire [1:0] c863_r0d;
  wire [1:0] c863_r1d;
  wire c863_a;
  wire [1:0] c862_r0d;
  wire [1:0] c862_r1d;
  wire c862_a;
  wire [1:0] c861_r0d;
  wire [1:0] c861_r1d;
  wire c861_a;
  wire [1:0] c860_r0d;
  wire [1:0] c860_r1d;
  wire c860_a;
  wire c859_r;
  wire c859_a;
  wire [31:0] c858_r0d;
  wire [31:0] c858_r1d;
  wire c858_a;
  wire [31:0] c857_r0d;
  wire [31:0] c857_r1d;
  wire c857_a;
  wire c856_r;
  wire c856_a;
  wire [31:0] c855_r0d;
  wire [31:0] c855_r1d;
  wire c855_a;
  wire c854_r;
  wire c854_a;
  wire [1:0] c853_r0d;
  wire [1:0] c853_r1d;
  wire c853_a;
  wire [1:0] c852_r0d;
  wire [1:0] c852_r1d;
  wire c852_a;
  wire [1:0] c851_r0d;
  wire [1:0] c851_r1d;
  wire c851_a;
  wire [1:0] c850_r0d;
  wire [1:0] c850_r1d;
  wire c850_a;
  wire c849_r;
  wire c849_a;
  wire [31:0] c848_r0d;
  wire [31:0] c848_r1d;
  wire c848_a;
  wire [31:0] c847_r0d;
  wire [31:0] c847_r1d;
  wire c847_a;
  wire c846_r;
  wire c846_a;
  wire [31:0] c845_r0d;
  wire [31:0] c845_r1d;
  wire c845_a;
  wire c844_r;
  wire c844_a;
  wire [33:0] c843_r0d;
  wire [33:0] c843_r1d;
  wire c843_a;
  wire [1:0] c842_r0d;
  wire [1:0] c842_r1d;
  wire c842_a;
  wire [1:0] c841_r0d;
  wire [1:0] c841_r1d;
  wire c841_a;
  wire [1:0] c840_r0d;
  wire [1:0] c840_r1d;
  wire c840_a;
  wire [1:0] c839_r0d;
  wire [1:0] c839_r1d;
  wire c839_a;
  wire [1:0] c838_r0d;
  wire [1:0] c838_r1d;
  wire c838_a;
  wire [1:0] c837_r0d;
  wire [1:0] c837_r1d;
  wire c837_a;
  wire [1:0] c836_r0d;
  wire [1:0] c836_r1d;
  wire c836_a;
  wire [34:0] c835_r0d;
  wire [34:0] c835_r1d;
  wire c835_a;
  wire c834_r;
  wire c834_a;
  wire [34:0] c833_r0d;
  wire [34:0] c833_r1d;
  wire c833_a;
  wire [34:0] c832_r0d;
  wire [34:0] c832_r1d;
  wire c832_a;
  wire c831_r;
  wire c831_a;
  wire [34:0] c830_r0d;
  wire [34:0] c830_r1d;
  wire c830_a;
  wire c829_r;
  wire c829_a;
  wire [1:0] c828_r0d;
  wire [1:0] c828_r1d;
  wire c828_a;
  wire [1:0] c827_r0d;
  wire [1:0] c827_r1d;
  wire c827_a;
  wire [1:0] c826_r0d;
  wire [1:0] c826_r1d;
  wire c826_a;
  wire [1:0] c825_r0d;
  wire [1:0] c825_r1d;
  wire c825_a;
  wire [35:0] c824_r0d;
  wire [35:0] c824_r1d;
  wire c824_a;
  wire c823_r;
  wire c823_a;
  wire [35:0] c822_r0d;
  wire [35:0] c822_r1d;
  wire c822_a;
  wire [35:0] c821_r0d;
  wire [35:0] c821_r1d;
  wire c821_a;
  wire c820_r;
  wire c820_a;
  wire [35:0] c819_r0d;
  wire [35:0] c819_r1d;
  wire c819_a;
  wire c818_r;
  wire c818_a;
  wire [34:0] c817_r0d;
  wire [34:0] c817_r1d;
  wire c817_a;
  wire c816_r0d;
  wire c816_r1d;
  wire c816_a;
  wire c815_r0d;
  wire c815_r1d;
  wire c815_a;
  wire [31:0] c814_r0d;
  wire [31:0] c814_r1d;
  wire c814_a;
  wire [31:0] c813_r0d;
  wire [31:0] c813_r1d;
  wire c813_a;
  wire [1:0] c812_r0d;
  wire [1:0] c812_r1d;
  wire c812_a;
  wire [1:0] c811_r0d;
  wire [1:0] c811_r1d;
  wire c811_a;
  wire [1:0] c810_r0d;
  wire [1:0] c810_r1d;
  wire c810_a;
  wire [1:0] c809_r0d;
  wire [1:0] c809_r1d;
  wire c809_a;
  wire [31:0] c808_r0d;
  wire [31:0] c808_r1d;
  wire c808_a;
  wire c807_r;
  wire c807_a;
  wire [31:0] c806_r0d;
  wire [31:0] c806_r1d;
  wire c806_a;
  wire [31:0] c805_r0d;
  wire [31:0] c805_r1d;
  wire c805_a;
  wire c804_r;
  wire c804_a;
  wire [31:0] c803_r0d;
  wire [31:0] c803_r1d;
  wire c803_a;
  wire c802_r;
  wire c802_a;
  wire [2:0] c801_r0d;
  wire [2:0] c801_r1d;
  wire c801_a;
  wire [34:0] c800_r0d;
  wire [34:0] c800_r1d;
  wire c800_a;
  wire [8:0] c799_r0d;
  wire [8:0] c799_r1d;
  wire c799_a;
  wire [8:0] c798_r0d;
  wire [8:0] c798_r1d;
  wire c798_a;
  wire [8:0] c797_r0d;
  wire [8:0] c797_r1d;
  wire c797_a;
  wire [8:0] c796_r0d;
  wire [8:0] c796_r1d;
  wire c796_a;
  wire [8:0] c795_r0d;
  wire [8:0] c795_r1d;
  wire c795_a;
  wire [8:0] c794_r0d;
  wire [8:0] c794_r1d;
  wire c794_a;
  wire [8:0] c793_r0d;
  wire [8:0] c793_r1d;
  wire c793_a;
  wire [8:0] c792_r0d;
  wire [8:0] c792_r1d;
  wire c792_a;
  wire [8:0] c791_r0d;
  wire [8:0] c791_r1d;
  wire c791_a;
  wire [8:0] c790_r0d;
  wire [8:0] c790_r1d;
  wire c790_a;
  wire [8:0] c789_r0d;
  wire [8:0] c789_r1d;
  wire c789_a;
  wire [34:0] c788_r0d;
  wire [34:0] c788_r1d;
  wire c788_a;
  wire c787_r;
  wire c787_a;
  wire [34:0] c786_r0d;
  wire [34:0] c786_r1d;
  wire c786_a;
  wire [34:0] c785_r0d;
  wire [34:0] c785_r1d;
  wire c785_a;
  wire c784_r;
  wire c784_a;
  wire [34:0] c783_r0d;
  wire [34:0] c783_r1d;
  wire c783_a;
  wire c782_r;
  wire c782_a;
  wire [34:0] c781_r0d;
  wire [34:0] c781_r1d;
  wire c781_a;
  wire c780_r;
  wire c780_a;
  wire [34:0] c779_r0d;
  wire [34:0] c779_r1d;
  wire c779_a;
  wire c778_r;
  wire c778_a;
  wire [34:0] c777_r0d;
  wire [34:0] c777_r1d;
  wire c777_a;
  wire c776_r;
  wire c776_a;
  wire [34:0] c775_r0d;
  wire [34:0] c775_r1d;
  wire c775_a;
  wire c774_r;
  wire c774_a;
  wire [34:0] c773_r0d;
  wire [34:0] c773_r1d;
  wire c773_a;
  wire c772_r;
  wire c772_a;
  wire [34:0] c771_r0d;
  wire [34:0] c771_r1d;
  wire c771_a;
  wire c770_r;
  wire c770_a;
  wire [34:0] c769_r0d;
  wire [34:0] c769_r1d;
  wire c769_a;
  wire c768_r;
  wire c768_a;
  wire [34:0] c767_r0d;
  wire [34:0] c767_r1d;
  wire c767_a;
  wire [34:0] c766_r0d;
  wire [34:0] c766_r1d;
  wire c766_a;
  wire [34:0] c765_r0d;
  wire [34:0] c765_r1d;
  wire c765_a;
  wire [2:0] c764_r0d;
  wire [2:0] c764_r1d;
  wire c764_a;
  wire [2:0] c763_r0d;
  wire [2:0] c763_r1d;
  wire c763_a;
  wire [2:0] c762_r0d;
  wire [2:0] c762_r1d;
  wire c762_a;
  wire [2:0] c761_r0d;
  wire [2:0] c761_r1d;
  wire c761_a;
  wire [2:0] c760_r0d;
  wire [2:0] c760_r1d;
  wire c760_a;
  wire [31:0] c759_r0d;
  wire [31:0] c759_r1d;
  wire c759_a;
  wire c758_r;
  wire c758_a;
  wire [31:0] c757_r0d;
  wire [31:0] c757_r1d;
  wire c757_a;
  wire [31:0] c756_r0d;
  wire [31:0] c756_r1d;
  wire c756_a;
  wire c755_r;
  wire c755_a;
  wire [31:0] c754_r0d;
  wire [31:0] c754_r1d;
  wire c754_a;
  wire c753_r;
  wire c753_a;
  wire [31:0] c752_r0d;
  wire [31:0] c752_r1d;
  wire c752_a;
  wire c751_r;
  wire c751_a;
  wire [2:0] c750_r0d;
  wire [2:0] c750_r1d;
  wire c750_a;
  wire [2:0] c749_r0d;
  wire [2:0] c749_r1d;
  wire c749_a;
  wire [2:0] c748_r0d;
  wire [2:0] c748_r1d;
  wire c748_a;
  wire [2:0] c747_r0d;
  wire [2:0] c747_r1d;
  wire c747_a;
  wire [2:0] c746_r0d;
  wire [2:0] c746_r1d;
  wire c746_a;
  wire [31:0] c745_r0d;
  wire [31:0] c745_r1d;
  wire c745_a;
  wire c744_r;
  wire c744_a;
  wire [31:0] c743_r0d;
  wire [31:0] c743_r1d;
  wire c743_a;
  wire [31:0] c742_r0d;
  wire [31:0] c742_r1d;
  wire c742_a;
  wire c741_r;
  wire c741_a;
  wire [31:0] c740_r0d;
  wire [31:0] c740_r1d;
  wire c740_a;
  wire c739_r;
  wire c739_a;
  wire [31:0] c738_r0d;
  wire [31:0] c738_r1d;
  wire c738_a;
  wire c737_r;
  wire c737_a;
  wire [2:0] c736_r0d;
  wire [2:0] c736_r1d;
  wire c736_a;
  wire [2:0] c735_r0d;
  wire [2:0] c735_r1d;
  wire c735_a;
  wire [2:0] c734_r0d;
  wire [2:0] c734_r1d;
  wire c734_a;
  wire [2:0] c733_r0d;
  wire [2:0] c733_r1d;
  wire c733_a;
  wire [2:0] c732_r0d;
  wire [2:0] c732_r1d;
  wire c732_a;
  wire c731_r0d;
  wire c731_r1d;
  wire c731_a;
  wire c730_r;
  wire c730_a;
  wire c729_r0d;
  wire c729_r1d;
  wire c729_a;
  wire c728_r0d;
  wire c728_r1d;
  wire c728_a;
  wire c727_r;
  wire c727_a;
  wire c726_r0d;
  wire c726_r1d;
  wire c726_a;
  wire c725_r;
  wire c725_a;
  wire c724_r0d;
  wire c724_r1d;
  wire c724_a;
  wire c723_r;
  wire c723_a;
  wire [34:0] c722_r0d;
  wire [34:0] c722_r1d;
  wire c722_a;
  wire [2:0] c721_r0d;
  wire [2:0] c721_r1d;
  wire c721_a;
  wire [2:0] c720_r0d;
  wire [2:0] c720_r1d;
  wire c720_a;
  wire [2:0] c719_r0d;
  wire [2:0] c719_r1d;
  wire c719_a;
  wire [2:0] c718_r0d;
  wire [2:0] c718_r1d;
  wire c718_a;
  wire [31:0] c717_r0d;
  wire [31:0] c717_r1d;
  wire c717_a;
  wire [3:0] c716_r0d;
  wire [3:0] c716_r1d;
  wire c716_a;
  wire [2:0] c715_r0d;
  wire [2:0] c715_r1d;
  wire c715_a;
  wire [2:0] c714_r0d;
  wire [2:0] c714_r1d;
  wire c714_a;
  wire [2:0] c713_r0d;
  wire [2:0] c713_r1d;
  wire c713_a;
  wire [2:0] c712_r0d;
  wire [2:0] c712_r1d;
  wire c712_a;
  wire c711_r0d;
  wire c711_r1d;
  wire c711_a;
  wire [1:0] c710_r0d;
  wire [1:0] c710_r1d;
  wire c710_a;
  wire [1:0] c709_r0d;
  wire [1:0] c709_r1d;
  wire c709_a;
  wire [1:0] c708_r0d;
  wire [1:0] c708_r1d;
  wire c708_a;
  wire [1:0] c707_r0d;
  wire [1:0] c707_r1d;
  wire c707_a;
  wire c706_r0d;
  wire c706_r1d;
  wire c706_a;
  wire c705_r;
  wire c705_a;
  wire c704_r0d;
  wire c704_r1d;
  wire c704_a;
  wire c703_r0d;
  wire c703_r1d;
  wire c703_a;
  wire c702_r;
  wire c702_a;
  wire c701_r0d;
  wire c701_r1d;
  wire c701_a;
  wire c700_r;
  wire c700_a;
  wire [1:0] c699_r0d;
  wire [1:0] c699_r1d;
  wire c699_a;
  wire [1:0] c698_r0d;
  wire [1:0] c698_r1d;
  wire c698_a;
  wire [1:0] c697_r0d;
  wire [1:0] c697_r1d;
  wire c697_a;
  wire [1:0] c696_r0d;
  wire [1:0] c696_r1d;
  wire c696_a;
  wire c695_r0d;
  wire c695_r1d;
  wire c695_a;
  wire c694_r;
  wire c694_a;
  wire c693_r0d;
  wire c693_r1d;
  wire c693_a;
  wire c692_r0d;
  wire c692_r1d;
  wire c692_a;
  wire c691_r;
  wire c691_a;
  wire c690_r0d;
  wire c690_r1d;
  wire c690_a;
  wire c689_r;
  wire c689_a;
  wire [31:0] c688_r0d;
  wire [31:0] c688_r1d;
  wire c688_a;
  wire [1:0] c687_r0d;
  wire [1:0] c687_r1d;
  wire c687_a;
  wire [1:0] c686_r0d;
  wire [1:0] c686_r1d;
  wire c686_a;
  wire [1:0] c685_r0d;
  wire [1:0] c685_r1d;
  wire c685_a;
  wire [1:0] c684_r0d;
  wire [1:0] c684_r1d;
  wire c684_a;
  wire [31:0] c683_r0d;
  wire [31:0] c683_r1d;
  wire c683_a;
  wire c682_r;
  wire c682_a;
  wire [31:0] c681_r0d;
  wire [31:0] c681_r1d;
  wire c681_a;
  wire [31:0] c680_r0d;
  wire [31:0] c680_r1d;
  wire c680_a;
  wire c679_r;
  wire c679_a;
  wire [31:0] c678_r0d;
  wire [31:0] c678_r1d;
  wire c678_a;
  wire c677_r;
  wire c677_a;
  wire [2:0] c676_r0d;
  wire [2:0] c676_r1d;
  wire c676_a;
  wire [2:0] c675_r0d;
  wire [2:0] c675_r1d;
  wire c675_a;
  wire [2:0] c674_r0d;
  wire [2:0] c674_r1d;
  wire c674_a;
  wire [2:0] c673_r0d;
  wire [2:0] c673_r1d;
  wire c673_a;
  wire [2:0] c672_r0d;
  wire [2:0] c672_r1d;
  wire c672_a;
  wire c671_r0d;
  wire c671_r1d;
  wire c671_a;
  wire c670_r;
  wire c670_a;
  wire c669_r0d;
  wire c669_r1d;
  wire c669_a;
  wire c668_r0d;
  wire c668_r1d;
  wire c668_a;
  wire c667_r;
  wire c667_a;
  wire c666_r0d;
  wire c666_r1d;
  wire c666_a;
  wire c665_r;
  wire c665_a;
  wire c664_r0d;
  wire c664_r1d;
  wire c664_a;
  wire c663_r;
  wire c663_a;
  wire [1:0] c662_r0d;
  wire [1:0] c662_r1d;
  wire c662_a;
  wire [1:0] c661_r0d;
  wire [1:0] c661_r1d;
  wire c661_a;
  wire [1:0] c660_r0d;
  wire [1:0] c660_r1d;
  wire c660_a;
  wire [1:0] c659_r0d;
  wire [1:0] c659_r1d;
  wire c659_a;
  wire c658_r0d;
  wire c658_r1d;
  wire c658_a;
  wire c657_r;
  wire c657_a;
  wire c656_r0d;
  wire c656_r1d;
  wire c656_a;
  wire c655_r0d;
  wire c655_r1d;
  wire c655_a;
  wire c654_r;
  wire c654_a;
  wire c653_r0d;
  wire c653_r1d;
  wire c653_a;
  wire c652_r;
  wire c652_a;
  wire c651_r0d;
  wire c651_r1d;
  wire c651_a;
  wire c650_r0d;
  wire c650_r1d;
  wire c650_a;
  wire c649_r;
  wire c649_a;
  wire c648_r;
  wire c648_a;
  wire c647_r;
  wire c647_a;
  wire c646_r;
  wire c646_a;
  wire c645_r;
  wire c645_a;
  wire c644_r;
  wire c644_a;
  wire c643_r0d;
  wire c643_r1d;
  wire c643_a;
  wire c642_r;
  wire c642_a;
  wire c641_r0d;
  wire c641_r1d;
  wire c641_a;
  wire c640_r;
  wire c640_a;
  wire c639_r;
  wire c639_a;
  wire c638_r;
  wire c638_a;
  wire c637_r;
  wire c637_a;
  wire c636_r;
  wire c636_a;
  wire [31:0] c635_r0d;
  wire [31:0] c635_r1d;
  wire c635_a;
  wire c634_r;
  wire c634_a;
  wire c633_r;
  wire c633_a;
  wire c632_r;
  wire c632_a;
  wire c631_r0d;
  wire c631_r1d;
  wire c631_a;
  wire c630_r;
  wire c630_a;
  wire c629_r0d;
  wire c629_r1d;
  wire c629_a;
  wire c628_r;
  wire c628_a;
  wire c627_r;
  wire c627_a;
  wire c626_r0d;
  wire c626_r1d;
  wire c626_a;
  wire c625_r;
  wire c625_a;
  wire c624_r;
  wire c624_a;
  wire [31:0] c623_r0d;
  wire [31:0] c623_r1d;
  wire c623_a;
  wire c622_r;
  wire c622_a;
  wire c621_r;
  wire c621_a;
  wire c620_r;
  wire c620_a;
  wire c619_r;
  wire c619_a;
  wire c618_r;
  wire c618_a;
  wire c617_r;
  wire c617_a;
  wire [31:0] c616_r0d;
  wire [31:0] c616_r1d;
  wire c616_a;
  wire c615_r;
  wire c615_a;
  wire [31:0] c614_r0d;
  wire [31:0] c614_r1d;
  wire c614_a;
  wire c613_r;
  wire c613_a;
  wire c612_r;
  wire c612_a;
  wire c611_r0d;
  wire c611_r1d;
  wire c611_a;
  wire c610_r;
  wire c610_a;
  wire c609_r;
  wire c609_a;
  wire c608_r0d;
  wire c608_r1d;
  wire c608_a;
  wire c607_r;
  wire c607_a;
  wire c606_r0d;
  wire c606_r1d;
  wire c606_a;
  wire c605_r;
  wire c605_a;
  wire c604_r;
  wire c604_a;
  wire c603_r0d;
  wire c603_r1d;
  wire c603_a;
  wire c602_r;
  wire c602_a;
  wire c601_r0d;
  wire c601_r1d;
  wire c601_a;
  wire c600_r;
  wire c600_a;
  wire c599_r;
  wire c599_a;
  wire [31:0] c598_r0d;
  wire [31:0] c598_r1d;
  wire c598_a;
  wire c597_r;
  wire c597_a;
  wire [31:0] c596_r0d;
  wire [31:0] c596_r1d;
  wire c596_a;
  wire c595_r0d;
  wire c595_r1d;
  wire c595_a;
  wire c594_r;
  wire c594_a;
  wire c593_r;
  wire c593_a;
  wire c592_r;
  wire c592_a;
  wire c591_r;
  wire c591_a;
  wire c590_r;
  wire c590_a;
  wire c589_r;
  wire c589_a;
  wire c588_r;
  wire c588_a;
  wire [2:0] c587_r0d;
  wire [2:0] c587_r1d;
  wire c587_a;
  wire c586_r;
  wire c586_a;
  wire c585_r0d;
  wire c585_r1d;
  wire c585_a;
  wire c584_r;
  wire c584_a;
  wire c583_r0d;
  wire c583_r1d;
  wire c583_a;
  wire c582_r;
  wire c582_a;
  wire c581_r;
  wire c581_a;
  wire c580_r;
  wire c580_a;
  wire c579_r0d;
  wire c579_r1d;
  wire c579_a;
  wire c578_r;
  wire c578_a;
  wire c577_r;
  wire c577_a;
  wire c576_r0d;
  wire c576_r1d;
  wire c576_a;
  wire c575_r;
  wire c575_a;
  wire c574_r;
  wire c574_a;
  wire c573_r;
  wire c573_a;
  wire c572_r;
  wire c572_a;
  wire c571_r;
  wire c571_a;
  wire [31:0] c570_r0d;
  wire [31:0] c570_r1d;
  wire c570_a;
  wire c569_r;
  wire c569_a;
  wire [31:0] c568_r0d;
  wire [31:0] c568_r1d;
  wire c568_a;
  wire c567_r;
  wire c567_a;
  wire c566_r;
  wire c566_a;
  wire c565_r;
  wire c565_a;
  wire c564_r;
  wire c564_a;
  wire [31:0] c563_r0d;
  wire [31:0] c563_r1d;
  wire c563_a;
  wire c562_r;
  wire c562_a;
  wire c561_r;
  wire c561_a;
  wire [2:0] c560_r0d;
  wire [2:0] c560_r1d;
  wire c560_a;
  wire c559_r;
  wire c559_a;
  wire c558_r;
  wire c558_a;
  wire c557_r;
  wire c557_a;
  wire c556_r;
  wire c556_a;
  wire c555_r;
  wire c555_a;
  wire [31:0] c554_r0d;
  wire [31:0] c554_r1d;
  wire c554_a;
  wire c553_r;
  wire c553_a;
  wire [31:0] c552_r0d;
  wire [31:0] c552_r1d;
  wire c552_a;
  wire c551_r;
  wire c551_a;
  wire [31:0] c550_r0d;
  wire [31:0] c550_r1d;
  wire c550_a;
  wire c549_r;
  wire c549_a;
  wire c548_r;
  wire c548_a;
  wire [2:0] c547_r0d;
  wire [2:0] c547_r1d;
  wire c547_a;
  wire c546_r;
  wire c546_a;
  wire c545_r;
  wire c545_a;
  wire [2:0] c544_r0d;
  wire [2:0] c544_r1d;
  wire c544_a;
  wire c543_r;
  wire c543_a;
  wire c542_r;
  wire c542_a;
  wire [31:0] c541_r0d;
  wire [31:0] c541_r1d;
  wire c541_a;
  wire c540_r;
  wire c540_a;
  wire c539_r;
  wire c539_a;
  wire [31:0] c538_r0d;
  wire [31:0] c538_r1d;
  wire c538_a;
  wire c537_r0d;
  wire c537_r1d;
  wire c537_a;
  wire c536_r;
  wire c536_a;
  wire c535_r;
  wire c535_a;
  wire c534_r;
  wire c534_a;
  wire c533_r;
  wire c533_a;
  wire c532_r;
  wire c532_a;
  wire c531_r;
  wire c531_a;
  wire c530_r;
  wire c530_a;
  wire c529_r;
  wire c529_a;
  wire [31:0] c528_r0d;
  wire [31:0] c528_r1d;
  wire c528_a;
  wire c527_r;
  wire c527_a;
  wire [31:0] c526_r0d;
  wire [31:0] c526_r1d;
  wire c526_a;
  wire c525_r;
  wire c525_a;
  wire [31:0] c524_r0d;
  wire [31:0] c524_r1d;
  wire c524_a;
  wire c523_r;
  wire c523_a;
  wire [2:0] c522_r0d;
  wire [2:0] c522_r1d;
  wire c522_a;
  wire c521_r;
  wire c521_a;
  wire c520_r;
  wire c520_a;
  wire c519_r;
  wire c519_a;
  wire c518_r0d;
  wire c518_r1d;
  wire c518_a;
  wire c517_r;
  wire c517_a;
  wire c516_r;
  wire c516_a;
  wire c515_r0d;
  wire c515_r1d;
  wire c515_a;
  wire c514_r;
  wire c514_a;
  wire c513_r;
  wire c513_a;
  wire [31:0] c512_r0d;
  wire [31:0] c512_r1d;
  wire c512_a;
  wire [34:0] c511_r0d;
  wire [34:0] c511_r1d;
  wire c511_a;
  wire c510_r;
  wire c510_a;
  wire c509_r;
  wire c509_a;
  wire c508_r;
  wire c508_a;
  wire c507_r;
  wire c507_a;
  wire c506_r;
  wire c506_a;
  wire [32:0] c505_r0d;
  wire [32:0] c505_r1d;
  wire c505_a;
  wire c504_r;
  wire c504_a;
  wire [31:0] c503_r0d;
  wire [31:0] c503_r1d;
  wire c503_a;
  wire c502_r0d;
  wire c502_r1d;
  wire c502_a;
  wire c501_r;
  wire c501_a;
  wire [35:0] c500_r0d;
  wire [35:0] c500_r1d;
  wire c500_a;
  wire c499_r;
  wire c499_a;
  wire c498_r;
  wire c498_a;
  wire [31:0] c497_r0d;
  wire [31:0] c497_r1d;
  wire c497_a;
  wire [34:0] c496_r0d;
  wire [34:0] c496_r1d;
  wire c496_a;
  wire c495_r;
  wire c495_a;
  wire c494_r;
  wire c494_a;
  wire c493_r;
  wire c493_a;
  wire c492_r;
  wire c492_a;
  wire [32:0] c491_r0d;
  wire [32:0] c491_r1d;
  wire c491_a;
  wire c490_r;
  wire c490_a;
  wire [31:0] c489_r0d;
  wire [31:0] c489_r1d;
  wire c489_a;
  wire c488_r0d;
  wire c488_r1d;
  wire c488_a;
  wire c487_r;
  wire c487_a;
  wire [35:0] c486_r0d;
  wire [35:0] c486_r1d;
  wire c486_a;
  wire c485_r;
  wire c485_a;
  wire c484_r;
  wire c484_a;
  wire [31:0] c483_r0d;
  wire [31:0] c483_r1d;
  wire c483_a;
  wire [34:0] c482_r0d;
  wire [34:0] c482_r1d;
  wire c482_a;
  wire c481_r;
  wire c481_a;
  wire [2:0] c480_r0d;
  wire [2:0] c480_r1d;
  wire c480_a;
  wire c479_r;
  wire c479_a;
  wire c478_r;
  wire c478_a;
  wire c477_r;
  wire c477_a;
  wire c476_r;
  wire c476_a;
  wire c475_r;
  wire c475_a;
  wire c474_r0d;
  wire c474_r1d;
  wire c474_a;
  wire c473_r;
  wire c473_a;
  wire c472_r;
  wire c472_a;
  wire [9:0] c471_r0d;
  wire [9:0] c471_r1d;
  wire c471_a;
  wire c470_r;
  wire c470_a;
  wire c469_r;
  wire c469_a;
  wire [9:0] c468_r0d;
  wire [9:0] c468_r1d;
  wire c468_a;
  wire c467_r;
  wire c467_a;
  wire c466_r;
  wire c466_a;
  wire c465_r;
  wire c465_a;
  wire [8:0] c464_r0d;
  wire [8:0] c464_r1d;
  wire c464_a;
  wire [9:0] c463_r0d;
  wire [9:0] c463_r1d;
  wire c463_a;
  wire c462_r;
  wire c462_a;
  wire c461_r;
  wire c461_a;
  wire c460_r0d;
  wire c460_r1d;
  wire c460_a;
  wire c459_r;
  wire c459_a;
  wire c458_r0d;
  wire c458_r1d;
  wire c458_a;
  wire c457_r;
  wire c457_a;
  wire c456_r0d;
  wire c456_r1d;
  wire c456_a;
  wire c455_r;
  wire c455_a;
  wire c454_r0d;
  wire c454_r1d;
  wire c454_a;
  wire c453_r;
  wire c453_a;
  wire [34:0] c452_r0d;
  wire [34:0] c452_r1d;
  wire c452_a;
  wire [34:0] c451_r0d;
  wire [34:0] c451_r1d;
  wire c451_a;
  wire c450_r0d;
  wire c450_r1d;
  wire c450_a;
  wire c449_r;
  wire c449_a;
  wire c448_r;
  wire c448_a;
  wire c447_r;
  wire c447_a;
  wire c446_r;
  wire c446_a;
  wire c445_r;
  wire c445_a;
  wire c444_r0d;
  wire c444_r1d;
  wire c444_a;
  wire c443_r;
  wire c443_a;
  wire c442_r;
  wire c442_a;
  wire c441_r;
  wire c441_a;
  wire c440_r0d;
  wire c440_r1d;
  wire c440_a;
  wire c439_r;
  wire c439_a;
  wire c438_r;
  wire c438_a;
  wire c437_r0d;
  wire c437_r1d;
  wire c437_a;
  wire [1:0] c436_r0d;
  wire [1:0] c436_r1d;
  wire c436_a;
  wire c435_r;
  wire c435_a;
  wire c434_r0d;
  wire c434_r1d;
  wire c434_a;
  wire c433_r0d;
  wire c433_r1d;
  wire c433_a;
  wire [32:0] c432_r0d;
  wire [32:0] c432_r1d;
  wire c432_a;
  wire c431_r0d;
  wire c431_r1d;
  wire c431_a;
  wire c430_r;
  wire c430_a;
  wire c429_r;
  wire c429_a;
  wire [31:0] c428_r0d;
  wire [31:0] c428_r1d;
  wire c428_a;
  wire c427_r;
  wire c427_a;
  wire c426_r0d;
  wire c426_r1d;
  wire c426_a;
  wire c425_r;
  wire c425_a;
  wire c424_r;
  wire c424_a;
  wire [31:0] c423_r0d;
  wire [31:0] c423_r1d;
  wire c423_a;
  wire c422_r;
  wire c422_a;
  wire c421_r;
  wire c421_a;
  wire [31:0] c420_r0d;
  wire [31:0] c420_r1d;
  wire c420_a;
  wire c419_r;
  wire c419_a;
  wire c418_r;
  wire c418_a;
  wire c417_r;
  wire c417_a;
  wire c416_r;
  wire c416_a;
  wire c415_r;
  wire c415_a;
  wire c414_r;
  wire c414_a;
  wire c413_r0d;
  wire c413_r1d;
  wire c413_a;
  wire c412_r;
  wire c412_a;
  wire [31:0] c411_r0d;
  wire [31:0] c411_r1d;
  wire c411_a;
  wire c410_r;
  wire c410_a;
  wire [31:0] c409_r0d;
  wire [31:0] c409_r1d;
  wire c409_a;
  wire c408_r;
  wire c408_a;
  wire c407_r;
  wire c407_a;
  wire c406_r0d;
  wire c406_r1d;
  wire c406_a;
  wire c405_r;
  wire c405_a;
  wire c404_r;
  wire c404_a;
  wire [31:0] c403_r0d;
  wire [31:0] c403_r1d;
  wire c403_a;
  wire c402_r;
  wire c402_a;
  wire c401_r;
  wire c401_a;
  wire [31:0] c400_r0d;
  wire [31:0] c400_r1d;
  wire c400_a;
  wire c399_r;
  wire c399_a;
  wire [30:0] c398_r0d;
  wire [30:0] c398_r1d;
  wire c398_a;
  wire c397_r;
  wire c397_a;
  wire c396_r0d;
  wire c396_r1d;
  wire c396_a;
  wire c395_r;
  wire c395_a;
  wire c394_r;
  wire c394_a;
  wire c393_r;
  wire c393_a;
  wire c392_r;
  wire c392_a;
  wire c391_r;
  wire c391_a;
  wire c390_r0d;
  wire c390_r1d;
  wire c390_a;
  wire c389_r;
  wire c389_a;
  wire c388_r;
  wire c388_a;
  wire c387_r0d;
  wire c387_r1d;
  wire c387_a;
  wire c386_r;
  wire c386_a;
  wire c385_r;
  wire c385_a;
  wire [31:0] c384_r0d;
  wire [31:0] c384_r1d;
  wire c384_a;
  wire c383_r0d;
  wire c383_r1d;
  wire c383_a;
  wire c382_r;
  wire c382_a;
  wire c381_r;
  wire c381_a;
  wire c380_r;
  wire c380_a;
  wire c379_r;
  wire c379_a;
  wire c378_r;
  wire c378_a;
  wire c377_r;
  wire c377_a;
  wire c376_r0d;
  wire c376_r1d;
  wire c376_a;
  wire c375_r;
  wire c375_a;
  wire [31:0] c374_r0d;
  wire [31:0] c374_r1d;
  wire c374_a;
  wire c373_r;
  wire c373_a;
  wire c372_r;
  wire c372_a;
  wire c371_r;
  wire c371_a;
  wire c370_r0d;
  wire c370_r1d;
  wire c370_a;
  wire [32:0] c369_r0d;
  wire [32:0] c369_r1d;
  wire c369_a;
  wire c368_r0d;
  wire c368_r1d;
  wire c368_a;
  wire c367_r;
  wire c367_a;
  wire c366_r;
  wire c366_a;
  wire [31:0] c365_r0d;
  wire [31:0] c365_r1d;
  wire c365_a;
  wire c364_r;
  wire c364_a;
  wire c363_r;
  wire c363_a;
  wire c362_r0d;
  wire c362_r1d;
  wire c362_a;
  wire c361_r;
  wire c361_a;
  wire c360_r;
  wire c360_a;
  wire c359_r0d;
  wire c359_r1d;
  wire c359_a;
  wire c358_r;
  wire c358_a;
  wire c357_r;
  wire c357_a;
  wire [31:0] c356_r0d;
  wire [31:0] c356_r1d;
  wire c356_a;
  wire c355_r;
  wire c355_a;
  wire c354_r0d;
  wire c354_r1d;
  wire c354_a;
  wire c353_r;
  wire c353_a;
  wire c352_r;
  wire c352_a;
  wire c351_r;
  wire c351_a;
  wire [31:0] c350_r0d;
  wire [31:0] c350_r1d;
  wire c350_a;
  wire c349_r;
  wire c349_a;
  wire c348_r;
  wire c348_a;
  wire [31:0] c347_r0d;
  wire [31:0] c347_r1d;
  wire c347_a;
  wire c346_r;
  wire c346_a;
  wire c345_r;
  wire c345_a;
  wire c344_r;
  wire c344_a;
  wire c343_r;
  wire c343_a;
  wire c342_r0d;
  wire c342_r1d;
  wire c342_a;
  wire c341_r;
  wire c341_a;
  wire c340_r;
  wire c340_a;
  wire c339_r;
  wire c339_a;
  wire [3:0] c338_r0d;
  wire [3:0] c338_r1d;
  wire c338_a;
  wire c337_r;
  wire c337_a;
  wire c336_r;
  wire c336_a;
  wire [35:0] c335_r0d;
  wire [35:0] c335_r1d;
  wire c335_a;
  wire c334_r;
  wire c334_a;
  wire c333_r;
  wire c333_a;
  wire [34:0] c332_r0d;
  wire [34:0] c332_r1d;
  wire c332_a;
  wire c331_r;
  wire c331_a;
  wire c330_r;
  wire c330_a;
  wire [35:0] c329_r0d;
  wire [35:0] c329_r1d;
  wire c329_a;
  wire c328_r;
  wire c328_a;
  wire c327_r;
  wire c327_a;
  wire [34:0] c326_r0d;
  wire [34:0] c326_r1d;
  wire c326_a;
  wire c325_r;
  wire c325_a;
  wire c324_r0d;
  wire c324_r1d;
  wire c324_a;
  wire [33:0] c323_r0d;
  wire [33:0] c323_r1d;
  wire c323_a;
  wire c322_r;
  wire c322_a;
  wire c321_r0d;
  wire c321_r1d;
  wire c321_a;
  wire c320_r;
  wire c320_a;
  wire [32:0] c319_r0d;
  wire [32:0] c319_r1d;
  wire c319_a;
  wire c318_r;
  wire c318_a;
  wire c317_r;
  wire c317_a;
  wire c316_r;
  wire c316_a;
  wire c315_r;
  wire c315_a;
  wire c314_r0d;
  wire c314_r1d;
  wire c314_a;
  wire c313_r;
  wire c313_a;
  wire c312_r0d;
  wire c312_r1d;
  wire c312_a;
  wire c311_r;
  wire c311_a;
  wire c310_r;
  wire c310_a;
  wire c309_r;
  wire c309_a;
  wire c308_r;
  wire c308_a;
  wire c307_r;
  wire c307_a;
  wire c306_r;
  wire c306_a;
  wire c305_r0d;
  wire c305_r1d;
  wire c305_a;
  wire c304_r;
  wire c304_a;
  wire [34:0] c303_r0d;
  wire [34:0] c303_r1d;
  wire c303_a;
  wire c302_r;
  wire c302_a;
  wire [34:0] c301_r0d;
  wire [34:0] c301_r1d;
  wire c301_a;
  wire c300_r;
  wire c300_a;
  wire c299_r;
  wire c299_a;
  wire c298_r;
  wire c298_a;
  wire [34:0] c297_r0d;
  wire [34:0] c297_r1d;
  wire c297_a;
  wire c296_r;
  wire c296_a;
  wire [2:0] c295_r0d;
  wire [2:0] c295_r1d;
  wire c295_a;
  wire c294_r;
  wire c294_a;
  wire [31:0] c293_r0d;
  wire [31:0] c293_r1d;
  wire c293_a;
  wire [35:0] c292_r0d;
  wire [35:0] c292_r1d;
  wire c292_a;
  wire c291_r;
  wire c291_a;
  wire c290_r;
  wire c290_a;
  wire [31:0] c289_r0d;
  wire [31:0] c289_r1d;
  wire c289_a;
  wire [34:0] c288_r0d;
  wire [34:0] c288_r1d;
  wire c288_a;
  wire c287_r;
  wire c287_a;
  wire c286_r;
  wire c286_a;
  wire [34:0] c285_r0d;
  wire [34:0] c285_r1d;
  wire c285_a;
  wire c284_r;
  wire c284_a;
  wire [1:0] c283_r0d;
  wire [1:0] c283_r1d;
  wire c283_a;
  wire [32:0] c282_r0d;
  wire [32:0] c282_r1d;
  wire c282_a;
  wire c281_r;
  wire c281_a;
  wire c280_r0d;
  wire c280_r1d;
  wire c280_a;
  wire c279_r;
  wire c279_a;
  wire [31:0] c278_r0d;
  wire [31:0] c278_r1d;
  wire c278_a;
  wire [35:0] c277_r0d;
  wire [35:0] c277_r1d;
  wire c277_a;
  wire c276_r;
  wire c276_a;
  wire c275_r;
  wire c275_a;
  wire [34:0] c274_r0d;
  wire [34:0] c274_r1d;
  wire c274_a;
  wire c273_r;
  wire c273_a;
  wire c272_r;
  wire c272_a;
  wire c271_r;
  wire c271_a;
  wire [34:0] c270_r0d;
  wire [34:0] c270_r1d;
  wire c270_a;
  wire c269_r;
  wire c269_a;
  wire c268_r;
  wire c268_a;
  wire [34:0] c267_r0d;
  wire [34:0] c267_r1d;
  wire c267_a;
  wire c266_r;
  wire c266_a;
  wire c265_r;
  wire c265_a;
  wire [34:0] c264_r0d;
  wire [34:0] c264_r1d;
  wire c264_a;
  wire c263_r;
  wire c263_a;
  wire c262_r;
  wire c262_a;
  wire [34:0] c261_r0d;
  wire [34:0] c261_r1d;
  wire c261_a;
  wire c260_r;
  wire c260_a;
  wire c259_r;
  wire c259_a;
  wire [34:0] c258_r0d;
  wire [34:0] c258_r1d;
  wire c258_a;
  wire c257_r;
  wire c257_a;
  wire c256_r;
  wire c256_a;
  wire [34:0] c255_r0d;
  wire [34:0] c255_r1d;
  wire c255_a;
  wire c254_r;
  wire c254_a;
  wire c253_r;
  wire c253_a;
  wire [34:0] c252_r0d;
  wire [34:0] c252_r1d;
  wire c252_a;
  wire c251_r;
  wire c251_a;
  wire c250_r;
  wire c250_a;
  wire [34:0] c249_r0d;
  wire [34:0] c249_r1d;
  wire c249_a;
  wire c248_r;
  wire c248_a;
  wire c247_r;
  wire c247_a;
  wire [3:0] c246_r0d;
  wire [3:0] c246_r1d;
  wire c246_a;
  wire [34:0] c245_r0d;
  wire [34:0] c245_r1d;
  wire c245_a;
  wire c244_r;
  wire c244_a;
  wire [3:0] c243_r0d;
  wire [3:0] c243_r1d;
  wire c243_a;
  wire c242_r;
  wire c242_a;
  wire c241_r;
  wire c241_a;
  wire c240_r0d;
  wire c240_r1d;
  wire c240_a;
  wire c239_r;
  wire c239_a;
  wire c238_r;
  wire c238_a;
  wire [34:0] c237_r0d;
  wire [34:0] c237_r1d;
  wire c237_a;
  wire c236_r;
  wire c236_a;
  wire [34:0] c235_r0d;
  wire [34:0] c235_r1d;
  wire c235_a;
  wire c234_r;
  wire c234_a;
  wire c233_r;
  wire c233_a;
  wire [34:0] c232_r0d;
  wire [34:0] c232_r1d;
  wire c232_a;
  wire c231_r;
  wire c231_a;
  wire [34:0] c230_r0d;
  wire [34:0] c230_r1d;
  wire c230_a;
  wire c229_r;
  wire c229_a;
  wire c228_r;
  wire c228_a;
  wire [34:0] c227_r0d;
  wire [34:0] c227_r1d;
  wire c227_a;
  wire c226_r;
  wire c226_a;
  wire c225_r;
  wire c225_a;
  wire [34:0] c224_r0d;
  wire [34:0] c224_r1d;
  wire c224_a;
  wire c223_r0d;
  wire c223_r1d;
  wire c223_a;
  wire c222_r;
  wire c222_a;
  wire c221_r;
  wire c221_a;
  wire c220_r0d;
  wire c220_r1d;
  wire c220_a;
  wire c219_r;
  wire c219_a;
  wire c218_r;
  wire c218_a;
  wire c217_r;
  wire c217_a;
  wire [34:0] c216_r0d;
  wire [34:0] c216_r1d;
  wire c216_a;
  wire [34:0] c215_r0d;
  wire [34:0] c215_r1d;
  wire c215_a;
  wire c214_r;
  wire c214_a;
  wire c213_r;
  wire c213_a;
  wire [34:0] c212_r0d;
  wire [34:0] c212_r1d;
  wire c212_a;
  wire [34:0] c211_r0d;
  wire [34:0] c211_r1d;
  wire c211_a;
  wire c210_r;
  wire c210_a;
  wire c209_r;
  wire c209_a;
  wire [34:0] c208_r0d;
  wire [34:0] c208_r1d;
  wire c208_a;
  wire [34:0] c207_r0d;
  wire [34:0] c207_r1d;
  wire c207_a;
  wire c206_r;
  wire c206_a;
  wire c205_r;
  wire c205_a;
  wire [34:0] c204_r0d;
  wire [34:0] c204_r1d;
  wire c204_a;
  wire [34:0] c203_r0d;
  wire [34:0] c203_r1d;
  wire c203_a;
  wire c202_r;
  wire c202_a;
  wire c201_r;
  wire c201_a;
  wire c200_r;
  wire c200_a;
  wire c199_r;
  wire c199_a;
  wire c198_r;
  wire c198_a;
  wire c197_r;
  wire c197_a;
  wire c196_r;
  wire c196_a;
  wire c195_r0d;
  wire c195_r1d;
  wire c195_a;
  wire c194_r;
  wire c194_a;
  wire c193_r0d;
  wire c193_r1d;
  wire c193_a;
  wire c192_r;
  wire c192_a;
  wire [34:0] c191_r0d;
  wire [34:0] c191_r1d;
  wire c191_a;
  wire c190_r;
  wire c190_a;
  wire [35:0] c189_r0d;
  wire [35:0] c189_r1d;
  wire c189_a;
  wire c188_r;
  wire c188_a;
  wire [34:0] c187_r0d;
  wire [34:0] c187_r1d;
  wire c187_a;
  wire c186_r;
  wire c186_a;
  wire c185_r;
  wire c185_a;
  wire [35:0] c184_r0d;
  wire [35:0] c184_r1d;
  wire c184_a;
  wire c183_r;
  wire c183_a;
  wire c182_r;
  wire c182_a;
  wire [34:0] c181_r0d;
  wire [34:0] c181_r1d;
  wire c181_a;
  wire c180_r;
  wire c180_a;
  wire c179_r;
  wire c179_a;
  wire c178_r;
  wire c178_a;
  wire [3:0] c177_r0d;
  wire [3:0] c177_r1d;
  wire c177_a;
  wire c176_r;
  wire c176_a;
  wire c175_r;
  wire c175_a;
  wire [34:0] c174_r0d;
  wire [34:0] c174_r1d;
  wire c174_a;
  wire c173_r;
  wire c173_a;
  wire c172_r;
  wire c172_a;
  wire [35:0] c171_r0d;
  wire [35:0] c171_r1d;
  wire c171_a;
  wire c170_r;
  wire c170_a;
  wire c169_r;
  wire c169_a;
  wire c168_r;
  wire c168_a;
  wire c167_r;
  wire c167_a;
  wire c166_r;
  wire c166_a;
  wire c165_r0d;
  wire c165_r1d;
  wire c165_a;
  wire c164_r;
  wire c164_a;
  wire [31:0] c163_r0d;
  wire [31:0] c163_r1d;
  wire c163_a;
  wire c162_r;
  wire c162_a;
  wire [34:0] c161_r0d;
  wire [34:0] c161_r1d;
  wire c161_a;
  wire c160_r;
  wire c160_a;
  wire c159_r0d;
  wire c159_r1d;
  wire c159_a;
  wire [33:0] c158_r0d;
  wire [33:0] c158_r1d;
  wire c158_a;
  wire c157_r;
  wire c157_a;
  wire c156_r0d;
  wire c156_r1d;
  wire c156_a;
  wire [32:0] c155_r0d;
  wire [32:0] c155_r1d;
  wire c155_a;
  wire c154_r;
  wire c154_a;
  wire [31:0] c153_r0d;
  wire [31:0] c153_r1d;
  wire c153_a;
  wire c152_r;
  wire c152_a;
  wire c151_r0d;
  wire c151_r1d;
  wire c151_a;
  wire c150_r;
  wire c150_a;
  wire c149_r0d;
  wire c149_r1d;
  wire c149_a;
  wire c148_r;
  wire c148_a;
  wire c147_r;
  wire c147_a;
  wire c146_r;
  wire c146_a;
  wire [31:0] c145_r0d;
  wire [31:0] c145_r1d;
  wire c145_a;
  wire c144_r;
  wire c144_a;
  wire c143_r;
  wire c143_a;
  wire [31:0] c142_r0d;
  wire [31:0] c142_r1d;
  wire c142_a;
  wire c141_r;
  wire c141_a;
  wire c140_r;
  wire c140_a;
  wire [34:0] c139_r0d;
  wire [34:0] c139_r1d;
  wire c139_a;
  wire c138_r;
  wire c138_a;
  wire [32:0] c137_r0d;
  wire [32:0] c137_r1d;
  wire c137_a;
  wire [1:0] c136_r0d;
  wire [1:0] c136_r1d;
  wire c136_a;
  wire c135_r;
  wire c135_a;
  wire c134_r;
  wire c134_a;
  wire c133_r;
  wire c133_a;
  wire [34:0] c132_r0d;
  wire [34:0] c132_r1d;
  wire c132_a;
  wire c131_r;
  wire c131_a;
  wire [33:0] c130_r0d;
  wire [33:0] c130_r1d;
  wire c130_a;
  wire c129_r0d;
  wire c129_r1d;
  wire c129_a;
  wire c128_r;
  wire c128_a;
  wire c127_r;
  wire c127_a;
  wire c126_r;
  wire c126_a;
  wire [34:0] c125_r0d;
  wire [34:0] c125_r1d;
  wire c125_a;
  wire c124_r;
  wire c124_a;
  wire c123_r;
  wire c123_a;
  wire c122_r0d;
  wire c122_r1d;
  wire c122_a;
  wire c121_r;
  wire c121_a;
  wire c120_r;
  wire c120_a;
  wire c119_r0d;
  wire c119_r1d;
  wire c119_a;
  wire c118_r;
  wire c118_a;
  wire [32:0] c117_r0d;
  wire [32:0] c117_r1d;
  wire c117_a;
  wire [32:0] c116_r0d;
  wire [32:0] c116_r1d;
  wire c116_a;
  wire [33:0] c115_r0d;
  wire [33:0] c115_r1d;
  wire c115_a;
  wire c114_r;
  wire c114_a;
  wire c113_r;
  wire c113_a;
  wire c112_r;
  wire c112_a;
  wire c111_r;
  wire c111_a;
  wire c110_r;
  wire c110_a;
  wire [33:0] c109_r0d;
  wire [33:0] c109_r1d;
  wire c109_a;
  wire c108_r;
  wire c108_a;
  wire c107_r;
  wire c107_a;
  wire c106_r;
  wire c106_a;
  wire c105_r0d;
  wire c105_r1d;
  wire c105_a;
  wire c104_r;
  wire c104_a;
  wire c103_r;
  wire c103_a;
  wire [31:0] c102_r0d;
  wire [31:0] c102_r1d;
  wire c102_a;
  wire c101_r;
  wire c101_a;
  wire c100_r;
  wire c100_a;
  wire c99_r;
  wire c99_a;
  wire c98_r;
  wire c98_a;
  wire c97_r;
  wire c97_a;
  wire [32:0] c96_r0d;
  wire [32:0] c96_r1d;
  wire c96_a;
  wire c95_r;
  wire c95_a;
  wire [32:0] c94_r0d;
  wire [32:0] c94_r1d;
  wire c94_a;
  wire c93_r;
  wire c93_a;
  wire [33:0] c92_r0d;
  wire [33:0] c92_r1d;
  wire c92_a;
  wire [65:0] c91_r0d;
  wire [65:0] c91_r1d;
  wire c91_a;
  wire c90_r;
  wire c90_a;
  wire [32:0] c89_r0d;
  wire [32:0] c89_r1d;
  wire c89_a;
  wire c88_r;
  wire c88_a;
  wire [32:0] c87_r0d;
  wire [32:0] c87_r1d;
  wire c87_a;
  wire c86_r;
  wire c86_a;
  wire c85_r;
  wire c85_a;
  wire c84_r;
  wire c84_a;
  wire c83_r;
  wire c83_a;
  wire c82_r;
  wire c82_a;
  wire c81_r;
  wire c81_a;
  wire c80_r0d;
  wire c80_r1d;
  wire c80_a;
  wire c79_r;
  wire c79_a;
  wire [31:0] c78_r0d;
  wire [31:0] c78_r1d;
  wire c78_a;
  wire c77_r;
  wire c77_a;
  wire [31:0] c76_r0d;
  wire [31:0] c76_r1d;
  wire c76_a;
  wire c75_r;
  wire c75_a;
  wire c74_r;
  wire c74_a;
  wire c73_r;
  wire c73_a;
  wire [32:0] c72_r0d;
  wire [32:0] c72_r1d;
  wire c72_a;
  wire c71_r;
  wire c71_a;
  wire [31:0] c70_r0d;
  wire [31:0] c70_r1d;
  wire c70_a;
  wire c69_r;
  wire c69_a;
  wire c68_r0d;
  wire c68_r1d;
  wire c68_a;
  wire c67_r;
  wire c67_a;
  wire c66_r;
  wire c66_a;
  wire [32:0] c65_r0d;
  wire [32:0] c65_r1d;
  wire c65_a;
  wire c64_r;
  wire c64_a;
  wire [31:0] c63_r0d;
  wire [31:0] c63_r1d;
  wire c63_a;
  wire c62_r;
  wire c62_a;
  wire c61_r0d;
  wire c61_r1d;
  wire c61_a;
  wire c60_r;
  wire c60_a;
  wire c59_r;
  wire c59_a;
  wire c58_r;
  wire c58_a;
  wire c57_r;
  wire c57_a;
  wire c56_r;
  wire c56_a;
  wire c55_r;
  wire c55_a;
  wire c54_r;
  wire c54_a;
  wire [34:0] c53_r0d;
  wire [34:0] c53_r1d;
  wire c53_a;
  wire c52_r;
  wire c52_a;
  wire [34:0] c51_r0d;
  wire [34:0] c51_r1d;
  wire c51_a;
  wire c50_r;
  wire c50_a;
  wire [34:0] c49_r0d;
  wire [34:0] c49_r1d;
  wire c49_a;
  wire c48_r;
  wire c48_a;
  wire c47_r;
  wire c47_a;
  wire c46_r;
  wire c46_a;
  wire [34:0] c45_r0d;
  wire [34:0] c45_r1d;
  wire c45_a;
  wire [69:0] c44_r0d;
  wire [69:0] c44_r1d;
  wire c44_a;
  wire [34:0] c43_r0d;
  wire [34:0] c43_r1d;
  wire c43_a;
  wire [69:0] c42_r0d;
  wire [69:0] c42_r1d;
  wire c42_a;
  wire c41_r;
  wire c41_a;
  wire [34:0] c40_r0d;
  wire [34:0] c40_r1d;
  wire c40_a;
  wire c39_r;
  wire c39_a;
  wire [34:0] c38_r0d;
  wire [34:0] c38_r1d;
  wire c38_a;
  wire [34:0] c37_r0d;
  wire [34:0] c37_r1d;
  wire c37_a;
  wire [69:0] c36_r0d;
  wire [69:0] c36_r1d;
  wire c36_a;
  wire [34:0] c35_r0d;
  wire [34:0] c35_r1d;
  wire c35_a;
  wire [69:0] c34_r0d;
  wire [69:0] c34_r1d;
  wire c34_a;
  wire c33_r;
  wire c33_a;
  wire [34:0] c32_r0d;
  wire [34:0] c32_r1d;
  wire c32_a;
  wire c31_r;
  wire c31_a;
  wire [34:0] c30_r0d;
  wire [34:0] c30_r1d;
  wire c30_a;
  wire [34:0] c29_r0d;
  wire [34:0] c29_r1d;
  wire c29_a;
  wire [69:0] c28_r0d;
  wire [69:0] c28_r1d;
  wire c28_a;
  wire c27_r;
  wire c27_a;
  wire [34:0] c26_r0d;
  wire [34:0] c26_r1d;
  wire c26_a;
  wire c25_r;
  wire c25_a;
  wire [34:0] c24_r0d;
  wire [34:0] c24_r1d;
  wire c24_a;
  wire c23_r;
  wire c23_a;
  wire c22_r;
  wire c22_a;
  wire [34:0] c21_r0d;
  wire [34:0] c21_r1d;
  wire c21_a;
  wire [69:0] c20_r0d;
  wire [69:0] c20_r1d;
  wire c20_a;
  wire c19_r;
  wire c19_a;
  wire [34:0] c18_r0d;
  wire [34:0] c18_r1d;
  wire c18_a;
  wire [34:0] c17_r0d;
  wire [34:0] c17_r1d;
  wire c17_a;
  wire [69:0] c16_r0d;
  wire [69:0] c16_r1d;
  wire c16_a;
  wire c15_r;
  wire c15_a;
  wire [34:0] c14_r0d;
  wire [34:0] c14_r1d;
  wire c14_a;
  wire c13_r;
  wire c13_a;
  wire [34:0] c12_r0d;
  wire [34:0] c12_r1d;
  wire c12_a;
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I0 (c883_r0d, c883_r1d, c883_a, c607_r, c607_a, c630_r, c630_a, initialise);
  BrzJ_l11__280_202_29 I1 (c879_r, c879_a, c882_r0d, c882_r1d, c882_a, c883_r0d, c883_r1d, c883_a, initialise);
  BrzM_2_2 I2 (c880_r0d, c880_r1d, c880_a, c881_r0d, c881_r1d, c881_a, c882_r0d, c882_r1d, c882_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I3 (c876_r, c876_a, c881_r0d, c881_r1d, c881_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I4 (c874_r, c874_a, c880_r0d, c880_r1d, c880_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I5 (c878_r0d, c878_r1d, c878_a, c879_r, c879_a, mN_0r0d, mN_0r1d, mN_0a, initialise);
  BrzM_1_2 I6 (c875_r0d, c875_r1d, c875_a, c877_r0d, c877_r1d, c877_a, c878_r0d, c878_r1d, c878_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I7 (c629_r0d, c629_r1d, c629_a, c876_r, c876_a, c877_r0d, c877_r1d, c877_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I8 (c606_r0d, c606_r1d, c606_a, c874_r, c874_a, c875_r0d, c875_r1d, c875_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I9 (c873_r0d, c873_r1d, c873_a, c602_r, c602_a, c627_r, c627_a, initialise);
  BrzJ_l11__280_202_29 I10 (c869_r, c869_a, c872_r0d, c872_r1d, c872_a, c873_r0d, c873_r1d, c873_a, initialise);
  BrzM_2_2 I11 (c870_r0d, c870_r1d, c870_a, c871_r0d, c871_r1d, c871_a, c872_r0d, c872_r1d, c872_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I12 (c866_r, c866_a, c871_r0d, c871_r1d, c871_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I13 (c864_r, c864_a, c870_r0d, c870_r1d, c870_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I14 (c868_r0d, c868_r1d, c868_a, c869_r, c869_a, mZ_0r0d, mZ_0r1d, mZ_0a, initialise);
  BrzM_1_2 I15 (c865_r0d, c865_r1d, c865_a, c867_r0d, c867_r1d, c867_a, c868_r0d, c868_r1d, c868_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I16 (c626_r0d, c626_r1d, c626_a, c866_r, c866_a, c867_r0d, c867_r1d, c867_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I17 (c601_r0d, c601_r1d, c601_a, c864_r, c864_a, c865_r0d, c865_r1d, c865_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I18 (c863_r0d, c863_r1d, c863_a, c597_r, c597_a, c624_r, c624_a, initialise);
  BrzJ_l11__280_202_29 I19 (c859_r, c859_a, c862_r0d, c862_r1d, c862_a, c863_r0d, c863_r1d, c863_a, initialise);
  BrzM_2_2 I20 (c860_r0d, c860_r1d, c860_a, c861_r0d, c861_r1d, c861_a, c862_r0d, c862_r1d, c862_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I21 (c856_r, c856_a, c861_r0d, c861_r1d, c861_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I22 (c854_r, c854_a, c860_r0d, c860_r1d, c860_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I23 (c858_r0d, c858_r1d, c858_a, c859_r, c859_a, mpL_0r0d, mpL_0r1d, mpL_0a, initialise);
  BrzM_32_2 I24 (c855_r0d, c855_r1d, c855_a, c857_r0d, c857_r1d, c857_a, c858_r0d, c858_r1d, c858_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I25 (c623_r0d, c623_r1d, c623_a, c856_r, c856_a, c857_r0d, c857_r1d, c857_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I26 (c596_r0d, c596_r1d, c596_a, c854_r, c854_a, c855_r0d, c855_r1d, c855_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I27 (c853_r0d, c853_r1d, c853_a, c615_r, c615_a, c636_r, c636_a, initialise);
  BrzJ_l11__280_202_29 I28 (c849_r, c849_a, c852_r0d, c852_r1d, c852_a, c853_r0d, c853_r1d, c853_a, initialise);
  BrzM_2_2 I29 (c850_r0d, c850_r1d, c850_a, c851_r0d, c851_r1d, c851_a, c852_r0d, c852_r1d, c852_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I30 (c846_r, c846_a, c851_r0d, c851_r1d, c851_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I31 (c844_r, c844_a, c850_r0d, c850_r1d, c850_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I32 (c848_r0d, c848_r1d, c848_a, c849_r, c849_a, mpH_0r0d, mpH_0r1d, mpH_0a, initialise);
  BrzM_32_2 I33 (c845_r0d, c845_r1d, c845_a, c847_r0d, c847_r1d, c847_a, c848_r0d, c848_r1d, c848_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I34 (c635_r0d, c635_r1d, c635_a, c846_r, c846_a, c847_r0d, c847_r1d, c847_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I35 (c614_r0d, c614_r1d, c614_a, c844_r, c844_a, c845_r0d, c845_r1d, c845_a, initialise);
  BrzS_34_l12__2832_202_29_l97__28_28_28_281_m69m I36 (c843_r0d, c843_r1d, c843_a, c554_r0d, c554_r1d, c554_a, c563_r0d, c563_r1d, c563_a, initialise);
  BrzJ_l12__2832_202_29 I37 (c_0r0d, c_0r1d, c_0a, c842_r0d, c842_r1d, c842_a, c843_r0d, c843_r1d, c843_a, initialise);
  BrzM_2_2 I38 (c840_r0d, c840_r1d, c840_a, c841_r0d, c841_r1d, c841_a, c842_r0d, c842_r1d, c842_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I39 (c565_r, c565_a, c841_r0d, c841_r1d, c841_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I40 (c556_r, c556_a, c840_r0d, c840_r1d, c840_a);
  BrzJ_l12__2832_200_29 I41 (b_0r0d, b_0r1d, b_0a, c574_r, c574_a, c570_r0d, c570_r1d, c570_a, initialise);
  BrzJ_l12__2832_200_29 I42 (a_0r0d, a_0r1d, a_0a, c573_r, c573_a, c568_r0d, c568_r1d, c568_a, initialise);
  BrzJ_l11__283_200_29 I43 (mType_0r0d, mType_0r1d, mType_0a, c592_r, c592_a, c587_r0d, c587_r1d, c587_a, initialise);
  BrzJ_l11__281_200_29 I44 (bypassH_0r0d, bypassH_0r1d, bypassH_0a, c591_r, c591_a, c585_r0d, c585_r1d, c585_a, initialise);
  BrzJ_l11__281_200_29 I45 (bypass_0r0d, bypass_0r1d, bypass_0a, c590_r, c590_a, c583_r0d, c583_r1d, c583_a, initialise);
  BrzJ_l12__2835_200_29 I46 (c835_r0d, c835_r1d, c835_a, c198_r, c198_a, c187_r0d, c187_r1d, c187_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I47 (c839_r0d, c839_r1d, c839_a, c485_r, c485_a, c499_r, c499_a, initialise);
  BrzJ_l11__280_202_29 I48 (c834_r, c834_a, c838_r0d, c838_r1d, c838_a, c839_r0d, c839_r1d, c839_a, initialise);
  BrzM_2_2 I49 (c836_r0d, c836_r1d, c836_a, c837_r0d, c837_r1d, c837_a, c838_r0d, c838_r1d, c838_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I50 (c831_r, c831_a, c837_r0d, c837_r1d, c837_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I51 (c829_r, c829_a, c836_r0d, c836_r1d, c836_a);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I52 (c833_r0d, c833_r1d, c833_a, c834_r, c834_a, c835_r0d, c835_r1d, c835_a, initialise);
  BrzM_35_2 I53 (c830_r0d, c830_r1d, c830_a, c832_r0d, c832_r1d, c832_a, c833_r0d, c833_r1d, c833_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I54 (c496_r0d, c496_r1d, c496_a, c831_r, c831_a, c832_r0d, c832_r1d, c832_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I55 (c482_r0d, c482_r1d, c482_a, c829_r, c829_a, c830_r0d, c830_r1d, c830_a, initialise);
  BrzJ_l12__2836_200_29 I56 (c824_r0d, c824_r1d, c824_a, c199_r, c199_a, c189_r0d, c189_r1d, c189_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I57 (c828_r0d, c828_r1d, c828_a, c493_r, c493_a, c507_r, c507_a, initialise);
  BrzJ_l11__280_202_29 I58 (c823_r, c823_a, c827_r0d, c827_r1d, c827_a, c828_r0d, c828_r1d, c828_a, initialise);
  BrzM_2_2 I59 (c825_r0d, c825_r1d, c825_a, c826_r0d, c826_r1d, c826_a, c827_r0d, c827_r1d, c827_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I60 (c820_r, c820_a, c826_r0d, c826_r1d, c826_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I61 (c818_r, c818_a, c825_r0d, c825_r1d, c825_a);
  BrzF_36_l32__28_280_200_29_20_280_2036_29__m44m I62 (c822_r0d, c822_r1d, c822_a, c823_r, c823_a, c824_r0d, c824_r1d, c824_a, initialise);
  BrzM_36_2 I63 (c819_r0d, c819_r1d, c819_a, c821_r0d, c821_r1d, c821_a, c822_r0d, c822_r1d, c822_a, initialise);
  BrzF_36_l32__28_280_200_29_20_280_2036_29__m44m I64 (c500_r0d, c500_r1d, c500_a, c820_r, c820_a, c821_r0d, c821_r1d, c821_a, initialise);
  BrzF_36_l32__28_280_200_29_20_280_2036_29__m44m I65 (c486_r0d, c486_r1d, c486_a, c818_r, c818_a, c819_r0d, c819_r1d, c819_a, initialise);
  BrzJ_l12__2835_200_29 I66 (c817_r0d, c817_r1d, c817_a, c200_r, c200_a, c191_r0d, c191_r1d, c191_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I67 (c511_r0d, c511_r1d, c511_a, c514_r, c514_a, c817_r0d, c817_r1d, c817_a, initialise);
  BrzJ_l11__281_200_29 I68 (c816_r0d, c816_r1d, c816_a, c201_r, c201_a, c193_r0d, c193_r1d, c193_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I69 (c515_r0d, c515_r1d, c515_a, c517_r, c517_a, c816_r0d, c816_r1d, c816_a, initialise);
  BrzJ_l11__281_200_29 I70 (c815_r0d, c815_r1d, c815_a, c202_r, c202_a, c195_r0d, c195_r1d, c195_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I71 (c518_r0d, c518_r1d, c518_a, c520_r, c520_a, c815_r0d, c815_r1d, c815_a, initialise);
  BrzJ_l12__2832_200_29 I72 (c814_r0d, c814_r1d, c814_a, c532_r, c532_a, c524_r0d, c524_r1d, c524_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I73 (c538_r0d, c538_r1d, c538_a, c540_r, c540_a, c814_r0d, c814_r1d, c814_a, initialise);
  BrzJ_l12__2832_200_29 I74 (c813_r0d, c813_r1d, c813_a, c533_r, c533_a, c526_r0d, c526_r1d, c526_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I75 (c541_r0d, c541_r1d, c541_a, c543_r, c543_a, c813_r0d, c813_r1d, c813_a, initialise);
  BrzJ_l12__2832_200_29 I76 (c808_r0d, c808_r1d, c808_a, c534_r, c534_a, c528_r0d, c528_r1d, c528_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I77 (c812_r0d, c812_r1d, c812_a, c551_r, c551_a, c553_r, c553_a, initialise);
  BrzJ_l11__280_202_29 I78 (c807_r, c807_a, c811_r0d, c811_r1d, c811_a, c812_r0d, c812_r1d, c812_a, initialise);
  BrzM_2_2 I79 (c809_r0d, c809_r1d, c809_a, c810_r0d, c810_r1d, c810_a, c811_r0d, c811_r1d, c811_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I80 (c804_r, c804_a, c810_r0d, c810_r1d, c810_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I81 (c802_r, c802_a, c809_r0d, c809_r1d, c809_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I82 (c806_r0d, c806_r1d, c806_a, c807_r, c807_a, c808_r0d, c808_r1d, c808_a, initialise);
  BrzM_32_2 I83 (c803_r0d, c803_r1d, c803_a, c805_r0d, c805_r1d, c805_a, c806_r0d, c806_r1d, c806_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I84 (c552_r0d, c552_r1d, c552_a, c804_r, c804_a, c805_r0d, c805_r1d, c805_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I85 (c550_r0d, c550_r1d, c550_a, c802_r, c802_a, c803_r0d, c803_r1d, c803_a, initialise);
  BrzJ_l11__283_200_29 I86 (c801_r0d, c801_r1d, c801_a, c531_r, c531_a, c522_r0d, c522_r1d, c522_a, initialise);
  BrzF_3_l31__28_280_200_29_20_280_203_29_29 I87 (c544_r0d, c544_r1d, c544_a, c546_r, c546_a, c801_r0d, c801_r1d, c801_a, initialise);
  BrzJ_l12__2835_200_29 I88 (c800_r0d, c800_r1d, c800_a, c56_r, c56_a, c49_r0d, c49_r1d, c49_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I89 (c224_r0d, c224_r1d, c224_a, c226_r, c226_a, c800_r0d, c800_r1d, c800_a, initialise);
  BrzJ_l12__2835_200_29 I90 (c788_r0d, c788_r1d, c788_a, c57_r, c57_a, c51_r0d, c51_r1d, c51_a, initialise);
  BrzS_9_l11__280_209_29_l424__28_28_28_281__m68m I91 (c799_r0d, c799_r1d, c799_a, c248_r, c248_a, c251_r, c251_a, c254_r, c254_a, c257_r, c257_a, c260_r, c260_a, c263_r, c263_a, c266_r, c266_a, c269_r, c269_a, c272_r, c272_a, initialise);
  BrzJ_l11__280_209_29 I92 (c787_r, c787_a, c798_r0d, c798_r1d, c798_a, c799_r0d, c799_r1d, c799_a, initialise);
  BrzM_9_9 I93 (c789_r0d, c789_r1d, c789_a, c790_r0d, c790_r1d, c790_a, c791_r0d, c791_r1d, c791_a, c792_r0d, c792_r1d, c792_a, c793_r0d, c793_r1d, c793_a, c794_r0d, c794_r1d, c794_a, c795_r0d, c795_r1d, c795_a, c796_r0d, c796_r1d, c796_a, c797_r0d, c797_r1d, c797_a, c798_r0d, c798_r1d, c798_a, initialise);
  BrzO_0_9_l25__28_28num_209_20256_29_29 I94 (c784_r, c784_a, c797_r0d, c797_r1d, c797_a);
  BrzO_0_9_l25__28_28num_209_20128_29_29 I95 (c782_r, c782_a, c796_r0d, c796_r1d, c796_a);
  BrzO_0_9_l24__28_28num_209_2064_29_29 I96 (c780_r, c780_a, c795_r0d, c795_r1d, c795_a);
  BrzO_0_9_l24__28_28num_209_2032_29_29 I97 (c778_r, c778_a, c794_r0d, c794_r1d, c794_a);
  BrzO_0_9_l24__28_28num_209_2016_29_29 I98 (c776_r, c776_a, c793_r0d, c793_r1d, c793_a);
  BrzO_0_9_l23__28_28num_209_208_29_29 I99 (c774_r, c774_a, c792_r0d, c792_r1d, c792_a);
  BrzO_0_9_l23__28_28num_209_204_29_29 I100 (c772_r, c772_a, c791_r0d, c791_r1d, c791_a);
  BrzO_0_9_l23__28_28num_209_202_29_29 I101 (c770_r, c770_a, c790_r0d, c790_r1d, c790_a);
  BrzO_0_9_l23__28_28num_209_201_29_29 I102 (c768_r, c768_a, c789_r0d, c789_r1d, c789_a);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I103 (c786_r0d, c786_r1d, c786_a, c787_r, c787_a, c788_r0d, c788_r1d, c788_a, initialise);
  BrzM_35_9 I104 (c769_r0d, c769_r1d, c769_a, c771_r0d, c771_r1d, c771_a, c773_r0d, c773_r1d, c773_a, c775_r0d, c775_r1d, c775_a, c777_r0d, c777_r1d, c777_a, c779_r0d, c779_r1d, c779_a, c781_r0d, c781_r1d, c781_a, c783_r0d, c783_r1d, c783_a, c785_r0d, c785_r1d, c785_a, c786_r0d, c786_r1d, c786_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I105 (c270_r0d, c270_r1d, c270_a, c784_r, c784_a, c785_r0d, c785_r1d, c785_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I106 (c267_r0d, c267_r1d, c267_a, c782_r, c782_a, c783_r0d, c783_r1d, c783_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I107 (c264_r0d, c264_r1d, c264_a, c780_r, c780_a, c781_r0d, c781_r1d, c781_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I108 (c261_r0d, c261_r1d, c261_a, c778_r, c778_a, c779_r0d, c779_r1d, c779_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I109 (c258_r0d, c258_r1d, c258_a, c776_r, c776_a, c777_r0d, c777_r1d, c777_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I110 (c255_r0d, c255_r1d, c255_a, c774_r, c774_a, c775_r0d, c775_r1d, c775_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I111 (c252_r0d, c252_r1d, c252_a, c772_r, c772_a, c773_r0d, c773_r1d, c773_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I112 (c249_r0d, c249_r1d, c249_a, c770_r, c770_a, c771_r0d, c771_r1d, c771_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I113 (c245_r0d, c245_r1d, c245_a, c768_r, c768_a, c769_r0d, c769_r1d, c769_a, initialise);
  BrzJ_l12__2835_200_29 I114 (c767_r0d, c767_r1d, c767_a, c58_r, c58_a, c53_r0d, c53_r1d, c53_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I115 (c227_r0d, c227_r1d, c227_a, c229_r, c229_a, c767_r0d, c767_r1d, c767_a, initialise);
  BrzJ_l12__2835_200_29 I116 (c766_r0d, c766_r1d, c766_a, c239_r, c239_a, c237_r0d, c237_r1d, c237_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I117 (c45_r0d, c45_r1d, c45_a, c47_r, c47_a, c766_r0d, c766_r1d, c766_a, initialise);
  BrzJ_l12__2835_200_29 I118 (c765_r0d, c765_r1d, c765_a, c234_r, c234_a, c232_r0d, c232_r1d, c232_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I119 (c21_r0d, c21_r1d, c21_a, c23_r, c23_a, c765_r0d, c765_r1d, c765_a, initialise);
  BrzJ_l12__2832_200_29 I120 (c759_r0d, c759_r1d, c759_a, c83_r, c83_a, c76_r0d, c76_r1d, c76_a, initialise);
  BrzS_3_l11__280_203_29_l141__28_28_28_281__m64m I121 (c764_r0d, c764_r1d, c764_a, c144_r, c144_a, c349_r, c349_a, c402_r, c402_a, initialise);
  BrzJ_l11__280_203_29 I122 (c758_r, c758_a, c763_r0d, c763_r1d, c763_a, c764_r0d, c764_r1d, c764_a, initialise);
  BrzM_3_3 I123 (c760_r0d, c760_r1d, c760_a, c761_r0d, c761_r1d, c761_a, c762_r0d, c762_r1d, c762_a, c763_r0d, c763_r1d, c763_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I124 (c755_r, c755_a, c762_r0d, c762_r1d, c762_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I125 (c753_r, c753_a, c761_r0d, c761_r1d, c761_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I126 (c751_r, c751_a, c760_r0d, c760_r1d, c760_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I127 (c757_r0d, c757_r1d, c757_a, c758_r, c758_a, c759_r0d, c759_r1d, c759_a, initialise);
  BrzM_32_3 I128 (c752_r0d, c752_r1d, c752_a, c754_r0d, c754_r1d, c754_a, c756_r0d, c756_r1d, c756_a, c757_r0d, c757_r1d, c757_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I129 (c400_r0d, c400_r1d, c400_a, c755_r, c755_a, c756_r0d, c756_r1d, c756_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I130 (c347_r0d, c347_r1d, c347_a, c753_r, c753_a, c754_r0d, c754_r1d, c754_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I131 (c142_r0d, c142_r1d, c142_a, c751_r, c751_a, c752_r0d, c752_r1d, c752_a, initialise);
  BrzJ_l12__2832_200_29 I132 (c745_r0d, c745_r1d, c745_a, c84_r, c84_a, c78_r0d, c78_r1d, c78_a, initialise);
  BrzS_3_l11__280_203_29_l141__28_28_28_281__m64m I133 (c750_r0d, c750_r1d, c750_a, c147_r, c147_a, c352_r, c352_a, c405_r, c405_a, initialise);
  BrzJ_l11__280_203_29 I134 (c744_r, c744_a, c749_r0d, c749_r1d, c749_a, c750_r0d, c750_r1d, c750_a, initialise);
  BrzM_3_3 I135 (c746_r0d, c746_r1d, c746_a, c747_r0d, c747_r1d, c747_a, c748_r0d, c748_r1d, c748_a, c749_r0d, c749_r1d, c749_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I136 (c741_r, c741_a, c748_r0d, c748_r1d, c748_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I137 (c739_r, c739_a, c747_r0d, c747_r1d, c747_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I138 (c737_r, c737_a, c746_r0d, c746_r1d, c746_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I139 (c743_r0d, c743_r1d, c743_a, c744_r, c744_a, c745_r0d, c745_r1d, c745_a, initialise);
  BrzM_32_3 I140 (c738_r0d, c738_r1d, c738_a, c740_r0d, c740_r1d, c740_a, c742_r0d, c742_r1d, c742_a, c743_r0d, c743_r1d, c743_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I141 (c403_r0d, c403_r1d, c403_a, c741_r, c741_a, c742_r0d, c742_r1d, c742_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I142 (c350_r0d, c350_r1d, c350_a, c739_r, c739_a, c740_r0d, c740_r1d, c740_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I143 (c145_r0d, c145_r1d, c145_a, c737_r, c737_a, c738_r0d, c738_r1d, c738_a, initialise);
  BrzJ_l11__281_200_29 I144 (c731_r0d, c731_r1d, c731_a, c85_r, c85_a, c80_r0d, c80_r1d, c80_a, initialise);
  BrzS_3_l11__280_203_29_l141__28_28_28_281__m64m I145 (c736_r0d, c736_r1d, c736_a, c150_r, c150_a, c355_r, c355_a, c408_r, c408_a, initialise);
  BrzJ_l11__280_203_29 I146 (c730_r, c730_a, c735_r0d, c735_r1d, c735_a, c736_r0d, c736_r1d, c736_a, initialise);
  BrzM_3_3 I147 (c732_r0d, c732_r1d, c732_a, c733_r0d, c733_r1d, c733_a, c734_r0d, c734_r1d, c734_a, c735_r0d, c735_r1d, c735_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I148 (c727_r, c727_a, c734_r0d, c734_r1d, c734_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I149 (c725_r, c725_a, c733_r0d, c733_r1d, c733_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I150 (c723_r, c723_a, c732_r0d, c732_r1d, c732_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I151 (c729_r0d, c729_r1d, c729_a, c730_r, c730_a, c731_r0d, c731_r1d, c731_a, initialise);
  BrzM_1_3 I152 (c724_r0d, c724_r1d, c724_a, c726_r0d, c726_r1d, c726_a, c728_r0d, c728_r1d, c728_a, c729_r0d, c729_r1d, c729_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I153 (c406_r0d, c406_r1d, c406_a, c727_r, c727_a, c728_r0d, c728_r1d, c728_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I154 (c354_r0d, c354_r1d, c354_a, c725_r, c725_a, c726_r0d, c726_r1d, c726_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I155 (c149_r0d, c149_r1d, c149_a, c723_r, c723_a, c724_r0d, c724_r1d, c724_a, initialise);
  BrzS_35_l12__2832_203_29_l144__28_28_28_28_m70m I156 (c722_r0d, c722_r1d, c722_a, c163_r0d, c163_r1d, c163_a, c374_r0d, c374_r1d, c374_a, c411_r0d, c411_r1d, c411_a, initialise);
  BrzJ_l12__2832_203_29 I157 (c717_r0d, c717_r1d, c717_a, c721_r0d, c721_r1d, c721_a, c722_r0d, c722_r1d, c722_a, initialise);
  BrzM_3_3 I158 (c718_r0d, c718_r1d, c718_a, c719_r0d, c719_r1d, c719_a, c720_r0d, c720_r1d, c720_a, c721_r0d, c721_r1d, c721_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I159 (c416_r, c416_a, c720_r0d, c720_r1d, c720_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I160 (c379_r, c379_a, c719_r0d, c719_r1d, c719_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I161 (c168_r, c168_a, c718_r0d, c718_r1d, c718_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I162 (c102_r0d, c102_r1d, c102_a, c104_r, c104_a, c717_r0d, c717_r1d, c717_a, initialise);
  BrzS_4_l11__281_203_29_l141__28_28_28_281__m67m I163 (c716_r0d, c716_r1d, c716_a, c165_r0d, c165_r1d, c165_a, c376_r0d, c376_r1d, c376_a, c413_r0d, c413_r1d, c413_a, initialise);
  BrzJ_l11__281_203_29 I164 (c711_r0d, c711_r1d, c711_a, c715_r0d, c715_r1d, c715_a, c716_r0d, c716_r1d, c716_a, initialise);
  BrzM_3_3 I165 (c712_r0d, c712_r1d, c712_a, c713_r0d, c713_r1d, c713_a, c714_r0d, c714_r1d, c714_a, c715_r0d, c715_r1d, c715_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I166 (c417_r, c417_a, c714_r0d, c714_r1d, c714_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I167 (c380_r, c380_a, c713_r0d, c713_r1d, c713_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I168 (c169_r, c169_a, c712_r0d, c712_r1d, c712_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I169 (c105_r0d, c105_r1d, c105_a, c107_r, c107_a, c711_r0d, c711_r1d, c711_a, initialise);
  BrzJ_l11__281_200_29 I170 (c706_r0d, c706_r1d, c706_a, c453_r, c453_a, c456_r0d, c456_r1d, c456_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I171 (c710_r0d, c710_r1d, c710_a, c221_r, c221_a, c343_r, c343_a, initialise);
  BrzJ_l11__280_202_29 I172 (c705_r, c705_a, c709_r0d, c709_r1d, c709_a, c710_r0d, c710_r1d, c710_a, initialise);
  BrzM_2_2 I173 (c707_r0d, c707_r1d, c707_a, c708_r0d, c708_r1d, c708_a, c709_r0d, c709_r1d, c709_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I174 (c702_r, c702_a, c708_r0d, c708_r1d, c708_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I175 (c700_r, c700_a, c707_r0d, c707_r1d, c707_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I176 (c704_r0d, c704_r1d, c704_a, c705_r, c705_a, c706_r0d, c706_r1d, c706_a, initialise);
  BrzM_1_2 I177 (c701_r0d, c701_r1d, c701_a, c703_r0d, c703_r1d, c703_a, c704_r0d, c704_r1d, c704_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I178 (c342_r0d, c342_r1d, c342_a, c702_r, c702_a, c703_r0d, c703_r1d, c703_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I179 (c220_r0d, c220_r1d, c220_a, c700_r, c700_a, c701_r0d, c701_r1d, c701_a, initialise);
  BrzJ_l11__281_200_29 I180 (c695_r0d, c695_r1d, c695_a, c316_r, c316_a, c314_r0d, c314_r1d, c314_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I181 (c699_r0d, c699_r1d, c699_a, c462_r, c462_a, c475_r, c475_a, initialise);
  BrzJ_l11__280_202_29 I182 (c694_r, c694_a, c698_r0d, c698_r1d, c698_a, c699_r0d, c699_r1d, c699_a, initialise);
  BrzM_2_2 I183 (c696_r0d, c696_r1d, c696_a, c697_r0d, c697_r1d, c697_a, c698_r0d, c698_r1d, c698_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I184 (c691_r, c691_a, c697_r0d, c697_r1d, c697_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I185 (c689_r, c689_a, c696_r0d, c696_r1d, c696_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I186 (c693_r0d, c693_r1d, c693_a, c694_r, c694_a, c695_r0d, c695_r1d, c695_a, initialise);
  BrzM_1_2 I187 (c690_r0d, c690_r1d, c690_a, c692_r0d, c692_r1d, c692_a, c693_r0d, c693_r1d, c693_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I188 (c474_r0d, c474_r1d, c474_a, c691_r, c691_a, c692_r0d, c692_r1d, c692_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I189 (c460_r0d, c460_r1d, c460_a, c689_r, c689_a, c690_r0d, c690_r1d, c690_a, initialise);
  BrzJ_l12__2832_200_29 I190 (c688_r0d, c688_r1d, c688_a, c618_r, c618_a, c616_r0d, c616_r1d, c616_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I191 (c420_r0d, c420_r1d, c420_a, c422_r, c422_a, c688_r0d, c688_r1d, c688_a, initialise);
  BrzJ_l12__2832_200_29 I192 (c683_r0d, c683_r1d, c683_a, c600_r, c600_a, c598_r0d, c598_r1d, c598_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I193 (c687_r0d, c687_r1d, c687_a, c386_r, c386_a, c425_r, c425_a, initialise);
  BrzJ_l11__280_202_29 I194 (c682_r, c682_a, c686_r0d, c686_r1d, c686_a, c687_r0d, c687_r1d, c687_a, initialise);
  BrzM_2_2 I195 (c684_r0d, c684_r1d, c684_a, c685_r0d, c685_r1d, c685_a, c686_r0d, c686_r1d, c686_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I196 (c679_r, c679_a, c685_r0d, c685_r1d, c685_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I197 (c677_r, c677_a, c684_r0d, c684_r1d, c684_a);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I198 (c681_r0d, c681_r1d, c681_a, c682_r, c682_a, c683_r0d, c683_r1d, c683_a, initialise);
  BrzM_32_2 I199 (c678_r0d, c678_r1d, c678_a, c680_r0d, c680_r1d, c680_a, c681_r0d, c681_r1d, c681_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I200 (c423_r0d, c423_r1d, c423_a, c679_r, c679_a, c680_r0d, c680_r1d, c680_a, initialise);
  BrzF_32_l32__28_280_200_29_20_280_2032_29__m40m I201 (c384_r0d, c384_r1d, c384_a, c677_r, c677_a, c678_r0d, c678_r1d, c678_a, initialise);
  BrzJ_l11__281_200_29 I202 (c671_r0d, c671_r1d, c671_a, c605_r, c605_a, c603_r0d, c603_r1d, c603_a, initialise);
  BrzS_3_l11__280_203_29_l141__28_28_28_281__m64m I203 (c676_r0d, c676_r1d, c676_a, c389_r, c389_a, c439_r, c439_a, c442_r, c442_a, initialise);
  BrzJ_l11__280_203_29 I204 (c670_r, c670_a, c675_r0d, c675_r1d, c675_a, c676_r0d, c676_r1d, c676_a, initialise);
  BrzM_3_3 I205 (c672_r0d, c672_r1d, c672_a, c673_r0d, c673_r1d, c673_a, c674_r0d, c674_r1d, c674_a, c675_r0d, c675_r1d, c675_a, initialise);
  BrzO_0_3_l23__28_28num_203_204_29_29 I206 (c667_r, c667_a, c674_r0d, c674_r1d, c674_a);
  BrzO_0_3_l23__28_28num_203_202_29_29 I207 (c665_r, c665_a, c673_r0d, c673_r1d, c673_a);
  BrzO_0_3_l23__28_28num_203_201_29_29 I208 (c663_r, c663_a, c672_r0d, c672_r1d, c672_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I209 (c669_r0d, c669_r1d, c669_a, c670_r, c670_a, c671_r0d, c671_r1d, c671_a, initialise);
  BrzM_1_3 I210 (c664_r0d, c664_r1d, c664_a, c666_r0d, c666_r1d, c666_a, c668_r0d, c668_r1d, c668_a, c669_r0d, c669_r1d, c669_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I211 (c440_r0d, c440_r1d, c440_a, c667_r, c667_a, c668_r0d, c668_r1d, c668_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I212 (c437_r0d, c437_r1d, c437_a, c665_r, c665_a, c666_r0d, c666_r1d, c666_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I213 (c387_r0d, c387_r1d, c387_a, c663_r, c663_a, c664_r0d, c664_r1d, c664_a, initialise);
  BrzJ_l11__281_200_29 I214 (c658_r0d, c658_r1d, c658_a, c610_r, c610_a, c608_r0d, c608_r1d, c608_a, initialise);
  BrzS_2_l11__280_202_29_l95__28_28_28_281_2_m62m I215 (c662_r0d, c662_r1d, c662_a, c392_r, c392_a, c446_r, c446_a, initialise);
  BrzJ_l11__280_202_29 I216 (c657_r, c657_a, c661_r0d, c661_r1d, c661_a, c662_r0d, c662_r1d, c662_a, initialise);
  BrzM_2_2 I217 (c659_r0d, c659_r1d, c659_a, c660_r0d, c660_r1d, c660_a, c661_r0d, c661_r1d, c661_a, initialise);
  BrzO_0_2_l23__28_28num_202_202_29_29 I218 (c654_r, c654_a, c660_r0d, c660_r1d, c660_a);
  BrzO_0_2_l23__28_28num_202_201_29_29 I219 (c652_r, c652_a, c659_r0d, c659_r1d, c659_a);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I220 (c656_r0d, c656_r1d, c656_a, c657_r, c657_a, c658_r0d, c658_r1d, c658_a, initialise);
  BrzM_1_2 I221 (c653_r0d, c653_r1d, c653_a, c655_r0d, c655_r1d, c655_a, c656_r0d, c656_r1d, c656_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I222 (c444_r0d, c444_r1d, c444_a, c654_r, c654_a, c655_r0d, c655_r1d, c655_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I223 (c390_r0d, c390_r1d, c390_a, c652_r, c652_a, c653_r0d, c653_r1d, c653_a, initialise);
  BrzJ_l11__281_200_29 I224 (c651_r0d, c651_r1d, c651_a, c646_r, c646_a, c641_r0d, c641_r1d, c641_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I225 (c579_r0d, c579_r1d, c579_a, c581_r, c581_a, c651_r0d, c651_r1d, c651_a, initialise);
  BrzJ_l11__281_200_29 I226 (c650_r0d, c650_r1d, c650_a, c647_r, c647_a, c643_r0d, c643_r1d, c643_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I227 (c576_r0d, c576_r1d, c576_a, c578_r, c578_a, c650_r0d, c650_r1d, c650_a, initialise);
  BrzF_0_l101__28_280_200_29_20_280_200_29_2_m37m I228 (go_0r, go_0a, c60_r, c60_a, c114_r, c114_a, c449_r, c449_a, c479_r, c479_a, c536_r, c536_a, c594_r, c594_a, c649_r, c649_a, initialise);
  BrzM_0_2 I229 (c649_r, c649_a, c640_r, c640_a, c648_r, c648_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I230 (c648_r, c648_a, c646_r, c646_a, c647_r, c647_a, initialise);
  BrzJ_l11__280_200_29 I231 (c642_r, c642_a, c644_r, c644_a, c645_r, c645_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I232 (c643_r0d, c643_r1d, c643_a, c644_r, c644_a, c645_r, c645_a, c595_r0d, c595_r1d, c595_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m72m I233 (c641_r0d, c641_r1d, c641_a, c642_r, c642_a, c612_r, c612_a, c632_r, c632_a, c611_r0d, c611_r1d, c611_a, c631_r0d, c631_r1d, c631_a, initialise);
  BrzM_0_2 I234 (c621_r, c621_a, c639_r, c639_a, c640_r, c640_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I235 (c595_r0d, c595_r1d, c595_a, c620_r, c620_a, c638_r, c638_a, initialise);
  BrzJ_l19__280_200_200_200_29 I236 (c624_r, c624_a, c627_r, c627_a, c630_r, c630_a, c637_r, c637_a, c639_r, c639_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I237 (c638_r, c638_a, c622_r, c622_a, c625_r, c625_a, c628_r, c628_a, c632_r, c632_a, initialise);
  BrzM_0_2 I238 (c633_r, c633_a, c636_r, c636_a, c637_r, c637_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I239 (c631_r0d, c631_r1d, c631_a, c633_r, c633_a, c634_r, c634_a, initialise);
  BrzO_0_32_l24__28_28num_2032_200_29_29 I240 (c634_r, c634_a, c635_r0d, c635_r1d, c635_a);
  BrzO_0_1_l23__28_28num_201_200_29_29 I241 (c628_r, c628_a, c629_r0d, c629_r1d, c629_a);
  BrzO_0_1_l23__28_28num_201_200_29_29 I242 (c625_r, c625_a, c626_r0d, c626_r1d, c626_a);
  BrzO_0_32_l24__28_28num_2032_200_29_29 I243 (c622_r, c622_a, c623_r0d, c623_r1d, c623_a);
  BrzJ_l19__280_200_200_200_29 I244 (c597_r, c597_a, c602_r, c602_a, c607_r, c607_a, c619_r, c619_a, c621_r, c621_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I245 (c620_r, c620_a, c600_r, c600_a, c605_r, c605_a, c610_r, c610_a, c612_r, c612_a, initialise);
  BrzM_0_2 I246 (c613_r, c613_a, c615_r, c615_a, c619_r, c619_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I247 (c611_r0d, c611_r1d, c611_a, c613_r, c613_a, c618_r, c618_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I248 (c616_r0d, c616_r1d, c616_a, c617_r, c617_a, c617_r, c617_a, c614_r0d, c614_r1d, c614_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I249 (c608_r0d, c608_r1d, c608_a, c609_r, c609_a, c609_r, c609_a, c606_r0d, c606_r1d, c606_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I250 (c603_r0d, c603_r1d, c603_a, c604_r, c604_a, c604_r, c604_a, c601_r0d, c601_r1d, c601_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I251 (c598_r0d, c598_r1d, c598_a, c599_r, c599_a, c599_r, c599_a, c596_r0d, c596_r1d, c596_a, initialise);
  BrzM_0_2 I252 (c594_r, c594_a, c582_r, c582_a, c593_r, c593_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I253 (c593_r, c593_a, c590_r, c590_a, c591_r, c591_a, c592_r, c592_a, initialise);
  BrzJ_l15__280_200_200_29 I254 (c584_r, c584_a, c586_r, c586_a, c588_r, c588_a, c589_r, c589_a, initialise);
  BrzV_3_l6__28_29_l23__28_28_280_203_29_29__m75m I255 (c587_r0d, c587_r1d, c587_a, c588_r, c588_a, c545_r, c545_a, c548_r, c548_a, c561_r, c561_a, c544_r0d, c544_r1d, c544_a, c547_r0d, c547_r1d, c547_a, c560_r0d, c560_r1d, c560_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I256 (c585_r0d, c585_r1d, c585_a, c586_r, c586_a, c580_r, c580_a, c579_r0d, c579_r1d, c579_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m72m I257 (c583_r0d, c583_r1d, c583_a, c584_r, c584_a, c572_r, c572_a, c577_r, c577_a, c537_r0d, c537_r1d, c537_a, c576_r0d, c576_r1d, c576_a, initialise);
  BrzJ_l15__280_200_200_29 I258 (c567_r, c567_a, c578_r, c578_a, c581_r, c581_a, c582_r, c582_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I259 (c589_r, c589_a, c575_r, c575_a, c577_r, c577_a, c580_r, c580_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I260 (c575_r, c575_a, c573_r, c573_a, c574_r, c574_a, initialise);
  BrzJ_l11__280_200_29 I261 (c569_r, c569_a, c571_r, c571_a, c572_r, c572_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I262 (c570_r0d, c570_r1d, c570_a, c571_r, c571_a, c542_r, c542_a, c541_r0d, c541_r1d, c541_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I263 (c568_r0d, c568_r1d, c568_a, c569_r, c569_a, c539_r, c539_a, c538_r0d, c538_r1d, c538_a, initialise);
  BrzM_0_2 I264 (c559_r, c559_a, c566_r, c566_a, c567_r, c567_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I265 (c537_r0d, c537_r1d, c537_a, c558_r, c558_a, c561_r, c561_a, initialise);
  BrzM_0_2 I266 (c562_r, c562_a, c564_r, c564_a, c566_r, c566_a, initialise);
  BrzS_3_l11__280_203_29_l137__28_28_28_280__m63m I267 (c560_r0d, c560_r1d, c560_a, c562_r, c562_a, c565_r, c565_a, initialise);
  BrzF_32_l17__28_280_200_29_29 I268 (c563_r0d, c563_r1d, c563_a, c564_r, c564_a, initialise);
  BrzJ_l19__280_200_200_200_29 I269 (c540_r, c540_a, c543_r, c543_a, c546_r, c546_a, c557_r, c557_a, c559_r, c559_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I270 (c558_r, c558_a, c539_r, c539_a, c542_r, c542_a, c545_r, c545_a, c548_r, c548_a, initialise);
  BrzM_0_2 I271 (c551_r, c551_a, c553_r, c553_a, c557_r, c557_a, initialise);
  BrzS_3_l11__280_203_29_l137__28_28_28_280__m63m I272 (c547_r0d, c547_r1d, c547_a, c549_r, c549_a, c556_r, c556_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I273 (c554_r0d, c554_r1d, c554_a, c555_r, c555_a, c555_r, c555_a, c552_r0d, c552_r1d, c552_a, initialise);
  BrzO_0_32_l24__28_28num_2032_200_29_29 I274 (c549_r, c549_a, c550_r0d, c550_r1d, c550_a);
  BrzM_0_2 I275 (c536_r, c536_a, c521_r, c521_a, c535_r, c535_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I276 (c535_r, c535_a, c531_r, c531_a, c532_r, c532_a, c533_r, c533_a, c534_r, c534_a, initialise);
  BrzJ_l19__280_200_200_200_29 I277 (c523_r, c523_a, c525_r, c525_a, c527_r, c527_a, c529_r, c529_a, c530_r, c530_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I278 (c528_r0d, c528_r1d, c528_a, c529_r, c529_a, c513_r, c513_a, c512_r0d, c512_r1d, c512_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m81m I279 (c526_r0d, c526_r1d, c526_a, c527_r, c527_a, c490_r, c490_a, c504_r, c504_a, c489_r0d, c489_r1d, c489_a, c503_r0d, c503_r1d, c503_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m81m I280 (c524_r0d, c524_r1d, c524_a, c525_r, c525_a, c484_r, c484_a, c498_r, c498_a, c483_r0d, c483_r1d, c483_a, c497_r0d, c497_r1d, c497_a, initialise);
  BrzV_3_l6__28_29_l23__28_28_280_203_29_29__m76m I281 (c522_r0d, c522_r1d, c522_a, c523_r, c523_a, c481_r, c481_a, c516_r, c516_a, c519_r, c519_a, c480_r0d, c480_r1d, c480_a, c515_r0d, c515_r1d, c515_a, c518_r0d, c518_r1d, c518_a, initialise);
  BrzJ_l19__280_200_200_200_29 I282 (c510_r, c510_a, c514_r, c514_a, c517_r, c517_a, c520_r, c520_a, c521_r, c521_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I283 (c530_r, c530_a, c481_r, c481_a, c513_r, c513_a, c516_r, c516_a, c519_r, c519_a, initialise);
  BrzO_32_35_l76__28_28num_203_200_29_20_28a_m51m I284 (c512_r0d, c512_r1d, c512_a, c511_r0d, c511_r1d, c511_a);
  BrzM_0_2 I285 (c495_r, c495_a, c509_r, c509_a, c510_r, c510_a, initialise);
  BrzS_3_l11__280_203_29_l151__28_28_28_281__m65m I286 (c480_r0d, c480_r1d, c480_a, c494_r, c494_a, c508_r, c508_a, initialise);
  BrzJ_l11__280_200_29 I287 (c499_r, c499_a, c507_r, c507_a, c509_r, c509_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I288 (c508_r, c508_a, c498_r, c498_a, c506_r, c506_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I289 (c506_r, c506_a, c501_r, c501_a, c504_r, c504_a, initialise);
  BrzO_33_36_l76__28_28num_203_200_29_20_28a_m54m I290 (c505_r0d, c505_r1d, c505_a, c500_r0d, c500_r1d, c500_a);
  BrzJ_l12__281_2032_29 I291 (c502_r0d, c502_r1d, c502_a, c503_r0d, c503_r1d, c503_a, c505_r0d, c505_r1d, c505_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I292 (c501_r, c501_a, c502_r0d, c502_r1d, c502_a);
  BrzO_32_35_l76__28_28num_203_200_29_20_28a_m51m I293 (c497_r0d, c497_r1d, c497_a, c496_r0d, c496_r1d, c496_a);
  BrzJ_l11__280_200_29 I294 (c485_r, c485_a, c493_r, c493_a, c495_r, c495_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I295 (c494_r, c494_a, c484_r, c484_a, c492_r, c492_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I296 (c492_r, c492_a, c487_r, c487_a, c490_r, c490_a, initialise);
  BrzO_33_36_l91__28_28app_203_20_280_2032_2_m53m I297 (c491_r0d, c491_r1d, c491_a, c486_r0d, c486_r1d, c486_a);
  BrzJ_l12__281_2032_29 I298 (c488_r0d, c488_r1d, c488_a, c489_r0d, c489_r1d, c489_a, c491_r0d, c491_r1d, c491_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I299 (c487_r, c487_a, c488_r0d, c488_r1d, c488_a);
  BrzO_32_35_l91__28_28app_203_20_280_2031_2_m50m I300 (c483_r0d, c483_r1d, c483_a, c482_r0d, c482_r1d, c482_a);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I301 (c454_r0d, c454_r1d, c454_a, c455_r, c455_a, c455_r, c455_a, c458_r0d, c458_r1d, c458_a, initialise);
  BrzV_10_l6__28_29_l45__28_28_280_2010_29_2_m79m I302 (c471_r0d, c471_r1d, c471_a, c468_r0d, c468_r1d, c468_a, c472_r, c472_a, c469_r, c469_a, c465_r, c465_a, c461_r, c461_a, c464_r0d, c464_r1d, c464_a, c460_r0d, c460_r1d, c460_a, initialise);
  BrzV_10_l6__28_29_l24__28_28_280_2010_29_2_m78m I303 (c463_r0d, c463_r1d, c463_a, c466_r, c466_a, c467_r, c467_a, c468_r0d, c468_r1d, c468_a, initialise);
  BrzM_0_2 I304 (c479_r, c479_a, c478_r, c478_a, c453_r, c453_a, initialise);
  BrzM_0_2 I305 (c469_r, c469_a, c477_r, c477_a, c478_r, c478_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I306 (c458_r0d, c458_r1d, c458_a, c459_r, c459_a, c476_r, c476_a, initialise);
  BrzJ_l11__280_200_29 I307 (c472_r, c472_a, c475_r, c475_a, c477_r, c477_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I308 (c476_r, c476_a, c470_r, c470_a, c473_r, c473_a, initialise);
  BrzO_0_1_l23__28_28num_201_201_29_29 I309 (c473_r, c473_a, c474_r0d, c474_r1d, c474_a);
  BrzO_0_10_l26__28_28num_2010_20256_29_29 I310 (c470_r, c470_a, c471_r0d, c471_r1d, c471_a);
  BrzJ_l11__280_200_29 I311 (c462_r, c462_a, c466_r, c466_a, c467_r, c467_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I312 (c459_r, c459_a, c461_r, c461_a, c465_r, c465_a, initialise);
  BrzO_9_10_l75__28_28num_201_200_29_20_28ap_m49m I313 (c464_r0d, c464_r1d, c464_a, c463_r0d, c463_r1d, c463_a);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I314 (c456_r0d, c456_r1d, c456_a, c457_r, c457_a, c457_r, c457_a, c454_r0d, c454_r1d, c454_a, initialise);
  BrzJ_l12__2835_200_29 I315 (c452_r0d, c452_r1d, c452_a, c308_r, c308_a, c301_r0d, c301_r1d, c301_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I316 (c230_r0d, c230_r1d, c230_a, c231_r, c231_a, c452_r0d, c452_r1d, c452_a, initialise);
  BrzJ_l12__2835_200_29 I317 (c451_r0d, c451_r1d, c451_a, c309_r, c309_a, c303_r0d, c303_r1d, c303_a, initialise);
  BrzF_35_l32__28_280_200_29_20_280_2035_29__m43m I318 (c235_r0d, c235_r1d, c235_a, c236_r, c236_a, c451_r0d, c451_r1d, c451_a, initialise);
  BrzJ_l11__281_200_29 I319 (c450_r0d, c450_r1d, c450_a, c310_r, c310_a, c305_r0d, c305_r1d, c305_a, initialise);
  BrzF_1_l31__28_280_200_29_20_280_201_29_29 I320 (c240_r0d, c240_r1d, c240_a, c242_r, c242_a, c450_r0d, c450_r1d, c450_a, initialise);
  BrzV_4_l6__28_29_l43__28_28_280_204_29_29__m77m I321 (c338_r0d, c338_r1d, c338_a, c177_r0d, c177_r1d, c177_a, c340_r, c340_a, c179_r, c179_a, c247_r, c247_a, c244_r, c244_a, c241_r, c241_a, c246_r0d, c246_r1d, c246_a, c243_r0d, c243_r1d, c243_a, c240_r0d, c240_r1d, c240_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m83m I322 (c409_r0d, c409_r1d, c409_a, c410_r, c410_a, c445_r, c445_a, c429_r, c429_a, c421_r, c421_a, c444_r0d, c444_r1d, c444_a, c428_r0d, c428_r1d, c428_a, c420_r0d, c420_r1d, c420_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m81m I323 (c356_r0d, c356_r1d, c356_a, c358_r, c358_a, c424_r, c424_a, c385_r, c385_a, c423_r0d, c423_r1d, c423_a, c384_r0d, c384_r1d, c384_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m90m I324 (c125_r0d, c125_r1d, c125_a, c127_r, c127_a, c250_r, c250_a, c205_r, c205_a, c249_r0d, c249_r1d, c249_a, c204_r0d, c204_r1d, c204_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m90m I325 (c132_r0d, c132_r1d, c132_a, c134_r, c134_a, c253_r, c253_a, c209_r, c209_a, c252_r0d, c252_r1d, c252_a, c208_r0d, c208_r1d, c208_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m90m I326 (c161_r0d, c161_r1d, c161_a, c162_r, c162_a, c256_r, c256_a, c213_r, c213_a, c255_r0d, c255_r1d, c255_a, c212_r0d, c212_r1d, c212_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m90m I327 (c139_r0d, c139_r1d, c139_a, c141_r, c141_a, c259_r, c259_a, c217_r, c217_a, c258_r0d, c258_r1d, c258_a, c216_r0d, c216_r1d, c216_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I328 (c203_r0d, c203_r1d, c203_a, c206_r, c206_a, c271_r, c271_a, c270_r0d, c270_r1d, c270_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I329 (c207_r0d, c207_r1d, c207_a, c210_r, c210_a, c268_r, c268_a, c267_r0d, c267_r1d, c267_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I330 (c211_r0d, c211_r1d, c211_a, c214_r, c214_a, c265_r, c265_a, c264_r0d, c264_r1d, c264_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I331 (c215_r0d, c215_r1d, c215_a, c218_r, c218_a, c262_r, c262_a, c261_r0d, c261_r1d, c261_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m92m I332 (c274_r0d, c274_r1d, c274_a, c276_r, c276_a, c404_r, c404_a, c325_r, c325_a, c322_r, c322_a, c320_r, c320_a, c403_r0d, c403_r1d, c403_a, c324_r0d, c324_r1d, c324_a, c321_r0d, c321_r1d, c321_a, c319_r0d, c319_r1d, c319_a, initialise);
  BrzV_36_l6__28_29_l24__28_28_280_2036_29_2_m96m I333 (c277_r0d, c277_r1d, c277_a, c287_r, c287_a, c351_r, c351_a, c330_r, c330_a, c350_r0d, c350_r1d, c350_a, c329_r0d, c329_r1d, c329_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m86m I334 (c288_r0d, c288_r1d, c288_a, c291_r, c291_a, c399_r, c399_a, c333_r, c333_a, c398_r0d, c398_r1d, c398_a, c332_r0d, c332_r1d, c332_a, initialise);
  BrzV_36_l6__28_29_l24__28_28_280_2036_29_2_m97m I335 (c292_r0d, c292_r1d, c292_a, c299_r, c299_a, c397_r, c397_a, c348_r, c348_a, c339_r, c339_a, c336_r, c336_a, c396_r0d, c396_r1d, c396_a, c347_r0d, c347_r1d, c347_a, c338_r0d, c338_r1d, c338_a, c335_r0d, c335_r1d, c335_a, initialise);
  BrzV_35_l6__28_29_l45__28_28_280_2035_29_2_m94m I336 (c332_r0d, c332_r1d, c332_a, c174_r0d, c174_r1d, c174_a, c334_r, c334_a, c176_r, c176_a, c225_r, c225_a, c224_r0d, c224_r1d, c224_a, initialise);
  BrzV_35_l6__28_29_l45__28_28_280_2035_29_2_m94m I337 (c326_r0d, c326_r1d, c326_a, c181_r0d, c181_r1d, c181_a, c328_r, c328_a, c182_r, c182_a, c228_r, c228_a, c227_r0d, c227_r1d, c227_a, initialise);
  BrzV_36_l6__28_29_l45__28_28_280_2036_29_2_m98m I338 (c329_r0d, c329_r1d, c329_a, c184_r0d, c184_r1d, c184_a, c331_r, c331_a, c185_r, c185_a, c279_r, c279_a, c278_r0d, c278_r1d, c278_a, initialise);
  BrzV_36_l6__28_29_l45__28_28_280_2036_29_2_m98m I339 (c335_r0d, c335_r1d, c335_a, c171_r0d, c171_r1d, c171_a, c337_r, c337_a, c173_r, c173_a, c294_r, c294_a, c293_r0d, c293_r1d, c293_a, initialise);
  BrzV_1_l6__28_29_l43__28_28_280_201_29_29__m74m I340 (c359_r0d, c359_r1d, c359_a, c312_r0d, c312_r1d, c312_a, c361_r, c361_a, c313_r, c313_a, c407_r, c407_a, c318_r, c318_a, c406_r0d, c406_r1d, c406_a, c223_r0d, c223_r1d, c223_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I341 (c119_r0d, c119_r1d, c119_a, c121_r, c121_a, c382_r, c382_a, c383_r0d, c383_r1d, c383_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I342 (c122_r0d, c122_r1d, c122_a, c124_r, c124_a, c427_r, c427_a, c426_r0d, c426_r1d, c426_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m73m I343 (c370_r0d, c370_r1d, c370_a, c372_r, c372_a, c441_r, c441_a, c435_r, c435_a, c388_r, c388_a, c440_r0d, c440_r1d, c440_a, c434_r0d, c434_r1d, c434_a, c387_r0d, c387_r1d, c387_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I344 (c362_r0d, c362_r1d, c362_a, c364_r, c364_a, c391_r, c391_a, c390_r0d, c390_r1d, c390_a, initialise);
  BrzM_0_2 I345 (c449_r, c449_a, c448_r, c448_a, c118_r, c118_a, initialise);
  BrzM_0_2 I346 (c394_r, c394_a, c447_r, c447_a, c448_r, c448_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I347 (c383_r0d, c383_r1d, c383_a, c393_r, c393_a, c395_r, c395_a, initialise);
  BrzJ_l19__280_200_200_200_29 I348 (c422_r, c422_a, c425_r, c425_a, c443_r, c443_a, c446_r, c446_a, c447_r, c447_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I349 (c419_r, c419_a, c421_r, c421_a, c424_r, c424_a, c427_r, c427_a, c445_r, c445_a, initialise);
  BrzM_0_2 I350 (c439_r, c439_a, c442_r, c442_a, c443_r, c443_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I351 (c426_r0d, c426_r1d, c426_a, c438_r, c438_a, c441_r, c441_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I352 (c438_r, c438_a, c429_r, c429_a, c430_r, c430_a, c435_r, c435_a, initialise);
  BrzO_2_1_l119__28_28app_201_20_280_200_201_m47m I353 (c436_r0d, c436_r1d, c436_a, c437_r0d, c437_r1d, c437_a);
  BrzJ_l11__281_201_29 I354 (c433_r0d, c433_r1d, c433_a, c434_r0d, c434_r1d, c434_a, c436_r0d, c436_r1d, c436_a, initialise);
  BrzO_33_1_l196__28_28app_201_20_280_200_20_m52m I355 (c432_r0d, c432_r1d, c432_a, c433_r0d, c433_r1d, c433_a);
  BrzJ_l12__2832_201_29 I356 (c428_r0d, c428_r1d, c428_a, c431_r0d, c431_r1d, c431_a, c432_r0d, c432_r1d, c432_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I357 (c430_r, c430_a, c431_r0d, c431_r1d, c431_a);
  BrzJ_l19__280_200_200_200_29 I358 (c402_r, c402_a, c405_r, c405_a, c408_r, c408_a, c410_r, c410_a, c419_r, c419_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I359 (c395_r, c395_a, c401_r, c401_a, c404_r, c404_a, c407_r, c407_a, c418_r, c418_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I360 (c418_r, c418_a, c416_r, c416_a, c417_r, c417_a, initialise);
  BrzJ_l11__280_200_29 I361 (c412_r, c412_a, c414_r, c414_a, c415_r, c415_a, initialise);
  BrzF_1_l17__28_280_200_29_29 I362 (c413_r0d, c413_r1d, c413_a, c414_r, c414_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I363 (c411_r0d, c411_r1d, c411_a, c412_r, c412_a, c415_r, c415_a, c409_r0d, c409_r1d, c409_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I364 (c401_r, c401_a, c397_r, c397_a, c399_r, c399_a, initialise);
  BrzJ_l12__281_2031_29 I365 (c396_r0d, c396_r1d, c396_a, c398_r0d, c398_r1d, c398_a, c400_r0d, c400_r1d, c400_a, initialise);
  BrzJ_l15__280_200_200_29 I366 (c386_r, c386_a, c389_r, c389_a, c392_r, c392_a, c394_r, c394_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I367 (c393_r, c393_a, c385_r, c385_a, c388_r, c388_a, c391_r, c391_a, initialise);
  BrzJ_l19__280_200_200_200_29 I368 (c349_r, c349_a, c352_r, c352_a, c355_r, c355_a, c373_r, c373_a, c382_r, c382_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I369 (c346_r, c346_a, c348_r, c348_a, c351_r, c351_a, c353_r, c353_a, c381_r, c381_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I370 (c381_r, c381_a, c379_r, c379_a, c380_r, c380_a, initialise);
  BrzJ_l11__280_200_29 I371 (c375_r, c375_a, c377_r, c377_a, c378_r, c378_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I372 (c376_r0d, c376_r1d, c376_a, c377_r, c377_a, c360_r, c360_a, c359_r0d, c359_r1d, c359_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m82m I373 (c374_r0d, c374_r1d, c374_a, c375_r, c375_a, c357_r, c357_a, c363_r, c363_a, c366_r, c366_a, c356_r0d, c356_r1d, c356_a, c362_r0d, c362_r1d, c362_a, c365_r0d, c365_r1d, c365_a, initialise);
  BrzJ_l19__280_200_200_200_29 I374 (c358_r, c358_a, c361_r, c361_a, c364_r, c364_a, c372_r, c372_a, c373_r, c373_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I375 (c378_r, c378_a, c357_r, c357_a, c360_r, c360_a, c363_r, c363_a, c371_r, c371_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I376 (c371_r, c371_a, c366_r, c366_a, c367_r, c367_a, initialise);
  BrzO_33_1_l196__28_28app_201_20_280_200_20_m52m I377 (c369_r0d, c369_r1d, c369_a, c370_r0d, c370_r1d, c370_a);
  BrzJ_l12__2832_201_29 I378 (c365_r0d, c365_r1d, c365_a, c368_r0d, c368_r1d, c368_a, c369_r0d, c369_r1d, c369_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I379 (c367_r, c367_a, c368_r0d, c368_r1d, c368_a);
  BrzO_0_1_l23__28_28num_201_200_29_29 I380 (c353_r, c353_a, c354_r0d, c354_r1d, c354_a);
  BrzM_0_2 I381 (c222_r, c222_a, c345_r, c345_a, c317_r, c317_a, initialise);
  BrzS_1_l11__280_201_29_l95__28_28_28_280_2_m61m I382 (c223_r0d, c223_r1d, c223_a, c346_r, c346_a, c344_r, c344_a, initialise);
  BrzJ_l27__280_200_200_200_200_200_29 I383 (c328_r, c328_a, c331_r, c331_a, c334_r, c334_a, c337_r, c337_a, c340_r, c340_a, c343_r, c343_a, c345_r, c345_a, initialise);
  BrzF_0_l87__28_280_200_29_20_280_200_29_20_m36m I384 (c344_r, c344_a, c327_r, c327_a, c330_r, c330_a, c333_r, c333_a, c336_r, c336_a, c339_r, c339_a, c341_r, c341_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I385 (c341_r, c341_a, c342_r0d, c342_r1d, c342_a);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I386 (c327_r, c327_a, c320_r, c320_a, c322_r, c322_a, c325_r, c325_a, initialise);
  BrzJ_l12__2834_201_29 I387 (c323_r0d, c323_r1d, c323_a, c324_r0d, c324_r1d, c324_a, c326_r0d, c326_r1d, c326_a, initialise);
  BrzJ_l12__2833_201_29 I388 (c319_r0d, c319_r1d, c319_a, c321_r0d, c321_r1d, c321_a, c323_r0d, c323_r1d, c323_a, initialise);
  BrzJ_l35__280_200_200_200_200_200_200_200__m45m I389 (c226_r, c226_a, c229_r, c229_a, c231_r, c231_a, c236_r, c236_a, c242_r, c242_a, c273_r, c273_a, c300_r, c300_a, c313_r, c313_a, c318_r, c318_a, initialise);
  BrzF_0_l115__28_280_200_29_20_280_200_29_2_m38m I390 (c317_r, c317_a, c225_r, c225_a, c228_r, c228_a, c234_r, c234_a, c239_r, c239_a, c241_r, c241_a, c244_r, c244_a, c311_r, c311_a, c316_r, c316_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I391 (c314_r0d, c314_r1d, c314_a, c315_r, c315_a, c315_r, c315_a, c312_r0d, c312_r1d, c312_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I392 (c311_r, c311_a, c308_r, c308_a, c309_r, c309_a, c310_r, c310_a, initialise);
  BrzJ_l15__280_200_200_29 I393 (c302_r, c302_a, c304_r, c304_a, c306_r, c306_a, c307_r, c307_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I394 (c305_r0d, c305_r1d, c305_a, c306_r, c306_a, c281_r, c281_a, c280_r0d, c280_r1d, c280_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m88m I395 (c303_r0d, c303_r1d, c303_a, c304_r, c304_a, c275_r, c275_a, c284_r, c284_a, c274_r0d, c274_r1d, c274_a, c283_r0d, c283_r1d, c283_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m93m I396 (c301_r0d, c301_r1d, c301_a, c302_r, c302_a, c290_r, c290_a, c296_r, c296_a, c289_r0d, c289_r1d, c289_a, c295_r0d, c295_r1d, c295_a, initialise);
  BrzJ_l19__280_200_200_200_29 I397 (c276_r, c276_a, c287_r, c287_a, c291_r, c291_a, c299_r, c299_a, c300_r, c300_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I398 (c307_r, c307_a, c275_r, c275_a, c286_r, c286_a, c290_r, c290_a, c298_r, c298_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I399 (c298_r, c298_a, c294_r, c294_a, c296_r, c296_a, initialise);
  BrzO_35_36_l76__28_28num_201_200_29_20_28a_m56m I400 (c297_r0d, c297_r1d, c297_a, c292_r0d, c292_r1d, c292_a);
  BrzJ_l12__2832_203_29 I401 (c293_r0d, c293_r1d, c293_a, c295_r0d, c295_r1d, c295_a, c297_r0d, c297_r1d, c297_a, initialise);
  BrzO_32_35_l91__28_28app_203_20_280_2031_2_m50m I402 (c289_r0d, c289_r1d, c289_a, c288_r0d, c288_r1d, c288_a);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I403 (c286_r, c286_a, c279_r, c279_a, c281_r, c281_a, c284_r, c284_a, initialise);
  BrzO_35_36_l76__28_28num_201_200_29_20_28a_m56m I404 (c285_r0d, c285_r1d, c285_a, c277_r0d, c277_r1d, c277_a);
  BrzJ_l12__2833_202_29 I405 (c282_r0d, c282_r1d, c282_a, c283_r0d, c283_r1d, c283_a, c285_r0d, c285_r1d, c285_a, initialise);
  BrzJ_l12__2832_201_29 I406 (c278_r0d, c278_r1d, c278_a, c280_r0d, c280_r1d, c280_a, c282_r0d, c282_r1d, c282_a, initialise);
  BrzM_0_9 I407 (c248_r, c248_a, c251_r, c251_a, c254_r, c254_a, c257_r, c257_a, c260_r, c260_a, c263_r, c263_a, c266_r, c266_a, c269_r, c269_a, c272_r, c272_a, c273_r, c273_a, initialise);
  BrzS_4_l11__280_204_29_l521__28_28_28_280__m66m I408 (c243_r0d, c243_r1d, c243_a, c247_r, c247_a, c250_r, c250_a, c253_r, c253_a, c256_r, c256_a, c259_r, c259_a, c262_r, c262_a, c265_r, c265_a, c268_r, c268_a, c271_r, c271_a, initialise);
  BrzO_4_35_l91__28_28app_2031_20_280_203_20_m48m I409 (c246_r0d, c246_r1d, c246_a, c245_r0d, c245_r1d, c245_a);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I410 (c237_r0d, c237_r1d, c237_a, c238_r, c238_a, c238_r, c238_a, c235_r0d, c235_r1d, c235_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I411 (c232_r0d, c232_r1d, c232_a, c233_r, c233_a, c233_r, c233_a, c230_r0d, c230_r1d, c230_a, initialise);
  BrzJ_l23__280_200_200_200_200_29 I412 (c206_r, c206_a, c210_r, c210_a, c214_r, c214_a, c218_r, c218_a, c221_r, c221_a, c222_r, c222_a, initialise);
  BrzF_0_l73__28_280_200_29_20_280_200_29_20_m35m I413 (c186_r, c186_a, c205_r, c205_a, c209_r, c209_a, c213_r, c213_a, c217_r, c217_a, c219_r, c219_a, initialise);
  BrzO_0_1_l23__28_28num_201_201_29_29 I414 (c219_r, c219_a, c220_r0d, c220_r1d, c220_a);
  BrzO_35_35_l34__28_28not_20_280_200_2035_2_m55m I415 (c216_r0d, c216_r1d, c216_a, c215_r0d, c215_r1d, c215_a);
  BrzO_35_35_l34__28_28not_20_280_200_2035_2_m55m I416 (c212_r0d, c212_r1d, c212_a, c211_r0d, c211_r1d, c211_a);
  BrzO_35_35_l34__28_28not_20_280_200_2035_2_m55m I417 (c208_r0d, c208_r1d, c208_a, c207_r0d, c207_r1d, c207_a);
  BrzO_35_35_l34__28_28not_20_280_200_2035_2_m55m I418 (c204_r0d, c204_r1d, c204_a, c203_r0d, c203_r1d, c203_a);
  BrzF_0_l73__28_280_200_29_20_280_200_29_20_m35m I419 (c118_r, c118_a, c198_r, c198_a, c199_r, c199_a, c200_r, c200_a, c201_r, c201_a, c202_r, c202_a, initialise);
  BrzJ_l23__280_200_200_200_200_29 I420 (c188_r, c188_a, c190_r, c190_a, c192_r, c192_a, c194_r, c194_a, c196_r, c196_a, c197_r, c197_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I421 (c195_r0d, c195_r1d, c195_a, c196_r, c196_a, c123_r, c123_a, c122_r0d, c122_r1d, c122_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I422 (c193_r0d, c193_r1d, c193_a, c194_r, c194_a, c120_r, c120_a, c119_r0d, c119_r1d, c119_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m87m I423 (c191_r0d, c191_r1d, c191_a, c192_r, c192_a, c175_r, c175_a, c174_r0d, c174_r1d, c174_a, initialise);
  BrzV_36_l6__28_29_l24__28_28_280_2036_29_2_m95m I424 (c189_r0d, c189_r1d, c189_a, c190_r, c190_a, c172_r, c172_a, c178_r, c178_a, c171_r0d, c171_r1d, c171_a, c177_r0d, c177_r1d, c177_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m89m I425 (c187_r0d, c187_r1d, c187_a, c188_r, c188_a, c126_r, c126_a, c131_r, c131_a, c138_r, c138_a, c143_r, c143_a, c146_r, c146_a, c152_r, c152_a, c160_r, c160_a, c125_r0d, c125_r1d, c125_a, c130_r0d, c130_r1d, c130_a, c137_r0d, c137_r1d, c137_a, c142_r0d, c142_r1d, c142_a, c145_r0d, c145_r1d, c145_a, c151_r0d, c151_r1d, c151_a, c159_r0d, c159_r1d, c159_a, initialise);
  BrzJ_l59__280_200_200_200_200_200_200_200__m46m I426 (c121_r, c121_a, c124_r, c124_a, c127_r, c127_a, c134_r, c134_a, c141_r, c141_a, c144_r, c144_a, c147_r, c147_a, c150_r, c150_a, c162_r, c162_a, c173_r, c173_a, c176_r, c176_a, c179_r, c179_a, c182_r, c182_a, c185_r, c185_a, c186_r, c186_a, initialise);
  BrzF_0_l199__28_280_200_29_20_280_200_29_2_m39m I427 (c197_r, c197_a, c120_r, c120_a, c123_r, c123_a, c126_r, c126_a, c133_r, c133_a, c140_r, c140_a, c143_r, c143_a, c146_r, c146_a, c148_r, c148_a, c170_r, c170_a, c172_r, c172_a, c175_r, c175_a, c178_r, c178_a, c180_r, c180_a, c183_r, c183_a, initialise);
  BrzO_0_36_l24__28_28num_2036_200_29_29 I428 (c183_r, c183_a, c184_r0d, c184_r1d, c184_a);
  BrzO_0_35_l24__28_28num_2035_200_29_29 I429 (c180_r, c180_a, c181_r0d, c181_r1d, c181_a);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I430 (c170_r, c170_a, c168_r, c168_a, c169_r, c169_a, initialise);
  BrzJ_l11__280_200_29 I431 (c164_r, c164_a, c166_r, c166_a, c167_r, c167_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m71m I432 (c165_r0d, c165_r1d, c165_a, c166_r, c166_a, c157_r, c157_a, c156_r0d, c156_r1d, c156_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I433 (c163_r0d, c163_r1d, c163_a, c164_r, c164_a, c154_r, c154_a, c153_r0d, c153_r1d, c153_a, initialise);
  BrzF_0_l59__28_280_200_29_20_280_200_29_20_m34m I434 (c167_r, c167_a, c152_r, c152_a, c154_r, c154_a, c157_r, c157_a, c160_r, c160_a, initialise);
  BrzJ_l12__2834_201_29 I435 (c158_r0d, c158_r1d, c158_a, c159_r0d, c159_r1d, c159_a, c161_r0d, c161_r1d, c161_a, initialise);
  BrzJ_l12__2833_201_29 I436 (c155_r0d, c155_r1d, c155_a, c156_r0d, c156_r1d, c156_a, c158_r0d, c158_r1d, c158_a, initialise);
  BrzJ_l12__281_2032_29 I437 (c151_r0d, c151_r1d, c151_a, c153_r0d, c153_r1d, c153_a, c155_r0d, c155_r1d, c155_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I438 (c148_r, c148_a, c149_r0d, c149_r1d, c149_a);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I439 (c140_r, c140_a, c135_r, c135_a, c138_r, c138_a, initialise);
  BrzJ_l12__282_2033_29 I440 (c136_r0d, c136_r1d, c136_a, c137_r0d, c137_r1d, c137_a, c139_r0d, c139_r1d, c139_a, initialise);
  BrzO_0_2_l23__28_28num_202_200_29_29 I441 (c135_r, c135_a, c136_r0d, c136_r1d, c136_a);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I442 (c133_r, c133_a, c128_r, c128_a, c131_r, c131_a, initialise);
  BrzJ_l12__281_2034_29 I443 (c129_r0d, c129_r1d, c129_a, c130_r0d, c130_r1d, c130_a, c132_r0d, c132_r1d, c132_a, initialise);
  BrzO_0_1_l23__28_28num_201_200_29_29 I444 (c128_r, c128_a, c129_r0d, c129_r1d, c129_a);
  BrzJ_l12__2833_200_29 I445 (c117_r0d, c117_r1d, c117_a, c99_r, c99_a, c94_r0d, c94_r1d, c94_a, initialise);
  BrzF_33_l32__28_280_200_29_20_280_2033_29__m41m I446 (c65_r0d, c65_r1d, c65_a, c67_r, c67_a, c117_r0d, c117_r1d, c117_a, initialise);
  BrzJ_l12__2833_200_29 I447 (c116_r0d, c116_r1d, c116_a, c100_r, c100_a, c96_r0d, c96_r1d, c96_a, initialise);
  BrzF_33_l32__28_280_200_29_20_280_2033_29__m41m I448 (c72_r0d, c72_r1d, c72_a, c74_r, c74_a, c116_r0d, c116_r1d, c116_a, initialise);
  BrzJ_l12__2834_200_29 I449 (c115_r0d, c115_r1d, c115_a, c111_r, c111_a, c109_r0d, c109_r1d, c109_a, initialise);
  BrzF_34_l32__28_280_200_29_20_280_2034_29__m42m I450 (c92_r0d, c92_r1d, c92_a, c93_r, c93_a, c115_r0d, c115_r1d, c115_a, initialise);
  BrzM_0_2 I451 (c114_r, c114_a, c113_r, c113_a, c112_r, c112_a, initialise);
  BrzJ_l15__280_200_200_29 I452 (c75_r, c75_a, c93_r, c93_a, c108_r, c108_a, c113_r, c113_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I453 (c112_r, c112_a, c86_r, c86_a, c101_r, c101_a, c111_r, c111_a, initialise);
  BrzV_34_l6__28_29_l24__28_28_280_2034_29_2_m85m I454 (c109_r0d, c109_r1d, c109_a, c110_r, c110_a, c103_r, c103_a, c106_r, c106_a, c102_r0d, c102_r1d, c102_a, c105_r0d, c105_r1d, c105_a, initialise);
  BrzJ_l11__280_200_29 I455 (c104_r, c104_a, c107_r, c107_a, c108_r, c108_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I456 (c110_r, c110_a, c103_r, c103_a, c106_r, c106_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I457 (c101_r, c101_a, c99_r, c99_a, c100_r, c100_a, initialise);
  BrzJ_l11__280_200_29 I458 (c95_r, c95_a, c97_r, c97_a, c98_r, c98_a, initialise);
  BrzV_33_l6__28_29_l24__28_28_280_2033_29_2_m84m I459 (c96_r0d, c96_r1d, c96_a, c97_r, c97_a, c90_r, c90_a, c89_r0d, c89_r1d, c89_a, initialise);
  BrzV_33_l6__28_29_l24__28_28_280_2033_29_2_m84m I460 (c94_r0d, c94_r1d, c94_a, c95_r, c95_a, c88_r, c88_a, c87_r0d, c87_r1d, c87_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I461 (c98_r, c98_a, c88_r, c88_a, c90_r, c90_a, initialise);
  BrzO_66_34_l270__28_28app_201_20_280_200_2_m57m I462 (c91_r0d, c91_r1d, c91_a, c92_r0d, c92_r1d, c92_a);
  BrzJ_l13__2833_2033_29 I463 (c87_r0d, c87_r1d, c87_a, c89_r0d, c89_r1d, c89_a, c91_r0d, c91_r1d, c91_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I464 (c86_r, c86_a, c83_r, c83_a, c84_r, c84_a, c85_r, c85_a, initialise);
  BrzJ_l15__280_200_200_29 I465 (c77_r, c77_a, c79_r, c79_a, c81_r, c81_a, c82_r, c82_a, initialise);
  BrzV_1_l6__28_29_l23__28_28_280_201_29_29__m72m I466 (c80_r0d, c80_r1d, c80_a, c81_r, c81_a, c62_r, c62_a, c69_r, c69_a, c61_r0d, c61_r1d, c61_a, c68_r0d, c68_r1d, c68_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I467 (c78_r0d, c78_r1d, c78_a, c79_r, c79_a, c71_r, c71_a, c70_r0d, c70_r1d, c70_a, initialise);
  BrzV_32_l6__28_29_l24__28_28_280_2032_29_2_m80m I468 (c76_r0d, c76_r1d, c76_a, c77_r, c77_a, c64_r, c64_a, c63_r0d, c63_r1d, c63_a, initialise);
  BrzJ_l11__280_200_29 I469 (c67_r, c67_a, c74_r, c74_a, c75_r, c75_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I470 (c82_r, c82_a, c66_r, c66_a, c73_r, c73_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I471 (c73_r, c73_a, c69_r, c69_a, c71_r, c71_a, initialise);
  BrzJ_l12__281_2032_29 I472 (c68_r0d, c68_r1d, c68_a, c70_r0d, c70_r1d, c70_a, c72_r0d, c72_r1d, c72_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I473 (c66_r, c66_a, c62_r, c62_a, c64_r, c64_a, initialise);
  BrzJ_l12__281_2032_29 I474 (c61_r0d, c61_r1d, c61_a, c63_r0d, c63_r1d, c63_a, c65_r0d, c65_r1d, c65_a, initialise);
  BrzM_0_2 I475 (c60_r, c60_a, c48_r, c48_a, c59_r, c59_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I476 (c59_r, c59_a, c56_r, c56_a, c57_r, c57_a, c58_r, c58_a, initialise);
  BrzJ_l15__280_200_200_29 I477 (c50_r, c50_a, c52_r, c52_a, c54_r, c54_a, c55_r, c55_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m91m I478 (c53_r0d, c53_r1d, c53_a, c54_r, c54_a, c19_r, c19_a, c31_r, c31_a, c39_r, c39_a, c18_r0d, c18_r1d, c18_a, c30_r0d, c30_r1d, c30_a, c38_r0d, c38_r1d, c38_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m91m I479 (c51_r0d, c51_r1d, c51_a, c52_r, c52_a, c15_r, c15_a, c27_r, c27_a, c41_r, c41_a, c14_r0d, c14_r1d, c14_a, c26_r0d, c26_r1d, c26_a, c40_r0d, c40_r1d, c40_a, initialise);
  BrzV_35_l6__28_29_l24__28_28_280_2035_29_2_m91m I480 (c49_r0d, c49_r1d, c49_a, c50_r, c50_a, c13_r, c13_a, c25_r, c25_a, c33_r, c33_a, c12_r0d, c12_r1d, c12_a, c24_r0d, c24_r1d, c24_a, c32_r0d, c32_r1d, c32_a, initialise);
  BrzJ_l11__280_200_29 I481 (c23_r, c23_a, c47_r, c47_a, c48_r, c48_a, initialise);
  BrzF_0_l31__28_280_200_29_20_280_200_29_29 I482 (c55_r, c55_a, c22_r, c22_a, c46_r, c46_a, initialise);
  BrzF_0_l87__28_280_200_29_20_280_200_29_20_m36m I483 (c46_r, c46_a, c25_r, c25_a, c27_r, c27_a, c31_r, c31_a, c33_r, c33_a, c39_r, c39_a, c41_r, c41_a, initialise);
  BrzO_70_35_l123__28_28app_201_20_280_200_2_m59m I484 (c44_r0d, c44_r1d, c44_a, c45_r0d, c45_r1d, c45_a);
  BrzJ_l13__2835_2035_29 I485 (c37_r0d, c37_r1d, c37_a, c43_r0d, c43_r1d, c43_a, c44_r0d, c44_r1d, c44_a, initialise);
  BrzO_70_35_l124__28_28app_201_20_280_200_2_m58m I486 (c42_r0d, c42_r1d, c42_a, c43_r0d, c43_r1d, c43_a);
  BrzJ_l13__2835_2035_29 I487 (c38_r0d, c38_r1d, c38_a, c40_r0d, c40_r1d, c40_a, c42_r0d, c42_r1d, c42_a, initialise);
  BrzO_70_35_l123__28_28app_201_20_280_200_2_m59m I488 (c36_r0d, c36_r1d, c36_a, c37_r0d, c37_r1d, c37_a);
  BrzJ_l13__2835_2035_29 I489 (c29_r0d, c29_r1d, c29_a, c35_r0d, c35_r1d, c35_a, c36_r0d, c36_r1d, c36_a, initialise);
  BrzO_70_35_l124__28_28app_201_20_280_200_2_m58m I490 (c34_r0d, c34_r1d, c34_a, c35_r0d, c35_r1d, c35_a);
  BrzJ_l13__2835_2035_29 I491 (c30_r0d, c30_r1d, c30_a, c32_r0d, c32_r1d, c32_a, c34_r0d, c34_r1d, c34_a, initialise);
  BrzO_70_35_l124__28_28app_201_20_280_200_2_m58m I492 (c28_r0d, c28_r1d, c28_a, c29_r0d, c29_r1d, c29_a);
  BrzJ_l13__2835_2035_29 I493 (c24_r0d, c24_r1d, c24_a, c26_r0d, c26_r1d, c26_a, c28_r0d, c28_r1d, c28_a, initialise);
  BrzF_0_l45__28_280_200_29_20_280_200_29_20_m33m I494 (c22_r, c22_a, c13_r, c13_a, c15_r, c15_a, c19_r, c19_a, initialise);
  BrzO_70_35_l124__28_28app_201_20_280_200_2_m60m I495 (c20_r0d, c20_r1d, c20_a, c21_r0d, c21_r1d, c21_a);
  BrzJ_l13__2835_2035_29 I496 (c17_r0d, c17_r1d, c17_a, c18_r0d, c18_r1d, c18_a, c20_r0d, c20_r1d, c20_a, initialise);
  BrzO_70_35_l124__28_28app_201_20_280_200_2_m60m I497 (c16_r0d, c16_r1d, c16_a, c17_r0d, c17_r1d, c17_a);
  BrzJ_l13__2835_2035_29 I498 (c12_r0d, c12_r1d, c12_a, c14_r0d, c14_r1d, c14_a, c16_r0d, c16_r1d, c16_a, initialise);
endmodule

