//
// by teak gui
//
// Generated on: Thu Oct 18 12:43:35 BST 2012
//


`timescale 1ns/1ps

// tko0m1_1nm1b0 TeakO [
//     (1,TeakOConstant 1 0)] [One 0,One 1]
module tko0m1_1nm1b0 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0, i_0r);
  GND I1 (o_0r1);
  BUFF I2 (i_0a, o_0a);
endmodule

// tkvdoFetchI1_wo0w1_ro0w1 TeakV "doFetchI" 1 [] [0] [0] [Many [1],Many [0],Many [0],Many [1]]
module tkvdoFetchI1_wo0w1_ro0w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input wg_0r0;
  input wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  input reset;
  wire wf_0;
  wire wt_0;
  wire df_0;
  wire dt_0;
  wire wc_0;
  wire wacks_0;
  wire wenr_0;
  wire wen_0;
  wire anyread_0;
  wire nreset_0;
  wire drlgf_0;
  wire drlgt_0;
  wire comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire conwgit_0;
  wire conwgif_0;
  wire conwig_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0, wenr_0, nreset_0);
  AND2 I2 (drlgf_0, wf_0, wen_0);
  AND2 I3 (drlgt_0, wt_0, wen_0);
  NOR2 I4 (df_0, dt_0, drlgt_0);
  NOR3 I5 (dt_0, df_0, drlgf_0, reset);
  AO22 I6 (wacks_0, drlgf_0, df_0, drlgt_0, dt_0);
  OR2 I7 (comp0_0, wg_0r0, wg_0r1);
  BUFF I8 (wc_0, comp0_0);
  AND2 I9 (conwgif_0, wg_0r0, conwig_0);
  AND2 I10 (conwgit_0, wg_0r1, conwig_0);
  BUFF I11 (conwigc_0, wc_0);
  AO22 I12 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I13 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I14 (wf_0, conwgif_0);
  BUFF I15 (wt_0, conwgit_0);
  BUFF I16 (wenr_0, wc_0);
  C2 I17 (wd_0r, conwig_0, wacks_0);
  AND2 I18 (rd_0r0, df_0, rg_0r);
  AND2 I19 (rd_0r1, dt_0, rg_0r);
  OR2 I20 (anyread_0, rg_0r, rg_0a);
  BUFF I21 (wg_0a, wd_0a);
  BUFF I22 (rg_0a, rd_0a);
endmodule

// tkm2x0b TeakM [Many [0,0],One 0]
module tkm2x0b (i_0r, i_0a, i_1r, i_1a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  output o_0r;
  input o_0a;
  input reset;
  wire nchosen_0;
  wire choice_0;
  wire choice_1;
  C2R I0 (choice_0, i_0r, nchosen_0, reset);
  C2R I1 (choice_1, i_1r, nchosen_0, reset);
  NOR2 I2 (nchosen_0, o_0r, o_0a);
  OR2 I3 (o_0r, choice_0, choice_1);
  C2R I4 (i_0a, choice_0, o_0a, reset);
  C2R I5 (i_1a, choice_1, o_0a, reset);
endmodule

// tkj1m1_0 TeakJ [Many [1,0],One 1]
module tkj1m1_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire joinf_0;
  wire joint_0;
  BUFF I0 (joinf_0, i_0r0);
  BUFF I1 (joint_0, i_0r1);
  BUFF I2 (icomplete_0, i_1r);
  C2 I3 (o_0r0, joinf_0, icomplete_0);
  C2 I4 (o_0r1, joint_0, icomplete_0);
  BUFF I5 (i_0a, o_0a);
  BUFF I6 (i_1a, o_0a);
endmodule

// tkf1mo0w0_o0w1 TeakF [0,0] [One 1,Many [0,1]]
module tkf1mo0w0_o0w1 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r0;
  output o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0, i_0r1);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_1r0, i_0r0);
  BUFF I3 (o_1r1, i_0r1);
  BUFF I4 (o_0r, icomplete_0);
  C3 I5 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tkm3x1b TeakM [Many [1,1,1],One 1]
module tkm3x1b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input i_1r0;
  input i_1r1;
  output i_1a;
  input i_2r0;
  input i_2r1;
  output i_2a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire gfint_0;
  wire gfint_1;
  wire gfint_2;
  wire gtint_0;
  wire gtint_1;
  wire gtint_2;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire nchosen_0;
  wire comp0_0;
  wire comp1_0;
  wire comp2_0;
  OR3 I0 (o_0r0, gfint_0, gfint_1, gfint_2);
  OR3 I1 (o_0r1, gtint_0, gtint_1, gtint_2);
  AND2 I2 (gtint_0, choice_0, i_0r1);
  AND2 I3 (gtint_1, choice_1, i_1r1);
  AND2 I4 (gtint_2, choice_2, i_2r1);
  AND2 I5 (gfint_0, choice_0, i_0r0);
  AND2 I6 (gfint_1, choice_1, i_1r0);
  AND2 I7 (gfint_2, choice_2, i_2r0);
  OR2 I8 (comp0_0, i_0r0, i_0r1);
  BUFF I9 (icomp_0, comp0_0);
  OR2 I10 (comp1_0, i_1r0, i_1r1);
  BUFF I11 (icomp_1, comp1_0);
  OR2 I12 (comp2_0, i_2r0, i_2r1);
  BUFF I13 (icomp_2, comp2_0);
  C2R I14 (choice_0, icomp_0, nchosen_0, reset);
  C2R I15 (choice_1, icomp_1, nchosen_0, reset);
  C2R I16 (choice_2, icomp_2, nchosen_0, reset);
  OR3 I17 (anychoice_0, choice_0, choice_1, choice_2);
  NOR2 I18 (nchosen_0, anychoice_0, o_0a);
  C2R I19 (i_0a, choice_0, o_0a, reset);
  C2R I20 (i_1a, choice_1, o_0a, reset);
  C2R I21 (i_2a, choice_2, o_0a, reset);
endmodule

// tko0m3_1nm3b1 TeakO [
//     (1,TeakOConstant 3 1)] [One 0,One 3]
module tko0m3_1nm3b1 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  GND I1 (o_0r0[0:0]);
  BUFF I2 (o_0r0[1:1], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  GND I4 (o_0r1[1:1]);
  GND I5 (o_0r1[2:2]);
  BUFF I6 (i_0a, o_0a);
endmodule

// tko0m3_1nm3b2 TeakO [
//     (1,TeakOConstant 3 2)] [One 0,One 3]
module tko0m3_1nm3b2 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[1:1], i_0r);
  GND I1 (o_0r0[1:1]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  GND I4 (o_0r1[0:0]);
  GND I5 (o_0r1[2:2]);
  BUFF I6 (i_0a, o_0a);
endmodule

// tko0m3_1nm3b4 TeakO [
//     (1,TeakOConstant 3 4)] [One 0,One 3]
module tko0m3_1nm3b4 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[2:2], i_0r);
  GND I1 (o_0r0[2:2]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  GND I4 (o_0r1[0:0]);
  GND I5 (o_0r1[1:1]);
  BUFF I6 (i_0a, o_0a);
endmodule

// tkm3x3b TeakM [Many [3,3,3],One 3]
module tkm3x3b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, o_0r0, o_0r1, o_0a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  input [2:0] i_1r0;
  input [2:0] i_1r1;
  output i_1a;
  input [2:0] i_2r0;
  input [2:0] i_2r1;
  output i_2a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire [2:0] gfint_0;
  wire [2:0] gfint_1;
  wire [2:0] gfint_2;
  wire [2:0] gtint_0;
  wire [2:0] gtint_1;
  wire [2:0] gtint_2;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire nchosen_0;
  wire [2:0] comp0_0;
  wire [2:0] comp1_0;
  wire [2:0] comp2_0;
  OR3 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  OR3 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  OR3 I2 (o_0r0[2:2], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  OR3 I3 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  OR3 I4 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  OR3 I5 (o_0r1[2:2], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  AND2 I6 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I7 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I8 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I9 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I10 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I11 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I12 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I13 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I14 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I15 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I16 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I17 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I18 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I19 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I20 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I21 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I22 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I23 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  OR2 I24 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I25 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I26 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I27 (icomp_0, comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  OR2 I28 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I29 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I30 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  C3 I31 (icomp_1, comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  OR2 I32 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I33 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I34 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  C3 I35 (icomp_2, comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C2R I36 (choice_0, icomp_0, nchosen_0, reset);
  C2R I37 (choice_1, icomp_1, nchosen_0, reset);
  C2R I38 (choice_2, icomp_2, nchosen_0, reset);
  OR3 I39 (anychoice_0, choice_0, choice_1, choice_2);
  NOR2 I40 (nchosen_0, anychoice_0, o_0a);
  C2R I41 (i_0a, choice_0, o_0a, reset);
  C2R I42 (i_1a, choice_1, o_0a, reset);
  C2R I43 (i_2a, choice_2, o_0a, reset);
endmodule

// tkj3m0_3 TeakJ [Many [0,3],One 3]
module tkj3m0_3 (i_0r, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  input [2:0] i_1r0;
  input [2:0] i_1r1;
  output i_1a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [2:0] joinf_0;
  wire [2:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_1r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_1r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_1r0[2:2]);
  BUFF I3 (joint_0[0:0], i_1r1[0:0]);
  BUFF I4 (joint_0[1:1], i_1r1[1:1]);
  BUFF I5 (joint_0[2:2], i_1r1[2:2]);
  BUFF I6 (icomplete_0, i_0r);
  C2 I7 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I8 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I9 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I10 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I11 (o_0r1[1:1], joint_0[1:1]);
  BUFF I12 (o_0r1[2:2], joint_0[2:2]);
  BUFF I13 (i_0a, o_0a);
  BUFF I14 (i_1a, o_0a);
endmodule

// tks3_o0w3_1o0w0_2o0w0_4o0w0 TeakS (0+:3) [([Imp 1 0],0),([Imp 2 0],0),([Imp 4 0],0)] [One 3,Many [0,
//   0,0]]
module tks3_o0w3_1o0w0_2o0w0_4o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire match2_0;
  wire [2:0] comp_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (match0_0, i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I2 (sel_1, match1_0);
  C3 I3 (match1_0, i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I4 (sel_2, match2_0);
  C3 I5 (match2_0, i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C2 I6 (gsel_0, sel_0, icomplete_0);
  C2 I7 (gsel_1, sel_1, icomplete_0);
  C2 I8 (gsel_2, sel_2, icomplete_0);
  OR2 I9 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I10 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I11 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I12 (icomplete_0, comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  BUFF I13 (o_0r, gsel_0);
  BUFF I14 (o_1r, gsel_1);
  BUFF I15 (o_2r, gsel_2);
  OR3 I16 (oack_0, o_0a, o_1a, o_2a);
  C2 I17 (i_0a, oack_0, icomplete_0);
endmodule

// tkr TeakR [One 0]
module tkr (o_0r, o_0a, reset);
  output o_0r;
  input o_0a;
  input reset;
  wire fb1_0;
  wire fb2_0;
  NOR2 I0 (fb1_0, reset, fb2_0);
  NOR2 I1 (fb2_0, o_0a, fb1_0);
  NOR2 I2 (o_0r, reset, fb1_0);
endmodule

// tko0m32_1nm32b0 TeakO [
//     (1,TeakOConstant 32 0)] [One 0,One 32]
module tko0m32_1nm32b0 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r);
  BUFF I1 (o_0r0[1:1], i_0r);
  BUFF I2 (o_0r0[2:2], i_0r);
  BUFF I3 (o_0r0[3:3], i_0r);
  BUFF I4 (o_0r0[4:4], i_0r);
  BUFF I5 (o_0r0[5:5], i_0r);
  BUFF I6 (o_0r0[6:6], i_0r);
  BUFF I7 (o_0r0[7:7], i_0r);
  BUFF I8 (o_0r0[8:8], i_0r);
  BUFF I9 (o_0r0[9:9], i_0r);
  BUFF I10 (o_0r0[10:10], i_0r);
  BUFF I11 (o_0r0[11:11], i_0r);
  BUFF I12 (o_0r0[12:12], i_0r);
  BUFF I13 (o_0r0[13:13], i_0r);
  BUFF I14 (o_0r0[14:14], i_0r);
  BUFF I15 (o_0r0[15:15], i_0r);
  BUFF I16 (o_0r0[16:16], i_0r);
  BUFF I17 (o_0r0[17:17], i_0r);
  BUFF I18 (o_0r0[18:18], i_0r);
  BUFF I19 (o_0r0[19:19], i_0r);
  BUFF I20 (o_0r0[20:20], i_0r);
  BUFF I21 (o_0r0[21:21], i_0r);
  BUFF I22 (o_0r0[22:22], i_0r);
  BUFF I23 (o_0r0[23:23], i_0r);
  BUFF I24 (o_0r0[24:24], i_0r);
  BUFF I25 (o_0r0[25:25], i_0r);
  BUFF I26 (o_0r0[26:26], i_0r);
  BUFF I27 (o_0r0[27:27], i_0r);
  BUFF I28 (o_0r0[28:28], i_0r);
  BUFF I29 (o_0r0[29:29], i_0r);
  BUFF I30 (o_0r0[30:30], i_0r);
  BUFF I31 (o_0r0[31:31], i_0r);
  GND I32 (o_0r1[0:0]);
  GND I33 (o_0r1[1:1]);
  GND I34 (o_0r1[2:2]);
  GND I35 (o_0r1[3:3]);
  GND I36 (o_0r1[4:4]);
  GND I37 (o_0r1[5:5]);
  GND I38 (o_0r1[6:6]);
  GND I39 (o_0r1[7:7]);
  GND I40 (o_0r1[8:8]);
  GND I41 (o_0r1[9:9]);
  GND I42 (o_0r1[10:10]);
  GND I43 (o_0r1[11:11]);
  GND I44 (o_0r1[12:12]);
  GND I45 (o_0r1[13:13]);
  GND I46 (o_0r1[14:14]);
  GND I47 (o_0r1[15:15]);
  GND I48 (o_0r1[16:16]);
  GND I49 (o_0r1[17:17]);
  GND I50 (o_0r1[18:18]);
  GND I51 (o_0r1[19:19]);
  GND I52 (o_0r1[20:20]);
  GND I53 (o_0r1[21:21]);
  GND I54 (o_0r1[22:22]);
  GND I55 (o_0r1[23:23]);
  GND I56 (o_0r1[24:24]);
  GND I57 (o_0r1[25:25]);
  GND I58 (o_0r1[26:26]);
  GND I59 (o_0r1[27:27]);
  GND I60 (o_0r1[28:28]);
  GND I61 (o_0r1[29:29]);
  GND I62 (o_0r1[30:30]);
  GND I63 (o_0r1[31:31]);
  BUFF I64 (i_0a, o_0a);
endmodule

// tko0m1_1nm1b1 TeakO [
//     (1,TeakOConstant 1 1)] [One 0,One 1]
module tko0m1_1nm1b1 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1, i_0r);
  GND I1 (o_0r0);
  BUFF I2 (i_0a, o_0a);
endmodule

// tkj0m0_0 TeakJ [Many [0,0],One 0]
module tkj0m0_0 (i_0r, i_0a, i_1r, i_1a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  output o_0r;
  input o_0a;
  input reset;
  C2 I0 (o_0r, i_0r, i_1r);
  BUFF I1 (i_0a, o_0a);
  BUFF I2 (i_1a, o_0a);
endmodule

// tkf0mo0w0_o0w0 TeakF [0,0] [One 0,Many [0,0]]
module tkf0mo0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  C2 I2 (i_0a, o_0a, o_1a);
endmodule

// tkvnewPc32_wo0w32_ro0w32 TeakV "newPc" 32 [] [0] [0] [Many [32],Many [0],Many [0],Many [32]]
module tkvnewPc32_wo0w32_ro0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I457 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I458 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I459 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I460 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I461 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I462 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I463 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I464 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I465 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I466 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I467 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I468 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I469 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I470 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I471 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I472 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I473 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I474 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I475 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I476 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I477 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I478 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I479 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I480 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I481 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I482 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I483 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I484 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I485 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I486 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I487 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  OR2 I488 (anyread_0, rg_0r, rg_0a);
  BUFF I489 (wg_0a, wd_0a);
  BUFF I490 (rg_0a, rd_0a);
endmodule

// tks1_o0w1_0o0w0_1o0w0 TeakS (0+:1) [([Imp 0 0],0),([Imp 1 0],0)] [One 1,Many [0,0]]
module tks1_o0w1_0o0w0_1o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire comp_0;
  BUFF I0 (sel_0, match0_0);
  BUFF I1 (match0_0, i_0r0);
  BUFF I2 (sel_1, match1_0);
  BUFF I3 (match1_0, i_0r1);
  C2 I4 (gsel_0, sel_0, icomplete_0);
  C2 I5 (gsel_1, sel_1, icomplete_0);
  OR2 I6 (comp_0, i_0r0, i_0r1);
  BUFF I7 (icomplete_0, comp_0);
  BUFF I8 (o_0r, gsel_0);
  BUFF I9 (o_1r, gsel_1);
  OR2 I10 (oack_0, o_0a, o_1a);
  C2 I11 (i_0a, oack_0, icomplete_0);
endmodule

// tkvdoFetch1_wo0w1_ro0w1 TeakV "doFetch" 1 [] [0] [0] [Many [1],Many [0],Many [0],Many [1]]
module tkvdoFetch1_wo0w1_ro0w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input wg_0r0;
  input wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  input reset;
  wire wf_0;
  wire wt_0;
  wire df_0;
  wire dt_0;
  wire wc_0;
  wire wacks_0;
  wire wenr_0;
  wire wen_0;
  wire anyread_0;
  wire nreset_0;
  wire drlgf_0;
  wire drlgt_0;
  wire comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire conwgit_0;
  wire conwgif_0;
  wire conwig_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0, wenr_0, nreset_0);
  AND2 I2 (drlgf_0, wf_0, wen_0);
  AND2 I3 (drlgt_0, wt_0, wen_0);
  NOR2 I4 (df_0, dt_0, drlgt_0);
  NOR3 I5 (dt_0, df_0, drlgf_0, reset);
  AO22 I6 (wacks_0, drlgf_0, df_0, drlgt_0, dt_0);
  OR2 I7 (comp0_0, wg_0r0, wg_0r1);
  BUFF I8 (wc_0, comp0_0);
  AND2 I9 (conwgif_0, wg_0r0, conwig_0);
  AND2 I10 (conwgit_0, wg_0r1, conwig_0);
  BUFF I11 (conwigc_0, wc_0);
  AO22 I12 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I13 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I14 (wf_0, conwgif_0);
  BUFF I15 (wt_0, conwgit_0);
  BUFF I16 (wenr_0, wc_0);
  C2 I17 (wd_0r, conwig_0, wacks_0);
  AND2 I18 (rd_0r0, df_0, rg_0r);
  AND2 I19 (rd_0r1, dt_0, rg_0r);
  OR2 I20 (anyread_0, rg_0r, rg_0a);
  BUFF I21 (wg_0a, wd_0a);
  BUFF I22 (rg_0a, rd_0a);
endmodule

// tkj33m32_1 TeakJ [Many [32,1],One 33]
module tkj33m32_1 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input i_1r0;
  input i_1r1;
  output i_1a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [32:0] joinf_0;
  wire [32:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joinf_0[32:32], i_1r0);
  BUFF I33 (joint_0[0:0], i_0r1[0:0]);
  BUFF I34 (joint_0[1:1], i_0r1[1:1]);
  BUFF I35 (joint_0[2:2], i_0r1[2:2]);
  BUFF I36 (joint_0[3:3], i_0r1[3:3]);
  BUFF I37 (joint_0[4:4], i_0r1[4:4]);
  BUFF I38 (joint_0[5:5], i_0r1[5:5]);
  BUFF I39 (joint_0[6:6], i_0r1[6:6]);
  BUFF I40 (joint_0[7:7], i_0r1[7:7]);
  BUFF I41 (joint_0[8:8], i_0r1[8:8]);
  BUFF I42 (joint_0[9:9], i_0r1[9:9]);
  BUFF I43 (joint_0[10:10], i_0r1[10:10]);
  BUFF I44 (joint_0[11:11], i_0r1[11:11]);
  BUFF I45 (joint_0[12:12], i_0r1[12:12]);
  BUFF I46 (joint_0[13:13], i_0r1[13:13]);
  BUFF I47 (joint_0[14:14], i_0r1[14:14]);
  BUFF I48 (joint_0[15:15], i_0r1[15:15]);
  BUFF I49 (joint_0[16:16], i_0r1[16:16]);
  BUFF I50 (joint_0[17:17], i_0r1[17:17]);
  BUFF I51 (joint_0[18:18], i_0r1[18:18]);
  BUFF I52 (joint_0[19:19], i_0r1[19:19]);
  BUFF I53 (joint_0[20:20], i_0r1[20:20]);
  BUFF I54 (joint_0[21:21], i_0r1[21:21]);
  BUFF I55 (joint_0[22:22], i_0r1[22:22]);
  BUFF I56 (joint_0[23:23], i_0r1[23:23]);
  BUFF I57 (joint_0[24:24], i_0r1[24:24]);
  BUFF I58 (joint_0[25:25], i_0r1[25:25]);
  BUFF I59 (joint_0[26:26], i_0r1[26:26]);
  BUFF I60 (joint_0[27:27], i_0r1[27:27]);
  BUFF I61 (joint_0[28:28], i_0r1[28:28]);
  BUFF I62 (joint_0[29:29], i_0r1[29:29]);
  BUFF I63 (joint_0[30:30], i_0r1[30:30]);
  BUFF I64 (joint_0[31:31], i_0r1[31:31]);
  BUFF I65 (joint_0[32:32], i_1r1);
  OR2 I66 (dcomplete_0, i_1r0, i_1r1);
  BUFF I67 (icomplete_0, dcomplete_0);
  C2 I68 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I69 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I70 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I71 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I72 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I73 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I74 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I75 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I76 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I77 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I78 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I79 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I80 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I81 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I82 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I83 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I84 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I85 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I86 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I87 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I88 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I89 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I90 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I91 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I92 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I93 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I94 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I95 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I96 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I97 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I98 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I99 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I100 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I101 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I102 (o_0r1[1:1], joint_0[1:1]);
  BUFF I103 (o_0r1[2:2], joint_0[2:2]);
  BUFF I104 (o_0r1[3:3], joint_0[3:3]);
  BUFF I105 (o_0r1[4:4], joint_0[4:4]);
  BUFF I106 (o_0r1[5:5], joint_0[5:5]);
  BUFF I107 (o_0r1[6:6], joint_0[6:6]);
  BUFF I108 (o_0r1[7:7], joint_0[7:7]);
  BUFF I109 (o_0r1[8:8], joint_0[8:8]);
  BUFF I110 (o_0r1[9:9], joint_0[9:9]);
  BUFF I111 (o_0r1[10:10], joint_0[10:10]);
  BUFF I112 (o_0r1[11:11], joint_0[11:11]);
  BUFF I113 (o_0r1[12:12], joint_0[12:12]);
  BUFF I114 (o_0r1[13:13], joint_0[13:13]);
  BUFF I115 (o_0r1[14:14], joint_0[14:14]);
  BUFF I116 (o_0r1[15:15], joint_0[15:15]);
  BUFF I117 (o_0r1[16:16], joint_0[16:16]);
  BUFF I118 (o_0r1[17:17], joint_0[17:17]);
  BUFF I119 (o_0r1[18:18], joint_0[18:18]);
  BUFF I120 (o_0r1[19:19], joint_0[19:19]);
  BUFF I121 (o_0r1[20:20], joint_0[20:20]);
  BUFF I122 (o_0r1[21:21], joint_0[21:21]);
  BUFF I123 (o_0r1[22:22], joint_0[22:22]);
  BUFF I124 (o_0r1[23:23], joint_0[23:23]);
  BUFF I125 (o_0r1[24:24], joint_0[24:24]);
  BUFF I126 (o_0r1[25:25], joint_0[25:25]);
  BUFF I127 (o_0r1[26:26], joint_0[26:26]);
  BUFF I128 (o_0r1[27:27], joint_0[27:27]);
  BUFF I129 (o_0r1[28:28], joint_0[28:28]);
  BUFF I130 (o_0r1[29:29], joint_0[29:29]);
  BUFF I131 (o_0r1[30:30], joint_0[30:30]);
  BUFF I132 (o_0r1[31:31], joint_0[31:31]);
  BUFF I133 (o_0r1[32:32], joint_0[32:32]);
  BUFF I134 (i_0a, o_0a);
  BUFF I135 (i_1a, o_0a);
endmodule

// tkj65m32_33 TeakJ [Many [32,33],One 65]
module tkj65m32_33 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [32:0] i_1r0;
  input [32:0] i_1r1;
  output i_1a;
  output [64:0] o_0r0;
  output [64:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [64:0] joinf_0;
  wire [64:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joinf_0[32:32], i_1r0[0:0]);
  BUFF I33 (joinf_0[33:33], i_1r0[1:1]);
  BUFF I34 (joinf_0[34:34], i_1r0[2:2]);
  BUFF I35 (joinf_0[35:35], i_1r0[3:3]);
  BUFF I36 (joinf_0[36:36], i_1r0[4:4]);
  BUFF I37 (joinf_0[37:37], i_1r0[5:5]);
  BUFF I38 (joinf_0[38:38], i_1r0[6:6]);
  BUFF I39 (joinf_0[39:39], i_1r0[7:7]);
  BUFF I40 (joinf_0[40:40], i_1r0[8:8]);
  BUFF I41 (joinf_0[41:41], i_1r0[9:9]);
  BUFF I42 (joinf_0[42:42], i_1r0[10:10]);
  BUFF I43 (joinf_0[43:43], i_1r0[11:11]);
  BUFF I44 (joinf_0[44:44], i_1r0[12:12]);
  BUFF I45 (joinf_0[45:45], i_1r0[13:13]);
  BUFF I46 (joinf_0[46:46], i_1r0[14:14]);
  BUFF I47 (joinf_0[47:47], i_1r0[15:15]);
  BUFF I48 (joinf_0[48:48], i_1r0[16:16]);
  BUFF I49 (joinf_0[49:49], i_1r0[17:17]);
  BUFF I50 (joinf_0[50:50], i_1r0[18:18]);
  BUFF I51 (joinf_0[51:51], i_1r0[19:19]);
  BUFF I52 (joinf_0[52:52], i_1r0[20:20]);
  BUFF I53 (joinf_0[53:53], i_1r0[21:21]);
  BUFF I54 (joinf_0[54:54], i_1r0[22:22]);
  BUFF I55 (joinf_0[55:55], i_1r0[23:23]);
  BUFF I56 (joinf_0[56:56], i_1r0[24:24]);
  BUFF I57 (joinf_0[57:57], i_1r0[25:25]);
  BUFF I58 (joinf_0[58:58], i_1r0[26:26]);
  BUFF I59 (joinf_0[59:59], i_1r0[27:27]);
  BUFF I60 (joinf_0[60:60], i_1r0[28:28]);
  BUFF I61 (joinf_0[61:61], i_1r0[29:29]);
  BUFF I62 (joinf_0[62:62], i_1r0[30:30]);
  BUFF I63 (joinf_0[63:63], i_1r0[31:31]);
  BUFF I64 (joinf_0[64:64], i_1r0[32:32]);
  BUFF I65 (joint_0[0:0], i_0r1[0:0]);
  BUFF I66 (joint_0[1:1], i_0r1[1:1]);
  BUFF I67 (joint_0[2:2], i_0r1[2:2]);
  BUFF I68 (joint_0[3:3], i_0r1[3:3]);
  BUFF I69 (joint_0[4:4], i_0r1[4:4]);
  BUFF I70 (joint_0[5:5], i_0r1[5:5]);
  BUFF I71 (joint_0[6:6], i_0r1[6:6]);
  BUFF I72 (joint_0[7:7], i_0r1[7:7]);
  BUFF I73 (joint_0[8:8], i_0r1[8:8]);
  BUFF I74 (joint_0[9:9], i_0r1[9:9]);
  BUFF I75 (joint_0[10:10], i_0r1[10:10]);
  BUFF I76 (joint_0[11:11], i_0r1[11:11]);
  BUFF I77 (joint_0[12:12], i_0r1[12:12]);
  BUFF I78 (joint_0[13:13], i_0r1[13:13]);
  BUFF I79 (joint_0[14:14], i_0r1[14:14]);
  BUFF I80 (joint_0[15:15], i_0r1[15:15]);
  BUFF I81 (joint_0[16:16], i_0r1[16:16]);
  BUFF I82 (joint_0[17:17], i_0r1[17:17]);
  BUFF I83 (joint_0[18:18], i_0r1[18:18]);
  BUFF I84 (joint_0[19:19], i_0r1[19:19]);
  BUFF I85 (joint_0[20:20], i_0r1[20:20]);
  BUFF I86 (joint_0[21:21], i_0r1[21:21]);
  BUFF I87 (joint_0[22:22], i_0r1[22:22]);
  BUFF I88 (joint_0[23:23], i_0r1[23:23]);
  BUFF I89 (joint_0[24:24], i_0r1[24:24]);
  BUFF I90 (joint_0[25:25], i_0r1[25:25]);
  BUFF I91 (joint_0[26:26], i_0r1[26:26]);
  BUFF I92 (joint_0[27:27], i_0r1[27:27]);
  BUFF I93 (joint_0[28:28], i_0r1[28:28]);
  BUFF I94 (joint_0[29:29], i_0r1[29:29]);
  BUFF I95 (joint_0[30:30], i_0r1[30:30]);
  BUFF I96 (joint_0[31:31], i_0r1[31:31]);
  BUFF I97 (joint_0[32:32], i_1r1[0:0]);
  BUFF I98 (joint_0[33:33], i_1r1[1:1]);
  BUFF I99 (joint_0[34:34], i_1r1[2:2]);
  BUFF I100 (joint_0[35:35], i_1r1[3:3]);
  BUFF I101 (joint_0[36:36], i_1r1[4:4]);
  BUFF I102 (joint_0[37:37], i_1r1[5:5]);
  BUFF I103 (joint_0[38:38], i_1r1[6:6]);
  BUFF I104 (joint_0[39:39], i_1r1[7:7]);
  BUFF I105 (joint_0[40:40], i_1r1[8:8]);
  BUFF I106 (joint_0[41:41], i_1r1[9:9]);
  BUFF I107 (joint_0[42:42], i_1r1[10:10]);
  BUFF I108 (joint_0[43:43], i_1r1[11:11]);
  BUFF I109 (joint_0[44:44], i_1r1[12:12]);
  BUFF I110 (joint_0[45:45], i_1r1[13:13]);
  BUFF I111 (joint_0[46:46], i_1r1[14:14]);
  BUFF I112 (joint_0[47:47], i_1r1[15:15]);
  BUFF I113 (joint_0[48:48], i_1r1[16:16]);
  BUFF I114 (joint_0[49:49], i_1r1[17:17]);
  BUFF I115 (joint_0[50:50], i_1r1[18:18]);
  BUFF I116 (joint_0[51:51], i_1r1[19:19]);
  BUFF I117 (joint_0[52:52], i_1r1[20:20]);
  BUFF I118 (joint_0[53:53], i_1r1[21:21]);
  BUFF I119 (joint_0[54:54], i_1r1[22:22]);
  BUFF I120 (joint_0[55:55], i_1r1[23:23]);
  BUFF I121 (joint_0[56:56], i_1r1[24:24]);
  BUFF I122 (joint_0[57:57], i_1r1[25:25]);
  BUFF I123 (joint_0[58:58], i_1r1[26:26]);
  BUFF I124 (joint_0[59:59], i_1r1[27:27]);
  BUFF I125 (joint_0[60:60], i_1r1[28:28]);
  BUFF I126 (joint_0[61:61], i_1r1[29:29]);
  BUFF I127 (joint_0[62:62], i_1r1[30:30]);
  BUFF I128 (joint_0[63:63], i_1r1[31:31]);
  BUFF I129 (joint_0[64:64], i_1r1[32:32]);
  OR2 I130 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I131 (icomplete_0, dcomplete_0);
  C2 I132 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I133 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I134 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I135 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I136 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I137 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I138 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I139 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I140 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I141 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I142 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I143 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I144 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I145 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I146 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I147 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I148 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I149 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I150 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I151 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I152 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I153 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I154 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I155 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I156 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I157 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I158 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I159 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I160 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I161 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I162 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I163 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I164 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I165 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I166 (o_0r0[33:33], joinf_0[33:33]);
  BUFF I167 (o_0r0[34:34], joinf_0[34:34]);
  BUFF I168 (o_0r0[35:35], joinf_0[35:35]);
  BUFF I169 (o_0r0[36:36], joinf_0[36:36]);
  BUFF I170 (o_0r0[37:37], joinf_0[37:37]);
  BUFF I171 (o_0r0[38:38], joinf_0[38:38]);
  BUFF I172 (o_0r0[39:39], joinf_0[39:39]);
  BUFF I173 (o_0r0[40:40], joinf_0[40:40]);
  BUFF I174 (o_0r0[41:41], joinf_0[41:41]);
  BUFF I175 (o_0r0[42:42], joinf_0[42:42]);
  BUFF I176 (o_0r0[43:43], joinf_0[43:43]);
  BUFF I177 (o_0r0[44:44], joinf_0[44:44]);
  BUFF I178 (o_0r0[45:45], joinf_0[45:45]);
  BUFF I179 (o_0r0[46:46], joinf_0[46:46]);
  BUFF I180 (o_0r0[47:47], joinf_0[47:47]);
  BUFF I181 (o_0r0[48:48], joinf_0[48:48]);
  BUFF I182 (o_0r0[49:49], joinf_0[49:49]);
  BUFF I183 (o_0r0[50:50], joinf_0[50:50]);
  BUFF I184 (o_0r0[51:51], joinf_0[51:51]);
  BUFF I185 (o_0r0[52:52], joinf_0[52:52]);
  BUFF I186 (o_0r0[53:53], joinf_0[53:53]);
  BUFF I187 (o_0r0[54:54], joinf_0[54:54]);
  BUFF I188 (o_0r0[55:55], joinf_0[55:55]);
  BUFF I189 (o_0r0[56:56], joinf_0[56:56]);
  BUFF I190 (o_0r0[57:57], joinf_0[57:57]);
  BUFF I191 (o_0r0[58:58], joinf_0[58:58]);
  BUFF I192 (o_0r0[59:59], joinf_0[59:59]);
  BUFF I193 (o_0r0[60:60], joinf_0[60:60]);
  BUFF I194 (o_0r0[61:61], joinf_0[61:61]);
  BUFF I195 (o_0r0[62:62], joinf_0[62:62]);
  BUFF I196 (o_0r0[63:63], joinf_0[63:63]);
  BUFF I197 (o_0r0[64:64], joinf_0[64:64]);
  BUFF I198 (o_0r1[1:1], joint_0[1:1]);
  BUFF I199 (o_0r1[2:2], joint_0[2:2]);
  BUFF I200 (o_0r1[3:3], joint_0[3:3]);
  BUFF I201 (o_0r1[4:4], joint_0[4:4]);
  BUFF I202 (o_0r1[5:5], joint_0[5:5]);
  BUFF I203 (o_0r1[6:6], joint_0[6:6]);
  BUFF I204 (o_0r1[7:7], joint_0[7:7]);
  BUFF I205 (o_0r1[8:8], joint_0[8:8]);
  BUFF I206 (o_0r1[9:9], joint_0[9:9]);
  BUFF I207 (o_0r1[10:10], joint_0[10:10]);
  BUFF I208 (o_0r1[11:11], joint_0[11:11]);
  BUFF I209 (o_0r1[12:12], joint_0[12:12]);
  BUFF I210 (o_0r1[13:13], joint_0[13:13]);
  BUFF I211 (o_0r1[14:14], joint_0[14:14]);
  BUFF I212 (o_0r1[15:15], joint_0[15:15]);
  BUFF I213 (o_0r1[16:16], joint_0[16:16]);
  BUFF I214 (o_0r1[17:17], joint_0[17:17]);
  BUFF I215 (o_0r1[18:18], joint_0[18:18]);
  BUFF I216 (o_0r1[19:19], joint_0[19:19]);
  BUFF I217 (o_0r1[20:20], joint_0[20:20]);
  BUFF I218 (o_0r1[21:21], joint_0[21:21]);
  BUFF I219 (o_0r1[22:22], joint_0[22:22]);
  BUFF I220 (o_0r1[23:23], joint_0[23:23]);
  BUFF I221 (o_0r1[24:24], joint_0[24:24]);
  BUFF I222 (o_0r1[25:25], joint_0[25:25]);
  BUFF I223 (o_0r1[26:26], joint_0[26:26]);
  BUFF I224 (o_0r1[27:27], joint_0[27:27]);
  BUFF I225 (o_0r1[28:28], joint_0[28:28]);
  BUFF I226 (o_0r1[29:29], joint_0[29:29]);
  BUFF I227 (o_0r1[30:30], joint_0[30:30]);
  BUFF I228 (o_0r1[31:31], joint_0[31:31]);
  BUFF I229 (o_0r1[32:32], joint_0[32:32]);
  BUFF I230 (o_0r1[33:33], joint_0[33:33]);
  BUFF I231 (o_0r1[34:34], joint_0[34:34]);
  BUFF I232 (o_0r1[35:35], joint_0[35:35]);
  BUFF I233 (o_0r1[36:36], joint_0[36:36]);
  BUFF I234 (o_0r1[37:37], joint_0[37:37]);
  BUFF I235 (o_0r1[38:38], joint_0[38:38]);
  BUFF I236 (o_0r1[39:39], joint_0[39:39]);
  BUFF I237 (o_0r1[40:40], joint_0[40:40]);
  BUFF I238 (o_0r1[41:41], joint_0[41:41]);
  BUFF I239 (o_0r1[42:42], joint_0[42:42]);
  BUFF I240 (o_0r1[43:43], joint_0[43:43]);
  BUFF I241 (o_0r1[44:44], joint_0[44:44]);
  BUFF I242 (o_0r1[45:45], joint_0[45:45]);
  BUFF I243 (o_0r1[46:46], joint_0[46:46]);
  BUFF I244 (o_0r1[47:47], joint_0[47:47]);
  BUFF I245 (o_0r1[48:48], joint_0[48:48]);
  BUFF I246 (o_0r1[49:49], joint_0[49:49]);
  BUFF I247 (o_0r1[50:50], joint_0[50:50]);
  BUFF I248 (o_0r1[51:51], joint_0[51:51]);
  BUFF I249 (o_0r1[52:52], joint_0[52:52]);
  BUFF I250 (o_0r1[53:53], joint_0[53:53]);
  BUFF I251 (o_0r1[54:54], joint_0[54:54]);
  BUFF I252 (o_0r1[55:55], joint_0[55:55]);
  BUFF I253 (o_0r1[56:56], joint_0[56:56]);
  BUFF I254 (o_0r1[57:57], joint_0[57:57]);
  BUFF I255 (o_0r1[58:58], joint_0[58:58]);
  BUFF I256 (o_0r1[59:59], joint_0[59:59]);
  BUFF I257 (o_0r1[60:60], joint_0[60:60]);
  BUFF I258 (o_0r1[61:61], joint_0[61:61]);
  BUFF I259 (o_0r1[62:62], joint_0[62:62]);
  BUFF I260 (o_0r1[63:63], joint_0[63:63]);
  BUFF I261 (o_0r1[64:64], joint_0[64:64]);
  BUFF I262 (i_0a, o_0a);
  BUFF I263 (i_1a, o_0a);
endmodule

// tkf0mo0w0_o0w0_o0w0 TeakF [0,0,0] [One 0,Many [0,0,0]]
module tkf0mo0w0_o0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  input reset;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  BUFF I2 (o_2r, i_0r);
  C3 I3 (i_0a, o_0a, o_1a, o_2a);
endmodule

// tkvfinst32_wo0w32_ro0w32 TeakV "finst" 32 [] [0] [0] [Many [32],Many [0],Many [0],Many [32]]
module tkvfinst32_wo0w32_ro0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I457 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I458 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I459 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I460 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I461 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I462 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I463 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I464 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I465 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I466 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I467 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I468 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I469 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I470 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I471 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I472 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I473 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I474 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I475 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I476 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I477 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I478 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I479 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I480 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I481 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I482 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I483 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I484 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I485 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I486 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I487 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  OR2 I488 (anyread_0, rg_0r, rg_0a);
  BUFF I489 (wg_0a, wd_0a);
  BUFF I490 (rg_0a, rd_0a);
endmodule

// tkj35m32_3 TeakJ [Many [32,3],One 35]
module tkj35m32_3 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [2:0] i_1r0;
  input [2:0] i_1r1;
  output i_1a;
  output [34:0] o_0r0;
  output [34:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [34:0] joinf_0;
  wire [34:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joinf_0[32:32], i_1r0[0:0]);
  BUFF I33 (joinf_0[33:33], i_1r0[1:1]);
  BUFF I34 (joinf_0[34:34], i_1r0[2:2]);
  BUFF I35 (joint_0[0:0], i_0r1[0:0]);
  BUFF I36 (joint_0[1:1], i_0r1[1:1]);
  BUFF I37 (joint_0[2:2], i_0r1[2:2]);
  BUFF I38 (joint_0[3:3], i_0r1[3:3]);
  BUFF I39 (joint_0[4:4], i_0r1[4:4]);
  BUFF I40 (joint_0[5:5], i_0r1[5:5]);
  BUFF I41 (joint_0[6:6], i_0r1[6:6]);
  BUFF I42 (joint_0[7:7], i_0r1[7:7]);
  BUFF I43 (joint_0[8:8], i_0r1[8:8]);
  BUFF I44 (joint_0[9:9], i_0r1[9:9]);
  BUFF I45 (joint_0[10:10], i_0r1[10:10]);
  BUFF I46 (joint_0[11:11], i_0r1[11:11]);
  BUFF I47 (joint_0[12:12], i_0r1[12:12]);
  BUFF I48 (joint_0[13:13], i_0r1[13:13]);
  BUFF I49 (joint_0[14:14], i_0r1[14:14]);
  BUFF I50 (joint_0[15:15], i_0r1[15:15]);
  BUFF I51 (joint_0[16:16], i_0r1[16:16]);
  BUFF I52 (joint_0[17:17], i_0r1[17:17]);
  BUFF I53 (joint_0[18:18], i_0r1[18:18]);
  BUFF I54 (joint_0[19:19], i_0r1[19:19]);
  BUFF I55 (joint_0[20:20], i_0r1[20:20]);
  BUFF I56 (joint_0[21:21], i_0r1[21:21]);
  BUFF I57 (joint_0[22:22], i_0r1[22:22]);
  BUFF I58 (joint_0[23:23], i_0r1[23:23]);
  BUFF I59 (joint_0[24:24], i_0r1[24:24]);
  BUFF I60 (joint_0[25:25], i_0r1[25:25]);
  BUFF I61 (joint_0[26:26], i_0r1[26:26]);
  BUFF I62 (joint_0[27:27], i_0r1[27:27]);
  BUFF I63 (joint_0[28:28], i_0r1[28:28]);
  BUFF I64 (joint_0[29:29], i_0r1[29:29]);
  BUFF I65 (joint_0[30:30], i_0r1[30:30]);
  BUFF I66 (joint_0[31:31], i_0r1[31:31]);
  BUFF I67 (joint_0[32:32], i_1r1[0:0]);
  BUFF I68 (joint_0[33:33], i_1r1[1:1]);
  BUFF I69 (joint_0[34:34], i_1r1[2:2]);
  OR2 I70 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I71 (icomplete_0, dcomplete_0);
  C2 I72 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I73 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I74 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I75 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I76 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I77 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I78 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I79 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I80 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I81 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I82 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I83 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I84 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I85 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I86 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I87 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I88 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I89 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I90 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I91 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I92 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I93 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I94 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I95 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I96 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I97 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I98 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I99 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I100 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I101 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I102 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I103 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I104 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I105 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I106 (o_0r0[33:33], joinf_0[33:33]);
  BUFF I107 (o_0r0[34:34], joinf_0[34:34]);
  BUFF I108 (o_0r1[1:1], joint_0[1:1]);
  BUFF I109 (o_0r1[2:2], joint_0[2:2]);
  BUFF I110 (o_0r1[3:3], joint_0[3:3]);
  BUFF I111 (o_0r1[4:4], joint_0[4:4]);
  BUFF I112 (o_0r1[5:5], joint_0[5:5]);
  BUFF I113 (o_0r1[6:6], joint_0[6:6]);
  BUFF I114 (o_0r1[7:7], joint_0[7:7]);
  BUFF I115 (o_0r1[8:8], joint_0[8:8]);
  BUFF I116 (o_0r1[9:9], joint_0[9:9]);
  BUFF I117 (o_0r1[10:10], joint_0[10:10]);
  BUFF I118 (o_0r1[11:11], joint_0[11:11]);
  BUFF I119 (o_0r1[12:12], joint_0[12:12]);
  BUFF I120 (o_0r1[13:13], joint_0[13:13]);
  BUFF I121 (o_0r1[14:14], joint_0[14:14]);
  BUFF I122 (o_0r1[15:15], joint_0[15:15]);
  BUFF I123 (o_0r1[16:16], joint_0[16:16]);
  BUFF I124 (o_0r1[17:17], joint_0[17:17]);
  BUFF I125 (o_0r1[18:18], joint_0[18:18]);
  BUFF I126 (o_0r1[19:19], joint_0[19:19]);
  BUFF I127 (o_0r1[20:20], joint_0[20:20]);
  BUFF I128 (o_0r1[21:21], joint_0[21:21]);
  BUFF I129 (o_0r1[22:22], joint_0[22:22]);
  BUFF I130 (o_0r1[23:23], joint_0[23:23]);
  BUFF I131 (o_0r1[24:24], joint_0[24:24]);
  BUFF I132 (o_0r1[25:25], joint_0[25:25]);
  BUFF I133 (o_0r1[26:26], joint_0[26:26]);
  BUFF I134 (o_0r1[27:27], joint_0[27:27]);
  BUFF I135 (o_0r1[28:28], joint_0[28:28]);
  BUFF I136 (o_0r1[29:29], joint_0[29:29]);
  BUFF I137 (o_0r1[30:30], joint_0[30:30]);
  BUFF I138 (o_0r1[31:31], joint_0[31:31]);
  BUFF I139 (o_0r1[32:32], joint_0[32:32]);
  BUFF I140 (o_0r1[33:33], joint_0[33:33]);
  BUFF I141 (o_0r1[34:34], joint_0[34:34]);
  BUFF I142 (i_0a, o_0a);
  BUFF I143 (i_1a, o_0a);
endmodule

// tko35m33_1api0w32b_2api32w3b_3nm1b0_4apt1o0w32bt3o0w1b_5nm30b0_6apt2o0w3bt5o0w30b_7addt4o0w33bt6o0w3
//   3b TeakO [
//     (1,TeakOAppend 1 [(0,0+:32)]),
//     (2,TeakOAppend 1 [(0,32+:3)]),
//     (3,TeakOConstant 1 0),
//     (4,TeakOAppend 1 [(1,0+:32),(3,0+:1)]),
//     (5,TeakOConstant 30 0),
//     (6,TeakOAppend 1 [(2,0+:3),(5,0+:30)]),
//     (7,TeakOp TeakOpAdd [(4,0+:33),(6,0+:33)])] [One 35,One 33]
module tko35m33_1api0w32b_2api32w3b_3nm1b0_4apt1o0w32bt3o0w1b_5nm30b0_6apt2o0w3bt5o0w30b_7addt4o0w33bt6o0w33b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [34:0] i_0r0;
  input [34:0] i_0r1;
  output i_0a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [34:0] gocomp_0;
  wire [11:0] simp371_0;
  wire [3:0] simp372_0;
  wire [1:0] simp373_0;
  wire [31:0] termf_1;
  wire [2:0] termf_2;
  wire termf_3;
  wire [32:0] termf_4;
  wire [29:0] termf_5;
  wire [32:0] termf_6;
  wire [31:0] termt_1;
  wire [2:0] termt_2;
  wire termt_3;
  wire [32:0] termt_4;
  wire [29:0] termt_5;
  wire [32:0] termt_6;
  wire [32:0] cf7__0;
  wire [32:0] ct7__0;
  wire [3:0] ha7__0;
  wire [7:0] fa7_1min_0;
  wire [1:0] simp2781_0;
  wire [1:0] simp2791_0;
  wire [7:0] fa7_2min_0;
  wire [1:0] simp2911_0;
  wire [1:0] simp2921_0;
  wire [7:0] fa7_3min_0;
  wire [1:0] simp3041_0;
  wire [1:0] simp3051_0;
  wire [7:0] fa7_4min_0;
  wire [1:0] simp3171_0;
  wire [1:0] simp3181_0;
  wire [7:0] fa7_5min_0;
  wire [1:0] simp3301_0;
  wire [1:0] simp3311_0;
  wire [7:0] fa7_6min_0;
  wire [1:0] simp3431_0;
  wire [1:0] simp3441_0;
  wire [7:0] fa7_7min_0;
  wire [1:0] simp3561_0;
  wire [1:0] simp3571_0;
  wire [7:0] fa7_8min_0;
  wire [1:0] simp3691_0;
  wire [1:0] simp3701_0;
  wire [7:0] fa7_9min_0;
  wire [1:0] simp3821_0;
  wire [1:0] simp3831_0;
  wire [7:0] fa7_10min_0;
  wire [1:0] simp3951_0;
  wire [1:0] simp3961_0;
  wire [7:0] fa7_11min_0;
  wire [1:0] simp4081_0;
  wire [1:0] simp4091_0;
  wire [7:0] fa7_12min_0;
  wire [1:0] simp4211_0;
  wire [1:0] simp4221_0;
  wire [7:0] fa7_13min_0;
  wire [1:0] simp4341_0;
  wire [1:0] simp4351_0;
  wire [7:0] fa7_14min_0;
  wire [1:0] simp4471_0;
  wire [1:0] simp4481_0;
  wire [7:0] fa7_15min_0;
  wire [1:0] simp4601_0;
  wire [1:0] simp4611_0;
  wire [7:0] fa7_16min_0;
  wire [1:0] simp4731_0;
  wire [1:0] simp4741_0;
  wire [7:0] fa7_17min_0;
  wire [1:0] simp4861_0;
  wire [1:0] simp4871_0;
  wire [7:0] fa7_18min_0;
  wire [1:0] simp4991_0;
  wire [1:0] simp5001_0;
  wire [7:0] fa7_19min_0;
  wire [1:0] simp5121_0;
  wire [1:0] simp5131_0;
  wire [7:0] fa7_20min_0;
  wire [1:0] simp5251_0;
  wire [1:0] simp5261_0;
  wire [7:0] fa7_21min_0;
  wire [1:0] simp5381_0;
  wire [1:0] simp5391_0;
  wire [7:0] fa7_22min_0;
  wire [1:0] simp5511_0;
  wire [1:0] simp5521_0;
  wire [7:0] fa7_23min_0;
  wire [1:0] simp5641_0;
  wire [1:0] simp5651_0;
  wire [7:0] fa7_24min_0;
  wire [1:0] simp5771_0;
  wire [1:0] simp5781_0;
  wire [7:0] fa7_25min_0;
  wire [1:0] simp5901_0;
  wire [1:0] simp5911_0;
  wire [7:0] fa7_26min_0;
  wire [1:0] simp6031_0;
  wire [1:0] simp6041_0;
  wire [7:0] fa7_27min_0;
  wire [1:0] simp6161_0;
  wire [1:0] simp6171_0;
  wire [7:0] fa7_28min_0;
  wire [1:0] simp6291_0;
  wire [1:0] simp6301_0;
  wire [7:0] fa7_29min_0;
  wire [1:0] simp6421_0;
  wire [1:0] simp6431_0;
  wire [7:0] fa7_30min_0;
  wire [1:0] simp6551_0;
  wire [1:0] simp6561_0;
  wire [7:0] fa7_31min_0;
  wire [1:0] simp6681_0;
  wire [1:0] simp6691_0;
  wire [7:0] fa7_32min_0;
  wire [1:0] simp6811_0;
  wire [1:0] simp6821_0;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I30 (gocomp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I31 (gocomp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I32 (gocomp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  OR2 I33 (gocomp_0[33:33], i_0r0[33:33], i_0r1[33:33]);
  OR2 I34 (gocomp_0[34:34], i_0r0[34:34], i_0r1[34:34]);
  C3 I35 (simp371_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  C3 I36 (simp371_0[1:1], gocomp_0[3:3], gocomp_0[4:4], gocomp_0[5:5]);
  C3 I37 (simp371_0[2:2], gocomp_0[6:6], gocomp_0[7:7], gocomp_0[8:8]);
  C3 I38 (simp371_0[3:3], gocomp_0[9:9], gocomp_0[10:10], gocomp_0[11:11]);
  C3 I39 (simp371_0[4:4], gocomp_0[12:12], gocomp_0[13:13], gocomp_0[14:14]);
  C3 I40 (simp371_0[5:5], gocomp_0[15:15], gocomp_0[16:16], gocomp_0[17:17]);
  C3 I41 (simp371_0[6:6], gocomp_0[18:18], gocomp_0[19:19], gocomp_0[20:20]);
  C3 I42 (simp371_0[7:7], gocomp_0[21:21], gocomp_0[22:22], gocomp_0[23:23]);
  C3 I43 (simp371_0[8:8], gocomp_0[24:24], gocomp_0[25:25], gocomp_0[26:26]);
  C3 I44 (simp371_0[9:9], gocomp_0[27:27], gocomp_0[28:28], gocomp_0[29:29]);
  C3 I45 (simp371_0[10:10], gocomp_0[30:30], gocomp_0[31:31], gocomp_0[32:32]);
  C2 I46 (simp371_0[11:11], gocomp_0[33:33], gocomp_0[34:34]);
  C3 I47 (simp372_0[0:0], simp371_0[0:0], simp371_0[1:1], simp371_0[2:2]);
  C3 I48 (simp372_0[1:1], simp371_0[3:3], simp371_0[4:4], simp371_0[5:5]);
  C3 I49 (simp372_0[2:2], simp371_0[6:6], simp371_0[7:7], simp371_0[8:8]);
  C3 I50 (simp372_0[3:3], simp371_0[9:9], simp371_0[10:10], simp371_0[11:11]);
  C3 I51 (simp373_0[0:0], simp372_0[0:0], simp372_0[1:1], simp372_0[2:2]);
  BUFF I52 (simp373_0[1:1], simp372_0[3:3]);
  C2 I53 (go_0, simp373_0[0:0], simp373_0[1:1]);
  BUFF I54 (termf_1[0:0], i_0r0[0:0]);
  BUFF I55 (termf_1[1:1], i_0r0[1:1]);
  BUFF I56 (termf_1[2:2], i_0r0[2:2]);
  BUFF I57 (termf_1[3:3], i_0r0[3:3]);
  BUFF I58 (termf_1[4:4], i_0r0[4:4]);
  BUFF I59 (termf_1[5:5], i_0r0[5:5]);
  BUFF I60 (termf_1[6:6], i_0r0[6:6]);
  BUFF I61 (termf_1[7:7], i_0r0[7:7]);
  BUFF I62 (termf_1[8:8], i_0r0[8:8]);
  BUFF I63 (termf_1[9:9], i_0r0[9:9]);
  BUFF I64 (termf_1[10:10], i_0r0[10:10]);
  BUFF I65 (termf_1[11:11], i_0r0[11:11]);
  BUFF I66 (termf_1[12:12], i_0r0[12:12]);
  BUFF I67 (termf_1[13:13], i_0r0[13:13]);
  BUFF I68 (termf_1[14:14], i_0r0[14:14]);
  BUFF I69 (termf_1[15:15], i_0r0[15:15]);
  BUFF I70 (termf_1[16:16], i_0r0[16:16]);
  BUFF I71 (termf_1[17:17], i_0r0[17:17]);
  BUFF I72 (termf_1[18:18], i_0r0[18:18]);
  BUFF I73 (termf_1[19:19], i_0r0[19:19]);
  BUFF I74 (termf_1[20:20], i_0r0[20:20]);
  BUFF I75 (termf_1[21:21], i_0r0[21:21]);
  BUFF I76 (termf_1[22:22], i_0r0[22:22]);
  BUFF I77 (termf_1[23:23], i_0r0[23:23]);
  BUFF I78 (termf_1[24:24], i_0r0[24:24]);
  BUFF I79 (termf_1[25:25], i_0r0[25:25]);
  BUFF I80 (termf_1[26:26], i_0r0[26:26]);
  BUFF I81 (termf_1[27:27], i_0r0[27:27]);
  BUFF I82 (termf_1[28:28], i_0r0[28:28]);
  BUFF I83 (termf_1[29:29], i_0r0[29:29]);
  BUFF I84 (termf_1[30:30], i_0r0[30:30]);
  BUFF I85 (termf_1[31:31], i_0r0[31:31]);
  BUFF I86 (termt_1[0:0], i_0r1[0:0]);
  BUFF I87 (termt_1[1:1], i_0r1[1:1]);
  BUFF I88 (termt_1[2:2], i_0r1[2:2]);
  BUFF I89 (termt_1[3:3], i_0r1[3:3]);
  BUFF I90 (termt_1[4:4], i_0r1[4:4]);
  BUFF I91 (termt_1[5:5], i_0r1[5:5]);
  BUFF I92 (termt_1[6:6], i_0r1[6:6]);
  BUFF I93 (termt_1[7:7], i_0r1[7:7]);
  BUFF I94 (termt_1[8:8], i_0r1[8:8]);
  BUFF I95 (termt_1[9:9], i_0r1[9:9]);
  BUFF I96 (termt_1[10:10], i_0r1[10:10]);
  BUFF I97 (termt_1[11:11], i_0r1[11:11]);
  BUFF I98 (termt_1[12:12], i_0r1[12:12]);
  BUFF I99 (termt_1[13:13], i_0r1[13:13]);
  BUFF I100 (termt_1[14:14], i_0r1[14:14]);
  BUFF I101 (termt_1[15:15], i_0r1[15:15]);
  BUFF I102 (termt_1[16:16], i_0r1[16:16]);
  BUFF I103 (termt_1[17:17], i_0r1[17:17]);
  BUFF I104 (termt_1[18:18], i_0r1[18:18]);
  BUFF I105 (termt_1[19:19], i_0r1[19:19]);
  BUFF I106 (termt_1[20:20], i_0r1[20:20]);
  BUFF I107 (termt_1[21:21], i_0r1[21:21]);
  BUFF I108 (termt_1[22:22], i_0r1[22:22]);
  BUFF I109 (termt_1[23:23], i_0r1[23:23]);
  BUFF I110 (termt_1[24:24], i_0r1[24:24]);
  BUFF I111 (termt_1[25:25], i_0r1[25:25]);
  BUFF I112 (termt_1[26:26], i_0r1[26:26]);
  BUFF I113 (termt_1[27:27], i_0r1[27:27]);
  BUFF I114 (termt_1[28:28], i_0r1[28:28]);
  BUFF I115 (termt_1[29:29], i_0r1[29:29]);
  BUFF I116 (termt_1[30:30], i_0r1[30:30]);
  BUFF I117 (termt_1[31:31], i_0r1[31:31]);
  BUFF I118 (termf_2[0:0], i_0r0[32:32]);
  BUFF I119 (termf_2[1:1], i_0r0[33:33]);
  BUFF I120 (termf_2[2:2], i_0r0[34:34]);
  BUFF I121 (termt_2[0:0], i_0r1[32:32]);
  BUFF I122 (termt_2[1:1], i_0r1[33:33]);
  BUFF I123 (termt_2[2:2], i_0r1[34:34]);
  BUFF I124 (termf_3, go_0);
  GND I125 (termt_3);
  BUFF I126 (termf_4[0:0], termf_1[0:0]);
  BUFF I127 (termf_4[1:1], termf_1[1:1]);
  BUFF I128 (termf_4[2:2], termf_1[2:2]);
  BUFF I129 (termf_4[3:3], termf_1[3:3]);
  BUFF I130 (termf_4[4:4], termf_1[4:4]);
  BUFF I131 (termf_4[5:5], termf_1[5:5]);
  BUFF I132 (termf_4[6:6], termf_1[6:6]);
  BUFF I133 (termf_4[7:7], termf_1[7:7]);
  BUFF I134 (termf_4[8:8], termf_1[8:8]);
  BUFF I135 (termf_4[9:9], termf_1[9:9]);
  BUFF I136 (termf_4[10:10], termf_1[10:10]);
  BUFF I137 (termf_4[11:11], termf_1[11:11]);
  BUFF I138 (termf_4[12:12], termf_1[12:12]);
  BUFF I139 (termf_4[13:13], termf_1[13:13]);
  BUFF I140 (termf_4[14:14], termf_1[14:14]);
  BUFF I141 (termf_4[15:15], termf_1[15:15]);
  BUFF I142 (termf_4[16:16], termf_1[16:16]);
  BUFF I143 (termf_4[17:17], termf_1[17:17]);
  BUFF I144 (termf_4[18:18], termf_1[18:18]);
  BUFF I145 (termf_4[19:19], termf_1[19:19]);
  BUFF I146 (termf_4[20:20], termf_1[20:20]);
  BUFF I147 (termf_4[21:21], termf_1[21:21]);
  BUFF I148 (termf_4[22:22], termf_1[22:22]);
  BUFF I149 (termf_4[23:23], termf_1[23:23]);
  BUFF I150 (termf_4[24:24], termf_1[24:24]);
  BUFF I151 (termf_4[25:25], termf_1[25:25]);
  BUFF I152 (termf_4[26:26], termf_1[26:26]);
  BUFF I153 (termf_4[27:27], termf_1[27:27]);
  BUFF I154 (termf_4[28:28], termf_1[28:28]);
  BUFF I155 (termf_4[29:29], termf_1[29:29]);
  BUFF I156 (termf_4[30:30], termf_1[30:30]);
  BUFF I157 (termf_4[31:31], termf_1[31:31]);
  BUFF I158 (termf_4[32:32], termf_3);
  BUFF I159 (termt_4[0:0], termt_1[0:0]);
  BUFF I160 (termt_4[1:1], termt_1[1:1]);
  BUFF I161 (termt_4[2:2], termt_1[2:2]);
  BUFF I162 (termt_4[3:3], termt_1[3:3]);
  BUFF I163 (termt_4[4:4], termt_1[4:4]);
  BUFF I164 (termt_4[5:5], termt_1[5:5]);
  BUFF I165 (termt_4[6:6], termt_1[6:6]);
  BUFF I166 (termt_4[7:7], termt_1[7:7]);
  BUFF I167 (termt_4[8:8], termt_1[8:8]);
  BUFF I168 (termt_4[9:9], termt_1[9:9]);
  BUFF I169 (termt_4[10:10], termt_1[10:10]);
  BUFF I170 (termt_4[11:11], termt_1[11:11]);
  BUFF I171 (termt_4[12:12], termt_1[12:12]);
  BUFF I172 (termt_4[13:13], termt_1[13:13]);
  BUFF I173 (termt_4[14:14], termt_1[14:14]);
  BUFF I174 (termt_4[15:15], termt_1[15:15]);
  BUFF I175 (termt_4[16:16], termt_1[16:16]);
  BUFF I176 (termt_4[17:17], termt_1[17:17]);
  BUFF I177 (termt_4[18:18], termt_1[18:18]);
  BUFF I178 (termt_4[19:19], termt_1[19:19]);
  BUFF I179 (termt_4[20:20], termt_1[20:20]);
  BUFF I180 (termt_4[21:21], termt_1[21:21]);
  BUFF I181 (termt_4[22:22], termt_1[22:22]);
  BUFF I182 (termt_4[23:23], termt_1[23:23]);
  BUFF I183 (termt_4[24:24], termt_1[24:24]);
  BUFF I184 (termt_4[25:25], termt_1[25:25]);
  BUFF I185 (termt_4[26:26], termt_1[26:26]);
  BUFF I186 (termt_4[27:27], termt_1[27:27]);
  BUFF I187 (termt_4[28:28], termt_1[28:28]);
  BUFF I188 (termt_4[29:29], termt_1[29:29]);
  BUFF I189 (termt_4[30:30], termt_1[30:30]);
  BUFF I190 (termt_4[31:31], termt_1[31:31]);
  BUFF I191 (termt_4[32:32], termt_3);
  BUFF I192 (termf_5[0:0], go_0);
  BUFF I193 (termf_5[1:1], go_0);
  BUFF I194 (termf_5[2:2], go_0);
  BUFF I195 (termf_5[3:3], go_0);
  BUFF I196 (termf_5[4:4], go_0);
  BUFF I197 (termf_5[5:5], go_0);
  BUFF I198 (termf_5[6:6], go_0);
  BUFF I199 (termf_5[7:7], go_0);
  BUFF I200 (termf_5[8:8], go_0);
  BUFF I201 (termf_5[9:9], go_0);
  BUFF I202 (termf_5[10:10], go_0);
  BUFF I203 (termf_5[11:11], go_0);
  BUFF I204 (termf_5[12:12], go_0);
  BUFF I205 (termf_5[13:13], go_0);
  BUFF I206 (termf_5[14:14], go_0);
  BUFF I207 (termf_5[15:15], go_0);
  BUFF I208 (termf_5[16:16], go_0);
  BUFF I209 (termf_5[17:17], go_0);
  BUFF I210 (termf_5[18:18], go_0);
  BUFF I211 (termf_5[19:19], go_0);
  BUFF I212 (termf_5[20:20], go_0);
  BUFF I213 (termf_5[21:21], go_0);
  BUFF I214 (termf_5[22:22], go_0);
  BUFF I215 (termf_5[23:23], go_0);
  BUFF I216 (termf_5[24:24], go_0);
  BUFF I217 (termf_5[25:25], go_0);
  BUFF I218 (termf_5[26:26], go_0);
  BUFF I219 (termf_5[27:27], go_0);
  BUFF I220 (termf_5[28:28], go_0);
  BUFF I221 (termf_5[29:29], go_0);
  GND I222 (termt_5[0:0]);
  GND I223 (termt_5[1:1]);
  GND I224 (termt_5[2:2]);
  GND I225 (termt_5[3:3]);
  GND I226 (termt_5[4:4]);
  GND I227 (termt_5[5:5]);
  GND I228 (termt_5[6:6]);
  GND I229 (termt_5[7:7]);
  GND I230 (termt_5[8:8]);
  GND I231 (termt_5[9:9]);
  GND I232 (termt_5[10:10]);
  GND I233 (termt_5[11:11]);
  GND I234 (termt_5[12:12]);
  GND I235 (termt_5[13:13]);
  GND I236 (termt_5[14:14]);
  GND I237 (termt_5[15:15]);
  GND I238 (termt_5[16:16]);
  GND I239 (termt_5[17:17]);
  GND I240 (termt_5[18:18]);
  GND I241 (termt_5[19:19]);
  GND I242 (termt_5[20:20]);
  GND I243 (termt_5[21:21]);
  GND I244 (termt_5[22:22]);
  GND I245 (termt_5[23:23]);
  GND I246 (termt_5[24:24]);
  GND I247 (termt_5[25:25]);
  GND I248 (termt_5[26:26]);
  GND I249 (termt_5[27:27]);
  GND I250 (termt_5[28:28]);
  GND I251 (termt_5[29:29]);
  BUFF I252 (termf_6[0:0], termf_2[0:0]);
  BUFF I253 (termf_6[1:1], termf_2[1:1]);
  BUFF I254 (termf_6[2:2], termf_2[2:2]);
  BUFF I255 (termf_6[3:3], termf_5[0:0]);
  BUFF I256 (termf_6[4:4], termf_5[1:1]);
  BUFF I257 (termf_6[5:5], termf_5[2:2]);
  BUFF I258 (termf_6[6:6], termf_5[3:3]);
  BUFF I259 (termf_6[7:7], termf_5[4:4]);
  BUFF I260 (termf_6[8:8], termf_5[5:5]);
  BUFF I261 (termf_6[9:9], termf_5[6:6]);
  BUFF I262 (termf_6[10:10], termf_5[7:7]);
  BUFF I263 (termf_6[11:11], termf_5[8:8]);
  BUFF I264 (termf_6[12:12], termf_5[9:9]);
  BUFF I265 (termf_6[13:13], termf_5[10:10]);
  BUFF I266 (termf_6[14:14], termf_5[11:11]);
  BUFF I267 (termf_6[15:15], termf_5[12:12]);
  BUFF I268 (termf_6[16:16], termf_5[13:13]);
  BUFF I269 (termf_6[17:17], termf_5[14:14]);
  BUFF I270 (termf_6[18:18], termf_5[15:15]);
  BUFF I271 (termf_6[19:19], termf_5[16:16]);
  BUFF I272 (termf_6[20:20], termf_5[17:17]);
  BUFF I273 (termf_6[21:21], termf_5[18:18]);
  BUFF I274 (termf_6[22:22], termf_5[19:19]);
  BUFF I275 (termf_6[23:23], termf_5[20:20]);
  BUFF I276 (termf_6[24:24], termf_5[21:21]);
  BUFF I277 (termf_6[25:25], termf_5[22:22]);
  BUFF I278 (termf_6[26:26], termf_5[23:23]);
  BUFF I279 (termf_6[27:27], termf_5[24:24]);
  BUFF I280 (termf_6[28:28], termf_5[25:25]);
  BUFF I281 (termf_6[29:29], termf_5[26:26]);
  BUFF I282 (termf_6[30:30], termf_5[27:27]);
  BUFF I283 (termf_6[31:31], termf_5[28:28]);
  BUFF I284 (termf_6[32:32], termf_5[29:29]);
  BUFF I285 (termt_6[0:0], termt_2[0:0]);
  BUFF I286 (termt_6[1:1], termt_2[1:1]);
  BUFF I287 (termt_6[2:2], termt_2[2:2]);
  BUFF I288 (termt_6[3:3], termt_5[0:0]);
  BUFF I289 (termt_6[4:4], termt_5[1:1]);
  BUFF I290 (termt_6[5:5], termt_5[2:2]);
  BUFF I291 (termt_6[6:6], termt_5[3:3]);
  BUFF I292 (termt_6[7:7], termt_5[4:4]);
  BUFF I293 (termt_6[8:8], termt_5[5:5]);
  BUFF I294 (termt_6[9:9], termt_5[6:6]);
  BUFF I295 (termt_6[10:10], termt_5[7:7]);
  BUFF I296 (termt_6[11:11], termt_5[8:8]);
  BUFF I297 (termt_6[12:12], termt_5[9:9]);
  BUFF I298 (termt_6[13:13], termt_5[10:10]);
  BUFF I299 (termt_6[14:14], termt_5[11:11]);
  BUFF I300 (termt_6[15:15], termt_5[12:12]);
  BUFF I301 (termt_6[16:16], termt_5[13:13]);
  BUFF I302 (termt_6[17:17], termt_5[14:14]);
  BUFF I303 (termt_6[18:18], termt_5[15:15]);
  BUFF I304 (termt_6[19:19], termt_5[16:16]);
  BUFF I305 (termt_6[20:20], termt_5[17:17]);
  BUFF I306 (termt_6[21:21], termt_5[18:18]);
  BUFF I307 (termt_6[22:22], termt_5[19:19]);
  BUFF I308 (termt_6[23:23], termt_5[20:20]);
  BUFF I309 (termt_6[24:24], termt_5[21:21]);
  BUFF I310 (termt_6[25:25], termt_5[22:22]);
  BUFF I311 (termt_6[26:26], termt_5[23:23]);
  BUFF I312 (termt_6[27:27], termt_5[24:24]);
  BUFF I313 (termt_6[28:28], termt_5[25:25]);
  BUFF I314 (termt_6[29:29], termt_5[26:26]);
  BUFF I315 (termt_6[30:30], termt_5[27:27]);
  BUFF I316 (termt_6[31:31], termt_5[28:28]);
  BUFF I317 (termt_6[32:32], termt_5[29:29]);
  C2 I318 (ha7__0[0:0], termf_6[0:0], termf_4[0:0]);
  C2 I319 (ha7__0[1:1], termf_6[0:0], termt_4[0:0]);
  C2 I320 (ha7__0[2:2], termt_6[0:0], termf_4[0:0]);
  C2 I321 (ha7__0[3:3], termt_6[0:0], termt_4[0:0]);
  OR3 I322 (cf7__0[0:0], ha7__0[0:0], ha7__0[1:1], ha7__0[2:2]);
  BUFF I323 (ct7__0[0:0], ha7__0[3:3]);
  OR2 I324 (o_0r0[0:0], ha7__0[0:0], ha7__0[3:3]);
  OR2 I325 (o_0r1[0:0], ha7__0[1:1], ha7__0[2:2]);
  C3 I326 (fa7_1min_0[0:0], cf7__0[0:0], termf_6[1:1], termf_4[1:1]);
  C3 I327 (fa7_1min_0[1:1], cf7__0[0:0], termf_6[1:1], termt_4[1:1]);
  C3 I328 (fa7_1min_0[2:2], cf7__0[0:0], termt_6[1:1], termf_4[1:1]);
  C3 I329 (fa7_1min_0[3:3], cf7__0[0:0], termt_6[1:1], termt_4[1:1]);
  C3 I330 (fa7_1min_0[4:4], ct7__0[0:0], termf_6[1:1], termf_4[1:1]);
  C3 I331 (fa7_1min_0[5:5], ct7__0[0:0], termf_6[1:1], termt_4[1:1]);
  C3 I332 (fa7_1min_0[6:6], ct7__0[0:0], termt_6[1:1], termf_4[1:1]);
  C3 I333 (fa7_1min_0[7:7], ct7__0[0:0], termt_6[1:1], termt_4[1:1]);
  NOR3 I334 (simp2781_0[0:0], fa7_1min_0[0:0], fa7_1min_0[3:3], fa7_1min_0[5:5]);
  INV I335 (simp2781_0[1:1], fa7_1min_0[6:6]);
  NAND2 I336 (o_0r0[1:1], simp2781_0[0:0], simp2781_0[1:1]);
  NOR3 I337 (simp2791_0[0:0], fa7_1min_0[1:1], fa7_1min_0[2:2], fa7_1min_0[4:4]);
  INV I338 (simp2791_0[1:1], fa7_1min_0[7:7]);
  NAND2 I339 (o_0r1[1:1], simp2791_0[0:0], simp2791_0[1:1]);
  AO222 I340 (ct7__0[1:1], termt_4[1:1], termt_6[1:1], termt_4[1:1], ct7__0[0:0], termt_6[1:1], ct7__0[0:0]);
  AO222 I341 (cf7__0[1:1], termf_4[1:1], termf_6[1:1], termf_4[1:1], cf7__0[0:0], termf_6[1:1], cf7__0[0:0]);
  C3 I342 (fa7_2min_0[0:0], cf7__0[1:1], termf_6[2:2], termf_4[2:2]);
  C3 I343 (fa7_2min_0[1:1], cf7__0[1:1], termf_6[2:2], termt_4[2:2]);
  C3 I344 (fa7_2min_0[2:2], cf7__0[1:1], termt_6[2:2], termf_4[2:2]);
  C3 I345 (fa7_2min_0[3:3], cf7__0[1:1], termt_6[2:2], termt_4[2:2]);
  C3 I346 (fa7_2min_0[4:4], ct7__0[1:1], termf_6[2:2], termf_4[2:2]);
  C3 I347 (fa7_2min_0[5:5], ct7__0[1:1], termf_6[2:2], termt_4[2:2]);
  C3 I348 (fa7_2min_0[6:6], ct7__0[1:1], termt_6[2:2], termf_4[2:2]);
  C3 I349 (fa7_2min_0[7:7], ct7__0[1:1], termt_6[2:2], termt_4[2:2]);
  NOR3 I350 (simp2911_0[0:0], fa7_2min_0[0:0], fa7_2min_0[3:3], fa7_2min_0[5:5]);
  INV I351 (simp2911_0[1:1], fa7_2min_0[6:6]);
  NAND2 I352 (o_0r0[2:2], simp2911_0[0:0], simp2911_0[1:1]);
  NOR3 I353 (simp2921_0[0:0], fa7_2min_0[1:1], fa7_2min_0[2:2], fa7_2min_0[4:4]);
  INV I354 (simp2921_0[1:1], fa7_2min_0[7:7]);
  NAND2 I355 (o_0r1[2:2], simp2921_0[0:0], simp2921_0[1:1]);
  AO222 I356 (ct7__0[2:2], termt_4[2:2], termt_6[2:2], termt_4[2:2], ct7__0[1:1], termt_6[2:2], ct7__0[1:1]);
  AO222 I357 (cf7__0[2:2], termf_4[2:2], termf_6[2:2], termf_4[2:2], cf7__0[1:1], termf_6[2:2], cf7__0[1:1]);
  C3 I358 (fa7_3min_0[0:0], cf7__0[2:2], termf_6[3:3], termf_4[3:3]);
  C3 I359 (fa7_3min_0[1:1], cf7__0[2:2], termf_6[3:3], termt_4[3:3]);
  C3 I360 (fa7_3min_0[2:2], cf7__0[2:2], termt_6[3:3], termf_4[3:3]);
  C3 I361 (fa7_3min_0[3:3], cf7__0[2:2], termt_6[3:3], termt_4[3:3]);
  C3 I362 (fa7_3min_0[4:4], ct7__0[2:2], termf_6[3:3], termf_4[3:3]);
  C3 I363 (fa7_3min_0[5:5], ct7__0[2:2], termf_6[3:3], termt_4[3:3]);
  C3 I364 (fa7_3min_0[6:6], ct7__0[2:2], termt_6[3:3], termf_4[3:3]);
  C3 I365 (fa7_3min_0[7:7], ct7__0[2:2], termt_6[3:3], termt_4[3:3]);
  NOR3 I366 (simp3041_0[0:0], fa7_3min_0[0:0], fa7_3min_0[3:3], fa7_3min_0[5:5]);
  INV I367 (simp3041_0[1:1], fa7_3min_0[6:6]);
  NAND2 I368 (o_0r0[3:3], simp3041_0[0:0], simp3041_0[1:1]);
  NOR3 I369 (simp3051_0[0:0], fa7_3min_0[1:1], fa7_3min_0[2:2], fa7_3min_0[4:4]);
  INV I370 (simp3051_0[1:1], fa7_3min_0[7:7]);
  NAND2 I371 (o_0r1[3:3], simp3051_0[0:0], simp3051_0[1:1]);
  AO222 I372 (ct7__0[3:3], termt_4[3:3], termt_6[3:3], termt_4[3:3], ct7__0[2:2], termt_6[3:3], ct7__0[2:2]);
  AO222 I373 (cf7__0[3:3], termf_4[3:3], termf_6[3:3], termf_4[3:3], cf7__0[2:2], termf_6[3:3], cf7__0[2:2]);
  C3 I374 (fa7_4min_0[0:0], cf7__0[3:3], termf_6[4:4], termf_4[4:4]);
  C3 I375 (fa7_4min_0[1:1], cf7__0[3:3], termf_6[4:4], termt_4[4:4]);
  C3 I376 (fa7_4min_0[2:2], cf7__0[3:3], termt_6[4:4], termf_4[4:4]);
  C3 I377 (fa7_4min_0[3:3], cf7__0[3:3], termt_6[4:4], termt_4[4:4]);
  C3 I378 (fa7_4min_0[4:4], ct7__0[3:3], termf_6[4:4], termf_4[4:4]);
  C3 I379 (fa7_4min_0[5:5], ct7__0[3:3], termf_6[4:4], termt_4[4:4]);
  C3 I380 (fa7_4min_0[6:6], ct7__0[3:3], termt_6[4:4], termf_4[4:4]);
  C3 I381 (fa7_4min_0[7:7], ct7__0[3:3], termt_6[4:4], termt_4[4:4]);
  NOR3 I382 (simp3171_0[0:0], fa7_4min_0[0:0], fa7_4min_0[3:3], fa7_4min_0[5:5]);
  INV I383 (simp3171_0[1:1], fa7_4min_0[6:6]);
  NAND2 I384 (o_0r0[4:4], simp3171_0[0:0], simp3171_0[1:1]);
  NOR3 I385 (simp3181_0[0:0], fa7_4min_0[1:1], fa7_4min_0[2:2], fa7_4min_0[4:4]);
  INV I386 (simp3181_0[1:1], fa7_4min_0[7:7]);
  NAND2 I387 (o_0r1[4:4], simp3181_0[0:0], simp3181_0[1:1]);
  AO222 I388 (ct7__0[4:4], termt_4[4:4], termt_6[4:4], termt_4[4:4], ct7__0[3:3], termt_6[4:4], ct7__0[3:3]);
  AO222 I389 (cf7__0[4:4], termf_4[4:4], termf_6[4:4], termf_4[4:4], cf7__0[3:3], termf_6[4:4], cf7__0[3:3]);
  C3 I390 (fa7_5min_0[0:0], cf7__0[4:4], termf_6[5:5], termf_4[5:5]);
  C3 I391 (fa7_5min_0[1:1], cf7__0[4:4], termf_6[5:5], termt_4[5:5]);
  C3 I392 (fa7_5min_0[2:2], cf7__0[4:4], termt_6[5:5], termf_4[5:5]);
  C3 I393 (fa7_5min_0[3:3], cf7__0[4:4], termt_6[5:5], termt_4[5:5]);
  C3 I394 (fa7_5min_0[4:4], ct7__0[4:4], termf_6[5:5], termf_4[5:5]);
  C3 I395 (fa7_5min_0[5:5], ct7__0[4:4], termf_6[5:5], termt_4[5:5]);
  C3 I396 (fa7_5min_0[6:6], ct7__0[4:4], termt_6[5:5], termf_4[5:5]);
  C3 I397 (fa7_5min_0[7:7], ct7__0[4:4], termt_6[5:5], termt_4[5:5]);
  NOR3 I398 (simp3301_0[0:0], fa7_5min_0[0:0], fa7_5min_0[3:3], fa7_5min_0[5:5]);
  INV I399 (simp3301_0[1:1], fa7_5min_0[6:6]);
  NAND2 I400 (o_0r0[5:5], simp3301_0[0:0], simp3301_0[1:1]);
  NOR3 I401 (simp3311_0[0:0], fa7_5min_0[1:1], fa7_5min_0[2:2], fa7_5min_0[4:4]);
  INV I402 (simp3311_0[1:1], fa7_5min_0[7:7]);
  NAND2 I403 (o_0r1[5:5], simp3311_0[0:0], simp3311_0[1:1]);
  AO222 I404 (ct7__0[5:5], termt_4[5:5], termt_6[5:5], termt_4[5:5], ct7__0[4:4], termt_6[5:5], ct7__0[4:4]);
  AO222 I405 (cf7__0[5:5], termf_4[5:5], termf_6[5:5], termf_4[5:5], cf7__0[4:4], termf_6[5:5], cf7__0[4:4]);
  C3 I406 (fa7_6min_0[0:0], cf7__0[5:5], termf_6[6:6], termf_4[6:6]);
  C3 I407 (fa7_6min_0[1:1], cf7__0[5:5], termf_6[6:6], termt_4[6:6]);
  C3 I408 (fa7_6min_0[2:2], cf7__0[5:5], termt_6[6:6], termf_4[6:6]);
  C3 I409 (fa7_6min_0[3:3], cf7__0[5:5], termt_6[6:6], termt_4[6:6]);
  C3 I410 (fa7_6min_0[4:4], ct7__0[5:5], termf_6[6:6], termf_4[6:6]);
  C3 I411 (fa7_6min_0[5:5], ct7__0[5:5], termf_6[6:6], termt_4[6:6]);
  C3 I412 (fa7_6min_0[6:6], ct7__0[5:5], termt_6[6:6], termf_4[6:6]);
  C3 I413 (fa7_6min_0[7:7], ct7__0[5:5], termt_6[6:6], termt_4[6:6]);
  NOR3 I414 (simp3431_0[0:0], fa7_6min_0[0:0], fa7_6min_0[3:3], fa7_6min_0[5:5]);
  INV I415 (simp3431_0[1:1], fa7_6min_0[6:6]);
  NAND2 I416 (o_0r0[6:6], simp3431_0[0:0], simp3431_0[1:1]);
  NOR3 I417 (simp3441_0[0:0], fa7_6min_0[1:1], fa7_6min_0[2:2], fa7_6min_0[4:4]);
  INV I418 (simp3441_0[1:1], fa7_6min_0[7:7]);
  NAND2 I419 (o_0r1[6:6], simp3441_0[0:0], simp3441_0[1:1]);
  AO222 I420 (ct7__0[6:6], termt_4[6:6], termt_6[6:6], termt_4[6:6], ct7__0[5:5], termt_6[6:6], ct7__0[5:5]);
  AO222 I421 (cf7__0[6:6], termf_4[6:6], termf_6[6:6], termf_4[6:6], cf7__0[5:5], termf_6[6:6], cf7__0[5:5]);
  C3 I422 (fa7_7min_0[0:0], cf7__0[6:6], termf_6[7:7], termf_4[7:7]);
  C3 I423 (fa7_7min_0[1:1], cf7__0[6:6], termf_6[7:7], termt_4[7:7]);
  C3 I424 (fa7_7min_0[2:2], cf7__0[6:6], termt_6[7:7], termf_4[7:7]);
  C3 I425 (fa7_7min_0[3:3], cf7__0[6:6], termt_6[7:7], termt_4[7:7]);
  C3 I426 (fa7_7min_0[4:4], ct7__0[6:6], termf_6[7:7], termf_4[7:7]);
  C3 I427 (fa7_7min_0[5:5], ct7__0[6:6], termf_6[7:7], termt_4[7:7]);
  C3 I428 (fa7_7min_0[6:6], ct7__0[6:6], termt_6[7:7], termf_4[7:7]);
  C3 I429 (fa7_7min_0[7:7], ct7__0[6:6], termt_6[7:7], termt_4[7:7]);
  NOR3 I430 (simp3561_0[0:0], fa7_7min_0[0:0], fa7_7min_0[3:3], fa7_7min_0[5:5]);
  INV I431 (simp3561_0[1:1], fa7_7min_0[6:6]);
  NAND2 I432 (o_0r0[7:7], simp3561_0[0:0], simp3561_0[1:1]);
  NOR3 I433 (simp3571_0[0:0], fa7_7min_0[1:1], fa7_7min_0[2:2], fa7_7min_0[4:4]);
  INV I434 (simp3571_0[1:1], fa7_7min_0[7:7]);
  NAND2 I435 (o_0r1[7:7], simp3571_0[0:0], simp3571_0[1:1]);
  AO222 I436 (ct7__0[7:7], termt_4[7:7], termt_6[7:7], termt_4[7:7], ct7__0[6:6], termt_6[7:7], ct7__0[6:6]);
  AO222 I437 (cf7__0[7:7], termf_4[7:7], termf_6[7:7], termf_4[7:7], cf7__0[6:6], termf_6[7:7], cf7__0[6:6]);
  C3 I438 (fa7_8min_0[0:0], cf7__0[7:7], termf_6[8:8], termf_4[8:8]);
  C3 I439 (fa7_8min_0[1:1], cf7__0[7:7], termf_6[8:8], termt_4[8:8]);
  C3 I440 (fa7_8min_0[2:2], cf7__0[7:7], termt_6[8:8], termf_4[8:8]);
  C3 I441 (fa7_8min_0[3:3], cf7__0[7:7], termt_6[8:8], termt_4[8:8]);
  C3 I442 (fa7_8min_0[4:4], ct7__0[7:7], termf_6[8:8], termf_4[8:8]);
  C3 I443 (fa7_8min_0[5:5], ct7__0[7:7], termf_6[8:8], termt_4[8:8]);
  C3 I444 (fa7_8min_0[6:6], ct7__0[7:7], termt_6[8:8], termf_4[8:8]);
  C3 I445 (fa7_8min_0[7:7], ct7__0[7:7], termt_6[8:8], termt_4[8:8]);
  NOR3 I446 (simp3691_0[0:0], fa7_8min_0[0:0], fa7_8min_0[3:3], fa7_8min_0[5:5]);
  INV I447 (simp3691_0[1:1], fa7_8min_0[6:6]);
  NAND2 I448 (o_0r0[8:8], simp3691_0[0:0], simp3691_0[1:1]);
  NOR3 I449 (simp3701_0[0:0], fa7_8min_0[1:1], fa7_8min_0[2:2], fa7_8min_0[4:4]);
  INV I450 (simp3701_0[1:1], fa7_8min_0[7:7]);
  NAND2 I451 (o_0r1[8:8], simp3701_0[0:0], simp3701_0[1:1]);
  AO222 I452 (ct7__0[8:8], termt_4[8:8], termt_6[8:8], termt_4[8:8], ct7__0[7:7], termt_6[8:8], ct7__0[7:7]);
  AO222 I453 (cf7__0[8:8], termf_4[8:8], termf_6[8:8], termf_4[8:8], cf7__0[7:7], termf_6[8:8], cf7__0[7:7]);
  C3 I454 (fa7_9min_0[0:0], cf7__0[8:8], termf_6[9:9], termf_4[9:9]);
  C3 I455 (fa7_9min_0[1:1], cf7__0[8:8], termf_6[9:9], termt_4[9:9]);
  C3 I456 (fa7_9min_0[2:2], cf7__0[8:8], termt_6[9:9], termf_4[9:9]);
  C3 I457 (fa7_9min_0[3:3], cf7__0[8:8], termt_6[9:9], termt_4[9:9]);
  C3 I458 (fa7_9min_0[4:4], ct7__0[8:8], termf_6[9:9], termf_4[9:9]);
  C3 I459 (fa7_9min_0[5:5], ct7__0[8:8], termf_6[9:9], termt_4[9:9]);
  C3 I460 (fa7_9min_0[6:6], ct7__0[8:8], termt_6[9:9], termf_4[9:9]);
  C3 I461 (fa7_9min_0[7:7], ct7__0[8:8], termt_6[9:9], termt_4[9:9]);
  NOR3 I462 (simp3821_0[0:0], fa7_9min_0[0:0], fa7_9min_0[3:3], fa7_9min_0[5:5]);
  INV I463 (simp3821_0[1:1], fa7_9min_0[6:6]);
  NAND2 I464 (o_0r0[9:9], simp3821_0[0:0], simp3821_0[1:1]);
  NOR3 I465 (simp3831_0[0:0], fa7_9min_0[1:1], fa7_9min_0[2:2], fa7_9min_0[4:4]);
  INV I466 (simp3831_0[1:1], fa7_9min_0[7:7]);
  NAND2 I467 (o_0r1[9:9], simp3831_0[0:0], simp3831_0[1:1]);
  AO222 I468 (ct7__0[9:9], termt_4[9:9], termt_6[9:9], termt_4[9:9], ct7__0[8:8], termt_6[9:9], ct7__0[8:8]);
  AO222 I469 (cf7__0[9:9], termf_4[9:9], termf_6[9:9], termf_4[9:9], cf7__0[8:8], termf_6[9:9], cf7__0[8:8]);
  C3 I470 (fa7_10min_0[0:0], cf7__0[9:9], termf_6[10:10], termf_4[10:10]);
  C3 I471 (fa7_10min_0[1:1], cf7__0[9:9], termf_6[10:10], termt_4[10:10]);
  C3 I472 (fa7_10min_0[2:2], cf7__0[9:9], termt_6[10:10], termf_4[10:10]);
  C3 I473 (fa7_10min_0[3:3], cf7__0[9:9], termt_6[10:10], termt_4[10:10]);
  C3 I474 (fa7_10min_0[4:4], ct7__0[9:9], termf_6[10:10], termf_4[10:10]);
  C3 I475 (fa7_10min_0[5:5], ct7__0[9:9], termf_6[10:10], termt_4[10:10]);
  C3 I476 (fa7_10min_0[6:6], ct7__0[9:9], termt_6[10:10], termf_4[10:10]);
  C3 I477 (fa7_10min_0[7:7], ct7__0[9:9], termt_6[10:10], termt_4[10:10]);
  NOR3 I478 (simp3951_0[0:0], fa7_10min_0[0:0], fa7_10min_0[3:3], fa7_10min_0[5:5]);
  INV I479 (simp3951_0[1:1], fa7_10min_0[6:6]);
  NAND2 I480 (o_0r0[10:10], simp3951_0[0:0], simp3951_0[1:1]);
  NOR3 I481 (simp3961_0[0:0], fa7_10min_0[1:1], fa7_10min_0[2:2], fa7_10min_0[4:4]);
  INV I482 (simp3961_0[1:1], fa7_10min_0[7:7]);
  NAND2 I483 (o_0r1[10:10], simp3961_0[0:0], simp3961_0[1:1]);
  AO222 I484 (ct7__0[10:10], termt_4[10:10], termt_6[10:10], termt_4[10:10], ct7__0[9:9], termt_6[10:10], ct7__0[9:9]);
  AO222 I485 (cf7__0[10:10], termf_4[10:10], termf_6[10:10], termf_4[10:10], cf7__0[9:9], termf_6[10:10], cf7__0[9:9]);
  C3 I486 (fa7_11min_0[0:0], cf7__0[10:10], termf_6[11:11], termf_4[11:11]);
  C3 I487 (fa7_11min_0[1:1], cf7__0[10:10], termf_6[11:11], termt_4[11:11]);
  C3 I488 (fa7_11min_0[2:2], cf7__0[10:10], termt_6[11:11], termf_4[11:11]);
  C3 I489 (fa7_11min_0[3:3], cf7__0[10:10], termt_6[11:11], termt_4[11:11]);
  C3 I490 (fa7_11min_0[4:4], ct7__0[10:10], termf_6[11:11], termf_4[11:11]);
  C3 I491 (fa7_11min_0[5:5], ct7__0[10:10], termf_6[11:11], termt_4[11:11]);
  C3 I492 (fa7_11min_0[6:6], ct7__0[10:10], termt_6[11:11], termf_4[11:11]);
  C3 I493 (fa7_11min_0[7:7], ct7__0[10:10], termt_6[11:11], termt_4[11:11]);
  NOR3 I494 (simp4081_0[0:0], fa7_11min_0[0:0], fa7_11min_0[3:3], fa7_11min_0[5:5]);
  INV I495 (simp4081_0[1:1], fa7_11min_0[6:6]);
  NAND2 I496 (o_0r0[11:11], simp4081_0[0:0], simp4081_0[1:1]);
  NOR3 I497 (simp4091_0[0:0], fa7_11min_0[1:1], fa7_11min_0[2:2], fa7_11min_0[4:4]);
  INV I498 (simp4091_0[1:1], fa7_11min_0[7:7]);
  NAND2 I499 (o_0r1[11:11], simp4091_0[0:0], simp4091_0[1:1]);
  AO222 I500 (ct7__0[11:11], termt_4[11:11], termt_6[11:11], termt_4[11:11], ct7__0[10:10], termt_6[11:11], ct7__0[10:10]);
  AO222 I501 (cf7__0[11:11], termf_4[11:11], termf_6[11:11], termf_4[11:11], cf7__0[10:10], termf_6[11:11], cf7__0[10:10]);
  C3 I502 (fa7_12min_0[0:0], cf7__0[11:11], termf_6[12:12], termf_4[12:12]);
  C3 I503 (fa7_12min_0[1:1], cf7__0[11:11], termf_6[12:12], termt_4[12:12]);
  C3 I504 (fa7_12min_0[2:2], cf7__0[11:11], termt_6[12:12], termf_4[12:12]);
  C3 I505 (fa7_12min_0[3:3], cf7__0[11:11], termt_6[12:12], termt_4[12:12]);
  C3 I506 (fa7_12min_0[4:4], ct7__0[11:11], termf_6[12:12], termf_4[12:12]);
  C3 I507 (fa7_12min_0[5:5], ct7__0[11:11], termf_6[12:12], termt_4[12:12]);
  C3 I508 (fa7_12min_0[6:6], ct7__0[11:11], termt_6[12:12], termf_4[12:12]);
  C3 I509 (fa7_12min_0[7:7], ct7__0[11:11], termt_6[12:12], termt_4[12:12]);
  NOR3 I510 (simp4211_0[0:0], fa7_12min_0[0:0], fa7_12min_0[3:3], fa7_12min_0[5:5]);
  INV I511 (simp4211_0[1:1], fa7_12min_0[6:6]);
  NAND2 I512 (o_0r0[12:12], simp4211_0[0:0], simp4211_0[1:1]);
  NOR3 I513 (simp4221_0[0:0], fa7_12min_0[1:1], fa7_12min_0[2:2], fa7_12min_0[4:4]);
  INV I514 (simp4221_0[1:1], fa7_12min_0[7:7]);
  NAND2 I515 (o_0r1[12:12], simp4221_0[0:0], simp4221_0[1:1]);
  AO222 I516 (ct7__0[12:12], termt_4[12:12], termt_6[12:12], termt_4[12:12], ct7__0[11:11], termt_6[12:12], ct7__0[11:11]);
  AO222 I517 (cf7__0[12:12], termf_4[12:12], termf_6[12:12], termf_4[12:12], cf7__0[11:11], termf_6[12:12], cf7__0[11:11]);
  C3 I518 (fa7_13min_0[0:0], cf7__0[12:12], termf_6[13:13], termf_4[13:13]);
  C3 I519 (fa7_13min_0[1:1], cf7__0[12:12], termf_6[13:13], termt_4[13:13]);
  C3 I520 (fa7_13min_0[2:2], cf7__0[12:12], termt_6[13:13], termf_4[13:13]);
  C3 I521 (fa7_13min_0[3:3], cf7__0[12:12], termt_6[13:13], termt_4[13:13]);
  C3 I522 (fa7_13min_0[4:4], ct7__0[12:12], termf_6[13:13], termf_4[13:13]);
  C3 I523 (fa7_13min_0[5:5], ct7__0[12:12], termf_6[13:13], termt_4[13:13]);
  C3 I524 (fa7_13min_0[6:6], ct7__0[12:12], termt_6[13:13], termf_4[13:13]);
  C3 I525 (fa7_13min_0[7:7], ct7__0[12:12], termt_6[13:13], termt_4[13:13]);
  NOR3 I526 (simp4341_0[0:0], fa7_13min_0[0:0], fa7_13min_0[3:3], fa7_13min_0[5:5]);
  INV I527 (simp4341_0[1:1], fa7_13min_0[6:6]);
  NAND2 I528 (o_0r0[13:13], simp4341_0[0:0], simp4341_0[1:1]);
  NOR3 I529 (simp4351_0[0:0], fa7_13min_0[1:1], fa7_13min_0[2:2], fa7_13min_0[4:4]);
  INV I530 (simp4351_0[1:1], fa7_13min_0[7:7]);
  NAND2 I531 (o_0r1[13:13], simp4351_0[0:0], simp4351_0[1:1]);
  AO222 I532 (ct7__0[13:13], termt_4[13:13], termt_6[13:13], termt_4[13:13], ct7__0[12:12], termt_6[13:13], ct7__0[12:12]);
  AO222 I533 (cf7__0[13:13], termf_4[13:13], termf_6[13:13], termf_4[13:13], cf7__0[12:12], termf_6[13:13], cf7__0[12:12]);
  C3 I534 (fa7_14min_0[0:0], cf7__0[13:13], termf_6[14:14], termf_4[14:14]);
  C3 I535 (fa7_14min_0[1:1], cf7__0[13:13], termf_6[14:14], termt_4[14:14]);
  C3 I536 (fa7_14min_0[2:2], cf7__0[13:13], termt_6[14:14], termf_4[14:14]);
  C3 I537 (fa7_14min_0[3:3], cf7__0[13:13], termt_6[14:14], termt_4[14:14]);
  C3 I538 (fa7_14min_0[4:4], ct7__0[13:13], termf_6[14:14], termf_4[14:14]);
  C3 I539 (fa7_14min_0[5:5], ct7__0[13:13], termf_6[14:14], termt_4[14:14]);
  C3 I540 (fa7_14min_0[6:6], ct7__0[13:13], termt_6[14:14], termf_4[14:14]);
  C3 I541 (fa7_14min_0[7:7], ct7__0[13:13], termt_6[14:14], termt_4[14:14]);
  NOR3 I542 (simp4471_0[0:0], fa7_14min_0[0:0], fa7_14min_0[3:3], fa7_14min_0[5:5]);
  INV I543 (simp4471_0[1:1], fa7_14min_0[6:6]);
  NAND2 I544 (o_0r0[14:14], simp4471_0[0:0], simp4471_0[1:1]);
  NOR3 I545 (simp4481_0[0:0], fa7_14min_0[1:1], fa7_14min_0[2:2], fa7_14min_0[4:4]);
  INV I546 (simp4481_0[1:1], fa7_14min_0[7:7]);
  NAND2 I547 (o_0r1[14:14], simp4481_0[0:0], simp4481_0[1:1]);
  AO222 I548 (ct7__0[14:14], termt_4[14:14], termt_6[14:14], termt_4[14:14], ct7__0[13:13], termt_6[14:14], ct7__0[13:13]);
  AO222 I549 (cf7__0[14:14], termf_4[14:14], termf_6[14:14], termf_4[14:14], cf7__0[13:13], termf_6[14:14], cf7__0[13:13]);
  C3 I550 (fa7_15min_0[0:0], cf7__0[14:14], termf_6[15:15], termf_4[15:15]);
  C3 I551 (fa7_15min_0[1:1], cf7__0[14:14], termf_6[15:15], termt_4[15:15]);
  C3 I552 (fa7_15min_0[2:2], cf7__0[14:14], termt_6[15:15], termf_4[15:15]);
  C3 I553 (fa7_15min_0[3:3], cf7__0[14:14], termt_6[15:15], termt_4[15:15]);
  C3 I554 (fa7_15min_0[4:4], ct7__0[14:14], termf_6[15:15], termf_4[15:15]);
  C3 I555 (fa7_15min_0[5:5], ct7__0[14:14], termf_6[15:15], termt_4[15:15]);
  C3 I556 (fa7_15min_0[6:6], ct7__0[14:14], termt_6[15:15], termf_4[15:15]);
  C3 I557 (fa7_15min_0[7:7], ct7__0[14:14], termt_6[15:15], termt_4[15:15]);
  NOR3 I558 (simp4601_0[0:0], fa7_15min_0[0:0], fa7_15min_0[3:3], fa7_15min_0[5:5]);
  INV I559 (simp4601_0[1:1], fa7_15min_0[6:6]);
  NAND2 I560 (o_0r0[15:15], simp4601_0[0:0], simp4601_0[1:1]);
  NOR3 I561 (simp4611_0[0:0], fa7_15min_0[1:1], fa7_15min_0[2:2], fa7_15min_0[4:4]);
  INV I562 (simp4611_0[1:1], fa7_15min_0[7:7]);
  NAND2 I563 (o_0r1[15:15], simp4611_0[0:0], simp4611_0[1:1]);
  AO222 I564 (ct7__0[15:15], termt_4[15:15], termt_6[15:15], termt_4[15:15], ct7__0[14:14], termt_6[15:15], ct7__0[14:14]);
  AO222 I565 (cf7__0[15:15], termf_4[15:15], termf_6[15:15], termf_4[15:15], cf7__0[14:14], termf_6[15:15], cf7__0[14:14]);
  C3 I566 (fa7_16min_0[0:0], cf7__0[15:15], termf_6[16:16], termf_4[16:16]);
  C3 I567 (fa7_16min_0[1:1], cf7__0[15:15], termf_6[16:16], termt_4[16:16]);
  C3 I568 (fa7_16min_0[2:2], cf7__0[15:15], termt_6[16:16], termf_4[16:16]);
  C3 I569 (fa7_16min_0[3:3], cf7__0[15:15], termt_6[16:16], termt_4[16:16]);
  C3 I570 (fa7_16min_0[4:4], ct7__0[15:15], termf_6[16:16], termf_4[16:16]);
  C3 I571 (fa7_16min_0[5:5], ct7__0[15:15], termf_6[16:16], termt_4[16:16]);
  C3 I572 (fa7_16min_0[6:6], ct7__0[15:15], termt_6[16:16], termf_4[16:16]);
  C3 I573 (fa7_16min_0[7:7], ct7__0[15:15], termt_6[16:16], termt_4[16:16]);
  NOR3 I574 (simp4731_0[0:0], fa7_16min_0[0:0], fa7_16min_0[3:3], fa7_16min_0[5:5]);
  INV I575 (simp4731_0[1:1], fa7_16min_0[6:6]);
  NAND2 I576 (o_0r0[16:16], simp4731_0[0:0], simp4731_0[1:1]);
  NOR3 I577 (simp4741_0[0:0], fa7_16min_0[1:1], fa7_16min_0[2:2], fa7_16min_0[4:4]);
  INV I578 (simp4741_0[1:1], fa7_16min_0[7:7]);
  NAND2 I579 (o_0r1[16:16], simp4741_0[0:0], simp4741_0[1:1]);
  AO222 I580 (ct7__0[16:16], termt_4[16:16], termt_6[16:16], termt_4[16:16], ct7__0[15:15], termt_6[16:16], ct7__0[15:15]);
  AO222 I581 (cf7__0[16:16], termf_4[16:16], termf_6[16:16], termf_4[16:16], cf7__0[15:15], termf_6[16:16], cf7__0[15:15]);
  C3 I582 (fa7_17min_0[0:0], cf7__0[16:16], termf_6[17:17], termf_4[17:17]);
  C3 I583 (fa7_17min_0[1:1], cf7__0[16:16], termf_6[17:17], termt_4[17:17]);
  C3 I584 (fa7_17min_0[2:2], cf7__0[16:16], termt_6[17:17], termf_4[17:17]);
  C3 I585 (fa7_17min_0[3:3], cf7__0[16:16], termt_6[17:17], termt_4[17:17]);
  C3 I586 (fa7_17min_0[4:4], ct7__0[16:16], termf_6[17:17], termf_4[17:17]);
  C3 I587 (fa7_17min_0[5:5], ct7__0[16:16], termf_6[17:17], termt_4[17:17]);
  C3 I588 (fa7_17min_0[6:6], ct7__0[16:16], termt_6[17:17], termf_4[17:17]);
  C3 I589 (fa7_17min_0[7:7], ct7__0[16:16], termt_6[17:17], termt_4[17:17]);
  NOR3 I590 (simp4861_0[0:0], fa7_17min_0[0:0], fa7_17min_0[3:3], fa7_17min_0[5:5]);
  INV I591 (simp4861_0[1:1], fa7_17min_0[6:6]);
  NAND2 I592 (o_0r0[17:17], simp4861_0[0:0], simp4861_0[1:1]);
  NOR3 I593 (simp4871_0[0:0], fa7_17min_0[1:1], fa7_17min_0[2:2], fa7_17min_0[4:4]);
  INV I594 (simp4871_0[1:1], fa7_17min_0[7:7]);
  NAND2 I595 (o_0r1[17:17], simp4871_0[0:0], simp4871_0[1:1]);
  AO222 I596 (ct7__0[17:17], termt_4[17:17], termt_6[17:17], termt_4[17:17], ct7__0[16:16], termt_6[17:17], ct7__0[16:16]);
  AO222 I597 (cf7__0[17:17], termf_4[17:17], termf_6[17:17], termf_4[17:17], cf7__0[16:16], termf_6[17:17], cf7__0[16:16]);
  C3 I598 (fa7_18min_0[0:0], cf7__0[17:17], termf_6[18:18], termf_4[18:18]);
  C3 I599 (fa7_18min_0[1:1], cf7__0[17:17], termf_6[18:18], termt_4[18:18]);
  C3 I600 (fa7_18min_0[2:2], cf7__0[17:17], termt_6[18:18], termf_4[18:18]);
  C3 I601 (fa7_18min_0[3:3], cf7__0[17:17], termt_6[18:18], termt_4[18:18]);
  C3 I602 (fa7_18min_0[4:4], ct7__0[17:17], termf_6[18:18], termf_4[18:18]);
  C3 I603 (fa7_18min_0[5:5], ct7__0[17:17], termf_6[18:18], termt_4[18:18]);
  C3 I604 (fa7_18min_0[6:6], ct7__0[17:17], termt_6[18:18], termf_4[18:18]);
  C3 I605 (fa7_18min_0[7:7], ct7__0[17:17], termt_6[18:18], termt_4[18:18]);
  NOR3 I606 (simp4991_0[0:0], fa7_18min_0[0:0], fa7_18min_0[3:3], fa7_18min_0[5:5]);
  INV I607 (simp4991_0[1:1], fa7_18min_0[6:6]);
  NAND2 I608 (o_0r0[18:18], simp4991_0[0:0], simp4991_0[1:1]);
  NOR3 I609 (simp5001_0[0:0], fa7_18min_0[1:1], fa7_18min_0[2:2], fa7_18min_0[4:4]);
  INV I610 (simp5001_0[1:1], fa7_18min_0[7:7]);
  NAND2 I611 (o_0r1[18:18], simp5001_0[0:0], simp5001_0[1:1]);
  AO222 I612 (ct7__0[18:18], termt_4[18:18], termt_6[18:18], termt_4[18:18], ct7__0[17:17], termt_6[18:18], ct7__0[17:17]);
  AO222 I613 (cf7__0[18:18], termf_4[18:18], termf_6[18:18], termf_4[18:18], cf7__0[17:17], termf_6[18:18], cf7__0[17:17]);
  C3 I614 (fa7_19min_0[0:0], cf7__0[18:18], termf_6[19:19], termf_4[19:19]);
  C3 I615 (fa7_19min_0[1:1], cf7__0[18:18], termf_6[19:19], termt_4[19:19]);
  C3 I616 (fa7_19min_0[2:2], cf7__0[18:18], termt_6[19:19], termf_4[19:19]);
  C3 I617 (fa7_19min_0[3:3], cf7__0[18:18], termt_6[19:19], termt_4[19:19]);
  C3 I618 (fa7_19min_0[4:4], ct7__0[18:18], termf_6[19:19], termf_4[19:19]);
  C3 I619 (fa7_19min_0[5:5], ct7__0[18:18], termf_6[19:19], termt_4[19:19]);
  C3 I620 (fa7_19min_0[6:6], ct7__0[18:18], termt_6[19:19], termf_4[19:19]);
  C3 I621 (fa7_19min_0[7:7], ct7__0[18:18], termt_6[19:19], termt_4[19:19]);
  NOR3 I622 (simp5121_0[0:0], fa7_19min_0[0:0], fa7_19min_0[3:3], fa7_19min_0[5:5]);
  INV I623 (simp5121_0[1:1], fa7_19min_0[6:6]);
  NAND2 I624 (o_0r0[19:19], simp5121_0[0:0], simp5121_0[1:1]);
  NOR3 I625 (simp5131_0[0:0], fa7_19min_0[1:1], fa7_19min_0[2:2], fa7_19min_0[4:4]);
  INV I626 (simp5131_0[1:1], fa7_19min_0[7:7]);
  NAND2 I627 (o_0r1[19:19], simp5131_0[0:0], simp5131_0[1:1]);
  AO222 I628 (ct7__0[19:19], termt_4[19:19], termt_6[19:19], termt_4[19:19], ct7__0[18:18], termt_6[19:19], ct7__0[18:18]);
  AO222 I629 (cf7__0[19:19], termf_4[19:19], termf_6[19:19], termf_4[19:19], cf7__0[18:18], termf_6[19:19], cf7__0[18:18]);
  C3 I630 (fa7_20min_0[0:0], cf7__0[19:19], termf_6[20:20], termf_4[20:20]);
  C3 I631 (fa7_20min_0[1:1], cf7__0[19:19], termf_6[20:20], termt_4[20:20]);
  C3 I632 (fa7_20min_0[2:2], cf7__0[19:19], termt_6[20:20], termf_4[20:20]);
  C3 I633 (fa7_20min_0[3:3], cf7__0[19:19], termt_6[20:20], termt_4[20:20]);
  C3 I634 (fa7_20min_0[4:4], ct7__0[19:19], termf_6[20:20], termf_4[20:20]);
  C3 I635 (fa7_20min_0[5:5], ct7__0[19:19], termf_6[20:20], termt_4[20:20]);
  C3 I636 (fa7_20min_0[6:6], ct7__0[19:19], termt_6[20:20], termf_4[20:20]);
  C3 I637 (fa7_20min_0[7:7], ct7__0[19:19], termt_6[20:20], termt_4[20:20]);
  NOR3 I638 (simp5251_0[0:0], fa7_20min_0[0:0], fa7_20min_0[3:3], fa7_20min_0[5:5]);
  INV I639 (simp5251_0[1:1], fa7_20min_0[6:6]);
  NAND2 I640 (o_0r0[20:20], simp5251_0[0:0], simp5251_0[1:1]);
  NOR3 I641 (simp5261_0[0:0], fa7_20min_0[1:1], fa7_20min_0[2:2], fa7_20min_0[4:4]);
  INV I642 (simp5261_0[1:1], fa7_20min_0[7:7]);
  NAND2 I643 (o_0r1[20:20], simp5261_0[0:0], simp5261_0[1:1]);
  AO222 I644 (ct7__0[20:20], termt_4[20:20], termt_6[20:20], termt_4[20:20], ct7__0[19:19], termt_6[20:20], ct7__0[19:19]);
  AO222 I645 (cf7__0[20:20], termf_4[20:20], termf_6[20:20], termf_4[20:20], cf7__0[19:19], termf_6[20:20], cf7__0[19:19]);
  C3 I646 (fa7_21min_0[0:0], cf7__0[20:20], termf_6[21:21], termf_4[21:21]);
  C3 I647 (fa7_21min_0[1:1], cf7__0[20:20], termf_6[21:21], termt_4[21:21]);
  C3 I648 (fa7_21min_0[2:2], cf7__0[20:20], termt_6[21:21], termf_4[21:21]);
  C3 I649 (fa7_21min_0[3:3], cf7__0[20:20], termt_6[21:21], termt_4[21:21]);
  C3 I650 (fa7_21min_0[4:4], ct7__0[20:20], termf_6[21:21], termf_4[21:21]);
  C3 I651 (fa7_21min_0[5:5], ct7__0[20:20], termf_6[21:21], termt_4[21:21]);
  C3 I652 (fa7_21min_0[6:6], ct7__0[20:20], termt_6[21:21], termf_4[21:21]);
  C3 I653 (fa7_21min_0[7:7], ct7__0[20:20], termt_6[21:21], termt_4[21:21]);
  NOR3 I654 (simp5381_0[0:0], fa7_21min_0[0:0], fa7_21min_0[3:3], fa7_21min_0[5:5]);
  INV I655 (simp5381_0[1:1], fa7_21min_0[6:6]);
  NAND2 I656 (o_0r0[21:21], simp5381_0[0:0], simp5381_0[1:1]);
  NOR3 I657 (simp5391_0[0:0], fa7_21min_0[1:1], fa7_21min_0[2:2], fa7_21min_0[4:4]);
  INV I658 (simp5391_0[1:1], fa7_21min_0[7:7]);
  NAND2 I659 (o_0r1[21:21], simp5391_0[0:0], simp5391_0[1:1]);
  AO222 I660 (ct7__0[21:21], termt_4[21:21], termt_6[21:21], termt_4[21:21], ct7__0[20:20], termt_6[21:21], ct7__0[20:20]);
  AO222 I661 (cf7__0[21:21], termf_4[21:21], termf_6[21:21], termf_4[21:21], cf7__0[20:20], termf_6[21:21], cf7__0[20:20]);
  C3 I662 (fa7_22min_0[0:0], cf7__0[21:21], termf_6[22:22], termf_4[22:22]);
  C3 I663 (fa7_22min_0[1:1], cf7__0[21:21], termf_6[22:22], termt_4[22:22]);
  C3 I664 (fa7_22min_0[2:2], cf7__0[21:21], termt_6[22:22], termf_4[22:22]);
  C3 I665 (fa7_22min_0[3:3], cf7__0[21:21], termt_6[22:22], termt_4[22:22]);
  C3 I666 (fa7_22min_0[4:4], ct7__0[21:21], termf_6[22:22], termf_4[22:22]);
  C3 I667 (fa7_22min_0[5:5], ct7__0[21:21], termf_6[22:22], termt_4[22:22]);
  C3 I668 (fa7_22min_0[6:6], ct7__0[21:21], termt_6[22:22], termf_4[22:22]);
  C3 I669 (fa7_22min_0[7:7], ct7__0[21:21], termt_6[22:22], termt_4[22:22]);
  NOR3 I670 (simp5511_0[0:0], fa7_22min_0[0:0], fa7_22min_0[3:3], fa7_22min_0[5:5]);
  INV I671 (simp5511_0[1:1], fa7_22min_0[6:6]);
  NAND2 I672 (o_0r0[22:22], simp5511_0[0:0], simp5511_0[1:1]);
  NOR3 I673 (simp5521_0[0:0], fa7_22min_0[1:1], fa7_22min_0[2:2], fa7_22min_0[4:4]);
  INV I674 (simp5521_0[1:1], fa7_22min_0[7:7]);
  NAND2 I675 (o_0r1[22:22], simp5521_0[0:0], simp5521_0[1:1]);
  AO222 I676 (ct7__0[22:22], termt_4[22:22], termt_6[22:22], termt_4[22:22], ct7__0[21:21], termt_6[22:22], ct7__0[21:21]);
  AO222 I677 (cf7__0[22:22], termf_4[22:22], termf_6[22:22], termf_4[22:22], cf7__0[21:21], termf_6[22:22], cf7__0[21:21]);
  C3 I678 (fa7_23min_0[0:0], cf7__0[22:22], termf_6[23:23], termf_4[23:23]);
  C3 I679 (fa7_23min_0[1:1], cf7__0[22:22], termf_6[23:23], termt_4[23:23]);
  C3 I680 (fa7_23min_0[2:2], cf7__0[22:22], termt_6[23:23], termf_4[23:23]);
  C3 I681 (fa7_23min_0[3:3], cf7__0[22:22], termt_6[23:23], termt_4[23:23]);
  C3 I682 (fa7_23min_0[4:4], ct7__0[22:22], termf_6[23:23], termf_4[23:23]);
  C3 I683 (fa7_23min_0[5:5], ct7__0[22:22], termf_6[23:23], termt_4[23:23]);
  C3 I684 (fa7_23min_0[6:6], ct7__0[22:22], termt_6[23:23], termf_4[23:23]);
  C3 I685 (fa7_23min_0[7:7], ct7__0[22:22], termt_6[23:23], termt_4[23:23]);
  NOR3 I686 (simp5641_0[0:0], fa7_23min_0[0:0], fa7_23min_0[3:3], fa7_23min_0[5:5]);
  INV I687 (simp5641_0[1:1], fa7_23min_0[6:6]);
  NAND2 I688 (o_0r0[23:23], simp5641_0[0:0], simp5641_0[1:1]);
  NOR3 I689 (simp5651_0[0:0], fa7_23min_0[1:1], fa7_23min_0[2:2], fa7_23min_0[4:4]);
  INV I690 (simp5651_0[1:1], fa7_23min_0[7:7]);
  NAND2 I691 (o_0r1[23:23], simp5651_0[0:0], simp5651_0[1:1]);
  AO222 I692 (ct7__0[23:23], termt_4[23:23], termt_6[23:23], termt_4[23:23], ct7__0[22:22], termt_6[23:23], ct7__0[22:22]);
  AO222 I693 (cf7__0[23:23], termf_4[23:23], termf_6[23:23], termf_4[23:23], cf7__0[22:22], termf_6[23:23], cf7__0[22:22]);
  C3 I694 (fa7_24min_0[0:0], cf7__0[23:23], termf_6[24:24], termf_4[24:24]);
  C3 I695 (fa7_24min_0[1:1], cf7__0[23:23], termf_6[24:24], termt_4[24:24]);
  C3 I696 (fa7_24min_0[2:2], cf7__0[23:23], termt_6[24:24], termf_4[24:24]);
  C3 I697 (fa7_24min_0[3:3], cf7__0[23:23], termt_6[24:24], termt_4[24:24]);
  C3 I698 (fa7_24min_0[4:4], ct7__0[23:23], termf_6[24:24], termf_4[24:24]);
  C3 I699 (fa7_24min_0[5:5], ct7__0[23:23], termf_6[24:24], termt_4[24:24]);
  C3 I700 (fa7_24min_0[6:6], ct7__0[23:23], termt_6[24:24], termf_4[24:24]);
  C3 I701 (fa7_24min_0[7:7], ct7__0[23:23], termt_6[24:24], termt_4[24:24]);
  NOR3 I702 (simp5771_0[0:0], fa7_24min_0[0:0], fa7_24min_0[3:3], fa7_24min_0[5:5]);
  INV I703 (simp5771_0[1:1], fa7_24min_0[6:6]);
  NAND2 I704 (o_0r0[24:24], simp5771_0[0:0], simp5771_0[1:1]);
  NOR3 I705 (simp5781_0[0:0], fa7_24min_0[1:1], fa7_24min_0[2:2], fa7_24min_0[4:4]);
  INV I706 (simp5781_0[1:1], fa7_24min_0[7:7]);
  NAND2 I707 (o_0r1[24:24], simp5781_0[0:0], simp5781_0[1:1]);
  AO222 I708 (ct7__0[24:24], termt_4[24:24], termt_6[24:24], termt_4[24:24], ct7__0[23:23], termt_6[24:24], ct7__0[23:23]);
  AO222 I709 (cf7__0[24:24], termf_4[24:24], termf_6[24:24], termf_4[24:24], cf7__0[23:23], termf_6[24:24], cf7__0[23:23]);
  C3 I710 (fa7_25min_0[0:0], cf7__0[24:24], termf_6[25:25], termf_4[25:25]);
  C3 I711 (fa7_25min_0[1:1], cf7__0[24:24], termf_6[25:25], termt_4[25:25]);
  C3 I712 (fa7_25min_0[2:2], cf7__0[24:24], termt_6[25:25], termf_4[25:25]);
  C3 I713 (fa7_25min_0[3:3], cf7__0[24:24], termt_6[25:25], termt_4[25:25]);
  C3 I714 (fa7_25min_0[4:4], ct7__0[24:24], termf_6[25:25], termf_4[25:25]);
  C3 I715 (fa7_25min_0[5:5], ct7__0[24:24], termf_6[25:25], termt_4[25:25]);
  C3 I716 (fa7_25min_0[6:6], ct7__0[24:24], termt_6[25:25], termf_4[25:25]);
  C3 I717 (fa7_25min_0[7:7], ct7__0[24:24], termt_6[25:25], termt_4[25:25]);
  NOR3 I718 (simp5901_0[0:0], fa7_25min_0[0:0], fa7_25min_0[3:3], fa7_25min_0[5:5]);
  INV I719 (simp5901_0[1:1], fa7_25min_0[6:6]);
  NAND2 I720 (o_0r0[25:25], simp5901_0[0:0], simp5901_0[1:1]);
  NOR3 I721 (simp5911_0[0:0], fa7_25min_0[1:1], fa7_25min_0[2:2], fa7_25min_0[4:4]);
  INV I722 (simp5911_0[1:1], fa7_25min_0[7:7]);
  NAND2 I723 (o_0r1[25:25], simp5911_0[0:0], simp5911_0[1:1]);
  AO222 I724 (ct7__0[25:25], termt_4[25:25], termt_6[25:25], termt_4[25:25], ct7__0[24:24], termt_6[25:25], ct7__0[24:24]);
  AO222 I725 (cf7__0[25:25], termf_4[25:25], termf_6[25:25], termf_4[25:25], cf7__0[24:24], termf_6[25:25], cf7__0[24:24]);
  C3 I726 (fa7_26min_0[0:0], cf7__0[25:25], termf_6[26:26], termf_4[26:26]);
  C3 I727 (fa7_26min_0[1:1], cf7__0[25:25], termf_6[26:26], termt_4[26:26]);
  C3 I728 (fa7_26min_0[2:2], cf7__0[25:25], termt_6[26:26], termf_4[26:26]);
  C3 I729 (fa7_26min_0[3:3], cf7__0[25:25], termt_6[26:26], termt_4[26:26]);
  C3 I730 (fa7_26min_0[4:4], ct7__0[25:25], termf_6[26:26], termf_4[26:26]);
  C3 I731 (fa7_26min_0[5:5], ct7__0[25:25], termf_6[26:26], termt_4[26:26]);
  C3 I732 (fa7_26min_0[6:6], ct7__0[25:25], termt_6[26:26], termf_4[26:26]);
  C3 I733 (fa7_26min_0[7:7], ct7__0[25:25], termt_6[26:26], termt_4[26:26]);
  NOR3 I734 (simp6031_0[0:0], fa7_26min_0[0:0], fa7_26min_0[3:3], fa7_26min_0[5:5]);
  INV I735 (simp6031_0[1:1], fa7_26min_0[6:6]);
  NAND2 I736 (o_0r0[26:26], simp6031_0[0:0], simp6031_0[1:1]);
  NOR3 I737 (simp6041_0[0:0], fa7_26min_0[1:1], fa7_26min_0[2:2], fa7_26min_0[4:4]);
  INV I738 (simp6041_0[1:1], fa7_26min_0[7:7]);
  NAND2 I739 (o_0r1[26:26], simp6041_0[0:0], simp6041_0[1:1]);
  AO222 I740 (ct7__0[26:26], termt_4[26:26], termt_6[26:26], termt_4[26:26], ct7__0[25:25], termt_6[26:26], ct7__0[25:25]);
  AO222 I741 (cf7__0[26:26], termf_4[26:26], termf_6[26:26], termf_4[26:26], cf7__0[25:25], termf_6[26:26], cf7__0[25:25]);
  C3 I742 (fa7_27min_0[0:0], cf7__0[26:26], termf_6[27:27], termf_4[27:27]);
  C3 I743 (fa7_27min_0[1:1], cf7__0[26:26], termf_6[27:27], termt_4[27:27]);
  C3 I744 (fa7_27min_0[2:2], cf7__0[26:26], termt_6[27:27], termf_4[27:27]);
  C3 I745 (fa7_27min_0[3:3], cf7__0[26:26], termt_6[27:27], termt_4[27:27]);
  C3 I746 (fa7_27min_0[4:4], ct7__0[26:26], termf_6[27:27], termf_4[27:27]);
  C3 I747 (fa7_27min_0[5:5], ct7__0[26:26], termf_6[27:27], termt_4[27:27]);
  C3 I748 (fa7_27min_0[6:6], ct7__0[26:26], termt_6[27:27], termf_4[27:27]);
  C3 I749 (fa7_27min_0[7:7], ct7__0[26:26], termt_6[27:27], termt_4[27:27]);
  NOR3 I750 (simp6161_0[0:0], fa7_27min_0[0:0], fa7_27min_0[3:3], fa7_27min_0[5:5]);
  INV I751 (simp6161_0[1:1], fa7_27min_0[6:6]);
  NAND2 I752 (o_0r0[27:27], simp6161_0[0:0], simp6161_0[1:1]);
  NOR3 I753 (simp6171_0[0:0], fa7_27min_0[1:1], fa7_27min_0[2:2], fa7_27min_0[4:4]);
  INV I754 (simp6171_0[1:1], fa7_27min_0[7:7]);
  NAND2 I755 (o_0r1[27:27], simp6171_0[0:0], simp6171_0[1:1]);
  AO222 I756 (ct7__0[27:27], termt_4[27:27], termt_6[27:27], termt_4[27:27], ct7__0[26:26], termt_6[27:27], ct7__0[26:26]);
  AO222 I757 (cf7__0[27:27], termf_4[27:27], termf_6[27:27], termf_4[27:27], cf7__0[26:26], termf_6[27:27], cf7__0[26:26]);
  C3 I758 (fa7_28min_0[0:0], cf7__0[27:27], termf_6[28:28], termf_4[28:28]);
  C3 I759 (fa7_28min_0[1:1], cf7__0[27:27], termf_6[28:28], termt_4[28:28]);
  C3 I760 (fa7_28min_0[2:2], cf7__0[27:27], termt_6[28:28], termf_4[28:28]);
  C3 I761 (fa7_28min_0[3:3], cf7__0[27:27], termt_6[28:28], termt_4[28:28]);
  C3 I762 (fa7_28min_0[4:4], ct7__0[27:27], termf_6[28:28], termf_4[28:28]);
  C3 I763 (fa7_28min_0[5:5], ct7__0[27:27], termf_6[28:28], termt_4[28:28]);
  C3 I764 (fa7_28min_0[6:6], ct7__0[27:27], termt_6[28:28], termf_4[28:28]);
  C3 I765 (fa7_28min_0[7:7], ct7__0[27:27], termt_6[28:28], termt_4[28:28]);
  NOR3 I766 (simp6291_0[0:0], fa7_28min_0[0:0], fa7_28min_0[3:3], fa7_28min_0[5:5]);
  INV I767 (simp6291_0[1:1], fa7_28min_0[6:6]);
  NAND2 I768 (o_0r0[28:28], simp6291_0[0:0], simp6291_0[1:1]);
  NOR3 I769 (simp6301_0[0:0], fa7_28min_0[1:1], fa7_28min_0[2:2], fa7_28min_0[4:4]);
  INV I770 (simp6301_0[1:1], fa7_28min_0[7:7]);
  NAND2 I771 (o_0r1[28:28], simp6301_0[0:0], simp6301_0[1:1]);
  AO222 I772 (ct7__0[28:28], termt_4[28:28], termt_6[28:28], termt_4[28:28], ct7__0[27:27], termt_6[28:28], ct7__0[27:27]);
  AO222 I773 (cf7__0[28:28], termf_4[28:28], termf_6[28:28], termf_4[28:28], cf7__0[27:27], termf_6[28:28], cf7__0[27:27]);
  C3 I774 (fa7_29min_0[0:0], cf7__0[28:28], termf_6[29:29], termf_4[29:29]);
  C3 I775 (fa7_29min_0[1:1], cf7__0[28:28], termf_6[29:29], termt_4[29:29]);
  C3 I776 (fa7_29min_0[2:2], cf7__0[28:28], termt_6[29:29], termf_4[29:29]);
  C3 I777 (fa7_29min_0[3:3], cf7__0[28:28], termt_6[29:29], termt_4[29:29]);
  C3 I778 (fa7_29min_0[4:4], ct7__0[28:28], termf_6[29:29], termf_4[29:29]);
  C3 I779 (fa7_29min_0[5:5], ct7__0[28:28], termf_6[29:29], termt_4[29:29]);
  C3 I780 (fa7_29min_0[6:6], ct7__0[28:28], termt_6[29:29], termf_4[29:29]);
  C3 I781 (fa7_29min_0[7:7], ct7__0[28:28], termt_6[29:29], termt_4[29:29]);
  NOR3 I782 (simp6421_0[0:0], fa7_29min_0[0:0], fa7_29min_0[3:3], fa7_29min_0[5:5]);
  INV I783 (simp6421_0[1:1], fa7_29min_0[6:6]);
  NAND2 I784 (o_0r0[29:29], simp6421_0[0:0], simp6421_0[1:1]);
  NOR3 I785 (simp6431_0[0:0], fa7_29min_0[1:1], fa7_29min_0[2:2], fa7_29min_0[4:4]);
  INV I786 (simp6431_0[1:1], fa7_29min_0[7:7]);
  NAND2 I787 (o_0r1[29:29], simp6431_0[0:0], simp6431_0[1:1]);
  AO222 I788 (ct7__0[29:29], termt_4[29:29], termt_6[29:29], termt_4[29:29], ct7__0[28:28], termt_6[29:29], ct7__0[28:28]);
  AO222 I789 (cf7__0[29:29], termf_4[29:29], termf_6[29:29], termf_4[29:29], cf7__0[28:28], termf_6[29:29], cf7__0[28:28]);
  C3 I790 (fa7_30min_0[0:0], cf7__0[29:29], termf_6[30:30], termf_4[30:30]);
  C3 I791 (fa7_30min_0[1:1], cf7__0[29:29], termf_6[30:30], termt_4[30:30]);
  C3 I792 (fa7_30min_0[2:2], cf7__0[29:29], termt_6[30:30], termf_4[30:30]);
  C3 I793 (fa7_30min_0[3:3], cf7__0[29:29], termt_6[30:30], termt_4[30:30]);
  C3 I794 (fa7_30min_0[4:4], ct7__0[29:29], termf_6[30:30], termf_4[30:30]);
  C3 I795 (fa7_30min_0[5:5], ct7__0[29:29], termf_6[30:30], termt_4[30:30]);
  C3 I796 (fa7_30min_0[6:6], ct7__0[29:29], termt_6[30:30], termf_4[30:30]);
  C3 I797 (fa7_30min_0[7:7], ct7__0[29:29], termt_6[30:30], termt_4[30:30]);
  NOR3 I798 (simp6551_0[0:0], fa7_30min_0[0:0], fa7_30min_0[3:3], fa7_30min_0[5:5]);
  INV I799 (simp6551_0[1:1], fa7_30min_0[6:6]);
  NAND2 I800 (o_0r0[30:30], simp6551_0[0:0], simp6551_0[1:1]);
  NOR3 I801 (simp6561_0[0:0], fa7_30min_0[1:1], fa7_30min_0[2:2], fa7_30min_0[4:4]);
  INV I802 (simp6561_0[1:1], fa7_30min_0[7:7]);
  NAND2 I803 (o_0r1[30:30], simp6561_0[0:0], simp6561_0[1:1]);
  AO222 I804 (ct7__0[30:30], termt_4[30:30], termt_6[30:30], termt_4[30:30], ct7__0[29:29], termt_6[30:30], ct7__0[29:29]);
  AO222 I805 (cf7__0[30:30], termf_4[30:30], termf_6[30:30], termf_4[30:30], cf7__0[29:29], termf_6[30:30], cf7__0[29:29]);
  C3 I806 (fa7_31min_0[0:0], cf7__0[30:30], termf_6[31:31], termf_4[31:31]);
  C3 I807 (fa7_31min_0[1:1], cf7__0[30:30], termf_6[31:31], termt_4[31:31]);
  C3 I808 (fa7_31min_0[2:2], cf7__0[30:30], termt_6[31:31], termf_4[31:31]);
  C3 I809 (fa7_31min_0[3:3], cf7__0[30:30], termt_6[31:31], termt_4[31:31]);
  C3 I810 (fa7_31min_0[4:4], ct7__0[30:30], termf_6[31:31], termf_4[31:31]);
  C3 I811 (fa7_31min_0[5:5], ct7__0[30:30], termf_6[31:31], termt_4[31:31]);
  C3 I812 (fa7_31min_0[6:6], ct7__0[30:30], termt_6[31:31], termf_4[31:31]);
  C3 I813 (fa7_31min_0[7:7], ct7__0[30:30], termt_6[31:31], termt_4[31:31]);
  NOR3 I814 (simp6681_0[0:0], fa7_31min_0[0:0], fa7_31min_0[3:3], fa7_31min_0[5:5]);
  INV I815 (simp6681_0[1:1], fa7_31min_0[6:6]);
  NAND2 I816 (o_0r0[31:31], simp6681_0[0:0], simp6681_0[1:1]);
  NOR3 I817 (simp6691_0[0:0], fa7_31min_0[1:1], fa7_31min_0[2:2], fa7_31min_0[4:4]);
  INV I818 (simp6691_0[1:1], fa7_31min_0[7:7]);
  NAND2 I819 (o_0r1[31:31], simp6691_0[0:0], simp6691_0[1:1]);
  AO222 I820 (ct7__0[31:31], termt_4[31:31], termt_6[31:31], termt_4[31:31], ct7__0[30:30], termt_6[31:31], ct7__0[30:30]);
  AO222 I821 (cf7__0[31:31], termf_4[31:31], termf_6[31:31], termf_4[31:31], cf7__0[30:30], termf_6[31:31], cf7__0[30:30]);
  C3 I822 (fa7_32min_0[0:0], cf7__0[31:31], termf_6[32:32], termf_4[32:32]);
  C3 I823 (fa7_32min_0[1:1], cf7__0[31:31], termf_6[32:32], termt_4[32:32]);
  C3 I824 (fa7_32min_0[2:2], cf7__0[31:31], termt_6[32:32], termf_4[32:32]);
  C3 I825 (fa7_32min_0[3:3], cf7__0[31:31], termt_6[32:32], termt_4[32:32]);
  C3 I826 (fa7_32min_0[4:4], ct7__0[31:31], termf_6[32:32], termf_4[32:32]);
  C3 I827 (fa7_32min_0[5:5], ct7__0[31:31], termf_6[32:32], termt_4[32:32]);
  C3 I828 (fa7_32min_0[6:6], ct7__0[31:31], termt_6[32:32], termf_4[32:32]);
  C3 I829 (fa7_32min_0[7:7], ct7__0[31:31], termt_6[32:32], termt_4[32:32]);
  NOR3 I830 (simp6811_0[0:0], fa7_32min_0[0:0], fa7_32min_0[3:3], fa7_32min_0[5:5]);
  INV I831 (simp6811_0[1:1], fa7_32min_0[6:6]);
  NAND2 I832 (o_0r0[32:32], simp6811_0[0:0], simp6811_0[1:1]);
  NOR3 I833 (simp6821_0[0:0], fa7_32min_0[1:1], fa7_32min_0[2:2], fa7_32min_0[4:4]);
  INV I834 (simp6821_0[1:1], fa7_32min_0[7:7]);
  NAND2 I835 (o_0r1[32:32], simp6821_0[0:0], simp6821_0[1:1]);
  AO222 I836 (ct7__0[32:32], termt_4[32:32], termt_6[32:32], termt_4[32:32], ct7__0[31:31], termt_6[32:32], ct7__0[31:31]);
  AO222 I837 (cf7__0[32:32], termf_4[32:32], termf_6[32:32], termf_4[32:32], cf7__0[31:31], termf_6[32:32], cf7__0[31:31]);
  BUFF I838 (i_0a, o_0a);
endmodule

// tkf33mo0w32 TeakF [0] [One 33,Many [32]]
module tkf33mo0w32 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [32:0] i_0r0;
  input [32:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  wire ucomplete_0;
  wire comp_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (comp_0, i_0r0[32:32], i_0r1[32:32]);
  BUFF I2 (ucomplete_0, comp_0);
  C2 I3 (acomplete_0, ucomplete_0, icomplete_0);
  C2 I4 (o_0r0[0:0], i_0r0[0:0], icomplete_0);
  BUFF I5 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I6 (o_0r0[2:2], i_0r0[2:2]);
  BUFF I7 (o_0r0[3:3], i_0r0[3:3]);
  BUFF I8 (o_0r0[4:4], i_0r0[4:4]);
  BUFF I9 (o_0r0[5:5], i_0r0[5:5]);
  BUFF I10 (o_0r0[6:6], i_0r0[6:6]);
  BUFF I11 (o_0r0[7:7], i_0r0[7:7]);
  BUFF I12 (o_0r0[8:8], i_0r0[8:8]);
  BUFF I13 (o_0r0[9:9], i_0r0[9:9]);
  BUFF I14 (o_0r0[10:10], i_0r0[10:10]);
  BUFF I15 (o_0r0[11:11], i_0r0[11:11]);
  BUFF I16 (o_0r0[12:12], i_0r0[12:12]);
  BUFF I17 (o_0r0[13:13], i_0r0[13:13]);
  BUFF I18 (o_0r0[14:14], i_0r0[14:14]);
  BUFF I19 (o_0r0[15:15], i_0r0[15:15]);
  BUFF I20 (o_0r0[16:16], i_0r0[16:16]);
  BUFF I21 (o_0r0[17:17], i_0r0[17:17]);
  BUFF I22 (o_0r0[18:18], i_0r0[18:18]);
  BUFF I23 (o_0r0[19:19], i_0r0[19:19]);
  BUFF I24 (o_0r0[20:20], i_0r0[20:20]);
  BUFF I25 (o_0r0[21:21], i_0r0[21:21]);
  BUFF I26 (o_0r0[22:22], i_0r0[22:22]);
  BUFF I27 (o_0r0[23:23], i_0r0[23:23]);
  BUFF I28 (o_0r0[24:24], i_0r0[24:24]);
  BUFF I29 (o_0r0[25:25], i_0r0[25:25]);
  BUFF I30 (o_0r0[26:26], i_0r0[26:26]);
  BUFF I31 (o_0r0[27:27], i_0r0[27:27]);
  BUFF I32 (o_0r0[28:28], i_0r0[28:28]);
  BUFF I33 (o_0r0[29:29], i_0r0[29:29]);
  BUFF I34 (o_0r0[30:30], i_0r0[30:30]);
  BUFF I35 (o_0r0[31:31], i_0r0[31:31]);
  C2 I36 (o_0r1[0:0], i_0r1[0:0], icomplete_0);
  BUFF I37 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I38 (o_0r1[2:2], i_0r1[2:2]);
  BUFF I39 (o_0r1[3:3], i_0r1[3:3]);
  BUFF I40 (o_0r1[4:4], i_0r1[4:4]);
  BUFF I41 (o_0r1[5:5], i_0r1[5:5]);
  BUFF I42 (o_0r1[6:6], i_0r1[6:6]);
  BUFF I43 (o_0r1[7:7], i_0r1[7:7]);
  BUFF I44 (o_0r1[8:8], i_0r1[8:8]);
  BUFF I45 (o_0r1[9:9], i_0r1[9:9]);
  BUFF I46 (o_0r1[10:10], i_0r1[10:10]);
  BUFF I47 (o_0r1[11:11], i_0r1[11:11]);
  BUFF I48 (o_0r1[12:12], i_0r1[12:12]);
  BUFF I49 (o_0r1[13:13], i_0r1[13:13]);
  BUFF I50 (o_0r1[14:14], i_0r1[14:14]);
  BUFF I51 (o_0r1[15:15], i_0r1[15:15]);
  BUFF I52 (o_0r1[16:16], i_0r1[16:16]);
  BUFF I53 (o_0r1[17:17], i_0r1[17:17]);
  BUFF I54 (o_0r1[18:18], i_0r1[18:18]);
  BUFF I55 (o_0r1[19:19], i_0r1[19:19]);
  BUFF I56 (o_0r1[20:20], i_0r1[20:20]);
  BUFF I57 (o_0r1[21:21], i_0r1[21:21]);
  BUFF I58 (o_0r1[22:22], i_0r1[22:22]);
  BUFF I59 (o_0r1[23:23], i_0r1[23:23]);
  BUFF I60 (o_0r1[24:24], i_0r1[24:24]);
  BUFF I61 (o_0r1[25:25], i_0r1[25:25]);
  BUFF I62 (o_0r1[26:26], i_0r1[26:26]);
  BUFF I63 (o_0r1[27:27], i_0r1[27:27]);
  BUFF I64 (o_0r1[28:28], i_0r1[28:28]);
  BUFF I65 (o_0r1[29:29], i_0r1[29:29]);
  BUFF I66 (o_0r1[30:30], i_0r1[30:30]);
  BUFF I67 (o_0r1[31:31], i_0r1[31:31]);
  C2 I68 (i_0a, acomplete_0, o_0a);
endmodule

// tkj0m0_0_0 TeakJ [Many [0,0,0],One 0]
module tkj0m0_0_0 (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  output o_0r;
  input o_0a;
  input reset;
  C3 I0 (o_0r, i_0r, i_1r, i_2r);
  BUFF I1 (i_0a, o_0a);
  BUFF I2 (i_1a, o_0a);
  BUFF I3 (i_2a, o_0a);
endmodule

// tko0m2_1nm2b1 TeakO [
//     (1,TeakOConstant 2 1)] [One 0,One 2]
module tko0m2_1nm2b1 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  GND I1 (o_0r0[0:0]);
  BUFF I2 (o_0r0[1:1], i_0r);
  GND I3 (o_0r1[1:1]);
  BUFF I4 (i_0a, o_0a);
endmodule

// tko0m2_1nm2b2 TeakO [
//     (1,TeakOConstant 2 2)] [One 0,One 2]
module tko0m2_1nm2b2 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[1:1], i_0r);
  GND I1 (o_0r0[1:1]);
  BUFF I2 (o_0r0[0:0], i_0r);
  GND I3 (o_0r1[0:0]);
  BUFF I4 (i_0a, o_0a);
endmodule

// tkm2x2b TeakM [Many [2,2],One 2]
module tkm2x2b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  input [1:0] i_1r0;
  input [1:0] i_1r1;
  output i_1a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  wire [1:0] gfint_0;
  wire [1:0] gfint_1;
  wire [1:0] gtint_0;
  wire [1:0] gtint_1;
  wire choice_0;
  wire choice_1;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire nchosen_0;
  wire [1:0] comp0_0;
  wire [1:0] comp1_0;
  OR2 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0]);
  OR2 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1]);
  OR2 I2 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0]);
  OR2 I3 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1]);
  AND2 I4 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I5 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I6 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I7 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I8 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I9 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I10 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I11 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  OR2 I12 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I13 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  C2 I14 (icomp_0, comp0_0[0:0], comp0_0[1:1]);
  OR2 I15 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I16 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  C2 I17 (icomp_1, comp1_0[0:0], comp1_0[1:1]);
  C2R I18 (choice_0, icomp_0, nchosen_0, reset);
  C2R I19 (choice_1, icomp_1, nchosen_0, reset);
  OR2 I20 (anychoice_0, choice_0, choice_1);
  NOR2 I21 (nchosen_0, anychoice_0, o_0a);
  C2R I22 (i_0a, choice_0, o_0a, reset);
  C2R I23 (i_1a, choice_1, o_0a, reset);
endmodule

// tkj2m0_2 TeakJ [Many [0,2],One 2]
module tkj2m0_2 (i_0r, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  input [1:0] i_1r0;
  input [1:0] i_1r1;
  output i_1a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [1:0] joinf_0;
  wire [1:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_1r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_1r0[1:1]);
  BUFF I2 (joint_0[0:0], i_1r1[0:0]);
  BUFF I3 (joint_0[1:1], i_1r1[1:1]);
  BUFF I4 (icomplete_0, i_0r);
  C2 I5 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I6 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I7 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I8 (o_0r1[1:1], joint_0[1:1]);
  BUFF I9 (i_0a, o_0a);
  BUFF I10 (i_1a, o_0a);
endmodule

// tks2_o0w2_1o0w0_2o0w0 TeakS (0+:2) [([Imp 1 0],0),([Imp 2 0],0)] [One 2,Many [0,0]]
module tks2_o0w2_1o0w0_2o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire [1:0] comp_0;
  BUFF I0 (sel_0, match0_0);
  C2 I1 (match0_0, i_0r1[0:0], i_0r0[1:1]);
  BUFF I2 (sel_1, match1_0);
  C2 I3 (match1_0, i_0r0[0:0], i_0r1[1:1]);
  C2 I4 (gsel_0, sel_0, icomplete_0);
  C2 I5 (gsel_1, sel_1, icomplete_0);
  OR2 I6 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I7 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  C2 I8 (icomplete_0, comp_0[0:0], comp_0[1:1]);
  BUFF I9 (o_0r, gsel_0);
  BUFF I10 (o_1r, gsel_1);
  OR2 I11 (oack_0, o_0a, o_1a);
  C2 I12 (i_0a, oack_0, icomplete_0);
endmodule

// tkvnewStream1_wo0w1_ro0w1 TeakV "newStream" 1 [] [0] [0] [Many [1],Many [0],Many [0],Many [1]]
module tkvnewStream1_wo0w1_ro0w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input wg_0r0;
  input wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  input reset;
  wire wf_0;
  wire wt_0;
  wire df_0;
  wire dt_0;
  wire wc_0;
  wire wacks_0;
  wire wenr_0;
  wire wen_0;
  wire anyread_0;
  wire nreset_0;
  wire drlgf_0;
  wire drlgt_0;
  wire comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire conwgit_0;
  wire conwgif_0;
  wire conwig_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0, wenr_0, nreset_0);
  AND2 I2 (drlgf_0, wf_0, wen_0);
  AND2 I3 (drlgt_0, wt_0, wen_0);
  NOR2 I4 (df_0, dt_0, drlgt_0);
  NOR3 I5 (dt_0, df_0, drlgf_0, reset);
  AO22 I6 (wacks_0, drlgf_0, df_0, drlgt_0, dt_0);
  OR2 I7 (comp0_0, wg_0r0, wg_0r1);
  BUFF I8 (wc_0, comp0_0);
  AND2 I9 (conwgif_0, wg_0r0, conwig_0);
  AND2 I10 (conwgit_0, wg_0r1, conwig_0);
  BUFF I11 (conwigc_0, wc_0);
  AO22 I12 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I13 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I14 (wf_0, conwgif_0);
  BUFF I15 (wt_0, conwgit_0);
  BUFF I16 (wenr_0, wc_0);
  C2 I17 (wd_0r, conwig_0, wacks_0);
  AND2 I18 (rd_0r0, df_0, rg_0r);
  AND2 I19 (rd_0r1, dt_0, rg_0r);
  OR2 I20 (anyread_0, rg_0r, rg_0a);
  BUFF I21 (wg_0a, wd_0a);
  BUFF I22 (rg_0a, rd_0a);
endmodule

// tkvpcTemp32_wo0w32_ro0w32 TeakV "pcTemp" 32 [] [0] [0] [Many [32],Many [0],Many [0],Many [32]]
module tkvpcTemp32_wo0w32_ro0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I457 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I458 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I459 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I460 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I461 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I462 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I463 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I464 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I465 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I466 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I467 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I468 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I469 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I470 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I471 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I472 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I473 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I474 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I475 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I476 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I477 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I478 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I479 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I480 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I481 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I482 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I483 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I484 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I485 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I486 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I487 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  OR2 I488 (anyread_0, rg_0r, rg_0a);
  BUFF I489 (wg_0a, wd_0a);
  BUFF I490 (rg_0a, rd_0a);
endmodule

// tkf32mo0w0_o0w32 TeakF [0,0] [One 32,Many [0,32]]
module tkf32mo0w0_o0w32 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [31:0] o_1r0;
  output [31:0] o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_1r0[0:0], i_0r0[0:0]);
  BUFF I3 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I4 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I5 (o_1r0[3:3], i_0r0[3:3]);
  BUFF I6 (o_1r0[4:4], i_0r0[4:4]);
  BUFF I7 (o_1r0[5:5], i_0r0[5:5]);
  BUFF I8 (o_1r0[6:6], i_0r0[6:6]);
  BUFF I9 (o_1r0[7:7], i_0r0[7:7]);
  BUFF I10 (o_1r0[8:8], i_0r0[8:8]);
  BUFF I11 (o_1r0[9:9], i_0r0[9:9]);
  BUFF I12 (o_1r0[10:10], i_0r0[10:10]);
  BUFF I13 (o_1r0[11:11], i_0r0[11:11]);
  BUFF I14 (o_1r0[12:12], i_0r0[12:12]);
  BUFF I15 (o_1r0[13:13], i_0r0[13:13]);
  BUFF I16 (o_1r0[14:14], i_0r0[14:14]);
  BUFF I17 (o_1r0[15:15], i_0r0[15:15]);
  BUFF I18 (o_1r0[16:16], i_0r0[16:16]);
  BUFF I19 (o_1r0[17:17], i_0r0[17:17]);
  BUFF I20 (o_1r0[18:18], i_0r0[18:18]);
  BUFF I21 (o_1r0[19:19], i_0r0[19:19]);
  BUFF I22 (o_1r0[20:20], i_0r0[20:20]);
  BUFF I23 (o_1r0[21:21], i_0r0[21:21]);
  BUFF I24 (o_1r0[22:22], i_0r0[22:22]);
  BUFF I25 (o_1r0[23:23], i_0r0[23:23]);
  BUFF I26 (o_1r0[24:24], i_0r0[24:24]);
  BUFF I27 (o_1r0[25:25], i_0r0[25:25]);
  BUFF I28 (o_1r0[26:26], i_0r0[26:26]);
  BUFF I29 (o_1r0[27:27], i_0r0[27:27]);
  BUFF I30 (o_1r0[28:28], i_0r0[28:28]);
  BUFF I31 (o_1r0[29:29], i_0r0[29:29]);
  BUFF I32 (o_1r0[30:30], i_0r0[30:30]);
  BUFF I33 (o_1r0[31:31], i_0r0[31:31]);
  BUFF I34 (o_1r1[0:0], i_0r1[0:0]);
  BUFF I35 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I36 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I37 (o_1r1[3:3], i_0r1[3:3]);
  BUFF I38 (o_1r1[4:4], i_0r1[4:4]);
  BUFF I39 (o_1r1[5:5], i_0r1[5:5]);
  BUFF I40 (o_1r1[6:6], i_0r1[6:6]);
  BUFF I41 (o_1r1[7:7], i_0r1[7:7]);
  BUFF I42 (o_1r1[8:8], i_0r1[8:8]);
  BUFF I43 (o_1r1[9:9], i_0r1[9:9]);
  BUFF I44 (o_1r1[10:10], i_0r1[10:10]);
  BUFF I45 (o_1r1[11:11], i_0r1[11:11]);
  BUFF I46 (o_1r1[12:12], i_0r1[12:12]);
  BUFF I47 (o_1r1[13:13], i_0r1[13:13]);
  BUFF I48 (o_1r1[14:14], i_0r1[14:14]);
  BUFF I49 (o_1r1[15:15], i_0r1[15:15]);
  BUFF I50 (o_1r1[16:16], i_0r1[16:16]);
  BUFF I51 (o_1r1[17:17], i_0r1[17:17]);
  BUFF I52 (o_1r1[18:18], i_0r1[18:18]);
  BUFF I53 (o_1r1[19:19], i_0r1[19:19]);
  BUFF I54 (o_1r1[20:20], i_0r1[20:20]);
  BUFF I55 (o_1r1[21:21], i_0r1[21:21]);
  BUFF I56 (o_1r1[22:22], i_0r1[22:22]);
  BUFF I57 (o_1r1[23:23], i_0r1[23:23]);
  BUFF I58 (o_1r1[24:24], i_0r1[24:24]);
  BUFF I59 (o_1r1[25:25], i_0r1[25:25]);
  BUFF I60 (o_1r1[26:26], i_0r1[26:26]);
  BUFF I61 (o_1r1[27:27], i_0r1[27:27]);
  BUFF I62 (o_1r1[28:28], i_0r1[28:28]);
  BUFF I63 (o_1r1[29:29], i_0r1[29:29]);
  BUFF I64 (o_1r1[30:30], i_0r1[30:30]);
  BUFF I65 (o_1r1[31:31], i_0r1[31:31]);
  BUFF I66 (o_0r, icomplete_0);
  C3 I67 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tkm3x32b TeakM [Many [32,32,32],One 32]
module tkm3x32b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  input [31:0] i_2r0;
  input [31:0] i_2r1;
  output i_2a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire [31:0] gfint_0;
  wire [31:0] gfint_1;
  wire [31:0] gfint_2;
  wire [31:0] gtint_0;
  wire [31:0] gtint_1;
  wire [31:0] gtint_2;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire nchosen_0;
  wire [31:0] comp0_0;
  wire [10:0] simp3031_0;
  wire [3:0] simp3032_0;
  wire [1:0] simp3033_0;
  wire [31:0] comp1_0;
  wire [10:0] simp3371_0;
  wire [3:0] simp3372_0;
  wire [1:0] simp3373_0;
  wire [31:0] comp2_0;
  wire [10:0] simp3711_0;
  wire [3:0] simp3712_0;
  wire [1:0] simp3713_0;
  OR3 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  OR3 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  OR3 I2 (o_0r0[2:2], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  OR3 I3 (o_0r0[3:3], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  OR3 I4 (o_0r0[4:4], gfint_0[4:4], gfint_1[4:4], gfint_2[4:4]);
  OR3 I5 (o_0r0[5:5], gfint_0[5:5], gfint_1[5:5], gfint_2[5:5]);
  OR3 I6 (o_0r0[6:6], gfint_0[6:6], gfint_1[6:6], gfint_2[6:6]);
  OR3 I7 (o_0r0[7:7], gfint_0[7:7], gfint_1[7:7], gfint_2[7:7]);
  OR3 I8 (o_0r0[8:8], gfint_0[8:8], gfint_1[8:8], gfint_2[8:8]);
  OR3 I9 (o_0r0[9:9], gfint_0[9:9], gfint_1[9:9], gfint_2[9:9]);
  OR3 I10 (o_0r0[10:10], gfint_0[10:10], gfint_1[10:10], gfint_2[10:10]);
  OR3 I11 (o_0r0[11:11], gfint_0[11:11], gfint_1[11:11], gfint_2[11:11]);
  OR3 I12 (o_0r0[12:12], gfint_0[12:12], gfint_1[12:12], gfint_2[12:12]);
  OR3 I13 (o_0r0[13:13], gfint_0[13:13], gfint_1[13:13], gfint_2[13:13]);
  OR3 I14 (o_0r0[14:14], gfint_0[14:14], gfint_1[14:14], gfint_2[14:14]);
  OR3 I15 (o_0r0[15:15], gfint_0[15:15], gfint_1[15:15], gfint_2[15:15]);
  OR3 I16 (o_0r0[16:16], gfint_0[16:16], gfint_1[16:16], gfint_2[16:16]);
  OR3 I17 (o_0r0[17:17], gfint_0[17:17], gfint_1[17:17], gfint_2[17:17]);
  OR3 I18 (o_0r0[18:18], gfint_0[18:18], gfint_1[18:18], gfint_2[18:18]);
  OR3 I19 (o_0r0[19:19], gfint_0[19:19], gfint_1[19:19], gfint_2[19:19]);
  OR3 I20 (o_0r0[20:20], gfint_0[20:20], gfint_1[20:20], gfint_2[20:20]);
  OR3 I21 (o_0r0[21:21], gfint_0[21:21], gfint_1[21:21], gfint_2[21:21]);
  OR3 I22 (o_0r0[22:22], gfint_0[22:22], gfint_1[22:22], gfint_2[22:22]);
  OR3 I23 (o_0r0[23:23], gfint_0[23:23], gfint_1[23:23], gfint_2[23:23]);
  OR3 I24 (o_0r0[24:24], gfint_0[24:24], gfint_1[24:24], gfint_2[24:24]);
  OR3 I25 (o_0r0[25:25], gfint_0[25:25], gfint_1[25:25], gfint_2[25:25]);
  OR3 I26 (o_0r0[26:26], gfint_0[26:26], gfint_1[26:26], gfint_2[26:26]);
  OR3 I27 (o_0r0[27:27], gfint_0[27:27], gfint_1[27:27], gfint_2[27:27]);
  OR3 I28 (o_0r0[28:28], gfint_0[28:28], gfint_1[28:28], gfint_2[28:28]);
  OR3 I29 (o_0r0[29:29], gfint_0[29:29], gfint_1[29:29], gfint_2[29:29]);
  OR3 I30 (o_0r0[30:30], gfint_0[30:30], gfint_1[30:30], gfint_2[30:30]);
  OR3 I31 (o_0r0[31:31], gfint_0[31:31], gfint_1[31:31], gfint_2[31:31]);
  OR3 I32 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  OR3 I33 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  OR3 I34 (o_0r1[2:2], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  OR3 I35 (o_0r1[3:3], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  OR3 I36 (o_0r1[4:4], gtint_0[4:4], gtint_1[4:4], gtint_2[4:4]);
  OR3 I37 (o_0r1[5:5], gtint_0[5:5], gtint_1[5:5], gtint_2[5:5]);
  OR3 I38 (o_0r1[6:6], gtint_0[6:6], gtint_1[6:6], gtint_2[6:6]);
  OR3 I39 (o_0r1[7:7], gtint_0[7:7], gtint_1[7:7], gtint_2[7:7]);
  OR3 I40 (o_0r1[8:8], gtint_0[8:8], gtint_1[8:8], gtint_2[8:8]);
  OR3 I41 (o_0r1[9:9], gtint_0[9:9], gtint_1[9:9], gtint_2[9:9]);
  OR3 I42 (o_0r1[10:10], gtint_0[10:10], gtint_1[10:10], gtint_2[10:10]);
  OR3 I43 (o_0r1[11:11], gtint_0[11:11], gtint_1[11:11], gtint_2[11:11]);
  OR3 I44 (o_0r1[12:12], gtint_0[12:12], gtint_1[12:12], gtint_2[12:12]);
  OR3 I45 (o_0r1[13:13], gtint_0[13:13], gtint_1[13:13], gtint_2[13:13]);
  OR3 I46 (o_0r1[14:14], gtint_0[14:14], gtint_1[14:14], gtint_2[14:14]);
  OR3 I47 (o_0r1[15:15], gtint_0[15:15], gtint_1[15:15], gtint_2[15:15]);
  OR3 I48 (o_0r1[16:16], gtint_0[16:16], gtint_1[16:16], gtint_2[16:16]);
  OR3 I49 (o_0r1[17:17], gtint_0[17:17], gtint_1[17:17], gtint_2[17:17]);
  OR3 I50 (o_0r1[18:18], gtint_0[18:18], gtint_1[18:18], gtint_2[18:18]);
  OR3 I51 (o_0r1[19:19], gtint_0[19:19], gtint_1[19:19], gtint_2[19:19]);
  OR3 I52 (o_0r1[20:20], gtint_0[20:20], gtint_1[20:20], gtint_2[20:20]);
  OR3 I53 (o_0r1[21:21], gtint_0[21:21], gtint_1[21:21], gtint_2[21:21]);
  OR3 I54 (o_0r1[22:22], gtint_0[22:22], gtint_1[22:22], gtint_2[22:22]);
  OR3 I55 (o_0r1[23:23], gtint_0[23:23], gtint_1[23:23], gtint_2[23:23]);
  OR3 I56 (o_0r1[24:24], gtint_0[24:24], gtint_1[24:24], gtint_2[24:24]);
  OR3 I57 (o_0r1[25:25], gtint_0[25:25], gtint_1[25:25], gtint_2[25:25]);
  OR3 I58 (o_0r1[26:26], gtint_0[26:26], gtint_1[26:26], gtint_2[26:26]);
  OR3 I59 (o_0r1[27:27], gtint_0[27:27], gtint_1[27:27], gtint_2[27:27]);
  OR3 I60 (o_0r1[28:28], gtint_0[28:28], gtint_1[28:28], gtint_2[28:28]);
  OR3 I61 (o_0r1[29:29], gtint_0[29:29], gtint_1[29:29], gtint_2[29:29]);
  OR3 I62 (o_0r1[30:30], gtint_0[30:30], gtint_1[30:30], gtint_2[30:30]);
  OR3 I63 (o_0r1[31:31], gtint_0[31:31], gtint_1[31:31], gtint_2[31:31]);
  AND2 I64 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I65 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I66 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I67 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I68 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I69 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I70 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I71 (gtint_0[7:7], choice_0, i_0r1[7:7]);
  AND2 I72 (gtint_0[8:8], choice_0, i_0r1[8:8]);
  AND2 I73 (gtint_0[9:9], choice_0, i_0r1[9:9]);
  AND2 I74 (gtint_0[10:10], choice_0, i_0r1[10:10]);
  AND2 I75 (gtint_0[11:11], choice_0, i_0r1[11:11]);
  AND2 I76 (gtint_0[12:12], choice_0, i_0r1[12:12]);
  AND2 I77 (gtint_0[13:13], choice_0, i_0r1[13:13]);
  AND2 I78 (gtint_0[14:14], choice_0, i_0r1[14:14]);
  AND2 I79 (gtint_0[15:15], choice_0, i_0r1[15:15]);
  AND2 I80 (gtint_0[16:16], choice_0, i_0r1[16:16]);
  AND2 I81 (gtint_0[17:17], choice_0, i_0r1[17:17]);
  AND2 I82 (gtint_0[18:18], choice_0, i_0r1[18:18]);
  AND2 I83 (gtint_0[19:19], choice_0, i_0r1[19:19]);
  AND2 I84 (gtint_0[20:20], choice_0, i_0r1[20:20]);
  AND2 I85 (gtint_0[21:21], choice_0, i_0r1[21:21]);
  AND2 I86 (gtint_0[22:22], choice_0, i_0r1[22:22]);
  AND2 I87 (gtint_0[23:23], choice_0, i_0r1[23:23]);
  AND2 I88 (gtint_0[24:24], choice_0, i_0r1[24:24]);
  AND2 I89 (gtint_0[25:25], choice_0, i_0r1[25:25]);
  AND2 I90 (gtint_0[26:26], choice_0, i_0r1[26:26]);
  AND2 I91 (gtint_0[27:27], choice_0, i_0r1[27:27]);
  AND2 I92 (gtint_0[28:28], choice_0, i_0r1[28:28]);
  AND2 I93 (gtint_0[29:29], choice_0, i_0r1[29:29]);
  AND2 I94 (gtint_0[30:30], choice_0, i_0r1[30:30]);
  AND2 I95 (gtint_0[31:31], choice_0, i_0r1[31:31]);
  AND2 I96 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I97 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I98 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I99 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I100 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I101 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I102 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I103 (gtint_1[7:7], choice_1, i_1r1[7:7]);
  AND2 I104 (gtint_1[8:8], choice_1, i_1r1[8:8]);
  AND2 I105 (gtint_1[9:9], choice_1, i_1r1[9:9]);
  AND2 I106 (gtint_1[10:10], choice_1, i_1r1[10:10]);
  AND2 I107 (gtint_1[11:11], choice_1, i_1r1[11:11]);
  AND2 I108 (gtint_1[12:12], choice_1, i_1r1[12:12]);
  AND2 I109 (gtint_1[13:13], choice_1, i_1r1[13:13]);
  AND2 I110 (gtint_1[14:14], choice_1, i_1r1[14:14]);
  AND2 I111 (gtint_1[15:15], choice_1, i_1r1[15:15]);
  AND2 I112 (gtint_1[16:16], choice_1, i_1r1[16:16]);
  AND2 I113 (gtint_1[17:17], choice_1, i_1r1[17:17]);
  AND2 I114 (gtint_1[18:18], choice_1, i_1r1[18:18]);
  AND2 I115 (gtint_1[19:19], choice_1, i_1r1[19:19]);
  AND2 I116 (gtint_1[20:20], choice_1, i_1r1[20:20]);
  AND2 I117 (gtint_1[21:21], choice_1, i_1r1[21:21]);
  AND2 I118 (gtint_1[22:22], choice_1, i_1r1[22:22]);
  AND2 I119 (gtint_1[23:23], choice_1, i_1r1[23:23]);
  AND2 I120 (gtint_1[24:24], choice_1, i_1r1[24:24]);
  AND2 I121 (gtint_1[25:25], choice_1, i_1r1[25:25]);
  AND2 I122 (gtint_1[26:26], choice_1, i_1r1[26:26]);
  AND2 I123 (gtint_1[27:27], choice_1, i_1r1[27:27]);
  AND2 I124 (gtint_1[28:28], choice_1, i_1r1[28:28]);
  AND2 I125 (gtint_1[29:29], choice_1, i_1r1[29:29]);
  AND2 I126 (gtint_1[30:30], choice_1, i_1r1[30:30]);
  AND2 I127 (gtint_1[31:31], choice_1, i_1r1[31:31]);
  AND2 I128 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I129 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I130 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I131 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AND2 I132 (gtint_2[4:4], choice_2, i_2r1[4:4]);
  AND2 I133 (gtint_2[5:5], choice_2, i_2r1[5:5]);
  AND2 I134 (gtint_2[6:6], choice_2, i_2r1[6:6]);
  AND2 I135 (gtint_2[7:7], choice_2, i_2r1[7:7]);
  AND2 I136 (gtint_2[8:8], choice_2, i_2r1[8:8]);
  AND2 I137 (gtint_2[9:9], choice_2, i_2r1[9:9]);
  AND2 I138 (gtint_2[10:10], choice_2, i_2r1[10:10]);
  AND2 I139 (gtint_2[11:11], choice_2, i_2r1[11:11]);
  AND2 I140 (gtint_2[12:12], choice_2, i_2r1[12:12]);
  AND2 I141 (gtint_2[13:13], choice_2, i_2r1[13:13]);
  AND2 I142 (gtint_2[14:14], choice_2, i_2r1[14:14]);
  AND2 I143 (gtint_2[15:15], choice_2, i_2r1[15:15]);
  AND2 I144 (gtint_2[16:16], choice_2, i_2r1[16:16]);
  AND2 I145 (gtint_2[17:17], choice_2, i_2r1[17:17]);
  AND2 I146 (gtint_2[18:18], choice_2, i_2r1[18:18]);
  AND2 I147 (gtint_2[19:19], choice_2, i_2r1[19:19]);
  AND2 I148 (gtint_2[20:20], choice_2, i_2r1[20:20]);
  AND2 I149 (gtint_2[21:21], choice_2, i_2r1[21:21]);
  AND2 I150 (gtint_2[22:22], choice_2, i_2r1[22:22]);
  AND2 I151 (gtint_2[23:23], choice_2, i_2r1[23:23]);
  AND2 I152 (gtint_2[24:24], choice_2, i_2r1[24:24]);
  AND2 I153 (gtint_2[25:25], choice_2, i_2r1[25:25]);
  AND2 I154 (gtint_2[26:26], choice_2, i_2r1[26:26]);
  AND2 I155 (gtint_2[27:27], choice_2, i_2r1[27:27]);
  AND2 I156 (gtint_2[28:28], choice_2, i_2r1[28:28]);
  AND2 I157 (gtint_2[29:29], choice_2, i_2r1[29:29]);
  AND2 I158 (gtint_2[30:30], choice_2, i_2r1[30:30]);
  AND2 I159 (gtint_2[31:31], choice_2, i_2r1[31:31]);
  AND2 I160 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I161 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I162 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I163 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I164 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I165 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I166 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I167 (gfint_0[7:7], choice_0, i_0r0[7:7]);
  AND2 I168 (gfint_0[8:8], choice_0, i_0r0[8:8]);
  AND2 I169 (gfint_0[9:9], choice_0, i_0r0[9:9]);
  AND2 I170 (gfint_0[10:10], choice_0, i_0r0[10:10]);
  AND2 I171 (gfint_0[11:11], choice_0, i_0r0[11:11]);
  AND2 I172 (gfint_0[12:12], choice_0, i_0r0[12:12]);
  AND2 I173 (gfint_0[13:13], choice_0, i_0r0[13:13]);
  AND2 I174 (gfint_0[14:14], choice_0, i_0r0[14:14]);
  AND2 I175 (gfint_0[15:15], choice_0, i_0r0[15:15]);
  AND2 I176 (gfint_0[16:16], choice_0, i_0r0[16:16]);
  AND2 I177 (gfint_0[17:17], choice_0, i_0r0[17:17]);
  AND2 I178 (gfint_0[18:18], choice_0, i_0r0[18:18]);
  AND2 I179 (gfint_0[19:19], choice_0, i_0r0[19:19]);
  AND2 I180 (gfint_0[20:20], choice_0, i_0r0[20:20]);
  AND2 I181 (gfint_0[21:21], choice_0, i_0r0[21:21]);
  AND2 I182 (gfint_0[22:22], choice_0, i_0r0[22:22]);
  AND2 I183 (gfint_0[23:23], choice_0, i_0r0[23:23]);
  AND2 I184 (gfint_0[24:24], choice_0, i_0r0[24:24]);
  AND2 I185 (gfint_0[25:25], choice_0, i_0r0[25:25]);
  AND2 I186 (gfint_0[26:26], choice_0, i_0r0[26:26]);
  AND2 I187 (gfint_0[27:27], choice_0, i_0r0[27:27]);
  AND2 I188 (gfint_0[28:28], choice_0, i_0r0[28:28]);
  AND2 I189 (gfint_0[29:29], choice_0, i_0r0[29:29]);
  AND2 I190 (gfint_0[30:30], choice_0, i_0r0[30:30]);
  AND2 I191 (gfint_0[31:31], choice_0, i_0r0[31:31]);
  AND2 I192 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I193 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I194 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I195 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I196 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I197 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I198 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I199 (gfint_1[7:7], choice_1, i_1r0[7:7]);
  AND2 I200 (gfint_1[8:8], choice_1, i_1r0[8:8]);
  AND2 I201 (gfint_1[9:9], choice_1, i_1r0[9:9]);
  AND2 I202 (gfint_1[10:10], choice_1, i_1r0[10:10]);
  AND2 I203 (gfint_1[11:11], choice_1, i_1r0[11:11]);
  AND2 I204 (gfint_1[12:12], choice_1, i_1r0[12:12]);
  AND2 I205 (gfint_1[13:13], choice_1, i_1r0[13:13]);
  AND2 I206 (gfint_1[14:14], choice_1, i_1r0[14:14]);
  AND2 I207 (gfint_1[15:15], choice_1, i_1r0[15:15]);
  AND2 I208 (gfint_1[16:16], choice_1, i_1r0[16:16]);
  AND2 I209 (gfint_1[17:17], choice_1, i_1r0[17:17]);
  AND2 I210 (gfint_1[18:18], choice_1, i_1r0[18:18]);
  AND2 I211 (gfint_1[19:19], choice_1, i_1r0[19:19]);
  AND2 I212 (gfint_1[20:20], choice_1, i_1r0[20:20]);
  AND2 I213 (gfint_1[21:21], choice_1, i_1r0[21:21]);
  AND2 I214 (gfint_1[22:22], choice_1, i_1r0[22:22]);
  AND2 I215 (gfint_1[23:23], choice_1, i_1r0[23:23]);
  AND2 I216 (gfint_1[24:24], choice_1, i_1r0[24:24]);
  AND2 I217 (gfint_1[25:25], choice_1, i_1r0[25:25]);
  AND2 I218 (gfint_1[26:26], choice_1, i_1r0[26:26]);
  AND2 I219 (gfint_1[27:27], choice_1, i_1r0[27:27]);
  AND2 I220 (gfint_1[28:28], choice_1, i_1r0[28:28]);
  AND2 I221 (gfint_1[29:29], choice_1, i_1r0[29:29]);
  AND2 I222 (gfint_1[30:30], choice_1, i_1r0[30:30]);
  AND2 I223 (gfint_1[31:31], choice_1, i_1r0[31:31]);
  AND2 I224 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I225 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I226 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I227 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AND2 I228 (gfint_2[4:4], choice_2, i_2r0[4:4]);
  AND2 I229 (gfint_2[5:5], choice_2, i_2r0[5:5]);
  AND2 I230 (gfint_2[6:6], choice_2, i_2r0[6:6]);
  AND2 I231 (gfint_2[7:7], choice_2, i_2r0[7:7]);
  AND2 I232 (gfint_2[8:8], choice_2, i_2r0[8:8]);
  AND2 I233 (gfint_2[9:9], choice_2, i_2r0[9:9]);
  AND2 I234 (gfint_2[10:10], choice_2, i_2r0[10:10]);
  AND2 I235 (gfint_2[11:11], choice_2, i_2r0[11:11]);
  AND2 I236 (gfint_2[12:12], choice_2, i_2r0[12:12]);
  AND2 I237 (gfint_2[13:13], choice_2, i_2r0[13:13]);
  AND2 I238 (gfint_2[14:14], choice_2, i_2r0[14:14]);
  AND2 I239 (gfint_2[15:15], choice_2, i_2r0[15:15]);
  AND2 I240 (gfint_2[16:16], choice_2, i_2r0[16:16]);
  AND2 I241 (gfint_2[17:17], choice_2, i_2r0[17:17]);
  AND2 I242 (gfint_2[18:18], choice_2, i_2r0[18:18]);
  AND2 I243 (gfint_2[19:19], choice_2, i_2r0[19:19]);
  AND2 I244 (gfint_2[20:20], choice_2, i_2r0[20:20]);
  AND2 I245 (gfint_2[21:21], choice_2, i_2r0[21:21]);
  AND2 I246 (gfint_2[22:22], choice_2, i_2r0[22:22]);
  AND2 I247 (gfint_2[23:23], choice_2, i_2r0[23:23]);
  AND2 I248 (gfint_2[24:24], choice_2, i_2r0[24:24]);
  AND2 I249 (gfint_2[25:25], choice_2, i_2r0[25:25]);
  AND2 I250 (gfint_2[26:26], choice_2, i_2r0[26:26]);
  AND2 I251 (gfint_2[27:27], choice_2, i_2r0[27:27]);
  AND2 I252 (gfint_2[28:28], choice_2, i_2r0[28:28]);
  AND2 I253 (gfint_2[29:29], choice_2, i_2r0[29:29]);
  AND2 I254 (gfint_2[30:30], choice_2, i_2r0[30:30]);
  AND2 I255 (gfint_2[31:31], choice_2, i_2r0[31:31]);
  OR2 I256 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I257 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I258 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I259 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I260 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I261 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I262 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I263 (comp0_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I264 (comp0_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I265 (comp0_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I266 (comp0_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I267 (comp0_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I268 (comp0_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I269 (comp0_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I270 (comp0_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I271 (comp0_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I272 (comp0_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I273 (comp0_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I274 (comp0_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I275 (comp0_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I276 (comp0_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I277 (comp0_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I278 (comp0_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I279 (comp0_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I280 (comp0_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I281 (comp0_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I282 (comp0_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I283 (comp0_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I284 (comp0_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I285 (comp0_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I286 (comp0_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I287 (comp0_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  C3 I288 (simp3031_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I289 (simp3031_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I290 (simp3031_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I291 (simp3031_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I292 (simp3031_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I293 (simp3031_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I294 (simp3031_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I295 (simp3031_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I296 (simp3031_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I297 (simp3031_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I298 (simp3031_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I299 (simp3032_0[0:0], simp3031_0[0:0], simp3031_0[1:1], simp3031_0[2:2]);
  C3 I300 (simp3032_0[1:1], simp3031_0[3:3], simp3031_0[4:4], simp3031_0[5:5]);
  C3 I301 (simp3032_0[2:2], simp3031_0[6:6], simp3031_0[7:7], simp3031_0[8:8]);
  C2 I302 (simp3032_0[3:3], simp3031_0[9:9], simp3031_0[10:10]);
  C3 I303 (simp3033_0[0:0], simp3032_0[0:0], simp3032_0[1:1], simp3032_0[2:2]);
  BUFF I304 (simp3033_0[1:1], simp3032_0[3:3]);
  C2 I305 (icomp_0, simp3033_0[0:0], simp3033_0[1:1]);
  OR2 I306 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I307 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I308 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I309 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I310 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I311 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I312 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  OR2 I313 (comp1_0[7:7], i_1r0[7:7], i_1r1[7:7]);
  OR2 I314 (comp1_0[8:8], i_1r0[8:8], i_1r1[8:8]);
  OR2 I315 (comp1_0[9:9], i_1r0[9:9], i_1r1[9:9]);
  OR2 I316 (comp1_0[10:10], i_1r0[10:10], i_1r1[10:10]);
  OR2 I317 (comp1_0[11:11], i_1r0[11:11], i_1r1[11:11]);
  OR2 I318 (comp1_0[12:12], i_1r0[12:12], i_1r1[12:12]);
  OR2 I319 (comp1_0[13:13], i_1r0[13:13], i_1r1[13:13]);
  OR2 I320 (comp1_0[14:14], i_1r0[14:14], i_1r1[14:14]);
  OR2 I321 (comp1_0[15:15], i_1r0[15:15], i_1r1[15:15]);
  OR2 I322 (comp1_0[16:16], i_1r0[16:16], i_1r1[16:16]);
  OR2 I323 (comp1_0[17:17], i_1r0[17:17], i_1r1[17:17]);
  OR2 I324 (comp1_0[18:18], i_1r0[18:18], i_1r1[18:18]);
  OR2 I325 (comp1_0[19:19], i_1r0[19:19], i_1r1[19:19]);
  OR2 I326 (comp1_0[20:20], i_1r0[20:20], i_1r1[20:20]);
  OR2 I327 (comp1_0[21:21], i_1r0[21:21], i_1r1[21:21]);
  OR2 I328 (comp1_0[22:22], i_1r0[22:22], i_1r1[22:22]);
  OR2 I329 (comp1_0[23:23], i_1r0[23:23], i_1r1[23:23]);
  OR2 I330 (comp1_0[24:24], i_1r0[24:24], i_1r1[24:24]);
  OR2 I331 (comp1_0[25:25], i_1r0[25:25], i_1r1[25:25]);
  OR2 I332 (comp1_0[26:26], i_1r0[26:26], i_1r1[26:26]);
  OR2 I333 (comp1_0[27:27], i_1r0[27:27], i_1r1[27:27]);
  OR2 I334 (comp1_0[28:28], i_1r0[28:28], i_1r1[28:28]);
  OR2 I335 (comp1_0[29:29], i_1r0[29:29], i_1r1[29:29]);
  OR2 I336 (comp1_0[30:30], i_1r0[30:30], i_1r1[30:30]);
  OR2 I337 (comp1_0[31:31], i_1r0[31:31], i_1r1[31:31]);
  C3 I338 (simp3371_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I339 (simp3371_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  C3 I340 (simp3371_0[2:2], comp1_0[6:6], comp1_0[7:7], comp1_0[8:8]);
  C3 I341 (simp3371_0[3:3], comp1_0[9:9], comp1_0[10:10], comp1_0[11:11]);
  C3 I342 (simp3371_0[4:4], comp1_0[12:12], comp1_0[13:13], comp1_0[14:14]);
  C3 I343 (simp3371_0[5:5], comp1_0[15:15], comp1_0[16:16], comp1_0[17:17]);
  C3 I344 (simp3371_0[6:6], comp1_0[18:18], comp1_0[19:19], comp1_0[20:20]);
  C3 I345 (simp3371_0[7:7], comp1_0[21:21], comp1_0[22:22], comp1_0[23:23]);
  C3 I346 (simp3371_0[8:8], comp1_0[24:24], comp1_0[25:25], comp1_0[26:26]);
  C3 I347 (simp3371_0[9:9], comp1_0[27:27], comp1_0[28:28], comp1_0[29:29]);
  C2 I348 (simp3371_0[10:10], comp1_0[30:30], comp1_0[31:31]);
  C3 I349 (simp3372_0[0:0], simp3371_0[0:0], simp3371_0[1:1], simp3371_0[2:2]);
  C3 I350 (simp3372_0[1:1], simp3371_0[3:3], simp3371_0[4:4], simp3371_0[5:5]);
  C3 I351 (simp3372_0[2:2], simp3371_0[6:6], simp3371_0[7:7], simp3371_0[8:8]);
  C2 I352 (simp3372_0[3:3], simp3371_0[9:9], simp3371_0[10:10]);
  C3 I353 (simp3373_0[0:0], simp3372_0[0:0], simp3372_0[1:1], simp3372_0[2:2]);
  BUFF I354 (simp3373_0[1:1], simp3372_0[3:3]);
  C2 I355 (icomp_1, simp3373_0[0:0], simp3373_0[1:1]);
  OR2 I356 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I357 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I358 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2 I359 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  OR2 I360 (comp2_0[4:4], i_2r0[4:4], i_2r1[4:4]);
  OR2 I361 (comp2_0[5:5], i_2r0[5:5], i_2r1[5:5]);
  OR2 I362 (comp2_0[6:6], i_2r0[6:6], i_2r1[6:6]);
  OR2 I363 (comp2_0[7:7], i_2r0[7:7], i_2r1[7:7]);
  OR2 I364 (comp2_0[8:8], i_2r0[8:8], i_2r1[8:8]);
  OR2 I365 (comp2_0[9:9], i_2r0[9:9], i_2r1[9:9]);
  OR2 I366 (comp2_0[10:10], i_2r0[10:10], i_2r1[10:10]);
  OR2 I367 (comp2_0[11:11], i_2r0[11:11], i_2r1[11:11]);
  OR2 I368 (comp2_0[12:12], i_2r0[12:12], i_2r1[12:12]);
  OR2 I369 (comp2_0[13:13], i_2r0[13:13], i_2r1[13:13]);
  OR2 I370 (comp2_0[14:14], i_2r0[14:14], i_2r1[14:14]);
  OR2 I371 (comp2_0[15:15], i_2r0[15:15], i_2r1[15:15]);
  OR2 I372 (comp2_0[16:16], i_2r0[16:16], i_2r1[16:16]);
  OR2 I373 (comp2_0[17:17], i_2r0[17:17], i_2r1[17:17]);
  OR2 I374 (comp2_0[18:18], i_2r0[18:18], i_2r1[18:18]);
  OR2 I375 (comp2_0[19:19], i_2r0[19:19], i_2r1[19:19]);
  OR2 I376 (comp2_0[20:20], i_2r0[20:20], i_2r1[20:20]);
  OR2 I377 (comp2_0[21:21], i_2r0[21:21], i_2r1[21:21]);
  OR2 I378 (comp2_0[22:22], i_2r0[22:22], i_2r1[22:22]);
  OR2 I379 (comp2_0[23:23], i_2r0[23:23], i_2r1[23:23]);
  OR2 I380 (comp2_0[24:24], i_2r0[24:24], i_2r1[24:24]);
  OR2 I381 (comp2_0[25:25], i_2r0[25:25], i_2r1[25:25]);
  OR2 I382 (comp2_0[26:26], i_2r0[26:26], i_2r1[26:26]);
  OR2 I383 (comp2_0[27:27], i_2r0[27:27], i_2r1[27:27]);
  OR2 I384 (comp2_0[28:28], i_2r0[28:28], i_2r1[28:28]);
  OR2 I385 (comp2_0[29:29], i_2r0[29:29], i_2r1[29:29]);
  OR2 I386 (comp2_0[30:30], i_2r0[30:30], i_2r1[30:30]);
  OR2 I387 (comp2_0[31:31], i_2r0[31:31], i_2r1[31:31]);
  C3 I388 (simp3711_0[0:0], comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C3 I389 (simp3711_0[1:1], comp2_0[3:3], comp2_0[4:4], comp2_0[5:5]);
  C3 I390 (simp3711_0[2:2], comp2_0[6:6], comp2_0[7:7], comp2_0[8:8]);
  C3 I391 (simp3711_0[3:3], comp2_0[9:9], comp2_0[10:10], comp2_0[11:11]);
  C3 I392 (simp3711_0[4:4], comp2_0[12:12], comp2_0[13:13], comp2_0[14:14]);
  C3 I393 (simp3711_0[5:5], comp2_0[15:15], comp2_0[16:16], comp2_0[17:17]);
  C3 I394 (simp3711_0[6:6], comp2_0[18:18], comp2_0[19:19], comp2_0[20:20]);
  C3 I395 (simp3711_0[7:7], comp2_0[21:21], comp2_0[22:22], comp2_0[23:23]);
  C3 I396 (simp3711_0[8:8], comp2_0[24:24], comp2_0[25:25], comp2_0[26:26]);
  C3 I397 (simp3711_0[9:9], comp2_0[27:27], comp2_0[28:28], comp2_0[29:29]);
  C2 I398 (simp3711_0[10:10], comp2_0[30:30], comp2_0[31:31]);
  C3 I399 (simp3712_0[0:0], simp3711_0[0:0], simp3711_0[1:1], simp3711_0[2:2]);
  C3 I400 (simp3712_0[1:1], simp3711_0[3:3], simp3711_0[4:4], simp3711_0[5:5]);
  C3 I401 (simp3712_0[2:2], simp3711_0[6:6], simp3711_0[7:7], simp3711_0[8:8]);
  C2 I402 (simp3712_0[3:3], simp3711_0[9:9], simp3711_0[10:10]);
  C3 I403 (simp3713_0[0:0], simp3712_0[0:0], simp3712_0[1:1], simp3712_0[2:2]);
  BUFF I404 (simp3713_0[1:1], simp3712_0[3:3]);
  C2 I405 (icomp_2, simp3713_0[0:0], simp3713_0[1:1]);
  C2R I406 (choice_0, icomp_0, nchosen_0, reset);
  C2R I407 (choice_1, icomp_1, nchosen_0, reset);
  C2R I408 (choice_2, icomp_2, nchosen_0, reset);
  OR3 I409 (anychoice_0, choice_0, choice_1, choice_2);
  NOR2 I410 (nchosen_0, anychoice_0, o_0a);
  C2R I411 (i_0a, choice_0, o_0a, reset);
  C2R I412 (i_1a, choice_1, o_0a, reset);
  C2R I413 (i_2a, choice_2, o_0a, reset);
endmodule

// tkvpc32_wo0w32_ro0w32o0w32o0w32 TeakV "pc" 32 [] [0] [0,0,0] [Many [32],Many [0],Many [0,0,0],Many [
//   32,32,32]]
module tkvpc32_wo0w32_ro0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp6001_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I521 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I522 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I523 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I524 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I525 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I526 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I527 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I528 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I529 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I530 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I531 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I532 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I533 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I534 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I535 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I536 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I537 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I538 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I539 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I540 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I541 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I542 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I543 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I544 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I545 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I546 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I547 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I548 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I549 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I550 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I551 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I552 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I553 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I554 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I555 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I556 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I557 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I558 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I559 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I560 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I561 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I562 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I563 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I564 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I565 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I566 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I567 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I568 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I569 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I570 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I571 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I572 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I573 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I574 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I575 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I576 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I577 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I578 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I579 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I580 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I581 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I582 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I583 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I608 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I609 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I610 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I611 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I612 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I613 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I614 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I615 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  NOR3 I616 (simp6001_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I617 (simp6001_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I618 (anyread_0, simp6001_0[0:0], simp6001_0[1:1]);
  BUFF I619 (wg_0a, wd_0a);
  BUFF I620 (rg_0a, rd_0a);
  BUFF I621 (rg_1a, rd_1a);
  BUFF I622 (rg_2a, rd_2a);
endmodule

// tkj32m32_0 TeakJ [Many [32,0],One 32]
module tkj32m32_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [31:0] joinf_0;
  wire [31:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joint_0[0:0], i_0r1[0:0]);
  BUFF I33 (joint_0[1:1], i_0r1[1:1]);
  BUFF I34 (joint_0[2:2], i_0r1[2:2]);
  BUFF I35 (joint_0[3:3], i_0r1[3:3]);
  BUFF I36 (joint_0[4:4], i_0r1[4:4]);
  BUFF I37 (joint_0[5:5], i_0r1[5:5]);
  BUFF I38 (joint_0[6:6], i_0r1[6:6]);
  BUFF I39 (joint_0[7:7], i_0r1[7:7]);
  BUFF I40 (joint_0[8:8], i_0r1[8:8]);
  BUFF I41 (joint_0[9:9], i_0r1[9:9]);
  BUFF I42 (joint_0[10:10], i_0r1[10:10]);
  BUFF I43 (joint_0[11:11], i_0r1[11:11]);
  BUFF I44 (joint_0[12:12], i_0r1[12:12]);
  BUFF I45 (joint_0[13:13], i_0r1[13:13]);
  BUFF I46 (joint_0[14:14], i_0r1[14:14]);
  BUFF I47 (joint_0[15:15], i_0r1[15:15]);
  BUFF I48 (joint_0[16:16], i_0r1[16:16]);
  BUFF I49 (joint_0[17:17], i_0r1[17:17]);
  BUFF I50 (joint_0[18:18], i_0r1[18:18]);
  BUFF I51 (joint_0[19:19], i_0r1[19:19]);
  BUFF I52 (joint_0[20:20], i_0r1[20:20]);
  BUFF I53 (joint_0[21:21], i_0r1[21:21]);
  BUFF I54 (joint_0[22:22], i_0r1[22:22]);
  BUFF I55 (joint_0[23:23], i_0r1[23:23]);
  BUFF I56 (joint_0[24:24], i_0r1[24:24]);
  BUFF I57 (joint_0[25:25], i_0r1[25:25]);
  BUFF I58 (joint_0[26:26], i_0r1[26:26]);
  BUFF I59 (joint_0[27:27], i_0r1[27:27]);
  BUFF I60 (joint_0[28:28], i_0r1[28:28]);
  BUFF I61 (joint_0[29:29], i_0r1[29:29]);
  BUFF I62 (joint_0[30:30], i_0r1[30:30]);
  BUFF I63 (joint_0[31:31], i_0r1[31:31]);
  BUFF I64 (icomplete_0, i_1r);
  C2 I65 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I66 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I67 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I68 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I69 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I70 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I71 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I72 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I73 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I74 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I75 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I76 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I77 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I78 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I79 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I80 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I81 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I82 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I83 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I84 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I85 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I86 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I87 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I88 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I89 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I90 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I91 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I92 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I93 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I94 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I95 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I96 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I97 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I98 (o_0r1[1:1], joint_0[1:1]);
  BUFF I99 (o_0r1[2:2], joint_0[2:2]);
  BUFF I100 (o_0r1[3:3], joint_0[3:3]);
  BUFF I101 (o_0r1[4:4], joint_0[4:4]);
  BUFF I102 (o_0r1[5:5], joint_0[5:5]);
  BUFF I103 (o_0r1[6:6], joint_0[6:6]);
  BUFF I104 (o_0r1[7:7], joint_0[7:7]);
  BUFF I105 (o_0r1[8:8], joint_0[8:8]);
  BUFF I106 (o_0r1[9:9], joint_0[9:9]);
  BUFF I107 (o_0r1[10:10], joint_0[10:10]);
  BUFF I108 (o_0r1[11:11], joint_0[11:11]);
  BUFF I109 (o_0r1[12:12], joint_0[12:12]);
  BUFF I110 (o_0r1[13:13], joint_0[13:13]);
  BUFF I111 (o_0r1[14:14], joint_0[14:14]);
  BUFF I112 (o_0r1[15:15], joint_0[15:15]);
  BUFF I113 (o_0r1[16:16], joint_0[16:16]);
  BUFF I114 (o_0r1[17:17], joint_0[17:17]);
  BUFF I115 (o_0r1[18:18], joint_0[18:18]);
  BUFF I116 (o_0r1[19:19], joint_0[19:19]);
  BUFF I117 (o_0r1[20:20], joint_0[20:20]);
  BUFF I118 (o_0r1[21:21], joint_0[21:21]);
  BUFF I119 (o_0r1[22:22], joint_0[22:22]);
  BUFF I120 (o_0r1[23:23], joint_0[23:23]);
  BUFF I121 (o_0r1[24:24], joint_0[24:24]);
  BUFF I122 (o_0r1[25:25], joint_0[25:25]);
  BUFF I123 (o_0r1[26:26], joint_0[26:26]);
  BUFF I124 (o_0r1[27:27], joint_0[27:27]);
  BUFF I125 (o_0r1[28:28], joint_0[28:28]);
  BUFF I126 (o_0r1[29:29], joint_0[29:29]);
  BUFF I127 (o_0r1[30:30], joint_0[30:30]);
  BUFF I128 (o_0r1[31:31], joint_0[31:31]);
  BUFF I129 (i_0a, o_0a);
  BUFF I130 (i_1a, o_0a);
endmodule

// tkf65mo0w0_o0w65 TeakF [0,0] [One 65,Many [0,65]]
module tkf65mo0w0_o0w65 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [64:0] i_0r0;
  input [64:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [64:0] o_1r0;
  output [64:0] o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_1r0[0:0], i_0r0[0:0]);
  BUFF I3 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I4 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I5 (o_1r0[3:3], i_0r0[3:3]);
  BUFF I6 (o_1r0[4:4], i_0r0[4:4]);
  BUFF I7 (o_1r0[5:5], i_0r0[5:5]);
  BUFF I8 (o_1r0[6:6], i_0r0[6:6]);
  BUFF I9 (o_1r0[7:7], i_0r0[7:7]);
  BUFF I10 (o_1r0[8:8], i_0r0[8:8]);
  BUFF I11 (o_1r0[9:9], i_0r0[9:9]);
  BUFF I12 (o_1r0[10:10], i_0r0[10:10]);
  BUFF I13 (o_1r0[11:11], i_0r0[11:11]);
  BUFF I14 (o_1r0[12:12], i_0r0[12:12]);
  BUFF I15 (o_1r0[13:13], i_0r0[13:13]);
  BUFF I16 (o_1r0[14:14], i_0r0[14:14]);
  BUFF I17 (o_1r0[15:15], i_0r0[15:15]);
  BUFF I18 (o_1r0[16:16], i_0r0[16:16]);
  BUFF I19 (o_1r0[17:17], i_0r0[17:17]);
  BUFF I20 (o_1r0[18:18], i_0r0[18:18]);
  BUFF I21 (o_1r0[19:19], i_0r0[19:19]);
  BUFF I22 (o_1r0[20:20], i_0r0[20:20]);
  BUFF I23 (o_1r0[21:21], i_0r0[21:21]);
  BUFF I24 (o_1r0[22:22], i_0r0[22:22]);
  BUFF I25 (o_1r0[23:23], i_0r0[23:23]);
  BUFF I26 (o_1r0[24:24], i_0r0[24:24]);
  BUFF I27 (o_1r0[25:25], i_0r0[25:25]);
  BUFF I28 (o_1r0[26:26], i_0r0[26:26]);
  BUFF I29 (o_1r0[27:27], i_0r0[27:27]);
  BUFF I30 (o_1r0[28:28], i_0r0[28:28]);
  BUFF I31 (o_1r0[29:29], i_0r0[29:29]);
  BUFF I32 (o_1r0[30:30], i_0r0[30:30]);
  BUFF I33 (o_1r0[31:31], i_0r0[31:31]);
  BUFF I34 (o_1r0[32:32], i_0r0[32:32]);
  BUFF I35 (o_1r0[33:33], i_0r0[33:33]);
  BUFF I36 (o_1r0[34:34], i_0r0[34:34]);
  BUFF I37 (o_1r0[35:35], i_0r0[35:35]);
  BUFF I38 (o_1r0[36:36], i_0r0[36:36]);
  BUFF I39 (o_1r0[37:37], i_0r0[37:37]);
  BUFF I40 (o_1r0[38:38], i_0r0[38:38]);
  BUFF I41 (o_1r0[39:39], i_0r0[39:39]);
  BUFF I42 (o_1r0[40:40], i_0r0[40:40]);
  BUFF I43 (o_1r0[41:41], i_0r0[41:41]);
  BUFF I44 (o_1r0[42:42], i_0r0[42:42]);
  BUFF I45 (o_1r0[43:43], i_0r0[43:43]);
  BUFF I46 (o_1r0[44:44], i_0r0[44:44]);
  BUFF I47 (o_1r0[45:45], i_0r0[45:45]);
  BUFF I48 (o_1r0[46:46], i_0r0[46:46]);
  BUFF I49 (o_1r0[47:47], i_0r0[47:47]);
  BUFF I50 (o_1r0[48:48], i_0r0[48:48]);
  BUFF I51 (o_1r0[49:49], i_0r0[49:49]);
  BUFF I52 (o_1r0[50:50], i_0r0[50:50]);
  BUFF I53 (o_1r0[51:51], i_0r0[51:51]);
  BUFF I54 (o_1r0[52:52], i_0r0[52:52]);
  BUFF I55 (o_1r0[53:53], i_0r0[53:53]);
  BUFF I56 (o_1r0[54:54], i_0r0[54:54]);
  BUFF I57 (o_1r0[55:55], i_0r0[55:55]);
  BUFF I58 (o_1r0[56:56], i_0r0[56:56]);
  BUFF I59 (o_1r0[57:57], i_0r0[57:57]);
  BUFF I60 (o_1r0[58:58], i_0r0[58:58]);
  BUFF I61 (o_1r0[59:59], i_0r0[59:59]);
  BUFF I62 (o_1r0[60:60], i_0r0[60:60]);
  BUFF I63 (o_1r0[61:61], i_0r0[61:61]);
  BUFF I64 (o_1r0[62:62], i_0r0[62:62]);
  BUFF I65 (o_1r0[63:63], i_0r0[63:63]);
  BUFF I66 (o_1r0[64:64], i_0r0[64:64]);
  BUFF I67 (o_1r1[0:0], i_0r1[0:0]);
  BUFF I68 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I69 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I70 (o_1r1[3:3], i_0r1[3:3]);
  BUFF I71 (o_1r1[4:4], i_0r1[4:4]);
  BUFF I72 (o_1r1[5:5], i_0r1[5:5]);
  BUFF I73 (o_1r1[6:6], i_0r1[6:6]);
  BUFF I74 (o_1r1[7:7], i_0r1[7:7]);
  BUFF I75 (o_1r1[8:8], i_0r1[8:8]);
  BUFF I76 (o_1r1[9:9], i_0r1[9:9]);
  BUFF I77 (o_1r1[10:10], i_0r1[10:10]);
  BUFF I78 (o_1r1[11:11], i_0r1[11:11]);
  BUFF I79 (o_1r1[12:12], i_0r1[12:12]);
  BUFF I80 (o_1r1[13:13], i_0r1[13:13]);
  BUFF I81 (o_1r1[14:14], i_0r1[14:14]);
  BUFF I82 (o_1r1[15:15], i_0r1[15:15]);
  BUFF I83 (o_1r1[16:16], i_0r1[16:16]);
  BUFF I84 (o_1r1[17:17], i_0r1[17:17]);
  BUFF I85 (o_1r1[18:18], i_0r1[18:18]);
  BUFF I86 (o_1r1[19:19], i_0r1[19:19]);
  BUFF I87 (o_1r1[20:20], i_0r1[20:20]);
  BUFF I88 (o_1r1[21:21], i_0r1[21:21]);
  BUFF I89 (o_1r1[22:22], i_0r1[22:22]);
  BUFF I90 (o_1r1[23:23], i_0r1[23:23]);
  BUFF I91 (o_1r1[24:24], i_0r1[24:24]);
  BUFF I92 (o_1r1[25:25], i_0r1[25:25]);
  BUFF I93 (o_1r1[26:26], i_0r1[26:26]);
  BUFF I94 (o_1r1[27:27], i_0r1[27:27]);
  BUFF I95 (o_1r1[28:28], i_0r1[28:28]);
  BUFF I96 (o_1r1[29:29], i_0r1[29:29]);
  BUFF I97 (o_1r1[30:30], i_0r1[30:30]);
  BUFF I98 (o_1r1[31:31], i_0r1[31:31]);
  BUFF I99 (o_1r1[32:32], i_0r1[32:32]);
  BUFF I100 (o_1r1[33:33], i_0r1[33:33]);
  BUFF I101 (o_1r1[34:34], i_0r1[34:34]);
  BUFF I102 (o_1r1[35:35], i_0r1[35:35]);
  BUFF I103 (o_1r1[36:36], i_0r1[36:36]);
  BUFF I104 (o_1r1[37:37], i_0r1[37:37]);
  BUFF I105 (o_1r1[38:38], i_0r1[38:38]);
  BUFF I106 (o_1r1[39:39], i_0r1[39:39]);
  BUFF I107 (o_1r1[40:40], i_0r1[40:40]);
  BUFF I108 (o_1r1[41:41], i_0r1[41:41]);
  BUFF I109 (o_1r1[42:42], i_0r1[42:42]);
  BUFF I110 (o_1r1[43:43], i_0r1[43:43]);
  BUFF I111 (o_1r1[44:44], i_0r1[44:44]);
  BUFF I112 (o_1r1[45:45], i_0r1[45:45]);
  BUFF I113 (o_1r1[46:46], i_0r1[46:46]);
  BUFF I114 (o_1r1[47:47], i_0r1[47:47]);
  BUFF I115 (o_1r1[48:48], i_0r1[48:48]);
  BUFF I116 (o_1r1[49:49], i_0r1[49:49]);
  BUFF I117 (o_1r1[50:50], i_0r1[50:50]);
  BUFF I118 (o_1r1[51:51], i_0r1[51:51]);
  BUFF I119 (o_1r1[52:52], i_0r1[52:52]);
  BUFF I120 (o_1r1[53:53], i_0r1[53:53]);
  BUFF I121 (o_1r1[54:54], i_0r1[54:54]);
  BUFF I122 (o_1r1[55:55], i_0r1[55:55]);
  BUFF I123 (o_1r1[56:56], i_0r1[56:56]);
  BUFF I124 (o_1r1[57:57], i_0r1[57:57]);
  BUFF I125 (o_1r1[58:58], i_0r1[58:58]);
  BUFF I126 (o_1r1[59:59], i_0r1[59:59]);
  BUFF I127 (o_1r1[60:60], i_0r1[60:60]);
  BUFF I128 (o_1r1[61:61], i_0r1[61:61]);
  BUFF I129 (o_1r1[62:62], i_0r1[62:62]);
  BUFF I130 (o_1r1[63:63], i_0r1[63:63]);
  BUFF I131 (o_1r1[64:64], i_0r1[64:64]);
  BUFF I132 (o_0r, icomplete_0);
  C3 I133 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tko0m4_1nm4b8 TeakO [
//     (1,TeakOConstant 4 8)] [One 0,One 4]
module tko0m4_1nm4b8 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[3:3], i_0r);
  GND I1 (o_0r0[3:3]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  GND I5 (o_0r1[0:0]);
  GND I6 (o_0r1[1:1]);
  GND I7 (o_0r1[2:2]);
  BUFF I8 (i_0a, o_0a);
endmodule

// tko1m1_1noti0w1b TeakO [
//     (1,TeakOp TeakOpNot [(0,0+:1)])] [One 1,One 1]
module tko1m1_1noti0w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1, i_0r0);
  BUFF I1 (o_0r0, i_0r1);
  BUFF I2 (i_0a, o_0a);
endmodule

// tkj3m1_1_1 TeakJ [Many [1,1,1],One 3]
module tkj3m1_1_1 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input i_1r0;
  input i_1r1;
  output i_1a;
  input i_2r0;
  input i_2r1;
  output i_2a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [2:0] joinf_0;
  wire [2:0] joint_0;
  wire dcomplete_0;
  wire dcomplete_1;
  BUFF I0 (joinf_0[0:0], i_0r0);
  BUFF I1 (joinf_0[1:1], i_1r0);
  BUFF I2 (joinf_0[2:2], i_2r0);
  BUFF I3 (joint_0[0:0], i_0r1);
  BUFF I4 (joint_0[1:1], i_1r1);
  BUFF I5 (joint_0[2:2], i_2r1);
  OR2 I6 (dcomplete_0, i_1r0, i_1r1);
  OR2 I7 (dcomplete_1, i_2r0, i_2r1);
  C2 I8 (icomplete_0, dcomplete_0, dcomplete_1);
  C2 I9 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I10 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I11 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I12 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I13 (o_0r1[1:1], joint_0[1:1]);
  BUFF I14 (o_0r1[2:2], joint_0[2:2]);
  BUFF I15 (i_0a, o_0a);
  BUFF I16 (i_1a, o_0a);
  BUFF I17 (i_2a, o_0a);
endmodule

// tko0m5_1nm5b0 TeakO [
//     (1,TeakOConstant 5 0)] [One 0,One 5]
module tko0m5_1nm5b0 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [4:0] o_0r0;
  output [4:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r);
  BUFF I1 (o_0r0[1:1], i_0r);
  BUFF I2 (o_0r0[2:2], i_0r);
  BUFF I3 (o_0r0[3:3], i_0r);
  BUFF I4 (o_0r0[4:4], i_0r);
  GND I5 (o_0r1[0:0]);
  GND I6 (o_0r1[1:1]);
  GND I7 (o_0r1[2:2]);
  GND I8 (o_0r1[3:3]);
  GND I9 (o_0r1[4:4]);
  BUFF I10 (i_0a, o_0a);
endmodule

// tkj15m5_5_5 TeakJ [Many [5,5,5],One 15]
module tkj15m5_5_5 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, o_0r0, o_0r1, o_0a, reset);
  input [4:0] i_0r0;
  input [4:0] i_0r1;
  output i_0a;
  input [4:0] i_1r0;
  input [4:0] i_1r1;
  output i_1a;
  input [4:0] i_2r0;
  input [4:0] i_2r1;
  output i_2a;
  output [14:0] o_0r0;
  output [14:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [14:0] joinf_0;
  wire [14:0] joint_0;
  wire dcomplete_0;
  wire dcomplete_1;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_1r0[0:0]);
  BUFF I6 (joinf_0[6:6], i_1r0[1:1]);
  BUFF I7 (joinf_0[7:7], i_1r0[2:2]);
  BUFF I8 (joinf_0[8:8], i_1r0[3:3]);
  BUFF I9 (joinf_0[9:9], i_1r0[4:4]);
  BUFF I10 (joinf_0[10:10], i_2r0[0:0]);
  BUFF I11 (joinf_0[11:11], i_2r0[1:1]);
  BUFF I12 (joinf_0[12:12], i_2r0[2:2]);
  BUFF I13 (joinf_0[13:13], i_2r0[3:3]);
  BUFF I14 (joinf_0[14:14], i_2r0[4:4]);
  BUFF I15 (joint_0[0:0], i_0r1[0:0]);
  BUFF I16 (joint_0[1:1], i_0r1[1:1]);
  BUFF I17 (joint_0[2:2], i_0r1[2:2]);
  BUFF I18 (joint_0[3:3], i_0r1[3:3]);
  BUFF I19 (joint_0[4:4], i_0r1[4:4]);
  BUFF I20 (joint_0[5:5], i_1r1[0:0]);
  BUFF I21 (joint_0[6:6], i_1r1[1:1]);
  BUFF I22 (joint_0[7:7], i_1r1[2:2]);
  BUFF I23 (joint_0[8:8], i_1r1[3:3]);
  BUFF I24 (joint_0[9:9], i_1r1[4:4]);
  BUFF I25 (joint_0[10:10], i_2r1[0:0]);
  BUFF I26 (joint_0[11:11], i_2r1[1:1]);
  BUFF I27 (joint_0[12:12], i_2r1[2:2]);
  BUFF I28 (joint_0[13:13], i_2r1[3:3]);
  BUFF I29 (joint_0[14:14], i_2r1[4:4]);
  OR2 I30 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  OR2 I31 (dcomplete_1, i_2r0[0:0], i_2r1[0:0]);
  C2 I32 (icomplete_0, dcomplete_0, dcomplete_1);
  C2 I33 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I34 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I35 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I36 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I37 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I38 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I39 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I40 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I41 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I42 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I43 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I44 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I45 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I46 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I47 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I48 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I49 (o_0r1[1:1], joint_0[1:1]);
  BUFF I50 (o_0r1[2:2], joint_0[2:2]);
  BUFF I51 (o_0r1[3:3], joint_0[3:3]);
  BUFF I52 (o_0r1[4:4], joint_0[4:4]);
  BUFF I53 (o_0r1[5:5], joint_0[5:5]);
  BUFF I54 (o_0r1[6:6], joint_0[6:6]);
  BUFF I55 (o_0r1[7:7], joint_0[7:7]);
  BUFF I56 (o_0r1[8:8], joint_0[8:8]);
  BUFF I57 (o_0r1[9:9], joint_0[9:9]);
  BUFF I58 (o_0r1[10:10], joint_0[10:10]);
  BUFF I59 (o_0r1[11:11], joint_0[11:11]);
  BUFF I60 (o_0r1[12:12], joint_0[12:12]);
  BUFF I61 (o_0r1[13:13], joint_0[13:13]);
  BUFF I62 (o_0r1[14:14], joint_0[14:14]);
  BUFF I63 (i_0a, o_0a);
  BUFF I64 (i_1a, o_0a);
  BUFF I65 (i_2a, o_0a);
endmodule

// tko13m32_1ap19xi12w1b_2api0w13bt1o0w19b TeakO [
//     (1,TeakOAppend 19 [(0,12+:1)]),
//     (2,TeakOAppend 1 [(0,0+:13),(1,0+:19)])] [One 13,One 32]
module tko13m32_1ap19xi12w1b_2api0w13bt1o0w19b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [12:0] i_0r0;
  input [12:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire [18:0] termf_1;
  wire [18:0] termt_1;
  BUFF I0 (termf_1[0:0], i_0r0[12:12]);
  BUFF I1 (termt_1[0:0], i_0r1[12:12]);
  BUFF I2 (termf_1[1:1], i_0r0[12:12]);
  BUFF I3 (termt_1[1:1], i_0r1[12:12]);
  BUFF I4 (termf_1[2:2], i_0r0[12:12]);
  BUFF I5 (termt_1[2:2], i_0r1[12:12]);
  BUFF I6 (termf_1[3:3], i_0r0[12:12]);
  BUFF I7 (termt_1[3:3], i_0r1[12:12]);
  BUFF I8 (termf_1[4:4], i_0r0[12:12]);
  BUFF I9 (termt_1[4:4], i_0r1[12:12]);
  BUFF I10 (termf_1[5:5], i_0r0[12:12]);
  BUFF I11 (termt_1[5:5], i_0r1[12:12]);
  BUFF I12 (termf_1[6:6], i_0r0[12:12]);
  BUFF I13 (termt_1[6:6], i_0r1[12:12]);
  BUFF I14 (termf_1[7:7], i_0r0[12:12]);
  BUFF I15 (termt_1[7:7], i_0r1[12:12]);
  BUFF I16 (termf_1[8:8], i_0r0[12:12]);
  BUFF I17 (termt_1[8:8], i_0r1[12:12]);
  BUFF I18 (termf_1[9:9], i_0r0[12:12]);
  BUFF I19 (termt_1[9:9], i_0r1[12:12]);
  BUFF I20 (termf_1[10:10], i_0r0[12:12]);
  BUFF I21 (termt_1[10:10], i_0r1[12:12]);
  BUFF I22 (termf_1[11:11], i_0r0[12:12]);
  BUFF I23 (termt_1[11:11], i_0r1[12:12]);
  BUFF I24 (termf_1[12:12], i_0r0[12:12]);
  BUFF I25 (termt_1[12:12], i_0r1[12:12]);
  BUFF I26 (termf_1[13:13], i_0r0[12:12]);
  BUFF I27 (termt_1[13:13], i_0r1[12:12]);
  BUFF I28 (termf_1[14:14], i_0r0[12:12]);
  BUFF I29 (termt_1[14:14], i_0r1[12:12]);
  BUFF I30 (termf_1[15:15], i_0r0[12:12]);
  BUFF I31 (termt_1[15:15], i_0r1[12:12]);
  BUFF I32 (termf_1[16:16], i_0r0[12:12]);
  BUFF I33 (termt_1[16:16], i_0r1[12:12]);
  BUFF I34 (termf_1[17:17], i_0r0[12:12]);
  BUFF I35 (termt_1[17:17], i_0r1[12:12]);
  BUFF I36 (termf_1[18:18], i_0r0[12:12]);
  BUFF I37 (termt_1[18:18], i_0r1[12:12]);
  BUFF I38 (o_0r0[0:0], i_0r0[0:0]);
  BUFF I39 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I40 (o_0r0[2:2], i_0r0[2:2]);
  BUFF I41 (o_0r0[3:3], i_0r0[3:3]);
  BUFF I42 (o_0r0[4:4], i_0r0[4:4]);
  BUFF I43 (o_0r0[5:5], i_0r0[5:5]);
  BUFF I44 (o_0r0[6:6], i_0r0[6:6]);
  BUFF I45 (o_0r0[7:7], i_0r0[7:7]);
  BUFF I46 (o_0r0[8:8], i_0r0[8:8]);
  BUFF I47 (o_0r0[9:9], i_0r0[9:9]);
  BUFF I48 (o_0r0[10:10], i_0r0[10:10]);
  BUFF I49 (o_0r0[11:11], i_0r0[11:11]);
  BUFF I50 (o_0r0[12:12], i_0r0[12:12]);
  BUFF I51 (o_0r0[13:13], termf_1[0:0]);
  BUFF I52 (o_0r0[14:14], termf_1[1:1]);
  BUFF I53 (o_0r0[15:15], termf_1[2:2]);
  BUFF I54 (o_0r0[16:16], termf_1[3:3]);
  BUFF I55 (o_0r0[17:17], termf_1[4:4]);
  BUFF I56 (o_0r0[18:18], termf_1[5:5]);
  BUFF I57 (o_0r0[19:19], termf_1[6:6]);
  BUFF I58 (o_0r0[20:20], termf_1[7:7]);
  BUFF I59 (o_0r0[21:21], termf_1[8:8]);
  BUFF I60 (o_0r0[22:22], termf_1[9:9]);
  BUFF I61 (o_0r0[23:23], termf_1[10:10]);
  BUFF I62 (o_0r0[24:24], termf_1[11:11]);
  BUFF I63 (o_0r0[25:25], termf_1[12:12]);
  BUFF I64 (o_0r0[26:26], termf_1[13:13]);
  BUFF I65 (o_0r0[27:27], termf_1[14:14]);
  BUFF I66 (o_0r0[28:28], termf_1[15:15]);
  BUFF I67 (o_0r0[29:29], termf_1[16:16]);
  BUFF I68 (o_0r0[30:30], termf_1[17:17]);
  BUFF I69 (o_0r0[31:31], termf_1[18:18]);
  BUFF I70 (o_0r1[0:0], i_0r1[0:0]);
  BUFF I71 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I72 (o_0r1[2:2], i_0r1[2:2]);
  BUFF I73 (o_0r1[3:3], i_0r1[3:3]);
  BUFF I74 (o_0r1[4:4], i_0r1[4:4]);
  BUFF I75 (o_0r1[5:5], i_0r1[5:5]);
  BUFF I76 (o_0r1[6:6], i_0r1[6:6]);
  BUFF I77 (o_0r1[7:7], i_0r1[7:7]);
  BUFF I78 (o_0r1[8:8], i_0r1[8:8]);
  BUFF I79 (o_0r1[9:9], i_0r1[9:9]);
  BUFF I80 (o_0r1[10:10], i_0r1[10:10]);
  BUFF I81 (o_0r1[11:11], i_0r1[11:11]);
  BUFF I82 (o_0r1[12:12], i_0r1[12:12]);
  BUFF I83 (o_0r1[13:13], termt_1[0:0]);
  BUFF I84 (o_0r1[14:14], termt_1[1:1]);
  BUFF I85 (o_0r1[15:15], termt_1[2:2]);
  BUFF I86 (o_0r1[16:16], termt_1[3:3]);
  BUFF I87 (o_0r1[17:17], termt_1[4:4]);
  BUFF I88 (o_0r1[18:18], termt_1[5:5]);
  BUFF I89 (o_0r1[19:19], termt_1[6:6]);
  BUFF I90 (o_0r1[20:20], termt_1[7:7]);
  BUFF I91 (o_0r1[21:21], termt_1[8:8]);
  BUFF I92 (o_0r1[22:22], termt_1[9:9]);
  BUFF I93 (o_0r1[23:23], termt_1[10:10]);
  BUFF I94 (o_0r1[24:24], termt_1[11:11]);
  BUFF I95 (o_0r1[25:25], termt_1[12:12]);
  BUFF I96 (o_0r1[26:26], termt_1[13:13]);
  BUFF I97 (o_0r1[27:27], termt_1[14:14]);
  BUFF I98 (o_0r1[28:28], termt_1[15:15]);
  BUFF I99 (o_0r1[29:29], termt_1[16:16]);
  BUFF I100 (o_0r1[30:30], termt_1[17:17]);
  BUFF I101 (o_0r1[31:31], termt_1[18:18]);
  BUFF I102 (i_0a, o_0a);
endmodule

// tko0m4_1nm4b7 TeakO [
//     (1,TeakOConstant 4 7)] [One 0,One 4]
module tko0m4_1nm4b7 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  BUFF I1 (o_0r1[1:1], i_0r);
  BUFF I2 (o_0r1[2:2], i_0r);
  GND I3 (o_0r0[0:0]);
  GND I4 (o_0r0[1:1]);
  GND I5 (o_0r0[2:2]);
  BUFF I6 (o_0r0[3:3], i_0r);
  GND I7 (o_0r1[3:3]);
  BUFF I8 (i_0a, o_0a);
endmodule

// tkj74m3_4_3_15_1_5_6_1_32_4 TeakJ [Many [3,4,3,15,1,5,6,1,32,4],One 74]
module tkj74m3_4_3_15_1_5_6_1_32_4 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, i_4r0, i_4r1, i_4a, i_5r0, i_5r1, i_5a, i_6r0, i_6r1, i_6a, i_7r0, i_7r1, i_7a, i_8r0, i_8r1, i_8a, i_9r0, i_9r1, i_9a, o_0r0, o_0r1, o_0a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  input [3:0] i_1r0;
  input [3:0] i_1r1;
  output i_1a;
  input [2:0] i_2r0;
  input [2:0] i_2r1;
  output i_2a;
  input [14:0] i_3r0;
  input [14:0] i_3r1;
  output i_3a;
  input i_4r0;
  input i_4r1;
  output i_4a;
  input [4:0] i_5r0;
  input [4:0] i_5r1;
  output i_5a;
  input [5:0] i_6r0;
  input [5:0] i_6r1;
  output i_6a;
  input i_7r0;
  input i_7r1;
  output i_7a;
  input [31:0] i_8r0;
  input [31:0] i_8r1;
  output i_8a;
  input [3:0] i_9r0;
  input [3:0] i_9r1;
  output i_9a;
  output [73:0] o_0r0;
  output [73:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [73:0] joinf_0;
  wire [73:0] joint_0;
  wire dcomplete_0;
  wire dcomplete_1;
  wire dcomplete_2;
  wire dcomplete_3;
  wire dcomplete_4;
  wire dcomplete_5;
  wire dcomplete_6;
  wire dcomplete_7;
  wire dcomplete_8;
  wire [2:0] simp1691_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_1r0[0:0]);
  BUFF I4 (joinf_0[4:4], i_1r0[1:1]);
  BUFF I5 (joinf_0[5:5], i_1r0[2:2]);
  BUFF I6 (joinf_0[6:6], i_1r0[3:3]);
  BUFF I7 (joinf_0[7:7], i_2r0[0:0]);
  BUFF I8 (joinf_0[8:8], i_2r0[1:1]);
  BUFF I9 (joinf_0[9:9], i_2r0[2:2]);
  BUFF I10 (joinf_0[10:10], i_3r0[0:0]);
  BUFF I11 (joinf_0[11:11], i_3r0[1:1]);
  BUFF I12 (joinf_0[12:12], i_3r0[2:2]);
  BUFF I13 (joinf_0[13:13], i_3r0[3:3]);
  BUFF I14 (joinf_0[14:14], i_3r0[4:4]);
  BUFF I15 (joinf_0[15:15], i_3r0[5:5]);
  BUFF I16 (joinf_0[16:16], i_3r0[6:6]);
  BUFF I17 (joinf_0[17:17], i_3r0[7:7]);
  BUFF I18 (joinf_0[18:18], i_3r0[8:8]);
  BUFF I19 (joinf_0[19:19], i_3r0[9:9]);
  BUFF I20 (joinf_0[20:20], i_3r0[10:10]);
  BUFF I21 (joinf_0[21:21], i_3r0[11:11]);
  BUFF I22 (joinf_0[22:22], i_3r0[12:12]);
  BUFF I23 (joinf_0[23:23], i_3r0[13:13]);
  BUFF I24 (joinf_0[24:24], i_3r0[14:14]);
  BUFF I25 (joinf_0[25:25], i_4r0);
  BUFF I26 (joinf_0[26:26], i_5r0[0:0]);
  BUFF I27 (joinf_0[27:27], i_5r0[1:1]);
  BUFF I28 (joinf_0[28:28], i_5r0[2:2]);
  BUFF I29 (joinf_0[29:29], i_5r0[3:3]);
  BUFF I30 (joinf_0[30:30], i_5r0[4:4]);
  BUFF I31 (joinf_0[31:31], i_6r0[0:0]);
  BUFF I32 (joinf_0[32:32], i_6r0[1:1]);
  BUFF I33 (joinf_0[33:33], i_6r0[2:2]);
  BUFF I34 (joinf_0[34:34], i_6r0[3:3]);
  BUFF I35 (joinf_0[35:35], i_6r0[4:4]);
  BUFF I36 (joinf_0[36:36], i_6r0[5:5]);
  BUFF I37 (joinf_0[37:37], i_7r0);
  BUFF I38 (joinf_0[38:38], i_8r0[0:0]);
  BUFF I39 (joinf_0[39:39], i_8r0[1:1]);
  BUFF I40 (joinf_0[40:40], i_8r0[2:2]);
  BUFF I41 (joinf_0[41:41], i_8r0[3:3]);
  BUFF I42 (joinf_0[42:42], i_8r0[4:4]);
  BUFF I43 (joinf_0[43:43], i_8r0[5:5]);
  BUFF I44 (joinf_0[44:44], i_8r0[6:6]);
  BUFF I45 (joinf_0[45:45], i_8r0[7:7]);
  BUFF I46 (joinf_0[46:46], i_8r0[8:8]);
  BUFF I47 (joinf_0[47:47], i_8r0[9:9]);
  BUFF I48 (joinf_0[48:48], i_8r0[10:10]);
  BUFF I49 (joinf_0[49:49], i_8r0[11:11]);
  BUFF I50 (joinf_0[50:50], i_8r0[12:12]);
  BUFF I51 (joinf_0[51:51], i_8r0[13:13]);
  BUFF I52 (joinf_0[52:52], i_8r0[14:14]);
  BUFF I53 (joinf_0[53:53], i_8r0[15:15]);
  BUFF I54 (joinf_0[54:54], i_8r0[16:16]);
  BUFF I55 (joinf_0[55:55], i_8r0[17:17]);
  BUFF I56 (joinf_0[56:56], i_8r0[18:18]);
  BUFF I57 (joinf_0[57:57], i_8r0[19:19]);
  BUFF I58 (joinf_0[58:58], i_8r0[20:20]);
  BUFF I59 (joinf_0[59:59], i_8r0[21:21]);
  BUFF I60 (joinf_0[60:60], i_8r0[22:22]);
  BUFF I61 (joinf_0[61:61], i_8r0[23:23]);
  BUFF I62 (joinf_0[62:62], i_8r0[24:24]);
  BUFF I63 (joinf_0[63:63], i_8r0[25:25]);
  BUFF I64 (joinf_0[64:64], i_8r0[26:26]);
  BUFF I65 (joinf_0[65:65], i_8r0[27:27]);
  BUFF I66 (joinf_0[66:66], i_8r0[28:28]);
  BUFF I67 (joinf_0[67:67], i_8r0[29:29]);
  BUFF I68 (joinf_0[68:68], i_8r0[30:30]);
  BUFF I69 (joinf_0[69:69], i_8r0[31:31]);
  BUFF I70 (joinf_0[70:70], i_9r0[0:0]);
  BUFF I71 (joinf_0[71:71], i_9r0[1:1]);
  BUFF I72 (joinf_0[72:72], i_9r0[2:2]);
  BUFF I73 (joinf_0[73:73], i_9r0[3:3]);
  BUFF I74 (joint_0[0:0], i_0r1[0:0]);
  BUFF I75 (joint_0[1:1], i_0r1[1:1]);
  BUFF I76 (joint_0[2:2], i_0r1[2:2]);
  BUFF I77 (joint_0[3:3], i_1r1[0:0]);
  BUFF I78 (joint_0[4:4], i_1r1[1:1]);
  BUFF I79 (joint_0[5:5], i_1r1[2:2]);
  BUFF I80 (joint_0[6:6], i_1r1[3:3]);
  BUFF I81 (joint_0[7:7], i_2r1[0:0]);
  BUFF I82 (joint_0[8:8], i_2r1[1:1]);
  BUFF I83 (joint_0[9:9], i_2r1[2:2]);
  BUFF I84 (joint_0[10:10], i_3r1[0:0]);
  BUFF I85 (joint_0[11:11], i_3r1[1:1]);
  BUFF I86 (joint_0[12:12], i_3r1[2:2]);
  BUFF I87 (joint_0[13:13], i_3r1[3:3]);
  BUFF I88 (joint_0[14:14], i_3r1[4:4]);
  BUFF I89 (joint_0[15:15], i_3r1[5:5]);
  BUFF I90 (joint_0[16:16], i_3r1[6:6]);
  BUFF I91 (joint_0[17:17], i_3r1[7:7]);
  BUFF I92 (joint_0[18:18], i_3r1[8:8]);
  BUFF I93 (joint_0[19:19], i_3r1[9:9]);
  BUFF I94 (joint_0[20:20], i_3r1[10:10]);
  BUFF I95 (joint_0[21:21], i_3r1[11:11]);
  BUFF I96 (joint_0[22:22], i_3r1[12:12]);
  BUFF I97 (joint_0[23:23], i_3r1[13:13]);
  BUFF I98 (joint_0[24:24], i_3r1[14:14]);
  BUFF I99 (joint_0[25:25], i_4r1);
  BUFF I100 (joint_0[26:26], i_5r1[0:0]);
  BUFF I101 (joint_0[27:27], i_5r1[1:1]);
  BUFF I102 (joint_0[28:28], i_5r1[2:2]);
  BUFF I103 (joint_0[29:29], i_5r1[3:3]);
  BUFF I104 (joint_0[30:30], i_5r1[4:4]);
  BUFF I105 (joint_0[31:31], i_6r1[0:0]);
  BUFF I106 (joint_0[32:32], i_6r1[1:1]);
  BUFF I107 (joint_0[33:33], i_6r1[2:2]);
  BUFF I108 (joint_0[34:34], i_6r1[3:3]);
  BUFF I109 (joint_0[35:35], i_6r1[4:4]);
  BUFF I110 (joint_0[36:36], i_6r1[5:5]);
  BUFF I111 (joint_0[37:37], i_7r1);
  BUFF I112 (joint_0[38:38], i_8r1[0:0]);
  BUFF I113 (joint_0[39:39], i_8r1[1:1]);
  BUFF I114 (joint_0[40:40], i_8r1[2:2]);
  BUFF I115 (joint_0[41:41], i_8r1[3:3]);
  BUFF I116 (joint_0[42:42], i_8r1[4:4]);
  BUFF I117 (joint_0[43:43], i_8r1[5:5]);
  BUFF I118 (joint_0[44:44], i_8r1[6:6]);
  BUFF I119 (joint_0[45:45], i_8r1[7:7]);
  BUFF I120 (joint_0[46:46], i_8r1[8:8]);
  BUFF I121 (joint_0[47:47], i_8r1[9:9]);
  BUFF I122 (joint_0[48:48], i_8r1[10:10]);
  BUFF I123 (joint_0[49:49], i_8r1[11:11]);
  BUFF I124 (joint_0[50:50], i_8r1[12:12]);
  BUFF I125 (joint_0[51:51], i_8r1[13:13]);
  BUFF I126 (joint_0[52:52], i_8r1[14:14]);
  BUFF I127 (joint_0[53:53], i_8r1[15:15]);
  BUFF I128 (joint_0[54:54], i_8r1[16:16]);
  BUFF I129 (joint_0[55:55], i_8r1[17:17]);
  BUFF I130 (joint_0[56:56], i_8r1[18:18]);
  BUFF I131 (joint_0[57:57], i_8r1[19:19]);
  BUFF I132 (joint_0[58:58], i_8r1[20:20]);
  BUFF I133 (joint_0[59:59], i_8r1[21:21]);
  BUFF I134 (joint_0[60:60], i_8r1[22:22]);
  BUFF I135 (joint_0[61:61], i_8r1[23:23]);
  BUFF I136 (joint_0[62:62], i_8r1[24:24]);
  BUFF I137 (joint_0[63:63], i_8r1[25:25]);
  BUFF I138 (joint_0[64:64], i_8r1[26:26]);
  BUFF I139 (joint_0[65:65], i_8r1[27:27]);
  BUFF I140 (joint_0[66:66], i_8r1[28:28]);
  BUFF I141 (joint_0[67:67], i_8r1[29:29]);
  BUFF I142 (joint_0[68:68], i_8r1[30:30]);
  BUFF I143 (joint_0[69:69], i_8r1[31:31]);
  BUFF I144 (joint_0[70:70], i_9r1[0:0]);
  BUFF I145 (joint_0[71:71], i_9r1[1:1]);
  BUFF I146 (joint_0[72:72], i_9r1[2:2]);
  BUFF I147 (joint_0[73:73], i_9r1[3:3]);
  OR2 I148 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  OR2 I149 (dcomplete_1, i_2r0[0:0], i_2r1[0:0]);
  OR2 I150 (dcomplete_2, i_3r0[0:0], i_3r1[0:0]);
  OR2 I151 (dcomplete_3, i_4r0, i_4r1);
  OR2 I152 (dcomplete_4, i_5r0[0:0], i_5r1[0:0]);
  OR2 I153 (dcomplete_5, i_6r0[0:0], i_6r1[0:0]);
  OR2 I154 (dcomplete_6, i_7r0, i_7r1);
  OR2 I155 (dcomplete_7, i_8r0[0:0], i_8r1[0:0]);
  OR2 I156 (dcomplete_8, i_9r0[0:0], i_9r1[0:0]);
  C3 I157 (simp1691_0[0:0], dcomplete_0, dcomplete_1, dcomplete_2);
  C3 I158 (simp1691_0[1:1], dcomplete_3, dcomplete_4, dcomplete_5);
  C3 I159 (simp1691_0[2:2], dcomplete_6, dcomplete_7, dcomplete_8);
  C3 I160 (icomplete_0, simp1691_0[0:0], simp1691_0[1:1], simp1691_0[2:2]);
  C2 I161 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I162 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I163 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I164 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I165 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I166 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I167 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I168 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I169 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I170 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I171 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I172 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I173 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I174 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I175 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I176 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I177 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I178 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I179 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I180 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I181 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I182 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I183 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I184 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I185 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I186 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I187 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I188 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I189 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I190 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I191 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I192 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I193 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I194 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I195 (o_0r0[33:33], joinf_0[33:33]);
  BUFF I196 (o_0r0[34:34], joinf_0[34:34]);
  BUFF I197 (o_0r0[35:35], joinf_0[35:35]);
  BUFF I198 (o_0r0[36:36], joinf_0[36:36]);
  BUFF I199 (o_0r0[37:37], joinf_0[37:37]);
  BUFF I200 (o_0r0[38:38], joinf_0[38:38]);
  BUFF I201 (o_0r0[39:39], joinf_0[39:39]);
  BUFF I202 (o_0r0[40:40], joinf_0[40:40]);
  BUFF I203 (o_0r0[41:41], joinf_0[41:41]);
  BUFF I204 (o_0r0[42:42], joinf_0[42:42]);
  BUFF I205 (o_0r0[43:43], joinf_0[43:43]);
  BUFF I206 (o_0r0[44:44], joinf_0[44:44]);
  BUFF I207 (o_0r0[45:45], joinf_0[45:45]);
  BUFF I208 (o_0r0[46:46], joinf_0[46:46]);
  BUFF I209 (o_0r0[47:47], joinf_0[47:47]);
  BUFF I210 (o_0r0[48:48], joinf_0[48:48]);
  BUFF I211 (o_0r0[49:49], joinf_0[49:49]);
  BUFF I212 (o_0r0[50:50], joinf_0[50:50]);
  BUFF I213 (o_0r0[51:51], joinf_0[51:51]);
  BUFF I214 (o_0r0[52:52], joinf_0[52:52]);
  BUFF I215 (o_0r0[53:53], joinf_0[53:53]);
  BUFF I216 (o_0r0[54:54], joinf_0[54:54]);
  BUFF I217 (o_0r0[55:55], joinf_0[55:55]);
  BUFF I218 (o_0r0[56:56], joinf_0[56:56]);
  BUFF I219 (o_0r0[57:57], joinf_0[57:57]);
  BUFF I220 (o_0r0[58:58], joinf_0[58:58]);
  BUFF I221 (o_0r0[59:59], joinf_0[59:59]);
  BUFF I222 (o_0r0[60:60], joinf_0[60:60]);
  BUFF I223 (o_0r0[61:61], joinf_0[61:61]);
  BUFF I224 (o_0r0[62:62], joinf_0[62:62]);
  BUFF I225 (o_0r0[63:63], joinf_0[63:63]);
  BUFF I226 (o_0r0[64:64], joinf_0[64:64]);
  BUFF I227 (o_0r0[65:65], joinf_0[65:65]);
  BUFF I228 (o_0r0[66:66], joinf_0[66:66]);
  BUFF I229 (o_0r0[67:67], joinf_0[67:67]);
  BUFF I230 (o_0r0[68:68], joinf_0[68:68]);
  BUFF I231 (o_0r0[69:69], joinf_0[69:69]);
  BUFF I232 (o_0r0[70:70], joinf_0[70:70]);
  BUFF I233 (o_0r0[71:71], joinf_0[71:71]);
  BUFF I234 (o_0r0[72:72], joinf_0[72:72]);
  BUFF I235 (o_0r0[73:73], joinf_0[73:73]);
  BUFF I236 (o_0r1[1:1], joint_0[1:1]);
  BUFF I237 (o_0r1[2:2], joint_0[2:2]);
  BUFF I238 (o_0r1[3:3], joint_0[3:3]);
  BUFF I239 (o_0r1[4:4], joint_0[4:4]);
  BUFF I240 (o_0r1[5:5], joint_0[5:5]);
  BUFF I241 (o_0r1[6:6], joint_0[6:6]);
  BUFF I242 (o_0r1[7:7], joint_0[7:7]);
  BUFF I243 (o_0r1[8:8], joint_0[8:8]);
  BUFF I244 (o_0r1[9:9], joint_0[9:9]);
  BUFF I245 (o_0r1[10:10], joint_0[10:10]);
  BUFF I246 (o_0r1[11:11], joint_0[11:11]);
  BUFF I247 (o_0r1[12:12], joint_0[12:12]);
  BUFF I248 (o_0r1[13:13], joint_0[13:13]);
  BUFF I249 (o_0r1[14:14], joint_0[14:14]);
  BUFF I250 (o_0r1[15:15], joint_0[15:15]);
  BUFF I251 (o_0r1[16:16], joint_0[16:16]);
  BUFF I252 (o_0r1[17:17], joint_0[17:17]);
  BUFF I253 (o_0r1[18:18], joint_0[18:18]);
  BUFF I254 (o_0r1[19:19], joint_0[19:19]);
  BUFF I255 (o_0r1[20:20], joint_0[20:20]);
  BUFF I256 (o_0r1[21:21], joint_0[21:21]);
  BUFF I257 (o_0r1[22:22], joint_0[22:22]);
  BUFF I258 (o_0r1[23:23], joint_0[23:23]);
  BUFF I259 (o_0r1[24:24], joint_0[24:24]);
  BUFF I260 (o_0r1[25:25], joint_0[25:25]);
  BUFF I261 (o_0r1[26:26], joint_0[26:26]);
  BUFF I262 (o_0r1[27:27], joint_0[27:27]);
  BUFF I263 (o_0r1[28:28], joint_0[28:28]);
  BUFF I264 (o_0r1[29:29], joint_0[29:29]);
  BUFF I265 (o_0r1[30:30], joint_0[30:30]);
  BUFF I266 (o_0r1[31:31], joint_0[31:31]);
  BUFF I267 (o_0r1[32:32], joint_0[32:32]);
  BUFF I268 (o_0r1[33:33], joint_0[33:33]);
  BUFF I269 (o_0r1[34:34], joint_0[34:34]);
  BUFF I270 (o_0r1[35:35], joint_0[35:35]);
  BUFF I271 (o_0r1[36:36], joint_0[36:36]);
  BUFF I272 (o_0r1[37:37], joint_0[37:37]);
  BUFF I273 (o_0r1[38:38], joint_0[38:38]);
  BUFF I274 (o_0r1[39:39], joint_0[39:39]);
  BUFF I275 (o_0r1[40:40], joint_0[40:40]);
  BUFF I276 (o_0r1[41:41], joint_0[41:41]);
  BUFF I277 (o_0r1[42:42], joint_0[42:42]);
  BUFF I278 (o_0r1[43:43], joint_0[43:43]);
  BUFF I279 (o_0r1[44:44], joint_0[44:44]);
  BUFF I280 (o_0r1[45:45], joint_0[45:45]);
  BUFF I281 (o_0r1[46:46], joint_0[46:46]);
  BUFF I282 (o_0r1[47:47], joint_0[47:47]);
  BUFF I283 (o_0r1[48:48], joint_0[48:48]);
  BUFF I284 (o_0r1[49:49], joint_0[49:49]);
  BUFF I285 (o_0r1[50:50], joint_0[50:50]);
  BUFF I286 (o_0r1[51:51], joint_0[51:51]);
  BUFF I287 (o_0r1[52:52], joint_0[52:52]);
  BUFF I288 (o_0r1[53:53], joint_0[53:53]);
  BUFF I289 (o_0r1[54:54], joint_0[54:54]);
  BUFF I290 (o_0r1[55:55], joint_0[55:55]);
  BUFF I291 (o_0r1[56:56], joint_0[56:56]);
  BUFF I292 (o_0r1[57:57], joint_0[57:57]);
  BUFF I293 (o_0r1[58:58], joint_0[58:58]);
  BUFF I294 (o_0r1[59:59], joint_0[59:59]);
  BUFF I295 (o_0r1[60:60], joint_0[60:60]);
  BUFF I296 (o_0r1[61:61], joint_0[61:61]);
  BUFF I297 (o_0r1[62:62], joint_0[62:62]);
  BUFF I298 (o_0r1[63:63], joint_0[63:63]);
  BUFF I299 (o_0r1[64:64], joint_0[64:64]);
  BUFF I300 (o_0r1[65:65], joint_0[65:65]);
  BUFF I301 (o_0r1[66:66], joint_0[66:66]);
  BUFF I302 (o_0r1[67:67], joint_0[67:67]);
  BUFF I303 (o_0r1[68:68], joint_0[68:68]);
  BUFF I304 (o_0r1[69:69], joint_0[69:69]);
  BUFF I305 (o_0r1[70:70], joint_0[70:70]);
  BUFF I306 (o_0r1[71:71], joint_0[71:71]);
  BUFF I307 (o_0r1[72:72], joint_0[72:72]);
  BUFF I308 (o_0r1[73:73], joint_0[73:73]);
  BUFF I309 (i_0a, o_0a);
  BUFF I310 (i_1a, o_0a);
  BUFF I311 (i_2a, o_0a);
  BUFF I312 (i_3a, o_0a);
  BUFF I313 (i_4a, o_0a);
  BUFF I314 (i_5a, o_0a);
  BUFF I315 (i_6a, o_0a);
  BUFF I316 (i_7a, o_0a);
  BUFF I317 (i_8a, o_0a);
  BUFF I318 (i_9a, o_0a);
endmodule

// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 TeakF [0,0,0,0,0,0,0,0,0,
//   0,0,0,0,0] [One 0,Many [0,0,0,0,0,0,0,0,0,0,0,0,0,0]]
module tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, o_5r, o_5a, o_6r, o_6a, o_7r, o_7a, o_8r, o_8a, o_9r, o_9a, o_10r, o_10a, o_11r, o_11a, o_12r, o_12a, o_13r, o_13a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  output o_7r;
  input o_7a;
  output o_8r;
  input o_8a;
  output o_9r;
  input o_9a;
  output o_10r;
  input o_10a;
  output o_11r;
  input o_11a;
  output o_12r;
  input o_12a;
  output o_13r;
  input o_13a;
  input reset;
  wire [4:0] simp11_0;
  wire [1:0] simp12_0;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  BUFF I2 (o_2r, i_0r);
  BUFF I3 (o_3r, i_0r);
  BUFF I4 (o_4r, i_0r);
  BUFF I5 (o_5r, i_0r);
  BUFF I6 (o_6r, i_0r);
  BUFF I7 (o_7r, i_0r);
  BUFF I8 (o_8r, i_0r);
  BUFF I9 (o_9r, i_0r);
  BUFF I10 (o_10r, i_0r);
  BUFF I11 (o_11r, i_0r);
  BUFF I12 (o_12r, i_0r);
  BUFF I13 (o_13r, i_0r);
  C3 I14 (simp11_0[0:0], o_0a, o_1a, o_2a);
  C3 I15 (simp11_0[1:1], o_3a, o_4a, o_5a);
  C3 I16 (simp11_0[2:2], o_6a, o_7a, o_8a);
  C3 I17 (simp11_0[3:3], o_9a, o_10a, o_11a);
  C2 I18 (simp11_0[4:4], o_12a, o_13a);
  C3 I19 (simp12_0[0:0], simp11_0[0:0], simp11_0[1:1], simp11_0[2:2]);
  C2 I20 (simp12_0[1:1], simp11_0[3:3], simp11_0[4:4]);
  C2 I21 (i_0a, simp12_0[0:0], simp12_0[1:1]);
endmodule

// tkvimmOrReg1_wo0w1_ro0w1 TeakV "immOrReg" 1 [] [0] [0] [Many [1],Many [0],Many [0],Many [1]]
module tkvimmOrReg1_wo0w1_ro0w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input wg_0r0;
  input wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  input reset;
  wire wf_0;
  wire wt_0;
  wire df_0;
  wire dt_0;
  wire wc_0;
  wire wacks_0;
  wire wenr_0;
  wire wen_0;
  wire anyread_0;
  wire nreset_0;
  wire drlgf_0;
  wire drlgt_0;
  wire comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire conwgit_0;
  wire conwgif_0;
  wire conwig_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0, wenr_0, nreset_0);
  AND2 I2 (drlgf_0, wf_0, wen_0);
  AND2 I3 (drlgt_0, wt_0, wen_0);
  NOR2 I4 (df_0, dt_0, drlgt_0);
  NOR3 I5 (dt_0, df_0, drlgf_0, reset);
  AO22 I6 (wacks_0, drlgf_0, df_0, drlgt_0, dt_0);
  OR2 I7 (comp0_0, wg_0r0, wg_0r1);
  BUFF I8 (wc_0, comp0_0);
  AND2 I9 (conwgif_0, wg_0r0, conwig_0);
  AND2 I10 (conwgit_0, wg_0r1, conwig_0);
  BUFF I11 (conwigc_0, wc_0);
  AO22 I12 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I13 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I14 (wf_0, conwgif_0);
  BUFF I15 (wt_0, conwgit_0);
  BUFF I16 (wenr_0, wc_0);
  C2 I17 (wd_0r, conwig_0, wacks_0);
  AND2 I18 (rd_0r0, df_0, rg_0r);
  AND2 I19 (rd_0r1, dt_0, rg_0r);
  OR2 I20 (anyread_0, rg_0r, rg_0a);
  BUFF I21 (wg_0a, wd_0a);
  BUFF I22 (rg_0a, rd_0a);
endmodule

// tks1_o0w1_1o0w0_0o0w0 TeakS (0+:1) [([Imp 1 0],0),([Imp 0 0],0)] [One 1,Many [0,0]]
module tks1_o0w1_1o0w0_0o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire comp_0;
  BUFF I0 (sel_0, match0_0);
  BUFF I1 (match0_0, i_0r1);
  BUFF I2 (sel_1, match1_0);
  BUFF I3 (match1_0, i_0r0);
  C2 I4 (gsel_0, sel_0, icomplete_0);
  C2 I5 (gsel_1, sel_1, icomplete_0);
  OR2 I6 (comp_0, i_0r0, i_0r1);
  BUFF I7 (icomplete_0, comp_0);
  BUFF I8 (o_0r, gsel_0);
  BUFF I9 (o_1r, gsel_1);
  OR2 I10 (oack_0, o_0a, o_1a);
  C2 I11 (i_0a, oack_0, icomplete_0);
endmodule

// tks6_o0w6_9c30mac30mbc30mdc30mec30mfc30m20m21m22m23m24m28m2cm30m31m32m33m34m35m36m37m38m3co0w0_0m1m2
//   m3m4m5m6m7m8mcm10m11m12m13m14m15m16m17m18m1cm25m26m27o0w0 TeakS (0+:6) [([Imp 9 48,Imp 10 48,Imp 11 
//   48,Imp 13 48,Imp 14 48,Imp 15 48,Imp 32 0,Imp 33 0,Imp 34 0,Imp 35 0,Imp 36 0,Imp 40 0,Imp 44 0,Imp 
//   48 0,Imp 49 0,Imp 50 0,Imp 51 0,Imp 52 0,Imp 53 0,Imp 54 0,Imp 55 0,Imp 56 0,Imp 60 0],0),([Imp 0 0,
//   Imp 1 0,Imp 2 0,Imp 3 0,Imp 4 0,Imp 5 0,Imp 6 0,Imp 7 0,Imp 8 0,Imp 12 0,Imp 16 0,Imp 17 0,Imp 18 0,
//   Imp 19 0,Imp 20 0,Imp 21 0,Imp 22 0,Imp 23 0,Imp 24 0,Imp 28 0,Imp 37 0,Imp 38 0,Imp 39 0],0)] [One 
//   6,Many [0,0]]
module tks6_o0w6_9c30mac30mbc30mdc30mec30mfc30m20m21m22m23m24m28m2cm30m31m32m33m34m35m36m37m38m3co0w0_0m1m2m3m4m5m6m7m8mcm10m11m12m13m14m15m16m17m18m1cm25m26m27o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input [5:0] i_0r0;
  input [5:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire [22:0] match0_0;
  wire [7:0] simp71_0;
  wire [2:0] simp72_0;
  wire [1:0] simp81_0;
  wire [1:0] simp91_0;
  wire [1:0] simp101_0;
  wire [1:0] simp111_0;
  wire [1:0] simp121_0;
  wire [1:0] simp131_0;
  wire [1:0] simp141_0;
  wire [1:0] simp151_0;
  wire [1:0] simp161_0;
  wire [1:0] simp171_0;
  wire [1:0] simp181_0;
  wire [1:0] simp191_0;
  wire [1:0] simp201_0;
  wire [1:0] simp211_0;
  wire [1:0] simp221_0;
  wire [1:0] simp231_0;
  wire [1:0] simp241_0;
  wire [1:0] simp251_0;
  wire [1:0] simp261_0;
  wire [1:0] simp271_0;
  wire [1:0] simp281_0;
  wire [1:0] simp291_0;
  wire [1:0] simp301_0;
  wire [22:0] match1_0;
  wire [7:0] simp321_0;
  wire [2:0] simp322_0;
  wire [1:0] simp331_0;
  wire [1:0] simp341_0;
  wire [1:0] simp351_0;
  wire [1:0] simp361_0;
  wire [1:0] simp371_0;
  wire [1:0] simp381_0;
  wire [1:0] simp391_0;
  wire [1:0] simp401_0;
  wire [1:0] simp411_0;
  wire [1:0] simp421_0;
  wire [1:0] simp431_0;
  wire [1:0] simp441_0;
  wire [1:0] simp451_0;
  wire [1:0] simp461_0;
  wire [1:0] simp471_0;
  wire [1:0] simp481_0;
  wire [1:0] simp491_0;
  wire [1:0] simp501_0;
  wire [1:0] simp511_0;
  wire [1:0] simp521_0;
  wire [1:0] simp531_0;
  wire [1:0] simp541_0;
  wire [1:0] simp551_0;
  wire [5:0] comp_0;
  wire [1:0] simp651_0;
  NOR3 I0 (simp71_0[0:0], match0_0[0:0], match0_0[1:1], match0_0[2:2]);
  NOR3 I1 (simp71_0[1:1], match0_0[3:3], match0_0[4:4], match0_0[5:5]);
  NOR3 I2 (simp71_0[2:2], match0_0[6:6], match0_0[7:7], match0_0[8:8]);
  NOR3 I3 (simp71_0[3:3], match0_0[9:9], match0_0[10:10], match0_0[11:11]);
  NOR3 I4 (simp71_0[4:4], match0_0[12:12], match0_0[13:13], match0_0[14:14]);
  NOR3 I5 (simp71_0[5:5], match0_0[15:15], match0_0[16:16], match0_0[17:17]);
  NOR3 I6 (simp71_0[6:6], match0_0[18:18], match0_0[19:19], match0_0[20:20]);
  NOR2 I7 (simp71_0[7:7], match0_0[21:21], match0_0[22:22]);
  NAND3 I8 (simp72_0[0:0], simp71_0[0:0], simp71_0[1:1], simp71_0[2:2]);
  NAND3 I9 (simp72_0[1:1], simp71_0[3:3], simp71_0[4:4], simp71_0[5:5]);
  NAND2 I10 (simp72_0[2:2], simp71_0[6:6], simp71_0[7:7]);
  OR3 I11 (sel_0, simp72_0[0:0], simp72_0[1:1], simp72_0[2:2]);
  C3 I12 (simp81_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I13 (simp81_0[1:1], i_0r1[3:3]);
  C2 I14 (match0_0[0:0], simp81_0[0:0], simp81_0[1:1]);
  C3 I15 (simp91_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I16 (simp91_0[1:1], i_0r1[3:3]);
  C2 I17 (match0_0[1:1], simp91_0[0:0], simp91_0[1:1]);
  C3 I18 (simp101_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I19 (simp101_0[1:1], i_0r1[3:3]);
  C2 I20 (match0_0[2:2], simp101_0[0:0], simp101_0[1:1]);
  C3 I21 (simp111_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I22 (simp111_0[1:1], i_0r1[3:3]);
  C2 I23 (match0_0[3:3], simp111_0[0:0], simp111_0[1:1]);
  C3 I24 (simp121_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I25 (simp121_0[1:1], i_0r1[3:3]);
  C2 I26 (match0_0[4:4], simp121_0[0:0], simp121_0[1:1]);
  C3 I27 (simp131_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I28 (simp131_0[1:1], i_0r1[3:3]);
  C2 I29 (match0_0[5:5], simp131_0[0:0], simp131_0[1:1]);
  C3 I30 (simp141_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I31 (simp141_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I32 (match0_0[6:6], simp141_0[0:0], simp141_0[1:1]);
  C3 I33 (simp151_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I34 (simp151_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I35 (match0_0[7:7], simp151_0[0:0], simp151_0[1:1]);
  C3 I36 (simp161_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I37 (simp161_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I38 (match0_0[8:8], simp161_0[0:0], simp161_0[1:1]);
  C3 I39 (simp171_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I40 (simp171_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I41 (match0_0[9:9], simp171_0[0:0], simp171_0[1:1]);
  C3 I42 (simp181_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I43 (simp181_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I44 (match0_0[10:10], simp181_0[0:0], simp181_0[1:1]);
  C3 I45 (simp191_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I46 (simp191_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I47 (match0_0[11:11], simp191_0[0:0], simp191_0[1:1]);
  C3 I48 (simp201_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I49 (simp201_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I50 (match0_0[12:12], simp201_0[0:0], simp201_0[1:1]);
  C3 I51 (simp211_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I52 (simp211_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I53 (match0_0[13:13], simp211_0[0:0], simp211_0[1:1]);
  C3 I54 (simp221_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I55 (simp221_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I56 (match0_0[14:14], simp221_0[0:0], simp221_0[1:1]);
  C3 I57 (simp231_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I58 (simp231_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I59 (match0_0[15:15], simp231_0[0:0], simp231_0[1:1]);
  C3 I60 (simp241_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I61 (simp241_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I62 (match0_0[16:16], simp241_0[0:0], simp241_0[1:1]);
  C3 I63 (simp251_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I64 (simp251_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I65 (match0_0[17:17], simp251_0[0:0], simp251_0[1:1]);
  C3 I66 (simp261_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I67 (simp261_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I68 (match0_0[18:18], simp261_0[0:0], simp261_0[1:1]);
  C3 I69 (simp271_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I70 (simp271_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I71 (match0_0[19:19], simp271_0[0:0], simp271_0[1:1]);
  C3 I72 (simp281_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I73 (simp281_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I74 (match0_0[20:20], simp281_0[0:0], simp281_0[1:1]);
  C3 I75 (simp291_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I76 (simp291_0[1:1], i_0r1[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I77 (match0_0[21:21], simp291_0[0:0], simp291_0[1:1]);
  C3 I78 (simp301_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I79 (simp301_0[1:1], i_0r1[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I80 (match0_0[22:22], simp301_0[0:0], simp301_0[1:1]);
  NOR3 I81 (simp321_0[0:0], match1_0[0:0], match1_0[1:1], match1_0[2:2]);
  NOR3 I82 (simp321_0[1:1], match1_0[3:3], match1_0[4:4], match1_0[5:5]);
  NOR3 I83 (simp321_0[2:2], match1_0[6:6], match1_0[7:7], match1_0[8:8]);
  NOR3 I84 (simp321_0[3:3], match1_0[9:9], match1_0[10:10], match1_0[11:11]);
  NOR3 I85 (simp321_0[4:4], match1_0[12:12], match1_0[13:13], match1_0[14:14]);
  NOR3 I86 (simp321_0[5:5], match1_0[15:15], match1_0[16:16], match1_0[17:17]);
  NOR3 I87 (simp321_0[6:6], match1_0[18:18], match1_0[19:19], match1_0[20:20]);
  NOR2 I88 (simp321_0[7:7], match1_0[21:21], match1_0[22:22]);
  NAND3 I89 (simp322_0[0:0], simp321_0[0:0], simp321_0[1:1], simp321_0[2:2]);
  NAND3 I90 (simp322_0[1:1], simp321_0[3:3], simp321_0[4:4], simp321_0[5:5]);
  NAND2 I91 (simp322_0[2:2], simp321_0[6:6], simp321_0[7:7]);
  OR3 I92 (sel_1, simp322_0[0:0], simp322_0[1:1], simp322_0[2:2]);
  C3 I93 (simp331_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I94 (simp331_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I95 (match1_0[0:0], simp331_0[0:0], simp331_0[1:1]);
  C3 I96 (simp341_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I97 (simp341_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I98 (match1_0[1:1], simp341_0[0:0], simp341_0[1:1]);
  C3 I99 (simp351_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I100 (simp351_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I101 (match1_0[2:2], simp351_0[0:0], simp351_0[1:1]);
  C3 I102 (simp361_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I103 (simp361_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I104 (match1_0[3:3], simp361_0[0:0], simp361_0[1:1]);
  C3 I105 (simp371_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I106 (simp371_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I107 (match1_0[4:4], simp371_0[0:0], simp371_0[1:1]);
  C3 I108 (simp381_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I109 (simp381_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I110 (match1_0[5:5], simp381_0[0:0], simp381_0[1:1]);
  C3 I111 (simp391_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I112 (simp391_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I113 (match1_0[6:6], simp391_0[0:0], simp391_0[1:1]);
  C3 I114 (simp401_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I115 (simp401_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I116 (match1_0[7:7], simp401_0[0:0], simp401_0[1:1]);
  C3 I117 (simp411_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I118 (simp411_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I119 (match1_0[8:8], simp411_0[0:0], simp411_0[1:1]);
  C3 I120 (simp421_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I121 (simp421_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I122 (match1_0[9:9], simp421_0[0:0], simp421_0[1:1]);
  C3 I123 (simp431_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I124 (simp431_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I125 (match1_0[10:10], simp431_0[0:0], simp431_0[1:1]);
  C3 I126 (simp441_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I127 (simp441_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I128 (match1_0[11:11], simp441_0[0:0], simp441_0[1:1]);
  C3 I129 (simp451_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I130 (simp451_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I131 (match1_0[12:12], simp451_0[0:0], simp451_0[1:1]);
  C3 I132 (simp461_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I133 (simp461_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I134 (match1_0[13:13], simp461_0[0:0], simp461_0[1:1]);
  C3 I135 (simp471_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I136 (simp471_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I137 (match1_0[14:14], simp471_0[0:0], simp471_0[1:1]);
  C3 I138 (simp481_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I139 (simp481_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I140 (match1_0[15:15], simp481_0[0:0], simp481_0[1:1]);
  C3 I141 (simp491_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I142 (simp491_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I143 (match1_0[16:16], simp491_0[0:0], simp491_0[1:1]);
  C3 I144 (simp501_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I145 (simp501_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I146 (match1_0[17:17], simp501_0[0:0], simp501_0[1:1]);
  C3 I147 (simp511_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I148 (simp511_0[1:1], i_0r1[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I149 (match1_0[18:18], simp511_0[0:0], simp511_0[1:1]);
  C3 I150 (simp521_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I151 (simp521_0[1:1], i_0r1[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I152 (match1_0[19:19], simp521_0[0:0], simp521_0[1:1]);
  C3 I153 (simp531_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I154 (simp531_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I155 (match1_0[20:20], simp531_0[0:0], simp531_0[1:1]);
  C3 I156 (simp541_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I157 (simp541_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I158 (match1_0[21:21], simp541_0[0:0], simp541_0[1:1]);
  C3 I159 (simp551_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I160 (simp551_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I161 (match1_0[22:22], simp551_0[0:0], simp551_0[1:1]);
  C2 I162 (gsel_0, sel_0, icomplete_0);
  C2 I163 (gsel_1, sel_1, icomplete_0);
  OR2 I164 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I165 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I166 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I167 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I168 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I169 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  C3 I170 (simp651_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I171 (simp651_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C2 I172 (icomplete_0, simp651_0[0:0], simp651_0[1:1]);
  BUFF I173 (o_0r, gsel_0);
  BUFF I174 (o_1r, gsel_1);
  OR2 I175 (oack_0, o_0a, o_1a);
  C2 I176 (i_0a, oack_0, icomplete_0);
endmodule

// tkm2x1b TeakM [Many [1,1],One 1]
module tkm2x1b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input i_1r0;
  input i_1r1;
  output i_1a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire gfint_0;
  wire gfint_1;
  wire gtint_0;
  wire gtint_1;
  wire choice_0;
  wire choice_1;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire nchosen_0;
  wire comp0_0;
  wire comp1_0;
  OR2 I0 (o_0r0, gfint_0, gfint_1);
  OR2 I1 (o_0r1, gtint_0, gtint_1);
  AND2 I2 (gtint_0, choice_0, i_0r1);
  AND2 I3 (gtint_1, choice_1, i_1r1);
  AND2 I4 (gfint_0, choice_0, i_0r0);
  AND2 I5 (gfint_1, choice_1, i_1r0);
  OR2 I6 (comp0_0, i_0r0, i_0r1);
  BUFF I7 (icomp_0, comp0_0);
  OR2 I8 (comp1_0, i_1r0, i_1r1);
  BUFF I9 (icomp_1, comp1_0);
  C2R I10 (choice_0, icomp_0, nchosen_0, reset);
  C2R I11 (choice_1, icomp_1, nchosen_0, reset);
  OR2 I12 (anychoice_0, choice_0, choice_1);
  NOR2 I13 (nchosen_0, anychoice_0, o_0a);
  C2R I14 (i_0a, choice_0, o_0a, reset);
  C2R I15 (i_1a, choice_1, o_0a, reset);
endmodule

// tks3_o0w3_0c4m1m2m3c4o0w0_5m6o0w0 TeakS (0+:3) [([Imp 0 4,Imp 1 0,Imp 2 0,Imp 3 4],0),([Imp 5 0,Imp 
//   6 0],0)] [One 3,Many [0,0]]
module tks3_o0w3_0c4m1m2m3c4o0w0_5m6o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire [3:0] match0_0;
  wire [1:0] simp71_0;
  wire [1:0] match1_0;
  wire [2:0] comp_0;
  NOR3 I0 (simp71_0[0:0], match0_0[0:0], match0_0[1:1], match0_0[2:2]);
  INV I1 (simp71_0[1:1], match0_0[3:3]);
  NAND2 I2 (sel_0, simp71_0[0:0], simp71_0[1:1]);
  C2 I3 (match0_0[0:0], i_0r0[0:0], i_0r0[1:1]);
  C3 I4 (match0_0[1:1], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I5 (match0_0[2:2], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C2 I6 (match0_0[3:3], i_0r1[0:0], i_0r1[1:1]);
  OR2 I7 (sel_1, match1_0[0:0], match1_0[1:1]);
  C3 I8 (match1_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I9 (match1_0[1:1], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  C2 I10 (gsel_0, sel_0, icomplete_0);
  C2 I11 (gsel_1, sel_1, icomplete_0);
  OR2 I12 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I13 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I14 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I15 (icomplete_0, comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  BUFF I16 (o_0r, gsel_0);
  BUFF I17 (o_1r, gsel_1);
  OR2 I18 (oack_0, o_0a, o_1a);
  C2 I19 (i_0a, oack_0, icomplete_0);
endmodule

// tks3_o0w3_1c6m2c4m4o0w0_0o0w0 TeakS (0+:3) [([Imp 1 6,Imp 2 4,Imp 4 0],0),([Imp 0 0],0)] [One 3,Many
//    [0,0]]
module tks3_o0w3_1c6m2c4m4o0w0_0o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire [2:0] match0_0;
  wire match1_0;
  wire [2:0] comp_0;
  OR3 I0 (sel_0, match0_0[0:0], match0_0[1:1], match0_0[2:2]);
  BUFF I1 (match0_0[0:0], i_0r1[0:0]);
  C2 I2 (match0_0[1:1], i_0r0[0:0], i_0r1[1:1]);
  C3 I3 (match0_0[2:2], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I4 (sel_1, match1_0);
  C3 I5 (match1_0, i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C2 I6 (gsel_0, sel_0, icomplete_0);
  C2 I7 (gsel_1, sel_1, icomplete_0);
  OR2 I8 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I9 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I10 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I11 (icomplete_0, comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  BUFF I12 (o_0r, gsel_0);
  BUFF I13 (o_1r, gsel_1);
  OR2 I14 (oack_0, o_0a, o_1a);
  C2 I15 (i_0a, oack_0, icomplete_0);
endmodule

// tkvstore1_wo0w1_ro0w1o0w1 TeakV "store" 1 [] [0] [0,0] [Many [1],Many [0],Many [0,0],Many [1,1]]
module tkvstore1_wo0w1_ro0w1o0w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, reset);
  input wg_0r0;
  input wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  output rd_1r0;
  output rd_1r1;
  input rd_1a;
  input reset;
  wire wf_0;
  wire wt_0;
  wire df_0;
  wire dt_0;
  wire wc_0;
  wire wacks_0;
  wire wenr_0;
  wire wen_0;
  wire anyread_0;
  wire nreset_0;
  wire drlgf_0;
  wire drlgt_0;
  wire comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire conwgit_0;
  wire conwgif_0;
  wire conwig_0;
  wire [1:0] simp401_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0, wenr_0, nreset_0);
  AND2 I2 (drlgf_0, wf_0, wen_0);
  AND2 I3 (drlgt_0, wt_0, wen_0);
  NOR2 I4 (df_0, dt_0, drlgt_0);
  NOR3 I5 (dt_0, df_0, drlgf_0, reset);
  AO22 I6 (wacks_0, drlgf_0, df_0, drlgt_0, dt_0);
  OR2 I7 (comp0_0, wg_0r0, wg_0r1);
  BUFF I8 (wc_0, comp0_0);
  AND2 I9 (conwgif_0, wg_0r0, conwig_0);
  AND2 I10 (conwgit_0, wg_0r1, conwig_0);
  BUFF I11 (conwigc_0, wc_0);
  AO22 I12 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I13 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I14 (wf_0, conwgif_0);
  BUFF I15 (wt_0, conwgit_0);
  BUFF I16 (wenr_0, wc_0);
  C2 I17 (wd_0r, conwig_0, wacks_0);
  AND2 I18 (rd_0r0, df_0, rg_0r);
  AND2 I19 (rd_1r0, df_0, rg_1r);
  AND2 I20 (rd_0r1, dt_0, rg_0r);
  AND2 I21 (rd_1r1, dt_0, rg_1r);
  NOR3 I22 (simp401_0[0:0], rg_0r, rg_1r, rg_0a);
  INV I23 (simp401_0[1:1], rg_1a);
  NAND2 I24 (anyread_0, simp401_0[0:0], simp401_0[1:1]);
  BUFF I25 (wg_0a, wd_0a);
  BUFF I26 (rg_0a, rd_0a);
  BUFF I27 (rg_1a, rd_1a);
endmodule

// tkvmemAccess4_wo0w4_ro0w4 TeakV "memAccess" 4 [] [0] [0] [Many [4],Many [0],Many [0],Many [4]]
module tkvmemAccess4_wo0w4_ro0w4 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [3:0] wg_0r0;
  input [3:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [3:0] rd_0r0;
  output [3:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [3:0] wf_0;
  wire [3:0] wt_0;
  wire [3:0] df_0;
  wire [3:0] dt_0;
  wire wc_0;
  wire [3:0] wacks_0;
  wire [3:0] wenr_0;
  wire [3:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [3:0] drlgf_0;
  wire [3:0] drlgt_0;
  wire [3:0] comp0_0;
  wire [1:0] simp421_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [3:0] conwgit_0;
  wire [3:0] conwgif_0;
  wire conwig_0;
  wire [1:0] simp711_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I6 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I7 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I8 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I9 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I10 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I11 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I12 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  NOR2 I13 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I14 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I15 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I16 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR3 I17 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I18 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I19 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I20 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  AO22 I21 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I22 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I23 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I24 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  OR2 I25 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I26 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I27 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I28 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  C3 I29 (simp421_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  BUFF I30 (simp421_0[1:1], comp0_0[3:3]);
  C2 I31 (wc_0, simp421_0[0:0], simp421_0[1:1]);
  AND2 I32 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I33 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I34 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I35 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I36 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I37 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I38 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I39 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  BUFF I40 (conwigc_0, wc_0);
  AO22 I41 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I42 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I43 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I44 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I45 (wenr_0[0:0], wc_0);
  BUFF I46 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I47 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I48 (wenr_0[1:1], wc_0);
  BUFF I49 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I50 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I51 (wenr_0[2:2], wc_0);
  BUFF I52 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I53 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I54 (wenr_0[3:3], wc_0);
  C3 I55 (simp711_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C2 I56 (simp711_0[1:1], wacks_0[2:2], wacks_0[3:3]);
  C2 I57 (wd_0r, simp711_0[0:0], simp711_0[1:1]);
  AND2 I58 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I59 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I60 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I61 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I62 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I63 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I64 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I65 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  OR2 I66 (anyread_0, rg_0r, rg_0a);
  BUFF I67 (wg_0a, wd_0a);
  BUFF I68 (rg_0a, rd_0a);
endmodule

// tkvinstKind3_wo0w3_ro0w3o0w3o0w3 TeakV "instKind" 3 [] [0] [0,0,0] [Many [3],Many [0],Many [0,0,0],M
//   any [3,3,3]]
module tkvinstKind3_wo0w3_ro0w3o0w3o0w3 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [2:0] wg_0r0;
  input [2:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [2:0] rd_0r0;
  output [2:0] rd_0r1;
  input rd_0a;
  output [2:0] rd_1r0;
  output [2:0] rd_1r1;
  input rd_1a;
  output [2:0] rd_2r0;
  output [2:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [2:0] wf_0;
  wire [2:0] wt_0;
  wire [2:0] df_0;
  wire [2:0] dt_0;
  wire wc_0;
  wire [2:0] wacks_0;
  wire [2:0] wenr_0;
  wire [2:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [2:0] drlgf_0;
  wire [2:0] drlgt_0;
  wire [2:0] comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [2:0] conwgit_0;
  wire [2:0] conwgif_0;
  wire conwig_0;
  wire [1:0] simp591_0;
  wire [1:0] simp781_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I5 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I6 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I7 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I8 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I9 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  NOR2 I10 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I11 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I12 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR3 I13 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I14 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I15 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  AO22 I16 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I17 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I18 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  OR2 I19 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I20 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I21 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  C3 I22 (wc_0, comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  AND2 I23 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I24 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I25 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I26 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I27 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I28 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  BUFF I29 (conwigc_0, wc_0);
  AO22 I30 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I31 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I32 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I33 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I34 (wenr_0[0:0], wc_0);
  BUFF I35 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I36 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I37 (wenr_0[1:1], wc_0);
  BUFF I38 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I39 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I40 (wenr_0[2:2], wc_0);
  C3 I41 (simp591_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  BUFF I42 (simp591_0[1:1], wacks_0[2:2]);
  C2 I43 (wd_0r, simp591_0[0:0], simp591_0[1:1]);
  AND2 I44 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I45 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I46 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I47 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I48 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I49 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I50 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I51 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I52 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I53 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I54 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I55 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I56 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I57 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I58 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I59 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I60 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I61 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  NOR3 I62 (simp781_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I63 (simp781_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I64 (anyread_0, simp781_0[0:0], simp781_0[1:1]);
  BUFF I65 (wg_0a, wd_0a);
  BUFF I66 (rg_0a, rd_0a);
  BUFF I67 (rg_1a, rd_1a);
  BUFF I68 (rg_2a, rd_2a);
endmodule

// tko0m3_1nm3b0 TeakO [
//     (1,TeakOConstant 3 0)] [One 0,One 3]
module tko0m3_1nm3b0 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r);
  BUFF I1 (o_0r0[1:1], i_0r);
  BUFF I2 (o_0r0[2:2], i_0r);
  GND I3 (o_0r1[0:0]);
  GND I4 (o_0r1[1:1]);
  GND I5 (o_0r1[2:2]);
  BUFF I6 (i_0a, o_0a);
endmodule

// tko0m3_1nm3b3 TeakO [
//     (1,TeakOConstant 3 3)] [One 0,One 3]
module tko0m3_1nm3b3 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  BUFF I1 (o_0r1[1:1], i_0r);
  GND I2 (o_0r0[0:0]);
  GND I3 (o_0r0[1:1]);
  BUFF I4 (o_0r0[2:2], i_0r);
  GND I5 (o_0r1[2:2]);
  BUFF I6 (i_0a, o_0a);
endmodule

// tko0m4_1nm4b3 TeakO [
//     (1,TeakOConstant 4 3)] [One 0,One 4]
module tko0m4_1nm4b3 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  BUFF I1 (o_0r1[1:1], i_0r);
  GND I2 (o_0r0[0:0]);
  GND I3 (o_0r0[1:1]);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  GND I6 (o_0r1[2:2]);
  GND I7 (o_0r1[3:3]);
  BUFF I8 (i_0a, o_0a);
endmodule

// tko0m4_1nm4b5 TeakO [
//     (1,TeakOConstant 4 5)] [One 0,One 4]
module tko0m4_1nm4b5 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  BUFF I1 (o_0r1[2:2], i_0r);
  GND I2 (o_0r0[0:0]);
  GND I3 (o_0r0[2:2]);
  BUFF I4 (o_0r0[1:1], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  GND I6 (o_0r1[1:1]);
  GND I7 (o_0r1[3:3]);
  BUFF I8 (i_0a, o_0a);
endmodule

// tko0m4_1nm4b6 TeakO [
//     (1,TeakOConstant 4 6)] [One 0,One 4]
module tko0m4_1nm4b6 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[1:1], i_0r);
  BUFF I1 (o_0r1[2:2], i_0r);
  GND I2 (o_0r0[1:1]);
  GND I3 (o_0r0[2:2]);
  BUFF I4 (o_0r0[0:0], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  GND I6 (o_0r1[0:0]);
  GND I7 (o_0r1[3:3]);
  BUFF I8 (i_0a, o_0a);
endmodule

// tko0m3_1nm3b5 TeakO [
//     (1,TeakOConstant 3 5)] [One 0,One 3]
module tko0m3_1nm3b5 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  BUFF I1 (o_0r1[2:2], i_0r);
  GND I2 (o_0r0[0:0]);
  GND I3 (o_0r0[2:2]);
  BUFF I4 (o_0r0[1:1], i_0r);
  GND I5 (o_0r1[1:1]);
  BUFF I6 (i_0a, o_0a);
endmodule

// tko0m4_1nm4b2 TeakO [
//     (1,TeakOConstant 4 2)] [One 0,One 4]
module tko0m4_1nm4b2 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[1:1], i_0r);
  GND I1 (o_0r0[1:1]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  GND I5 (o_0r1[0:0]);
  GND I6 (o_0r1[2:2]);
  GND I7 (o_0r1[3:3]);
  BUFF I8 (i_0a, o_0a);
endmodule

// tko0m4_1nm4b4 TeakO [
//     (1,TeakOConstant 4 4)] [One 0,One 4]
module tko0m4_1nm4b4 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[2:2], i_0r);
  GND I1 (o_0r0[2:2]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  GND I5 (o_0r1[0:0]);
  GND I6 (o_0r1[1:1]);
  GND I7 (o_0r1[3:3]);
  BUFF I8 (i_0a, o_0a);
endmodule

// tko0m4_1nm4bb TeakO [
//     (1,TeakOConstant 4 11)] [One 0,One 4]
module tko0m4_1nm4bb (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  BUFF I1 (o_0r1[1:1], i_0r);
  BUFF I2 (o_0r1[3:3], i_0r);
  GND I3 (o_0r0[0:0]);
  GND I4 (o_0r0[1:1]);
  GND I5 (o_0r0[3:3]);
  BUFF I6 (o_0r0[2:2], i_0r);
  GND I7 (o_0r1[2:2]);
  BUFF I8 (i_0a, o_0a);
endmodule

// tko0m4_1nm4bd TeakO [
//     (1,TeakOConstant 4 13)] [One 0,One 4]
module tko0m4_1nm4bd (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  BUFF I1 (o_0r1[2:2], i_0r);
  BUFF I2 (o_0r1[3:3], i_0r);
  GND I3 (o_0r0[0:0]);
  GND I4 (o_0r0[2:2]);
  GND I5 (o_0r0[3:3]);
  BUFF I6 (o_0r0[1:1], i_0r);
  GND I7 (o_0r1[1:1]);
  BUFF I8 (i_0a, o_0a);
endmodule

// tks6_o0w6_8c30mbc30mcc30mdc30mec30mfc30m10c20m11c20m12c20m13c20m14c20m15c20m16c20m17c20m19c20m1ac20m
//   20m21m22m23m24m25m26m27m29m2ao0w0_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0_9o0w0_ao0w0 TeakS 
//   (0+:6) [([Imp 8 48,Imp 11 48,Imp 12 48,Imp 13 48,Imp 14 48,Imp 15 48,Imp 16 32,Imp 17 32,Imp 18 32,I
//   mp 19 32,Imp 20 32,Imp 21 32,Imp 22 32,Imp 23 32,Imp 25 32,Imp 26 32,Imp 32 0,Imp 33 0,Imp 34 0,Imp 
//   35 0,Imp 36 0,Imp 37 0,Imp 38 0,Imp 39 0,Imp 41 0,Imp 42 0],0),([Imp 0 0],0),([Imp 1 0],0),([Imp 2 0
//   ],0),([Imp 3 0],0),([Imp 4 0],0),([Imp 5 0],0),([Imp 6 0],0),([Imp 7 0],0),([Imp 9 0],0),([Imp 10 0]
//   ,0)] [One 6,Many [0,0,0,0,0,0,0,0,0,0,0]]
module tks6_o0w6_8c30mbc30mcc30mdc30mec30mfc30m10c20m11c20m12c20m13c20m14c20m15c20m16c20m17c20m19c20m1ac20m20m21m22m23m24m25m26m27m29m2ao0w0_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0_9o0w0_ao0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, o_5r, o_5a, o_6r, o_6a, o_7r, o_7a, o_8r, o_8a, o_9r, o_9a, o_10r, o_10a, reset);
  input [5:0] i_0r0;
  input [5:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  output o_7r;
  input o_7a;
  output o_8r;
  input o_8a;
  output o_9r;
  input o_9a;
  output o_10r;
  input o_10a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire sel_4;
  wire sel_5;
  wire sel_6;
  wire sel_7;
  wire sel_8;
  wire sel_9;
  wire sel_10;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire gsel_4;
  wire gsel_5;
  wire gsel_6;
  wire gsel_7;
  wire gsel_8;
  wire gsel_9;
  wire gsel_10;
  wire oack_0;
  wire [25:0] match0_0;
  wire [8:0] simp251_0;
  wire [2:0] simp252_0;
  wire [1:0] simp261_0;
  wire [1:0] simp271_0;
  wire [1:0] simp281_0;
  wire [1:0] simp291_0;
  wire [1:0] simp301_0;
  wire [1:0] simp311_0;
  wire [1:0] simp321_0;
  wire [1:0] simp331_0;
  wire [1:0] simp341_0;
  wire [1:0] simp351_0;
  wire [1:0] simp361_0;
  wire [1:0] simp371_0;
  wire [1:0] simp381_0;
  wire [1:0] simp391_0;
  wire [1:0] simp401_0;
  wire [1:0] simp411_0;
  wire [1:0] simp421_0;
  wire [1:0] simp431_0;
  wire [1:0] simp441_0;
  wire [1:0] simp451_0;
  wire [1:0] simp461_0;
  wire [1:0] simp471_0;
  wire [1:0] simp481_0;
  wire [1:0] simp491_0;
  wire [1:0] simp501_0;
  wire [1:0] simp511_0;
  wire match1_0;
  wire [1:0] simp541_0;
  wire match2_0;
  wire [1:0] simp571_0;
  wire match3_0;
  wire [1:0] simp601_0;
  wire match4_0;
  wire [1:0] simp631_0;
  wire match5_0;
  wire [1:0] simp661_0;
  wire match6_0;
  wire [1:0] simp691_0;
  wire match7_0;
  wire [1:0] simp721_0;
  wire match8_0;
  wire [1:0] simp751_0;
  wire match9_0;
  wire [1:0] simp781_0;
  wire match10_0;
  wire [1:0] simp811_0;
  wire [5:0] comp_0;
  wire [1:0] simp1001_0;
  wire [3:0] simp1121_0;
  wire [1:0] simp1122_0;
  NOR3 I0 (simp251_0[0:0], match0_0[0:0], match0_0[1:1], match0_0[2:2]);
  NOR3 I1 (simp251_0[1:1], match0_0[3:3], match0_0[4:4], match0_0[5:5]);
  NOR3 I2 (simp251_0[2:2], match0_0[6:6], match0_0[7:7], match0_0[8:8]);
  NOR3 I3 (simp251_0[3:3], match0_0[9:9], match0_0[10:10], match0_0[11:11]);
  NOR3 I4 (simp251_0[4:4], match0_0[12:12], match0_0[13:13], match0_0[14:14]);
  NOR3 I5 (simp251_0[5:5], match0_0[15:15], match0_0[16:16], match0_0[17:17]);
  NOR3 I6 (simp251_0[6:6], match0_0[18:18], match0_0[19:19], match0_0[20:20]);
  NOR3 I7 (simp251_0[7:7], match0_0[21:21], match0_0[22:22], match0_0[23:23]);
  NOR2 I8 (simp251_0[8:8], match0_0[24:24], match0_0[25:25]);
  NAND3 I9 (simp252_0[0:0], simp251_0[0:0], simp251_0[1:1], simp251_0[2:2]);
  NAND3 I10 (simp252_0[1:1], simp251_0[3:3], simp251_0[4:4], simp251_0[5:5]);
  NAND3 I11 (simp252_0[2:2], simp251_0[6:6], simp251_0[7:7], simp251_0[8:8]);
  OR3 I12 (sel_0, simp252_0[0:0], simp252_0[1:1], simp252_0[2:2]);
  C3 I13 (simp261_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I14 (simp261_0[1:1], i_0r1[3:3]);
  C2 I15 (match0_0[0:0], simp261_0[0:0], simp261_0[1:1]);
  C3 I16 (simp271_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I17 (simp271_0[1:1], i_0r1[3:3]);
  C2 I18 (match0_0[1:1], simp271_0[0:0], simp271_0[1:1]);
  C3 I19 (simp281_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I20 (simp281_0[1:1], i_0r1[3:3]);
  C2 I21 (match0_0[2:2], simp281_0[0:0], simp281_0[1:1]);
  C3 I22 (simp291_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I23 (simp291_0[1:1], i_0r1[3:3]);
  C2 I24 (match0_0[3:3], simp291_0[0:0], simp291_0[1:1]);
  C3 I25 (simp301_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I26 (simp301_0[1:1], i_0r1[3:3]);
  C2 I27 (match0_0[4:4], simp301_0[0:0], simp301_0[1:1]);
  C3 I28 (simp311_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I29 (simp311_0[1:1], i_0r1[3:3]);
  C2 I30 (match0_0[5:5], simp311_0[0:0], simp311_0[1:1]);
  C3 I31 (simp321_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C2 I32 (simp321_0[1:1], i_0r0[3:3], i_0r1[4:4]);
  C2 I33 (match0_0[6:6], simp321_0[0:0], simp321_0[1:1]);
  C3 I34 (simp331_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C2 I35 (simp331_0[1:1], i_0r0[3:3], i_0r1[4:4]);
  C2 I36 (match0_0[7:7], simp331_0[0:0], simp331_0[1:1]);
  C3 I37 (simp341_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C2 I38 (simp341_0[1:1], i_0r0[3:3], i_0r1[4:4]);
  C2 I39 (match0_0[8:8], simp341_0[0:0], simp341_0[1:1]);
  C3 I40 (simp351_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  C2 I41 (simp351_0[1:1], i_0r0[3:3], i_0r1[4:4]);
  C2 I42 (match0_0[9:9], simp351_0[0:0], simp351_0[1:1]);
  C3 I43 (simp361_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C2 I44 (simp361_0[1:1], i_0r0[3:3], i_0r1[4:4]);
  C2 I45 (match0_0[10:10], simp361_0[0:0], simp361_0[1:1]);
  C3 I46 (simp371_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  C2 I47 (simp371_0[1:1], i_0r0[3:3], i_0r1[4:4]);
  C2 I48 (match0_0[11:11], simp371_0[0:0], simp371_0[1:1]);
  C3 I49 (simp381_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  C2 I50 (simp381_0[1:1], i_0r0[3:3], i_0r1[4:4]);
  C2 I51 (match0_0[12:12], simp381_0[0:0], simp381_0[1:1]);
  C3 I52 (simp391_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  C2 I53 (simp391_0[1:1], i_0r0[3:3], i_0r1[4:4]);
  C2 I54 (match0_0[13:13], simp391_0[0:0], simp391_0[1:1]);
  C3 I55 (simp401_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C2 I56 (simp401_0[1:1], i_0r1[3:3], i_0r1[4:4]);
  C2 I57 (match0_0[14:14], simp401_0[0:0], simp401_0[1:1]);
  C3 I58 (simp411_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C2 I59 (simp411_0[1:1], i_0r1[3:3], i_0r1[4:4]);
  C2 I60 (match0_0[15:15], simp411_0[0:0], simp411_0[1:1]);
  C3 I61 (simp421_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I62 (simp421_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I63 (match0_0[16:16], simp421_0[0:0], simp421_0[1:1]);
  C3 I64 (simp431_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I65 (simp431_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I66 (match0_0[17:17], simp431_0[0:0], simp431_0[1:1]);
  C3 I67 (simp441_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I68 (simp441_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I69 (match0_0[18:18], simp441_0[0:0], simp441_0[1:1]);
  C3 I70 (simp451_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I71 (simp451_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I72 (match0_0[19:19], simp451_0[0:0], simp451_0[1:1]);
  C3 I73 (simp461_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I74 (simp461_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I75 (match0_0[20:20], simp461_0[0:0], simp461_0[1:1]);
  C3 I76 (simp471_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I77 (simp471_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I78 (match0_0[21:21], simp471_0[0:0], simp471_0[1:1]);
  C3 I79 (simp481_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I80 (simp481_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I81 (match0_0[22:22], simp481_0[0:0], simp481_0[1:1]);
  C3 I82 (simp491_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I83 (simp491_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I84 (match0_0[23:23], simp491_0[0:0], simp491_0[1:1]);
  C3 I85 (simp501_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I86 (simp501_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I87 (match0_0[24:24], simp501_0[0:0], simp501_0[1:1]);
  C3 I88 (simp511_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I89 (simp511_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I90 (match0_0[25:25], simp511_0[0:0], simp511_0[1:1]);
  BUFF I91 (sel_1, match1_0);
  C3 I92 (simp541_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I93 (simp541_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I94 (match1_0, simp541_0[0:0], simp541_0[1:1]);
  BUFF I95 (sel_2, match2_0);
  C3 I96 (simp571_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I97 (simp571_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I98 (match2_0, simp571_0[0:0], simp571_0[1:1]);
  BUFF I99 (sel_3, match3_0);
  C3 I100 (simp601_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I101 (simp601_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I102 (match3_0, simp601_0[0:0], simp601_0[1:1]);
  BUFF I103 (sel_4, match4_0);
  C3 I104 (simp631_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I105 (simp631_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I106 (match4_0, simp631_0[0:0], simp631_0[1:1]);
  BUFF I107 (sel_5, match5_0);
  C3 I108 (simp661_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I109 (simp661_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I110 (match5_0, simp661_0[0:0], simp661_0[1:1]);
  BUFF I111 (sel_6, match6_0);
  C3 I112 (simp691_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I113 (simp691_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I114 (match6_0, simp691_0[0:0], simp691_0[1:1]);
  BUFF I115 (sel_7, match7_0);
  C3 I116 (simp721_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I117 (simp721_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I118 (match7_0, simp721_0[0:0], simp721_0[1:1]);
  BUFF I119 (sel_8, match8_0);
  C3 I120 (simp751_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I121 (simp751_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I122 (match8_0, simp751_0[0:0], simp751_0[1:1]);
  BUFF I123 (sel_9, match9_0);
  C3 I124 (simp781_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I125 (simp781_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I126 (match9_0, simp781_0[0:0], simp781_0[1:1]);
  BUFF I127 (sel_10, match10_0);
  C3 I128 (simp811_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I129 (simp811_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I130 (match10_0, simp811_0[0:0], simp811_0[1:1]);
  C2 I131 (gsel_0, sel_0, icomplete_0);
  C2 I132 (gsel_1, sel_1, icomplete_0);
  C2 I133 (gsel_2, sel_2, icomplete_0);
  C2 I134 (gsel_3, sel_3, icomplete_0);
  C2 I135 (gsel_4, sel_4, icomplete_0);
  C2 I136 (gsel_5, sel_5, icomplete_0);
  C2 I137 (gsel_6, sel_6, icomplete_0);
  C2 I138 (gsel_7, sel_7, icomplete_0);
  C2 I139 (gsel_8, sel_8, icomplete_0);
  C2 I140 (gsel_9, sel_9, icomplete_0);
  C2 I141 (gsel_10, sel_10, icomplete_0);
  OR2 I142 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I143 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I144 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I145 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I146 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I147 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  C3 I148 (simp1001_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I149 (simp1001_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C2 I150 (icomplete_0, simp1001_0[0:0], simp1001_0[1:1]);
  BUFF I151 (o_0r, gsel_0);
  BUFF I152 (o_1r, gsel_1);
  BUFF I153 (o_2r, gsel_2);
  BUFF I154 (o_3r, gsel_3);
  BUFF I155 (o_4r, gsel_4);
  BUFF I156 (o_5r, gsel_5);
  BUFF I157 (o_6r, gsel_6);
  BUFF I158 (o_7r, gsel_7);
  BUFF I159 (o_8r, gsel_8);
  BUFF I160 (o_9r, gsel_9);
  BUFF I161 (o_10r, gsel_10);
  NOR3 I162 (simp1121_0[0:0], o_0a, o_1a, o_2a);
  NOR3 I163 (simp1121_0[1:1], o_3a, o_4a, o_5a);
  NOR3 I164 (simp1121_0[2:2], o_6a, o_7a, o_8a);
  NOR2 I165 (simp1121_0[3:3], o_9a, o_10a);
  NAND3 I166 (simp1122_0[0:0], simp1121_0[0:0], simp1121_0[1:1], simp1121_0[2:2]);
  INV I167 (simp1122_0[1:1], simp1121_0[3:3]);
  OR2 I168 (oack_0, simp1122_0[0:0], simp1122_0[1:1]);
  C2 I169 (i_0a, oack_0, icomplete_0);
endmodule

// tkm11x0b TeakM [Many [0,0,0,0,0,0,0,0,0,0,0],One 0]
module tkm11x0b (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, i_3r, i_3a, i_4r, i_4a, i_5r, i_5a, i_6r, i_6a, i_7r, i_7a, i_8r, i_8a, i_9r, i_9a, i_10r, i_10a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  input i_4r;
  output i_4a;
  input i_5r;
  output i_5a;
  input i_6r;
  output i_6a;
  input i_7r;
  output i_7a;
  input i_8r;
  output i_8a;
  input i_9r;
  output i_9a;
  input i_10r;
  output i_10a;
  output o_0r;
  input o_0a;
  input reset;
  wire nchosen_0;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire choice_4;
  wire choice_5;
  wire choice_6;
  wire choice_7;
  wire choice_8;
  wire choice_9;
  wire choice_10;
  wire [3:0] simp241_0;
  wire [1:0] simp242_0;
  C2R I0 (choice_0, i_0r, nchosen_0, reset);
  C2R I1 (choice_1, i_1r, nchosen_0, reset);
  C2R I2 (choice_2, i_2r, nchosen_0, reset);
  C2R I3 (choice_3, i_3r, nchosen_0, reset);
  C2R I4 (choice_4, i_4r, nchosen_0, reset);
  C2R I5 (choice_5, i_5r, nchosen_0, reset);
  C2R I6 (choice_6, i_6r, nchosen_0, reset);
  C2R I7 (choice_7, i_7r, nchosen_0, reset);
  C2R I8 (choice_8, i_8r, nchosen_0, reset);
  C2R I9 (choice_9, i_9r, nchosen_0, reset);
  C2R I10 (choice_10, i_10r, nchosen_0, reset);
  NOR2 I11 (nchosen_0, o_0r, o_0a);
  NOR3 I12 (simp241_0[0:0], choice_0, choice_1, choice_2);
  NOR3 I13 (simp241_0[1:1], choice_3, choice_4, choice_5);
  NOR3 I14 (simp241_0[2:2], choice_6, choice_7, choice_8);
  NOR2 I15 (simp241_0[3:3], choice_9, choice_10);
  NAND3 I16 (simp242_0[0:0], simp241_0[0:0], simp241_0[1:1], simp241_0[2:2]);
  INV I17 (simp242_0[1:1], simp241_0[3:3]);
  OR2 I18 (o_0r, simp242_0[0:0], simp242_0[1:1]);
  C2R I19 (i_0a, choice_0, o_0a, reset);
  C2R I20 (i_1a, choice_1, o_0a, reset);
  C2R I21 (i_2a, choice_2, o_0a, reset);
  C2R I22 (i_3a, choice_3, o_0a, reset);
  C2R I23 (i_4a, choice_4, o_0a, reset);
  C2R I24 (i_5a, choice_5, o_0a, reset);
  C2R I25 (i_6a, choice_6, o_0a, reset);
  C2R I26 (i_7a, choice_7, o_0a, reset);
  C2R I27 (i_8a, choice_8, o_0a, reset);
  C2R I28 (i_9a, choice_9, o_0a, reset);
  C2R I29 (i_10a, choice_10, o_0a, reset);
endmodule

// tkf3mo0w0_o0w3 TeakF [0,0] [One 3,Many [0,3]]
module tkf3mo0w0_o0w3 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [2:0] o_1r0;
  output [2:0] o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_1r0[0:0], i_0r0[0:0]);
  BUFF I3 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I4 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I5 (o_1r1[0:0], i_0r1[0:0]);
  BUFF I6 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I7 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I8 (o_0r, icomplete_0);
  C3 I9 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tkm11x3b TeakM [Many [3,3,3,3,3,3,3,3,3,3,3],One 3]
module tkm11x3b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, i_4r0, i_4r1, i_4a, i_5r0, i_5r1, i_5a, i_6r0, i_6r1, i_6a, i_7r0, i_7r1, i_7a, i_8r0, i_8r1, i_8a, i_9r0, i_9r1, i_9a, i_10r0, i_10r1, i_10a, o_0r0, o_0r1, o_0a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  input [2:0] i_1r0;
  input [2:0] i_1r1;
  output i_1a;
  input [2:0] i_2r0;
  input [2:0] i_2r1;
  output i_2a;
  input [2:0] i_3r0;
  input [2:0] i_3r1;
  output i_3a;
  input [2:0] i_4r0;
  input [2:0] i_4r1;
  output i_4a;
  input [2:0] i_5r0;
  input [2:0] i_5r1;
  output i_5a;
  input [2:0] i_6r0;
  input [2:0] i_6r1;
  output i_6a;
  input [2:0] i_7r0;
  input [2:0] i_7r1;
  output i_7a;
  input [2:0] i_8r0;
  input [2:0] i_8r1;
  output i_8a;
  input [2:0] i_9r0;
  input [2:0] i_9r1;
  output i_9a;
  input [2:0] i_10r0;
  input [2:0] i_10r1;
  output i_10a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire [2:0] gfint_0;
  wire [2:0] gfint_1;
  wire [2:0] gfint_2;
  wire [2:0] gfint_3;
  wire [2:0] gfint_4;
  wire [2:0] gfint_5;
  wire [2:0] gfint_6;
  wire [2:0] gfint_7;
  wire [2:0] gfint_8;
  wire [2:0] gfint_9;
  wire [2:0] gfint_10;
  wire [2:0] gtint_0;
  wire [2:0] gtint_1;
  wire [2:0] gtint_2;
  wire [2:0] gtint_3;
  wire [2:0] gtint_4;
  wire [2:0] gtint_5;
  wire [2:0] gtint_6;
  wire [2:0] gtint_7;
  wire [2:0] gtint_8;
  wire [2:0] gtint_9;
  wire [2:0] gtint_10;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire choice_4;
  wire choice_5;
  wire choice_6;
  wire choice_7;
  wire choice_8;
  wire choice_9;
  wire choice_10;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire icomp_3;
  wire icomp_4;
  wire icomp_5;
  wire icomp_6;
  wire icomp_7;
  wire icomp_8;
  wire icomp_9;
  wire icomp_10;
  wire nchosen_0;
  wire [3:0] simp461_0;
  wire [1:0] simp462_0;
  wire [3:0] simp471_0;
  wire [1:0] simp472_0;
  wire [3:0] simp481_0;
  wire [1:0] simp482_0;
  wire [3:0] simp491_0;
  wire [1:0] simp492_0;
  wire [3:0] simp501_0;
  wire [1:0] simp502_0;
  wire [3:0] simp511_0;
  wire [1:0] simp512_0;
  wire [2:0] comp0_0;
  wire [2:0] comp1_0;
  wire [2:0] comp2_0;
  wire [2:0] comp3_0;
  wire [2:0] comp4_0;
  wire [2:0] comp5_0;
  wire [2:0] comp6_0;
  wire [2:0] comp7_0;
  wire [2:0] comp8_0;
  wire [2:0] comp9_0;
  wire [2:0] comp10_0;
  wire [3:0] simp1841_0;
  wire [1:0] simp1842_0;
  NOR3 I0 (simp461_0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  NOR3 I1 (simp461_0[1:1], gfint_3[0:0], gfint_4[0:0], gfint_5[0:0]);
  NOR3 I2 (simp461_0[2:2], gfint_6[0:0], gfint_7[0:0], gfint_8[0:0]);
  NOR2 I3 (simp461_0[3:3], gfint_9[0:0], gfint_10[0:0]);
  NAND3 I4 (simp462_0[0:0], simp461_0[0:0], simp461_0[1:1], simp461_0[2:2]);
  INV I5 (simp462_0[1:1], simp461_0[3:3]);
  OR2 I6 (o_0r0[0:0], simp462_0[0:0], simp462_0[1:1]);
  NOR3 I7 (simp471_0[0:0], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  NOR3 I8 (simp471_0[1:1], gfint_3[1:1], gfint_4[1:1], gfint_5[1:1]);
  NOR3 I9 (simp471_0[2:2], gfint_6[1:1], gfint_7[1:1], gfint_8[1:1]);
  NOR2 I10 (simp471_0[3:3], gfint_9[1:1], gfint_10[1:1]);
  NAND3 I11 (simp472_0[0:0], simp471_0[0:0], simp471_0[1:1], simp471_0[2:2]);
  INV I12 (simp472_0[1:1], simp471_0[3:3]);
  OR2 I13 (o_0r0[1:1], simp472_0[0:0], simp472_0[1:1]);
  NOR3 I14 (simp481_0[0:0], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  NOR3 I15 (simp481_0[1:1], gfint_3[2:2], gfint_4[2:2], gfint_5[2:2]);
  NOR3 I16 (simp481_0[2:2], gfint_6[2:2], gfint_7[2:2], gfint_8[2:2]);
  NOR2 I17 (simp481_0[3:3], gfint_9[2:2], gfint_10[2:2]);
  NAND3 I18 (simp482_0[0:0], simp481_0[0:0], simp481_0[1:1], simp481_0[2:2]);
  INV I19 (simp482_0[1:1], simp481_0[3:3]);
  OR2 I20 (o_0r0[2:2], simp482_0[0:0], simp482_0[1:1]);
  NOR3 I21 (simp491_0[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  NOR3 I22 (simp491_0[1:1], gtint_3[0:0], gtint_4[0:0], gtint_5[0:0]);
  NOR3 I23 (simp491_0[2:2], gtint_6[0:0], gtint_7[0:0], gtint_8[0:0]);
  NOR2 I24 (simp491_0[3:3], gtint_9[0:0], gtint_10[0:0]);
  NAND3 I25 (simp492_0[0:0], simp491_0[0:0], simp491_0[1:1], simp491_0[2:2]);
  INV I26 (simp492_0[1:1], simp491_0[3:3]);
  OR2 I27 (o_0r1[0:0], simp492_0[0:0], simp492_0[1:1]);
  NOR3 I28 (simp501_0[0:0], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  NOR3 I29 (simp501_0[1:1], gtint_3[1:1], gtint_4[1:1], gtint_5[1:1]);
  NOR3 I30 (simp501_0[2:2], gtint_6[1:1], gtint_7[1:1], gtint_8[1:1]);
  NOR2 I31 (simp501_0[3:3], gtint_9[1:1], gtint_10[1:1]);
  NAND3 I32 (simp502_0[0:0], simp501_0[0:0], simp501_0[1:1], simp501_0[2:2]);
  INV I33 (simp502_0[1:1], simp501_0[3:3]);
  OR2 I34 (o_0r1[1:1], simp502_0[0:0], simp502_0[1:1]);
  NOR3 I35 (simp511_0[0:0], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  NOR3 I36 (simp511_0[1:1], gtint_3[2:2], gtint_4[2:2], gtint_5[2:2]);
  NOR3 I37 (simp511_0[2:2], gtint_6[2:2], gtint_7[2:2], gtint_8[2:2]);
  NOR2 I38 (simp511_0[3:3], gtint_9[2:2], gtint_10[2:2]);
  NAND3 I39 (simp512_0[0:0], simp511_0[0:0], simp511_0[1:1], simp511_0[2:2]);
  INV I40 (simp512_0[1:1], simp511_0[3:3]);
  OR2 I41 (o_0r1[2:2], simp512_0[0:0], simp512_0[1:1]);
  AND2 I42 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I43 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I44 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I45 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I46 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I47 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I48 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I49 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I50 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I51 (gtint_3[0:0], choice_3, i_3r1[0:0]);
  AND2 I52 (gtint_3[1:1], choice_3, i_3r1[1:1]);
  AND2 I53 (gtint_3[2:2], choice_3, i_3r1[2:2]);
  AND2 I54 (gtint_4[0:0], choice_4, i_4r1[0:0]);
  AND2 I55 (gtint_4[1:1], choice_4, i_4r1[1:1]);
  AND2 I56 (gtint_4[2:2], choice_4, i_4r1[2:2]);
  AND2 I57 (gtint_5[0:0], choice_5, i_5r1[0:0]);
  AND2 I58 (gtint_5[1:1], choice_5, i_5r1[1:1]);
  AND2 I59 (gtint_5[2:2], choice_5, i_5r1[2:2]);
  AND2 I60 (gtint_6[0:0], choice_6, i_6r1[0:0]);
  AND2 I61 (gtint_6[1:1], choice_6, i_6r1[1:1]);
  AND2 I62 (gtint_6[2:2], choice_6, i_6r1[2:2]);
  AND2 I63 (gtint_7[0:0], choice_7, i_7r1[0:0]);
  AND2 I64 (gtint_7[1:1], choice_7, i_7r1[1:1]);
  AND2 I65 (gtint_7[2:2], choice_7, i_7r1[2:2]);
  AND2 I66 (gtint_8[0:0], choice_8, i_8r1[0:0]);
  AND2 I67 (gtint_8[1:1], choice_8, i_8r1[1:1]);
  AND2 I68 (gtint_8[2:2], choice_8, i_8r1[2:2]);
  AND2 I69 (gtint_9[0:0], choice_9, i_9r1[0:0]);
  AND2 I70 (gtint_9[1:1], choice_9, i_9r1[1:1]);
  AND2 I71 (gtint_9[2:2], choice_9, i_9r1[2:2]);
  AND2 I72 (gtint_10[0:0], choice_10, i_10r1[0:0]);
  AND2 I73 (gtint_10[1:1], choice_10, i_10r1[1:1]);
  AND2 I74 (gtint_10[2:2], choice_10, i_10r1[2:2]);
  AND2 I75 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I76 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I77 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I78 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I79 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I80 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I81 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I82 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I83 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I84 (gfint_3[0:0], choice_3, i_3r0[0:0]);
  AND2 I85 (gfint_3[1:1], choice_3, i_3r0[1:1]);
  AND2 I86 (gfint_3[2:2], choice_3, i_3r0[2:2]);
  AND2 I87 (gfint_4[0:0], choice_4, i_4r0[0:0]);
  AND2 I88 (gfint_4[1:1], choice_4, i_4r0[1:1]);
  AND2 I89 (gfint_4[2:2], choice_4, i_4r0[2:2]);
  AND2 I90 (gfint_5[0:0], choice_5, i_5r0[0:0]);
  AND2 I91 (gfint_5[1:1], choice_5, i_5r0[1:1]);
  AND2 I92 (gfint_5[2:2], choice_5, i_5r0[2:2]);
  AND2 I93 (gfint_6[0:0], choice_6, i_6r0[0:0]);
  AND2 I94 (gfint_6[1:1], choice_6, i_6r0[1:1]);
  AND2 I95 (gfint_6[2:2], choice_6, i_6r0[2:2]);
  AND2 I96 (gfint_7[0:0], choice_7, i_7r0[0:0]);
  AND2 I97 (gfint_7[1:1], choice_7, i_7r0[1:1]);
  AND2 I98 (gfint_7[2:2], choice_7, i_7r0[2:2]);
  AND2 I99 (gfint_8[0:0], choice_8, i_8r0[0:0]);
  AND2 I100 (gfint_8[1:1], choice_8, i_8r0[1:1]);
  AND2 I101 (gfint_8[2:2], choice_8, i_8r0[2:2]);
  AND2 I102 (gfint_9[0:0], choice_9, i_9r0[0:0]);
  AND2 I103 (gfint_9[1:1], choice_9, i_9r0[1:1]);
  AND2 I104 (gfint_9[2:2], choice_9, i_9r0[2:2]);
  AND2 I105 (gfint_10[0:0], choice_10, i_10r0[0:0]);
  AND2 I106 (gfint_10[1:1], choice_10, i_10r0[1:1]);
  AND2 I107 (gfint_10[2:2], choice_10, i_10r0[2:2]);
  OR2 I108 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I109 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I110 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I111 (icomp_0, comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  OR2 I112 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I113 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I114 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  C3 I115 (icomp_1, comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  OR2 I116 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I117 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I118 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  C3 I119 (icomp_2, comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  OR2 I120 (comp3_0[0:0], i_3r0[0:0], i_3r1[0:0]);
  OR2 I121 (comp3_0[1:1], i_3r0[1:1], i_3r1[1:1]);
  OR2 I122 (comp3_0[2:2], i_3r0[2:2], i_3r1[2:2]);
  C3 I123 (icomp_3, comp3_0[0:0], comp3_0[1:1], comp3_0[2:2]);
  OR2 I124 (comp4_0[0:0], i_4r0[0:0], i_4r1[0:0]);
  OR2 I125 (comp4_0[1:1], i_4r0[1:1], i_4r1[1:1]);
  OR2 I126 (comp4_0[2:2], i_4r0[2:2], i_4r1[2:2]);
  C3 I127 (icomp_4, comp4_0[0:0], comp4_0[1:1], comp4_0[2:2]);
  OR2 I128 (comp5_0[0:0], i_5r0[0:0], i_5r1[0:0]);
  OR2 I129 (comp5_0[1:1], i_5r0[1:1], i_5r1[1:1]);
  OR2 I130 (comp5_0[2:2], i_5r0[2:2], i_5r1[2:2]);
  C3 I131 (icomp_5, comp5_0[0:0], comp5_0[1:1], comp5_0[2:2]);
  OR2 I132 (comp6_0[0:0], i_6r0[0:0], i_6r1[0:0]);
  OR2 I133 (comp6_0[1:1], i_6r0[1:1], i_6r1[1:1]);
  OR2 I134 (comp6_0[2:2], i_6r0[2:2], i_6r1[2:2]);
  C3 I135 (icomp_6, comp6_0[0:0], comp6_0[1:1], comp6_0[2:2]);
  OR2 I136 (comp7_0[0:0], i_7r0[0:0], i_7r1[0:0]);
  OR2 I137 (comp7_0[1:1], i_7r0[1:1], i_7r1[1:1]);
  OR2 I138 (comp7_0[2:2], i_7r0[2:2], i_7r1[2:2]);
  C3 I139 (icomp_7, comp7_0[0:0], comp7_0[1:1], comp7_0[2:2]);
  OR2 I140 (comp8_0[0:0], i_8r0[0:0], i_8r1[0:0]);
  OR2 I141 (comp8_0[1:1], i_8r0[1:1], i_8r1[1:1]);
  OR2 I142 (comp8_0[2:2], i_8r0[2:2], i_8r1[2:2]);
  C3 I143 (icomp_8, comp8_0[0:0], comp8_0[1:1], comp8_0[2:2]);
  OR2 I144 (comp9_0[0:0], i_9r0[0:0], i_9r1[0:0]);
  OR2 I145 (comp9_0[1:1], i_9r0[1:1], i_9r1[1:1]);
  OR2 I146 (comp9_0[2:2], i_9r0[2:2], i_9r1[2:2]);
  C3 I147 (icomp_9, comp9_0[0:0], comp9_0[1:1], comp9_0[2:2]);
  OR2 I148 (comp10_0[0:0], i_10r0[0:0], i_10r1[0:0]);
  OR2 I149 (comp10_0[1:1], i_10r0[1:1], i_10r1[1:1]);
  OR2 I150 (comp10_0[2:2], i_10r0[2:2], i_10r1[2:2]);
  C3 I151 (icomp_10, comp10_0[0:0], comp10_0[1:1], comp10_0[2:2]);
  C2R I152 (choice_0, icomp_0, nchosen_0, reset);
  C2R I153 (choice_1, icomp_1, nchosen_0, reset);
  C2R I154 (choice_2, icomp_2, nchosen_0, reset);
  C2R I155 (choice_3, icomp_3, nchosen_0, reset);
  C2R I156 (choice_4, icomp_4, nchosen_0, reset);
  C2R I157 (choice_5, icomp_5, nchosen_0, reset);
  C2R I158 (choice_6, icomp_6, nchosen_0, reset);
  C2R I159 (choice_7, icomp_7, nchosen_0, reset);
  C2R I160 (choice_8, icomp_8, nchosen_0, reset);
  C2R I161 (choice_9, icomp_9, nchosen_0, reset);
  C2R I162 (choice_10, icomp_10, nchosen_0, reset);
  NOR3 I163 (simp1841_0[0:0], choice_0, choice_1, choice_2);
  NOR3 I164 (simp1841_0[1:1], choice_3, choice_4, choice_5);
  NOR3 I165 (simp1841_0[2:2], choice_6, choice_7, choice_8);
  NOR2 I166 (simp1841_0[3:3], choice_9, choice_10);
  NAND3 I167 (simp1842_0[0:0], simp1841_0[0:0], simp1841_0[1:1], simp1841_0[2:2]);
  INV I168 (simp1842_0[1:1], simp1841_0[3:3]);
  OR2 I169 (anychoice_0, simp1842_0[0:0], simp1842_0[1:1]);
  NOR2 I170 (nchosen_0, anychoice_0, o_0a);
  C2R I171 (i_0a, choice_0, o_0a, reset);
  C2R I172 (i_1a, choice_1, o_0a, reset);
  C2R I173 (i_2a, choice_2, o_0a, reset);
  C2R I174 (i_3a, choice_3, o_0a, reset);
  C2R I175 (i_4a, choice_4, o_0a, reset);
  C2R I176 (i_5a, choice_5, o_0a, reset);
  C2R I177 (i_6a, choice_6, o_0a, reset);
  C2R I178 (i_7a, choice_7, o_0a, reset);
  C2R I179 (i_8a, choice_8, o_0a, reset);
  C2R I180 (i_9a, choice_9, o_0a, reset);
  C2R I181 (i_10a, choice_10, o_0a, reset);
endmodule

// tko0m11_1nm11b1 TeakO [
//     (1,TeakOConstant 11 1)] [One 0,One 11]
module tko0m11_1nm11b1 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [10:0] o_0r0;
  output [10:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  GND I1 (o_0r0[0:0]);
  BUFF I2 (o_0r0[1:1], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  BUFF I6 (o_0r0[5:5], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  BUFF I8 (o_0r0[7:7], i_0r);
  BUFF I9 (o_0r0[8:8], i_0r);
  BUFF I10 (o_0r0[9:9], i_0r);
  BUFF I11 (o_0r0[10:10], i_0r);
  GND I12 (o_0r1[1:1]);
  GND I13 (o_0r1[2:2]);
  GND I14 (o_0r1[3:3]);
  GND I15 (o_0r1[4:4]);
  GND I16 (o_0r1[5:5]);
  GND I17 (o_0r1[6:6]);
  GND I18 (o_0r1[7:7]);
  GND I19 (o_0r1[8:8]);
  GND I20 (o_0r1[9:9]);
  GND I21 (o_0r1[10:10]);
  BUFF I22 (i_0a, o_0a);
endmodule

// tko0m11_1nm11b2 TeakO [
//     (1,TeakOConstant 11 2)] [One 0,One 11]
module tko0m11_1nm11b2 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [10:0] o_0r0;
  output [10:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[1:1], i_0r);
  GND I1 (o_0r0[1:1]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  BUFF I6 (o_0r0[5:5], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  BUFF I8 (o_0r0[7:7], i_0r);
  BUFF I9 (o_0r0[8:8], i_0r);
  BUFF I10 (o_0r0[9:9], i_0r);
  BUFF I11 (o_0r0[10:10], i_0r);
  GND I12 (o_0r1[0:0]);
  GND I13 (o_0r1[2:2]);
  GND I14 (o_0r1[3:3]);
  GND I15 (o_0r1[4:4]);
  GND I16 (o_0r1[5:5]);
  GND I17 (o_0r1[6:6]);
  GND I18 (o_0r1[7:7]);
  GND I19 (o_0r1[8:8]);
  GND I20 (o_0r1[9:9]);
  GND I21 (o_0r1[10:10]);
  BUFF I22 (i_0a, o_0a);
endmodule

// tko0m11_1nm11b4 TeakO [
//     (1,TeakOConstant 11 4)] [One 0,One 11]
module tko0m11_1nm11b4 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [10:0] o_0r0;
  output [10:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[2:2], i_0r);
  GND I1 (o_0r0[2:2]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  BUFF I6 (o_0r0[5:5], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  BUFF I8 (o_0r0[7:7], i_0r);
  BUFF I9 (o_0r0[8:8], i_0r);
  BUFF I10 (o_0r0[9:9], i_0r);
  BUFF I11 (o_0r0[10:10], i_0r);
  GND I12 (o_0r1[0:0]);
  GND I13 (o_0r1[1:1]);
  GND I14 (o_0r1[3:3]);
  GND I15 (o_0r1[4:4]);
  GND I16 (o_0r1[5:5]);
  GND I17 (o_0r1[6:6]);
  GND I18 (o_0r1[7:7]);
  GND I19 (o_0r1[8:8]);
  GND I20 (o_0r1[9:9]);
  GND I21 (o_0r1[10:10]);
  BUFF I22 (i_0a, o_0a);
endmodule

// tko0m11_1nm11b8 TeakO [
//     (1,TeakOConstant 11 8)] [One 0,One 11]
module tko0m11_1nm11b8 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [10:0] o_0r0;
  output [10:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[3:3], i_0r);
  GND I1 (o_0r0[3:3]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  BUFF I6 (o_0r0[5:5], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  BUFF I8 (o_0r0[7:7], i_0r);
  BUFF I9 (o_0r0[8:8], i_0r);
  BUFF I10 (o_0r0[9:9], i_0r);
  BUFF I11 (o_0r0[10:10], i_0r);
  GND I12 (o_0r1[0:0]);
  GND I13 (o_0r1[1:1]);
  GND I14 (o_0r1[2:2]);
  GND I15 (o_0r1[4:4]);
  GND I16 (o_0r1[5:5]);
  GND I17 (o_0r1[6:6]);
  GND I18 (o_0r1[7:7]);
  GND I19 (o_0r1[8:8]);
  GND I20 (o_0r1[9:9]);
  GND I21 (o_0r1[10:10]);
  BUFF I22 (i_0a, o_0a);
endmodule

// tko0m11_1nm11b10 TeakO [
//     (1,TeakOConstant 11 16)] [One 0,One 11]
module tko0m11_1nm11b10 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [10:0] o_0r0;
  output [10:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[4:4], i_0r);
  GND I1 (o_0r0[4:4]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  BUFF I6 (o_0r0[5:5], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  BUFF I8 (o_0r0[7:7], i_0r);
  BUFF I9 (o_0r0[8:8], i_0r);
  BUFF I10 (o_0r0[9:9], i_0r);
  BUFF I11 (o_0r0[10:10], i_0r);
  GND I12 (o_0r1[0:0]);
  GND I13 (o_0r1[1:1]);
  GND I14 (o_0r1[2:2]);
  GND I15 (o_0r1[3:3]);
  GND I16 (o_0r1[5:5]);
  GND I17 (o_0r1[6:6]);
  GND I18 (o_0r1[7:7]);
  GND I19 (o_0r1[8:8]);
  GND I20 (o_0r1[9:9]);
  GND I21 (o_0r1[10:10]);
  BUFF I22 (i_0a, o_0a);
endmodule

// tko0m11_1nm11b20 TeakO [
//     (1,TeakOConstant 11 32)] [One 0,One 11]
module tko0m11_1nm11b20 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [10:0] o_0r0;
  output [10:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[5:5], i_0r);
  GND I1 (o_0r0[5:5]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  BUFF I6 (o_0r0[4:4], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  BUFF I8 (o_0r0[7:7], i_0r);
  BUFF I9 (o_0r0[8:8], i_0r);
  BUFF I10 (o_0r0[9:9], i_0r);
  BUFF I11 (o_0r0[10:10], i_0r);
  GND I12 (o_0r1[0:0]);
  GND I13 (o_0r1[1:1]);
  GND I14 (o_0r1[2:2]);
  GND I15 (o_0r1[3:3]);
  GND I16 (o_0r1[4:4]);
  GND I17 (o_0r1[6:6]);
  GND I18 (o_0r1[7:7]);
  GND I19 (o_0r1[8:8]);
  GND I20 (o_0r1[9:9]);
  GND I21 (o_0r1[10:10]);
  BUFF I22 (i_0a, o_0a);
endmodule

// tko0m11_1nm11b40 TeakO [
//     (1,TeakOConstant 11 64)] [One 0,One 11]
module tko0m11_1nm11b40 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [10:0] o_0r0;
  output [10:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[6:6], i_0r);
  GND I1 (o_0r0[6:6]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  BUFF I6 (o_0r0[4:4], i_0r);
  BUFF I7 (o_0r0[5:5], i_0r);
  BUFF I8 (o_0r0[7:7], i_0r);
  BUFF I9 (o_0r0[8:8], i_0r);
  BUFF I10 (o_0r0[9:9], i_0r);
  BUFF I11 (o_0r0[10:10], i_0r);
  GND I12 (o_0r1[0:0]);
  GND I13 (o_0r1[1:1]);
  GND I14 (o_0r1[2:2]);
  GND I15 (o_0r1[3:3]);
  GND I16 (o_0r1[4:4]);
  GND I17 (o_0r1[5:5]);
  GND I18 (o_0r1[7:7]);
  GND I19 (o_0r1[8:8]);
  GND I20 (o_0r1[9:9]);
  GND I21 (o_0r1[10:10]);
  BUFF I22 (i_0a, o_0a);
endmodule

// tko0m11_1nm11b80 TeakO [
//     (1,TeakOConstant 11 128)] [One 0,One 11]
module tko0m11_1nm11b80 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [10:0] o_0r0;
  output [10:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[7:7], i_0r);
  GND I1 (o_0r0[7:7]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  BUFF I6 (o_0r0[4:4], i_0r);
  BUFF I7 (o_0r0[5:5], i_0r);
  BUFF I8 (o_0r0[6:6], i_0r);
  BUFF I9 (o_0r0[8:8], i_0r);
  BUFF I10 (o_0r0[9:9], i_0r);
  BUFF I11 (o_0r0[10:10], i_0r);
  GND I12 (o_0r1[0:0]);
  GND I13 (o_0r1[1:1]);
  GND I14 (o_0r1[2:2]);
  GND I15 (o_0r1[3:3]);
  GND I16 (o_0r1[4:4]);
  GND I17 (o_0r1[5:5]);
  GND I18 (o_0r1[6:6]);
  GND I19 (o_0r1[8:8]);
  GND I20 (o_0r1[9:9]);
  GND I21 (o_0r1[10:10]);
  BUFF I22 (i_0a, o_0a);
endmodule

// tko0m11_1nm11b100 TeakO [
//     (1,TeakOConstant 11 256)] [One 0,One 11]
module tko0m11_1nm11b100 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [10:0] o_0r0;
  output [10:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[8:8], i_0r);
  GND I1 (o_0r0[8:8]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  BUFF I6 (o_0r0[4:4], i_0r);
  BUFF I7 (o_0r0[5:5], i_0r);
  BUFF I8 (o_0r0[6:6], i_0r);
  BUFF I9 (o_0r0[7:7], i_0r);
  BUFF I10 (o_0r0[9:9], i_0r);
  BUFF I11 (o_0r0[10:10], i_0r);
  GND I12 (o_0r1[0:0]);
  GND I13 (o_0r1[1:1]);
  GND I14 (o_0r1[2:2]);
  GND I15 (o_0r1[3:3]);
  GND I16 (o_0r1[4:4]);
  GND I17 (o_0r1[5:5]);
  GND I18 (o_0r1[6:6]);
  GND I19 (o_0r1[7:7]);
  GND I20 (o_0r1[9:9]);
  GND I21 (o_0r1[10:10]);
  BUFF I22 (i_0a, o_0a);
endmodule

// tko0m11_1nm11b200 TeakO [
//     (1,TeakOConstant 11 512)] [One 0,One 11]
module tko0m11_1nm11b200 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [10:0] o_0r0;
  output [10:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[9:9], i_0r);
  GND I1 (o_0r0[9:9]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  BUFF I6 (o_0r0[4:4], i_0r);
  BUFF I7 (o_0r0[5:5], i_0r);
  BUFF I8 (o_0r0[6:6], i_0r);
  BUFF I9 (o_0r0[7:7], i_0r);
  BUFF I10 (o_0r0[8:8], i_0r);
  BUFF I11 (o_0r0[10:10], i_0r);
  GND I12 (o_0r1[0:0]);
  GND I13 (o_0r1[1:1]);
  GND I14 (o_0r1[2:2]);
  GND I15 (o_0r1[3:3]);
  GND I16 (o_0r1[4:4]);
  GND I17 (o_0r1[5:5]);
  GND I18 (o_0r1[6:6]);
  GND I19 (o_0r1[7:7]);
  GND I20 (o_0r1[8:8]);
  GND I21 (o_0r1[10:10]);
  BUFF I22 (i_0a, o_0a);
endmodule

// tko0m11_1nm11b400 TeakO [
//     (1,TeakOConstant 11 1024)] [One 0,One 11]
module tko0m11_1nm11b400 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [10:0] o_0r0;
  output [10:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[10:10], i_0r);
  GND I1 (o_0r0[10:10]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  BUFF I6 (o_0r0[4:4], i_0r);
  BUFF I7 (o_0r0[5:5], i_0r);
  BUFF I8 (o_0r0[6:6], i_0r);
  BUFF I9 (o_0r0[7:7], i_0r);
  BUFF I10 (o_0r0[8:8], i_0r);
  BUFF I11 (o_0r0[9:9], i_0r);
  GND I12 (o_0r1[0:0]);
  GND I13 (o_0r1[1:1]);
  GND I14 (o_0r1[2:2]);
  GND I15 (o_0r1[3:3]);
  GND I16 (o_0r1[4:4]);
  GND I17 (o_0r1[5:5]);
  GND I18 (o_0r1[6:6]);
  GND I19 (o_0r1[7:7]);
  GND I20 (o_0r1[8:8]);
  GND I21 (o_0r1[9:9]);
  BUFF I22 (i_0a, o_0a);
endmodule

// tkm11x11b TeakM [Many [11,11,11,11,11,11,11,11,11,11,11],One 11]
module tkm11x11b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, i_4r0, i_4r1, i_4a, i_5r0, i_5r1, i_5a, i_6r0, i_6r1, i_6a, i_7r0, i_7r1, i_7a, i_8r0, i_8r1, i_8a, i_9r0, i_9r1, i_9a, i_10r0, i_10r1, i_10a, o_0r0, o_0r1, o_0a, reset);
  input [10:0] i_0r0;
  input [10:0] i_0r1;
  output i_0a;
  input [10:0] i_1r0;
  input [10:0] i_1r1;
  output i_1a;
  input [10:0] i_2r0;
  input [10:0] i_2r1;
  output i_2a;
  input [10:0] i_3r0;
  input [10:0] i_3r1;
  output i_3a;
  input [10:0] i_4r0;
  input [10:0] i_4r1;
  output i_4a;
  input [10:0] i_5r0;
  input [10:0] i_5r1;
  output i_5a;
  input [10:0] i_6r0;
  input [10:0] i_6r1;
  output i_6a;
  input [10:0] i_7r0;
  input [10:0] i_7r1;
  output i_7a;
  input [10:0] i_8r0;
  input [10:0] i_8r1;
  output i_8a;
  input [10:0] i_9r0;
  input [10:0] i_9r1;
  output i_9a;
  input [10:0] i_10r0;
  input [10:0] i_10r1;
  output i_10a;
  output [10:0] o_0r0;
  output [10:0] o_0r1;
  input o_0a;
  input reset;
  wire [10:0] gfint_0;
  wire [10:0] gfint_1;
  wire [10:0] gfint_2;
  wire [10:0] gfint_3;
  wire [10:0] gfint_4;
  wire [10:0] gfint_5;
  wire [10:0] gfint_6;
  wire [10:0] gfint_7;
  wire [10:0] gfint_8;
  wire [10:0] gfint_9;
  wire [10:0] gfint_10;
  wire [10:0] gtint_0;
  wire [10:0] gtint_1;
  wire [10:0] gtint_2;
  wire [10:0] gtint_3;
  wire [10:0] gtint_4;
  wire [10:0] gtint_5;
  wire [10:0] gtint_6;
  wire [10:0] gtint_7;
  wire [10:0] gtint_8;
  wire [10:0] gtint_9;
  wire [10:0] gtint_10;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire choice_4;
  wire choice_5;
  wire choice_6;
  wire choice_7;
  wire choice_8;
  wire choice_9;
  wire choice_10;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire icomp_3;
  wire icomp_4;
  wire icomp_5;
  wire icomp_6;
  wire icomp_7;
  wire icomp_8;
  wire icomp_9;
  wire icomp_10;
  wire nchosen_0;
  wire [3:0] simp461_0;
  wire [1:0] simp462_0;
  wire [3:0] simp471_0;
  wire [1:0] simp472_0;
  wire [3:0] simp481_0;
  wire [1:0] simp482_0;
  wire [3:0] simp491_0;
  wire [1:0] simp492_0;
  wire [3:0] simp501_0;
  wire [1:0] simp502_0;
  wire [3:0] simp511_0;
  wire [1:0] simp512_0;
  wire [3:0] simp521_0;
  wire [1:0] simp522_0;
  wire [3:0] simp531_0;
  wire [1:0] simp532_0;
  wire [3:0] simp541_0;
  wire [1:0] simp542_0;
  wire [3:0] simp551_0;
  wire [1:0] simp552_0;
  wire [3:0] simp561_0;
  wire [1:0] simp562_0;
  wire [3:0] simp571_0;
  wire [1:0] simp572_0;
  wire [3:0] simp581_0;
  wire [1:0] simp582_0;
  wire [3:0] simp591_0;
  wire [1:0] simp592_0;
  wire [3:0] simp601_0;
  wire [1:0] simp602_0;
  wire [3:0] simp611_0;
  wire [1:0] simp612_0;
  wire [3:0] simp621_0;
  wire [1:0] simp622_0;
  wire [3:0] simp631_0;
  wire [1:0] simp632_0;
  wire [3:0] simp641_0;
  wire [1:0] simp642_0;
  wire [3:0] simp651_0;
  wire [1:0] simp652_0;
  wire [3:0] simp661_0;
  wire [1:0] simp662_0;
  wire [3:0] simp671_0;
  wire [1:0] simp672_0;
  wire [10:0] comp0_0;
  wire [3:0] simp3221_0;
  wire [1:0] simp3222_0;
  wire [10:0] comp1_0;
  wire [3:0] simp3351_0;
  wire [1:0] simp3352_0;
  wire [10:0] comp2_0;
  wire [3:0] simp3481_0;
  wire [1:0] simp3482_0;
  wire [10:0] comp3_0;
  wire [3:0] simp3611_0;
  wire [1:0] simp3612_0;
  wire [10:0] comp4_0;
  wire [3:0] simp3741_0;
  wire [1:0] simp3742_0;
  wire [10:0] comp5_0;
  wire [3:0] simp3871_0;
  wire [1:0] simp3872_0;
  wire [10:0] comp6_0;
  wire [3:0] simp4001_0;
  wire [1:0] simp4002_0;
  wire [10:0] comp7_0;
  wire [3:0] simp4131_0;
  wire [1:0] simp4132_0;
  wire [10:0] comp8_0;
  wire [3:0] simp4261_0;
  wire [1:0] simp4262_0;
  wire [10:0] comp9_0;
  wire [3:0] simp4391_0;
  wire [1:0] simp4392_0;
  wire [10:0] comp10_0;
  wire [3:0] simp4521_0;
  wire [1:0] simp4522_0;
  wire [3:0] simp4641_0;
  wire [1:0] simp4642_0;
  NOR3 I0 (simp461_0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  NOR3 I1 (simp461_0[1:1], gfint_3[0:0], gfint_4[0:0], gfint_5[0:0]);
  NOR3 I2 (simp461_0[2:2], gfint_6[0:0], gfint_7[0:0], gfint_8[0:0]);
  NOR2 I3 (simp461_0[3:3], gfint_9[0:0], gfint_10[0:0]);
  NAND3 I4 (simp462_0[0:0], simp461_0[0:0], simp461_0[1:1], simp461_0[2:2]);
  INV I5 (simp462_0[1:1], simp461_0[3:3]);
  OR2 I6 (o_0r0[0:0], simp462_0[0:0], simp462_0[1:1]);
  NOR3 I7 (simp471_0[0:0], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  NOR3 I8 (simp471_0[1:1], gfint_3[1:1], gfint_4[1:1], gfint_5[1:1]);
  NOR3 I9 (simp471_0[2:2], gfint_6[1:1], gfint_7[1:1], gfint_8[1:1]);
  NOR2 I10 (simp471_0[3:3], gfint_9[1:1], gfint_10[1:1]);
  NAND3 I11 (simp472_0[0:0], simp471_0[0:0], simp471_0[1:1], simp471_0[2:2]);
  INV I12 (simp472_0[1:1], simp471_0[3:3]);
  OR2 I13 (o_0r0[1:1], simp472_0[0:0], simp472_0[1:1]);
  NOR3 I14 (simp481_0[0:0], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  NOR3 I15 (simp481_0[1:1], gfint_3[2:2], gfint_4[2:2], gfint_5[2:2]);
  NOR3 I16 (simp481_0[2:2], gfint_6[2:2], gfint_7[2:2], gfint_8[2:2]);
  NOR2 I17 (simp481_0[3:3], gfint_9[2:2], gfint_10[2:2]);
  NAND3 I18 (simp482_0[0:0], simp481_0[0:0], simp481_0[1:1], simp481_0[2:2]);
  INV I19 (simp482_0[1:1], simp481_0[3:3]);
  OR2 I20 (o_0r0[2:2], simp482_0[0:0], simp482_0[1:1]);
  NOR3 I21 (simp491_0[0:0], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  NOR3 I22 (simp491_0[1:1], gfint_3[3:3], gfint_4[3:3], gfint_5[3:3]);
  NOR3 I23 (simp491_0[2:2], gfint_6[3:3], gfint_7[3:3], gfint_8[3:3]);
  NOR2 I24 (simp491_0[3:3], gfint_9[3:3], gfint_10[3:3]);
  NAND3 I25 (simp492_0[0:0], simp491_0[0:0], simp491_0[1:1], simp491_0[2:2]);
  INV I26 (simp492_0[1:1], simp491_0[3:3]);
  OR2 I27 (o_0r0[3:3], simp492_0[0:0], simp492_0[1:1]);
  NOR3 I28 (simp501_0[0:0], gfint_0[4:4], gfint_1[4:4], gfint_2[4:4]);
  NOR3 I29 (simp501_0[1:1], gfint_3[4:4], gfint_4[4:4], gfint_5[4:4]);
  NOR3 I30 (simp501_0[2:2], gfint_6[4:4], gfint_7[4:4], gfint_8[4:4]);
  NOR2 I31 (simp501_0[3:3], gfint_9[4:4], gfint_10[4:4]);
  NAND3 I32 (simp502_0[0:0], simp501_0[0:0], simp501_0[1:1], simp501_0[2:2]);
  INV I33 (simp502_0[1:1], simp501_0[3:3]);
  OR2 I34 (o_0r0[4:4], simp502_0[0:0], simp502_0[1:1]);
  NOR3 I35 (simp511_0[0:0], gfint_0[5:5], gfint_1[5:5], gfint_2[5:5]);
  NOR3 I36 (simp511_0[1:1], gfint_3[5:5], gfint_4[5:5], gfint_5[5:5]);
  NOR3 I37 (simp511_0[2:2], gfint_6[5:5], gfint_7[5:5], gfint_8[5:5]);
  NOR2 I38 (simp511_0[3:3], gfint_9[5:5], gfint_10[5:5]);
  NAND3 I39 (simp512_0[0:0], simp511_0[0:0], simp511_0[1:1], simp511_0[2:2]);
  INV I40 (simp512_0[1:1], simp511_0[3:3]);
  OR2 I41 (o_0r0[5:5], simp512_0[0:0], simp512_0[1:1]);
  NOR3 I42 (simp521_0[0:0], gfint_0[6:6], gfint_1[6:6], gfint_2[6:6]);
  NOR3 I43 (simp521_0[1:1], gfint_3[6:6], gfint_4[6:6], gfint_5[6:6]);
  NOR3 I44 (simp521_0[2:2], gfint_6[6:6], gfint_7[6:6], gfint_8[6:6]);
  NOR2 I45 (simp521_0[3:3], gfint_9[6:6], gfint_10[6:6]);
  NAND3 I46 (simp522_0[0:0], simp521_0[0:0], simp521_0[1:1], simp521_0[2:2]);
  INV I47 (simp522_0[1:1], simp521_0[3:3]);
  OR2 I48 (o_0r0[6:6], simp522_0[0:0], simp522_0[1:1]);
  NOR3 I49 (simp531_0[0:0], gfint_0[7:7], gfint_1[7:7], gfint_2[7:7]);
  NOR3 I50 (simp531_0[1:1], gfint_3[7:7], gfint_4[7:7], gfint_5[7:7]);
  NOR3 I51 (simp531_0[2:2], gfint_6[7:7], gfint_7[7:7], gfint_8[7:7]);
  NOR2 I52 (simp531_0[3:3], gfint_9[7:7], gfint_10[7:7]);
  NAND3 I53 (simp532_0[0:0], simp531_0[0:0], simp531_0[1:1], simp531_0[2:2]);
  INV I54 (simp532_0[1:1], simp531_0[3:3]);
  OR2 I55 (o_0r0[7:7], simp532_0[0:0], simp532_0[1:1]);
  NOR3 I56 (simp541_0[0:0], gfint_0[8:8], gfint_1[8:8], gfint_2[8:8]);
  NOR3 I57 (simp541_0[1:1], gfint_3[8:8], gfint_4[8:8], gfint_5[8:8]);
  NOR3 I58 (simp541_0[2:2], gfint_6[8:8], gfint_7[8:8], gfint_8[8:8]);
  NOR2 I59 (simp541_0[3:3], gfint_9[8:8], gfint_10[8:8]);
  NAND3 I60 (simp542_0[0:0], simp541_0[0:0], simp541_0[1:1], simp541_0[2:2]);
  INV I61 (simp542_0[1:1], simp541_0[3:3]);
  OR2 I62 (o_0r0[8:8], simp542_0[0:0], simp542_0[1:1]);
  NOR3 I63 (simp551_0[0:0], gfint_0[9:9], gfint_1[9:9], gfint_2[9:9]);
  NOR3 I64 (simp551_0[1:1], gfint_3[9:9], gfint_4[9:9], gfint_5[9:9]);
  NOR3 I65 (simp551_0[2:2], gfint_6[9:9], gfint_7[9:9], gfint_8[9:9]);
  NOR2 I66 (simp551_0[3:3], gfint_9[9:9], gfint_10[9:9]);
  NAND3 I67 (simp552_0[0:0], simp551_0[0:0], simp551_0[1:1], simp551_0[2:2]);
  INV I68 (simp552_0[1:1], simp551_0[3:3]);
  OR2 I69 (o_0r0[9:9], simp552_0[0:0], simp552_0[1:1]);
  NOR3 I70 (simp561_0[0:0], gfint_0[10:10], gfint_1[10:10], gfint_2[10:10]);
  NOR3 I71 (simp561_0[1:1], gfint_3[10:10], gfint_4[10:10], gfint_5[10:10]);
  NOR3 I72 (simp561_0[2:2], gfint_6[10:10], gfint_7[10:10], gfint_8[10:10]);
  NOR2 I73 (simp561_0[3:3], gfint_9[10:10], gfint_10[10:10]);
  NAND3 I74 (simp562_0[0:0], simp561_0[0:0], simp561_0[1:1], simp561_0[2:2]);
  INV I75 (simp562_0[1:1], simp561_0[3:3]);
  OR2 I76 (o_0r0[10:10], simp562_0[0:0], simp562_0[1:1]);
  NOR3 I77 (simp571_0[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  NOR3 I78 (simp571_0[1:1], gtint_3[0:0], gtint_4[0:0], gtint_5[0:0]);
  NOR3 I79 (simp571_0[2:2], gtint_6[0:0], gtint_7[0:0], gtint_8[0:0]);
  NOR2 I80 (simp571_0[3:3], gtint_9[0:0], gtint_10[0:0]);
  NAND3 I81 (simp572_0[0:0], simp571_0[0:0], simp571_0[1:1], simp571_0[2:2]);
  INV I82 (simp572_0[1:1], simp571_0[3:3]);
  OR2 I83 (o_0r1[0:0], simp572_0[0:0], simp572_0[1:1]);
  NOR3 I84 (simp581_0[0:0], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  NOR3 I85 (simp581_0[1:1], gtint_3[1:1], gtint_4[1:1], gtint_5[1:1]);
  NOR3 I86 (simp581_0[2:2], gtint_6[1:1], gtint_7[1:1], gtint_8[1:1]);
  NOR2 I87 (simp581_0[3:3], gtint_9[1:1], gtint_10[1:1]);
  NAND3 I88 (simp582_0[0:0], simp581_0[0:0], simp581_0[1:1], simp581_0[2:2]);
  INV I89 (simp582_0[1:1], simp581_0[3:3]);
  OR2 I90 (o_0r1[1:1], simp582_0[0:0], simp582_0[1:1]);
  NOR3 I91 (simp591_0[0:0], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  NOR3 I92 (simp591_0[1:1], gtint_3[2:2], gtint_4[2:2], gtint_5[2:2]);
  NOR3 I93 (simp591_0[2:2], gtint_6[2:2], gtint_7[2:2], gtint_8[2:2]);
  NOR2 I94 (simp591_0[3:3], gtint_9[2:2], gtint_10[2:2]);
  NAND3 I95 (simp592_0[0:0], simp591_0[0:0], simp591_0[1:1], simp591_0[2:2]);
  INV I96 (simp592_0[1:1], simp591_0[3:3]);
  OR2 I97 (o_0r1[2:2], simp592_0[0:0], simp592_0[1:1]);
  NOR3 I98 (simp601_0[0:0], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  NOR3 I99 (simp601_0[1:1], gtint_3[3:3], gtint_4[3:3], gtint_5[3:3]);
  NOR3 I100 (simp601_0[2:2], gtint_6[3:3], gtint_7[3:3], gtint_8[3:3]);
  NOR2 I101 (simp601_0[3:3], gtint_9[3:3], gtint_10[3:3]);
  NAND3 I102 (simp602_0[0:0], simp601_0[0:0], simp601_0[1:1], simp601_0[2:2]);
  INV I103 (simp602_0[1:1], simp601_0[3:3]);
  OR2 I104 (o_0r1[3:3], simp602_0[0:0], simp602_0[1:1]);
  NOR3 I105 (simp611_0[0:0], gtint_0[4:4], gtint_1[4:4], gtint_2[4:4]);
  NOR3 I106 (simp611_0[1:1], gtint_3[4:4], gtint_4[4:4], gtint_5[4:4]);
  NOR3 I107 (simp611_0[2:2], gtint_6[4:4], gtint_7[4:4], gtint_8[4:4]);
  NOR2 I108 (simp611_0[3:3], gtint_9[4:4], gtint_10[4:4]);
  NAND3 I109 (simp612_0[0:0], simp611_0[0:0], simp611_0[1:1], simp611_0[2:2]);
  INV I110 (simp612_0[1:1], simp611_0[3:3]);
  OR2 I111 (o_0r1[4:4], simp612_0[0:0], simp612_0[1:1]);
  NOR3 I112 (simp621_0[0:0], gtint_0[5:5], gtint_1[5:5], gtint_2[5:5]);
  NOR3 I113 (simp621_0[1:1], gtint_3[5:5], gtint_4[5:5], gtint_5[5:5]);
  NOR3 I114 (simp621_0[2:2], gtint_6[5:5], gtint_7[5:5], gtint_8[5:5]);
  NOR2 I115 (simp621_0[3:3], gtint_9[5:5], gtint_10[5:5]);
  NAND3 I116 (simp622_0[0:0], simp621_0[0:0], simp621_0[1:1], simp621_0[2:2]);
  INV I117 (simp622_0[1:1], simp621_0[3:3]);
  OR2 I118 (o_0r1[5:5], simp622_0[0:0], simp622_0[1:1]);
  NOR3 I119 (simp631_0[0:0], gtint_0[6:6], gtint_1[6:6], gtint_2[6:6]);
  NOR3 I120 (simp631_0[1:1], gtint_3[6:6], gtint_4[6:6], gtint_5[6:6]);
  NOR3 I121 (simp631_0[2:2], gtint_6[6:6], gtint_7[6:6], gtint_8[6:6]);
  NOR2 I122 (simp631_0[3:3], gtint_9[6:6], gtint_10[6:6]);
  NAND3 I123 (simp632_0[0:0], simp631_0[0:0], simp631_0[1:1], simp631_0[2:2]);
  INV I124 (simp632_0[1:1], simp631_0[3:3]);
  OR2 I125 (o_0r1[6:6], simp632_0[0:0], simp632_0[1:1]);
  NOR3 I126 (simp641_0[0:0], gtint_0[7:7], gtint_1[7:7], gtint_2[7:7]);
  NOR3 I127 (simp641_0[1:1], gtint_3[7:7], gtint_4[7:7], gtint_5[7:7]);
  NOR3 I128 (simp641_0[2:2], gtint_6[7:7], gtint_7[7:7], gtint_8[7:7]);
  NOR2 I129 (simp641_0[3:3], gtint_9[7:7], gtint_10[7:7]);
  NAND3 I130 (simp642_0[0:0], simp641_0[0:0], simp641_0[1:1], simp641_0[2:2]);
  INV I131 (simp642_0[1:1], simp641_0[3:3]);
  OR2 I132 (o_0r1[7:7], simp642_0[0:0], simp642_0[1:1]);
  NOR3 I133 (simp651_0[0:0], gtint_0[8:8], gtint_1[8:8], gtint_2[8:8]);
  NOR3 I134 (simp651_0[1:1], gtint_3[8:8], gtint_4[8:8], gtint_5[8:8]);
  NOR3 I135 (simp651_0[2:2], gtint_6[8:8], gtint_7[8:8], gtint_8[8:8]);
  NOR2 I136 (simp651_0[3:3], gtint_9[8:8], gtint_10[8:8]);
  NAND3 I137 (simp652_0[0:0], simp651_0[0:0], simp651_0[1:1], simp651_0[2:2]);
  INV I138 (simp652_0[1:1], simp651_0[3:3]);
  OR2 I139 (o_0r1[8:8], simp652_0[0:0], simp652_0[1:1]);
  NOR3 I140 (simp661_0[0:0], gtint_0[9:9], gtint_1[9:9], gtint_2[9:9]);
  NOR3 I141 (simp661_0[1:1], gtint_3[9:9], gtint_4[9:9], gtint_5[9:9]);
  NOR3 I142 (simp661_0[2:2], gtint_6[9:9], gtint_7[9:9], gtint_8[9:9]);
  NOR2 I143 (simp661_0[3:3], gtint_9[9:9], gtint_10[9:9]);
  NAND3 I144 (simp662_0[0:0], simp661_0[0:0], simp661_0[1:1], simp661_0[2:2]);
  INV I145 (simp662_0[1:1], simp661_0[3:3]);
  OR2 I146 (o_0r1[9:9], simp662_0[0:0], simp662_0[1:1]);
  NOR3 I147 (simp671_0[0:0], gtint_0[10:10], gtint_1[10:10], gtint_2[10:10]);
  NOR3 I148 (simp671_0[1:1], gtint_3[10:10], gtint_4[10:10], gtint_5[10:10]);
  NOR3 I149 (simp671_0[2:2], gtint_6[10:10], gtint_7[10:10], gtint_8[10:10]);
  NOR2 I150 (simp671_0[3:3], gtint_9[10:10], gtint_10[10:10]);
  NAND3 I151 (simp672_0[0:0], simp671_0[0:0], simp671_0[1:1], simp671_0[2:2]);
  INV I152 (simp672_0[1:1], simp671_0[3:3]);
  OR2 I153 (o_0r1[10:10], simp672_0[0:0], simp672_0[1:1]);
  AND2 I154 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I155 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I156 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I157 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I158 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I159 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I160 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I161 (gtint_0[7:7], choice_0, i_0r1[7:7]);
  AND2 I162 (gtint_0[8:8], choice_0, i_0r1[8:8]);
  AND2 I163 (gtint_0[9:9], choice_0, i_0r1[9:9]);
  AND2 I164 (gtint_0[10:10], choice_0, i_0r1[10:10]);
  AND2 I165 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I166 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I167 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I168 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I169 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I170 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I171 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I172 (gtint_1[7:7], choice_1, i_1r1[7:7]);
  AND2 I173 (gtint_1[8:8], choice_1, i_1r1[8:8]);
  AND2 I174 (gtint_1[9:9], choice_1, i_1r1[9:9]);
  AND2 I175 (gtint_1[10:10], choice_1, i_1r1[10:10]);
  AND2 I176 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I177 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I178 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I179 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AND2 I180 (gtint_2[4:4], choice_2, i_2r1[4:4]);
  AND2 I181 (gtint_2[5:5], choice_2, i_2r1[5:5]);
  AND2 I182 (gtint_2[6:6], choice_2, i_2r1[6:6]);
  AND2 I183 (gtint_2[7:7], choice_2, i_2r1[7:7]);
  AND2 I184 (gtint_2[8:8], choice_2, i_2r1[8:8]);
  AND2 I185 (gtint_2[9:9], choice_2, i_2r1[9:9]);
  AND2 I186 (gtint_2[10:10], choice_2, i_2r1[10:10]);
  AND2 I187 (gtint_3[0:0], choice_3, i_3r1[0:0]);
  AND2 I188 (gtint_3[1:1], choice_3, i_3r1[1:1]);
  AND2 I189 (gtint_3[2:2], choice_3, i_3r1[2:2]);
  AND2 I190 (gtint_3[3:3], choice_3, i_3r1[3:3]);
  AND2 I191 (gtint_3[4:4], choice_3, i_3r1[4:4]);
  AND2 I192 (gtint_3[5:5], choice_3, i_3r1[5:5]);
  AND2 I193 (gtint_3[6:6], choice_3, i_3r1[6:6]);
  AND2 I194 (gtint_3[7:7], choice_3, i_3r1[7:7]);
  AND2 I195 (gtint_3[8:8], choice_3, i_3r1[8:8]);
  AND2 I196 (gtint_3[9:9], choice_3, i_3r1[9:9]);
  AND2 I197 (gtint_3[10:10], choice_3, i_3r1[10:10]);
  AND2 I198 (gtint_4[0:0], choice_4, i_4r1[0:0]);
  AND2 I199 (gtint_4[1:1], choice_4, i_4r1[1:1]);
  AND2 I200 (gtint_4[2:2], choice_4, i_4r1[2:2]);
  AND2 I201 (gtint_4[3:3], choice_4, i_4r1[3:3]);
  AND2 I202 (gtint_4[4:4], choice_4, i_4r1[4:4]);
  AND2 I203 (gtint_4[5:5], choice_4, i_4r1[5:5]);
  AND2 I204 (gtint_4[6:6], choice_4, i_4r1[6:6]);
  AND2 I205 (gtint_4[7:7], choice_4, i_4r1[7:7]);
  AND2 I206 (gtint_4[8:8], choice_4, i_4r1[8:8]);
  AND2 I207 (gtint_4[9:9], choice_4, i_4r1[9:9]);
  AND2 I208 (gtint_4[10:10], choice_4, i_4r1[10:10]);
  AND2 I209 (gtint_5[0:0], choice_5, i_5r1[0:0]);
  AND2 I210 (gtint_5[1:1], choice_5, i_5r1[1:1]);
  AND2 I211 (gtint_5[2:2], choice_5, i_5r1[2:2]);
  AND2 I212 (gtint_5[3:3], choice_5, i_5r1[3:3]);
  AND2 I213 (gtint_5[4:4], choice_5, i_5r1[4:4]);
  AND2 I214 (gtint_5[5:5], choice_5, i_5r1[5:5]);
  AND2 I215 (gtint_5[6:6], choice_5, i_5r1[6:6]);
  AND2 I216 (gtint_5[7:7], choice_5, i_5r1[7:7]);
  AND2 I217 (gtint_5[8:8], choice_5, i_5r1[8:8]);
  AND2 I218 (gtint_5[9:9], choice_5, i_5r1[9:9]);
  AND2 I219 (gtint_5[10:10], choice_5, i_5r1[10:10]);
  AND2 I220 (gtint_6[0:0], choice_6, i_6r1[0:0]);
  AND2 I221 (gtint_6[1:1], choice_6, i_6r1[1:1]);
  AND2 I222 (gtint_6[2:2], choice_6, i_6r1[2:2]);
  AND2 I223 (gtint_6[3:3], choice_6, i_6r1[3:3]);
  AND2 I224 (gtint_6[4:4], choice_6, i_6r1[4:4]);
  AND2 I225 (gtint_6[5:5], choice_6, i_6r1[5:5]);
  AND2 I226 (gtint_6[6:6], choice_6, i_6r1[6:6]);
  AND2 I227 (gtint_6[7:7], choice_6, i_6r1[7:7]);
  AND2 I228 (gtint_6[8:8], choice_6, i_6r1[8:8]);
  AND2 I229 (gtint_6[9:9], choice_6, i_6r1[9:9]);
  AND2 I230 (gtint_6[10:10], choice_6, i_6r1[10:10]);
  AND2 I231 (gtint_7[0:0], choice_7, i_7r1[0:0]);
  AND2 I232 (gtint_7[1:1], choice_7, i_7r1[1:1]);
  AND2 I233 (gtint_7[2:2], choice_7, i_7r1[2:2]);
  AND2 I234 (gtint_7[3:3], choice_7, i_7r1[3:3]);
  AND2 I235 (gtint_7[4:4], choice_7, i_7r1[4:4]);
  AND2 I236 (gtint_7[5:5], choice_7, i_7r1[5:5]);
  AND2 I237 (gtint_7[6:6], choice_7, i_7r1[6:6]);
  AND2 I238 (gtint_7[7:7], choice_7, i_7r1[7:7]);
  AND2 I239 (gtint_7[8:8], choice_7, i_7r1[8:8]);
  AND2 I240 (gtint_7[9:9], choice_7, i_7r1[9:9]);
  AND2 I241 (gtint_7[10:10], choice_7, i_7r1[10:10]);
  AND2 I242 (gtint_8[0:0], choice_8, i_8r1[0:0]);
  AND2 I243 (gtint_8[1:1], choice_8, i_8r1[1:1]);
  AND2 I244 (gtint_8[2:2], choice_8, i_8r1[2:2]);
  AND2 I245 (gtint_8[3:3], choice_8, i_8r1[3:3]);
  AND2 I246 (gtint_8[4:4], choice_8, i_8r1[4:4]);
  AND2 I247 (gtint_8[5:5], choice_8, i_8r1[5:5]);
  AND2 I248 (gtint_8[6:6], choice_8, i_8r1[6:6]);
  AND2 I249 (gtint_8[7:7], choice_8, i_8r1[7:7]);
  AND2 I250 (gtint_8[8:8], choice_8, i_8r1[8:8]);
  AND2 I251 (gtint_8[9:9], choice_8, i_8r1[9:9]);
  AND2 I252 (gtint_8[10:10], choice_8, i_8r1[10:10]);
  AND2 I253 (gtint_9[0:0], choice_9, i_9r1[0:0]);
  AND2 I254 (gtint_9[1:1], choice_9, i_9r1[1:1]);
  AND2 I255 (gtint_9[2:2], choice_9, i_9r1[2:2]);
  AND2 I256 (gtint_9[3:3], choice_9, i_9r1[3:3]);
  AND2 I257 (gtint_9[4:4], choice_9, i_9r1[4:4]);
  AND2 I258 (gtint_9[5:5], choice_9, i_9r1[5:5]);
  AND2 I259 (gtint_9[6:6], choice_9, i_9r1[6:6]);
  AND2 I260 (gtint_9[7:7], choice_9, i_9r1[7:7]);
  AND2 I261 (gtint_9[8:8], choice_9, i_9r1[8:8]);
  AND2 I262 (gtint_9[9:9], choice_9, i_9r1[9:9]);
  AND2 I263 (gtint_9[10:10], choice_9, i_9r1[10:10]);
  AND2 I264 (gtint_10[0:0], choice_10, i_10r1[0:0]);
  AND2 I265 (gtint_10[1:1], choice_10, i_10r1[1:1]);
  AND2 I266 (gtint_10[2:2], choice_10, i_10r1[2:2]);
  AND2 I267 (gtint_10[3:3], choice_10, i_10r1[3:3]);
  AND2 I268 (gtint_10[4:4], choice_10, i_10r1[4:4]);
  AND2 I269 (gtint_10[5:5], choice_10, i_10r1[5:5]);
  AND2 I270 (gtint_10[6:6], choice_10, i_10r1[6:6]);
  AND2 I271 (gtint_10[7:7], choice_10, i_10r1[7:7]);
  AND2 I272 (gtint_10[8:8], choice_10, i_10r1[8:8]);
  AND2 I273 (gtint_10[9:9], choice_10, i_10r1[9:9]);
  AND2 I274 (gtint_10[10:10], choice_10, i_10r1[10:10]);
  AND2 I275 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I276 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I277 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I278 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I279 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I280 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I281 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I282 (gfint_0[7:7], choice_0, i_0r0[7:7]);
  AND2 I283 (gfint_0[8:8], choice_0, i_0r0[8:8]);
  AND2 I284 (gfint_0[9:9], choice_0, i_0r0[9:9]);
  AND2 I285 (gfint_0[10:10], choice_0, i_0r0[10:10]);
  AND2 I286 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I287 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I288 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I289 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I290 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I291 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I292 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I293 (gfint_1[7:7], choice_1, i_1r0[7:7]);
  AND2 I294 (gfint_1[8:8], choice_1, i_1r0[8:8]);
  AND2 I295 (gfint_1[9:9], choice_1, i_1r0[9:9]);
  AND2 I296 (gfint_1[10:10], choice_1, i_1r0[10:10]);
  AND2 I297 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I298 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I299 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I300 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AND2 I301 (gfint_2[4:4], choice_2, i_2r0[4:4]);
  AND2 I302 (gfint_2[5:5], choice_2, i_2r0[5:5]);
  AND2 I303 (gfint_2[6:6], choice_2, i_2r0[6:6]);
  AND2 I304 (gfint_2[7:7], choice_2, i_2r0[7:7]);
  AND2 I305 (gfint_2[8:8], choice_2, i_2r0[8:8]);
  AND2 I306 (gfint_2[9:9], choice_2, i_2r0[9:9]);
  AND2 I307 (gfint_2[10:10], choice_2, i_2r0[10:10]);
  AND2 I308 (gfint_3[0:0], choice_3, i_3r0[0:0]);
  AND2 I309 (gfint_3[1:1], choice_3, i_3r0[1:1]);
  AND2 I310 (gfint_3[2:2], choice_3, i_3r0[2:2]);
  AND2 I311 (gfint_3[3:3], choice_3, i_3r0[3:3]);
  AND2 I312 (gfint_3[4:4], choice_3, i_3r0[4:4]);
  AND2 I313 (gfint_3[5:5], choice_3, i_3r0[5:5]);
  AND2 I314 (gfint_3[6:6], choice_3, i_3r0[6:6]);
  AND2 I315 (gfint_3[7:7], choice_3, i_3r0[7:7]);
  AND2 I316 (gfint_3[8:8], choice_3, i_3r0[8:8]);
  AND2 I317 (gfint_3[9:9], choice_3, i_3r0[9:9]);
  AND2 I318 (gfint_3[10:10], choice_3, i_3r0[10:10]);
  AND2 I319 (gfint_4[0:0], choice_4, i_4r0[0:0]);
  AND2 I320 (gfint_4[1:1], choice_4, i_4r0[1:1]);
  AND2 I321 (gfint_4[2:2], choice_4, i_4r0[2:2]);
  AND2 I322 (gfint_4[3:3], choice_4, i_4r0[3:3]);
  AND2 I323 (gfint_4[4:4], choice_4, i_4r0[4:4]);
  AND2 I324 (gfint_4[5:5], choice_4, i_4r0[5:5]);
  AND2 I325 (gfint_4[6:6], choice_4, i_4r0[6:6]);
  AND2 I326 (gfint_4[7:7], choice_4, i_4r0[7:7]);
  AND2 I327 (gfint_4[8:8], choice_4, i_4r0[8:8]);
  AND2 I328 (gfint_4[9:9], choice_4, i_4r0[9:9]);
  AND2 I329 (gfint_4[10:10], choice_4, i_4r0[10:10]);
  AND2 I330 (gfint_5[0:0], choice_5, i_5r0[0:0]);
  AND2 I331 (gfint_5[1:1], choice_5, i_5r0[1:1]);
  AND2 I332 (gfint_5[2:2], choice_5, i_5r0[2:2]);
  AND2 I333 (gfint_5[3:3], choice_5, i_5r0[3:3]);
  AND2 I334 (gfint_5[4:4], choice_5, i_5r0[4:4]);
  AND2 I335 (gfint_5[5:5], choice_5, i_5r0[5:5]);
  AND2 I336 (gfint_5[6:6], choice_5, i_5r0[6:6]);
  AND2 I337 (gfint_5[7:7], choice_5, i_5r0[7:7]);
  AND2 I338 (gfint_5[8:8], choice_5, i_5r0[8:8]);
  AND2 I339 (gfint_5[9:9], choice_5, i_5r0[9:9]);
  AND2 I340 (gfint_5[10:10], choice_5, i_5r0[10:10]);
  AND2 I341 (gfint_6[0:0], choice_6, i_6r0[0:0]);
  AND2 I342 (gfint_6[1:1], choice_6, i_6r0[1:1]);
  AND2 I343 (gfint_6[2:2], choice_6, i_6r0[2:2]);
  AND2 I344 (gfint_6[3:3], choice_6, i_6r0[3:3]);
  AND2 I345 (gfint_6[4:4], choice_6, i_6r0[4:4]);
  AND2 I346 (gfint_6[5:5], choice_6, i_6r0[5:5]);
  AND2 I347 (gfint_6[6:6], choice_6, i_6r0[6:6]);
  AND2 I348 (gfint_6[7:7], choice_6, i_6r0[7:7]);
  AND2 I349 (gfint_6[8:8], choice_6, i_6r0[8:8]);
  AND2 I350 (gfint_6[9:9], choice_6, i_6r0[9:9]);
  AND2 I351 (gfint_6[10:10], choice_6, i_6r0[10:10]);
  AND2 I352 (gfint_7[0:0], choice_7, i_7r0[0:0]);
  AND2 I353 (gfint_7[1:1], choice_7, i_7r0[1:1]);
  AND2 I354 (gfint_7[2:2], choice_7, i_7r0[2:2]);
  AND2 I355 (gfint_7[3:3], choice_7, i_7r0[3:3]);
  AND2 I356 (gfint_7[4:4], choice_7, i_7r0[4:4]);
  AND2 I357 (gfint_7[5:5], choice_7, i_7r0[5:5]);
  AND2 I358 (gfint_7[6:6], choice_7, i_7r0[6:6]);
  AND2 I359 (gfint_7[7:7], choice_7, i_7r0[7:7]);
  AND2 I360 (gfint_7[8:8], choice_7, i_7r0[8:8]);
  AND2 I361 (gfint_7[9:9], choice_7, i_7r0[9:9]);
  AND2 I362 (gfint_7[10:10], choice_7, i_7r0[10:10]);
  AND2 I363 (gfint_8[0:0], choice_8, i_8r0[0:0]);
  AND2 I364 (gfint_8[1:1], choice_8, i_8r0[1:1]);
  AND2 I365 (gfint_8[2:2], choice_8, i_8r0[2:2]);
  AND2 I366 (gfint_8[3:3], choice_8, i_8r0[3:3]);
  AND2 I367 (gfint_8[4:4], choice_8, i_8r0[4:4]);
  AND2 I368 (gfint_8[5:5], choice_8, i_8r0[5:5]);
  AND2 I369 (gfint_8[6:6], choice_8, i_8r0[6:6]);
  AND2 I370 (gfint_8[7:7], choice_8, i_8r0[7:7]);
  AND2 I371 (gfint_8[8:8], choice_8, i_8r0[8:8]);
  AND2 I372 (gfint_8[9:9], choice_8, i_8r0[9:9]);
  AND2 I373 (gfint_8[10:10], choice_8, i_8r0[10:10]);
  AND2 I374 (gfint_9[0:0], choice_9, i_9r0[0:0]);
  AND2 I375 (gfint_9[1:1], choice_9, i_9r0[1:1]);
  AND2 I376 (gfint_9[2:2], choice_9, i_9r0[2:2]);
  AND2 I377 (gfint_9[3:3], choice_9, i_9r0[3:3]);
  AND2 I378 (gfint_9[4:4], choice_9, i_9r0[4:4]);
  AND2 I379 (gfint_9[5:5], choice_9, i_9r0[5:5]);
  AND2 I380 (gfint_9[6:6], choice_9, i_9r0[6:6]);
  AND2 I381 (gfint_9[7:7], choice_9, i_9r0[7:7]);
  AND2 I382 (gfint_9[8:8], choice_9, i_9r0[8:8]);
  AND2 I383 (gfint_9[9:9], choice_9, i_9r0[9:9]);
  AND2 I384 (gfint_9[10:10], choice_9, i_9r0[10:10]);
  AND2 I385 (gfint_10[0:0], choice_10, i_10r0[0:0]);
  AND2 I386 (gfint_10[1:1], choice_10, i_10r0[1:1]);
  AND2 I387 (gfint_10[2:2], choice_10, i_10r0[2:2]);
  AND2 I388 (gfint_10[3:3], choice_10, i_10r0[3:3]);
  AND2 I389 (gfint_10[4:4], choice_10, i_10r0[4:4]);
  AND2 I390 (gfint_10[5:5], choice_10, i_10r0[5:5]);
  AND2 I391 (gfint_10[6:6], choice_10, i_10r0[6:6]);
  AND2 I392 (gfint_10[7:7], choice_10, i_10r0[7:7]);
  AND2 I393 (gfint_10[8:8], choice_10, i_10r0[8:8]);
  AND2 I394 (gfint_10[9:9], choice_10, i_10r0[9:9]);
  AND2 I395 (gfint_10[10:10], choice_10, i_10r0[10:10]);
  OR2 I396 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I397 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I398 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I399 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I400 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I401 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I402 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I403 (comp0_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I404 (comp0_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I405 (comp0_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I406 (comp0_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  C3 I407 (simp3221_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I408 (simp3221_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I409 (simp3221_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C2 I410 (simp3221_0[3:3], comp0_0[9:9], comp0_0[10:10]);
  C3 I411 (simp3222_0[0:0], simp3221_0[0:0], simp3221_0[1:1], simp3221_0[2:2]);
  BUFF I412 (simp3222_0[1:1], simp3221_0[3:3]);
  C2 I413 (icomp_0, simp3222_0[0:0], simp3222_0[1:1]);
  OR2 I414 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I415 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I416 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I417 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I418 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I419 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I420 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  OR2 I421 (comp1_0[7:7], i_1r0[7:7], i_1r1[7:7]);
  OR2 I422 (comp1_0[8:8], i_1r0[8:8], i_1r1[8:8]);
  OR2 I423 (comp1_0[9:9], i_1r0[9:9], i_1r1[9:9]);
  OR2 I424 (comp1_0[10:10], i_1r0[10:10], i_1r1[10:10]);
  C3 I425 (simp3351_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I426 (simp3351_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  C3 I427 (simp3351_0[2:2], comp1_0[6:6], comp1_0[7:7], comp1_0[8:8]);
  C2 I428 (simp3351_0[3:3], comp1_0[9:9], comp1_0[10:10]);
  C3 I429 (simp3352_0[0:0], simp3351_0[0:0], simp3351_0[1:1], simp3351_0[2:2]);
  BUFF I430 (simp3352_0[1:1], simp3351_0[3:3]);
  C2 I431 (icomp_1, simp3352_0[0:0], simp3352_0[1:1]);
  OR2 I432 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I433 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I434 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2 I435 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  OR2 I436 (comp2_0[4:4], i_2r0[4:4], i_2r1[4:4]);
  OR2 I437 (comp2_0[5:5], i_2r0[5:5], i_2r1[5:5]);
  OR2 I438 (comp2_0[6:6], i_2r0[6:6], i_2r1[6:6]);
  OR2 I439 (comp2_0[7:7], i_2r0[7:7], i_2r1[7:7]);
  OR2 I440 (comp2_0[8:8], i_2r0[8:8], i_2r1[8:8]);
  OR2 I441 (comp2_0[9:9], i_2r0[9:9], i_2r1[9:9]);
  OR2 I442 (comp2_0[10:10], i_2r0[10:10], i_2r1[10:10]);
  C3 I443 (simp3481_0[0:0], comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C3 I444 (simp3481_0[1:1], comp2_0[3:3], comp2_0[4:4], comp2_0[5:5]);
  C3 I445 (simp3481_0[2:2], comp2_0[6:6], comp2_0[7:7], comp2_0[8:8]);
  C2 I446 (simp3481_0[3:3], comp2_0[9:9], comp2_0[10:10]);
  C3 I447 (simp3482_0[0:0], simp3481_0[0:0], simp3481_0[1:1], simp3481_0[2:2]);
  BUFF I448 (simp3482_0[1:1], simp3481_0[3:3]);
  C2 I449 (icomp_2, simp3482_0[0:0], simp3482_0[1:1]);
  OR2 I450 (comp3_0[0:0], i_3r0[0:0], i_3r1[0:0]);
  OR2 I451 (comp3_0[1:1], i_3r0[1:1], i_3r1[1:1]);
  OR2 I452 (comp3_0[2:2], i_3r0[2:2], i_3r1[2:2]);
  OR2 I453 (comp3_0[3:3], i_3r0[3:3], i_3r1[3:3]);
  OR2 I454 (comp3_0[4:4], i_3r0[4:4], i_3r1[4:4]);
  OR2 I455 (comp3_0[5:5], i_3r0[5:5], i_3r1[5:5]);
  OR2 I456 (comp3_0[6:6], i_3r0[6:6], i_3r1[6:6]);
  OR2 I457 (comp3_0[7:7], i_3r0[7:7], i_3r1[7:7]);
  OR2 I458 (comp3_0[8:8], i_3r0[8:8], i_3r1[8:8]);
  OR2 I459 (comp3_0[9:9], i_3r0[9:9], i_3r1[9:9]);
  OR2 I460 (comp3_0[10:10], i_3r0[10:10], i_3r1[10:10]);
  C3 I461 (simp3611_0[0:0], comp3_0[0:0], comp3_0[1:1], comp3_0[2:2]);
  C3 I462 (simp3611_0[1:1], comp3_0[3:3], comp3_0[4:4], comp3_0[5:5]);
  C3 I463 (simp3611_0[2:2], comp3_0[6:6], comp3_0[7:7], comp3_0[8:8]);
  C2 I464 (simp3611_0[3:3], comp3_0[9:9], comp3_0[10:10]);
  C3 I465 (simp3612_0[0:0], simp3611_0[0:0], simp3611_0[1:1], simp3611_0[2:2]);
  BUFF I466 (simp3612_0[1:1], simp3611_0[3:3]);
  C2 I467 (icomp_3, simp3612_0[0:0], simp3612_0[1:1]);
  OR2 I468 (comp4_0[0:0], i_4r0[0:0], i_4r1[0:0]);
  OR2 I469 (comp4_0[1:1], i_4r0[1:1], i_4r1[1:1]);
  OR2 I470 (comp4_0[2:2], i_4r0[2:2], i_4r1[2:2]);
  OR2 I471 (comp4_0[3:3], i_4r0[3:3], i_4r1[3:3]);
  OR2 I472 (comp4_0[4:4], i_4r0[4:4], i_4r1[4:4]);
  OR2 I473 (comp4_0[5:5], i_4r0[5:5], i_4r1[5:5]);
  OR2 I474 (comp4_0[6:6], i_4r0[6:6], i_4r1[6:6]);
  OR2 I475 (comp4_0[7:7], i_4r0[7:7], i_4r1[7:7]);
  OR2 I476 (comp4_0[8:8], i_4r0[8:8], i_4r1[8:8]);
  OR2 I477 (comp4_0[9:9], i_4r0[9:9], i_4r1[9:9]);
  OR2 I478 (comp4_0[10:10], i_4r0[10:10], i_4r1[10:10]);
  C3 I479 (simp3741_0[0:0], comp4_0[0:0], comp4_0[1:1], comp4_0[2:2]);
  C3 I480 (simp3741_0[1:1], comp4_0[3:3], comp4_0[4:4], comp4_0[5:5]);
  C3 I481 (simp3741_0[2:2], comp4_0[6:6], comp4_0[7:7], comp4_0[8:8]);
  C2 I482 (simp3741_0[3:3], comp4_0[9:9], comp4_0[10:10]);
  C3 I483 (simp3742_0[0:0], simp3741_0[0:0], simp3741_0[1:1], simp3741_0[2:2]);
  BUFF I484 (simp3742_0[1:1], simp3741_0[3:3]);
  C2 I485 (icomp_4, simp3742_0[0:0], simp3742_0[1:1]);
  OR2 I486 (comp5_0[0:0], i_5r0[0:0], i_5r1[0:0]);
  OR2 I487 (comp5_0[1:1], i_5r0[1:1], i_5r1[1:1]);
  OR2 I488 (comp5_0[2:2], i_5r0[2:2], i_5r1[2:2]);
  OR2 I489 (comp5_0[3:3], i_5r0[3:3], i_5r1[3:3]);
  OR2 I490 (comp5_0[4:4], i_5r0[4:4], i_5r1[4:4]);
  OR2 I491 (comp5_0[5:5], i_5r0[5:5], i_5r1[5:5]);
  OR2 I492 (comp5_0[6:6], i_5r0[6:6], i_5r1[6:6]);
  OR2 I493 (comp5_0[7:7], i_5r0[7:7], i_5r1[7:7]);
  OR2 I494 (comp5_0[8:8], i_5r0[8:8], i_5r1[8:8]);
  OR2 I495 (comp5_0[9:9], i_5r0[9:9], i_5r1[9:9]);
  OR2 I496 (comp5_0[10:10], i_5r0[10:10], i_5r1[10:10]);
  C3 I497 (simp3871_0[0:0], comp5_0[0:0], comp5_0[1:1], comp5_0[2:2]);
  C3 I498 (simp3871_0[1:1], comp5_0[3:3], comp5_0[4:4], comp5_0[5:5]);
  C3 I499 (simp3871_0[2:2], comp5_0[6:6], comp5_0[7:7], comp5_0[8:8]);
  C2 I500 (simp3871_0[3:3], comp5_0[9:9], comp5_0[10:10]);
  C3 I501 (simp3872_0[0:0], simp3871_0[0:0], simp3871_0[1:1], simp3871_0[2:2]);
  BUFF I502 (simp3872_0[1:1], simp3871_0[3:3]);
  C2 I503 (icomp_5, simp3872_0[0:0], simp3872_0[1:1]);
  OR2 I504 (comp6_0[0:0], i_6r0[0:0], i_6r1[0:0]);
  OR2 I505 (comp6_0[1:1], i_6r0[1:1], i_6r1[1:1]);
  OR2 I506 (comp6_0[2:2], i_6r0[2:2], i_6r1[2:2]);
  OR2 I507 (comp6_0[3:3], i_6r0[3:3], i_6r1[3:3]);
  OR2 I508 (comp6_0[4:4], i_6r0[4:4], i_6r1[4:4]);
  OR2 I509 (comp6_0[5:5], i_6r0[5:5], i_6r1[5:5]);
  OR2 I510 (comp6_0[6:6], i_6r0[6:6], i_6r1[6:6]);
  OR2 I511 (comp6_0[7:7], i_6r0[7:7], i_6r1[7:7]);
  OR2 I512 (comp6_0[8:8], i_6r0[8:8], i_6r1[8:8]);
  OR2 I513 (comp6_0[9:9], i_6r0[9:9], i_6r1[9:9]);
  OR2 I514 (comp6_0[10:10], i_6r0[10:10], i_6r1[10:10]);
  C3 I515 (simp4001_0[0:0], comp6_0[0:0], comp6_0[1:1], comp6_0[2:2]);
  C3 I516 (simp4001_0[1:1], comp6_0[3:3], comp6_0[4:4], comp6_0[5:5]);
  C3 I517 (simp4001_0[2:2], comp6_0[6:6], comp6_0[7:7], comp6_0[8:8]);
  C2 I518 (simp4001_0[3:3], comp6_0[9:9], comp6_0[10:10]);
  C3 I519 (simp4002_0[0:0], simp4001_0[0:0], simp4001_0[1:1], simp4001_0[2:2]);
  BUFF I520 (simp4002_0[1:1], simp4001_0[3:3]);
  C2 I521 (icomp_6, simp4002_0[0:0], simp4002_0[1:1]);
  OR2 I522 (comp7_0[0:0], i_7r0[0:0], i_7r1[0:0]);
  OR2 I523 (comp7_0[1:1], i_7r0[1:1], i_7r1[1:1]);
  OR2 I524 (comp7_0[2:2], i_7r0[2:2], i_7r1[2:2]);
  OR2 I525 (comp7_0[3:3], i_7r0[3:3], i_7r1[3:3]);
  OR2 I526 (comp7_0[4:4], i_7r0[4:4], i_7r1[4:4]);
  OR2 I527 (comp7_0[5:5], i_7r0[5:5], i_7r1[5:5]);
  OR2 I528 (comp7_0[6:6], i_7r0[6:6], i_7r1[6:6]);
  OR2 I529 (comp7_0[7:7], i_7r0[7:7], i_7r1[7:7]);
  OR2 I530 (comp7_0[8:8], i_7r0[8:8], i_7r1[8:8]);
  OR2 I531 (comp7_0[9:9], i_7r0[9:9], i_7r1[9:9]);
  OR2 I532 (comp7_0[10:10], i_7r0[10:10], i_7r1[10:10]);
  C3 I533 (simp4131_0[0:0], comp7_0[0:0], comp7_0[1:1], comp7_0[2:2]);
  C3 I534 (simp4131_0[1:1], comp7_0[3:3], comp7_0[4:4], comp7_0[5:5]);
  C3 I535 (simp4131_0[2:2], comp7_0[6:6], comp7_0[7:7], comp7_0[8:8]);
  C2 I536 (simp4131_0[3:3], comp7_0[9:9], comp7_0[10:10]);
  C3 I537 (simp4132_0[0:0], simp4131_0[0:0], simp4131_0[1:1], simp4131_0[2:2]);
  BUFF I538 (simp4132_0[1:1], simp4131_0[3:3]);
  C2 I539 (icomp_7, simp4132_0[0:0], simp4132_0[1:1]);
  OR2 I540 (comp8_0[0:0], i_8r0[0:0], i_8r1[0:0]);
  OR2 I541 (comp8_0[1:1], i_8r0[1:1], i_8r1[1:1]);
  OR2 I542 (comp8_0[2:2], i_8r0[2:2], i_8r1[2:2]);
  OR2 I543 (comp8_0[3:3], i_8r0[3:3], i_8r1[3:3]);
  OR2 I544 (comp8_0[4:4], i_8r0[4:4], i_8r1[4:4]);
  OR2 I545 (comp8_0[5:5], i_8r0[5:5], i_8r1[5:5]);
  OR2 I546 (comp8_0[6:6], i_8r0[6:6], i_8r1[6:6]);
  OR2 I547 (comp8_0[7:7], i_8r0[7:7], i_8r1[7:7]);
  OR2 I548 (comp8_0[8:8], i_8r0[8:8], i_8r1[8:8]);
  OR2 I549 (comp8_0[9:9], i_8r0[9:9], i_8r1[9:9]);
  OR2 I550 (comp8_0[10:10], i_8r0[10:10], i_8r1[10:10]);
  C3 I551 (simp4261_0[0:0], comp8_0[0:0], comp8_0[1:1], comp8_0[2:2]);
  C3 I552 (simp4261_0[1:1], comp8_0[3:3], comp8_0[4:4], comp8_0[5:5]);
  C3 I553 (simp4261_0[2:2], comp8_0[6:6], comp8_0[7:7], comp8_0[8:8]);
  C2 I554 (simp4261_0[3:3], comp8_0[9:9], comp8_0[10:10]);
  C3 I555 (simp4262_0[0:0], simp4261_0[0:0], simp4261_0[1:1], simp4261_0[2:2]);
  BUFF I556 (simp4262_0[1:1], simp4261_0[3:3]);
  C2 I557 (icomp_8, simp4262_0[0:0], simp4262_0[1:1]);
  OR2 I558 (comp9_0[0:0], i_9r0[0:0], i_9r1[0:0]);
  OR2 I559 (comp9_0[1:1], i_9r0[1:1], i_9r1[1:1]);
  OR2 I560 (comp9_0[2:2], i_9r0[2:2], i_9r1[2:2]);
  OR2 I561 (comp9_0[3:3], i_9r0[3:3], i_9r1[3:3]);
  OR2 I562 (comp9_0[4:4], i_9r0[4:4], i_9r1[4:4]);
  OR2 I563 (comp9_0[5:5], i_9r0[5:5], i_9r1[5:5]);
  OR2 I564 (comp9_0[6:6], i_9r0[6:6], i_9r1[6:6]);
  OR2 I565 (comp9_0[7:7], i_9r0[7:7], i_9r1[7:7]);
  OR2 I566 (comp9_0[8:8], i_9r0[8:8], i_9r1[8:8]);
  OR2 I567 (comp9_0[9:9], i_9r0[9:9], i_9r1[9:9]);
  OR2 I568 (comp9_0[10:10], i_9r0[10:10], i_9r1[10:10]);
  C3 I569 (simp4391_0[0:0], comp9_0[0:0], comp9_0[1:1], comp9_0[2:2]);
  C3 I570 (simp4391_0[1:1], comp9_0[3:3], comp9_0[4:4], comp9_0[5:5]);
  C3 I571 (simp4391_0[2:2], comp9_0[6:6], comp9_0[7:7], comp9_0[8:8]);
  C2 I572 (simp4391_0[3:3], comp9_0[9:9], comp9_0[10:10]);
  C3 I573 (simp4392_0[0:0], simp4391_0[0:0], simp4391_0[1:1], simp4391_0[2:2]);
  BUFF I574 (simp4392_0[1:1], simp4391_0[3:3]);
  C2 I575 (icomp_9, simp4392_0[0:0], simp4392_0[1:1]);
  OR2 I576 (comp10_0[0:0], i_10r0[0:0], i_10r1[0:0]);
  OR2 I577 (comp10_0[1:1], i_10r0[1:1], i_10r1[1:1]);
  OR2 I578 (comp10_0[2:2], i_10r0[2:2], i_10r1[2:2]);
  OR2 I579 (comp10_0[3:3], i_10r0[3:3], i_10r1[3:3]);
  OR2 I580 (comp10_0[4:4], i_10r0[4:4], i_10r1[4:4]);
  OR2 I581 (comp10_0[5:5], i_10r0[5:5], i_10r1[5:5]);
  OR2 I582 (comp10_0[6:6], i_10r0[6:6], i_10r1[6:6]);
  OR2 I583 (comp10_0[7:7], i_10r0[7:7], i_10r1[7:7]);
  OR2 I584 (comp10_0[8:8], i_10r0[8:8], i_10r1[8:8]);
  OR2 I585 (comp10_0[9:9], i_10r0[9:9], i_10r1[9:9]);
  OR2 I586 (comp10_0[10:10], i_10r0[10:10], i_10r1[10:10]);
  C3 I587 (simp4521_0[0:0], comp10_0[0:0], comp10_0[1:1], comp10_0[2:2]);
  C3 I588 (simp4521_0[1:1], comp10_0[3:3], comp10_0[4:4], comp10_0[5:5]);
  C3 I589 (simp4521_0[2:2], comp10_0[6:6], comp10_0[7:7], comp10_0[8:8]);
  C2 I590 (simp4521_0[3:3], comp10_0[9:9], comp10_0[10:10]);
  C3 I591 (simp4522_0[0:0], simp4521_0[0:0], simp4521_0[1:1], simp4521_0[2:2]);
  BUFF I592 (simp4522_0[1:1], simp4521_0[3:3]);
  C2 I593 (icomp_10, simp4522_0[0:0], simp4522_0[1:1]);
  C2R I594 (choice_0, icomp_0, nchosen_0, reset);
  C2R I595 (choice_1, icomp_1, nchosen_0, reset);
  C2R I596 (choice_2, icomp_2, nchosen_0, reset);
  C2R I597 (choice_3, icomp_3, nchosen_0, reset);
  C2R I598 (choice_4, icomp_4, nchosen_0, reset);
  C2R I599 (choice_5, icomp_5, nchosen_0, reset);
  C2R I600 (choice_6, icomp_6, nchosen_0, reset);
  C2R I601 (choice_7, icomp_7, nchosen_0, reset);
  C2R I602 (choice_8, icomp_8, nchosen_0, reset);
  C2R I603 (choice_9, icomp_9, nchosen_0, reset);
  C2R I604 (choice_10, icomp_10, nchosen_0, reset);
  NOR3 I605 (simp4641_0[0:0], choice_0, choice_1, choice_2);
  NOR3 I606 (simp4641_0[1:1], choice_3, choice_4, choice_5);
  NOR3 I607 (simp4641_0[2:2], choice_6, choice_7, choice_8);
  NOR2 I608 (simp4641_0[3:3], choice_9, choice_10);
  NAND3 I609 (simp4642_0[0:0], simp4641_0[0:0], simp4641_0[1:1], simp4641_0[2:2]);
  INV I610 (simp4642_0[1:1], simp4641_0[3:3]);
  OR2 I611 (anychoice_0, simp4642_0[0:0], simp4642_0[1:1]);
  NOR2 I612 (nchosen_0, anychoice_0, o_0a);
  C2R I613 (i_0a, choice_0, o_0a, reset);
  C2R I614 (i_1a, choice_1, o_0a, reset);
  C2R I615 (i_2a, choice_2, o_0a, reset);
  C2R I616 (i_3a, choice_3, o_0a, reset);
  C2R I617 (i_4a, choice_4, o_0a, reset);
  C2R I618 (i_5a, choice_5, o_0a, reset);
  C2R I619 (i_6a, choice_6, o_0a, reset);
  C2R I620 (i_7a, choice_7, o_0a, reset);
  C2R I621 (i_8a, choice_8, o_0a, reset);
  C2R I622 (i_9a, choice_9, o_0a, reset);
  C2R I623 (i_10a, choice_10, o_0a, reset);
endmodule

// tkj11m0_11 TeakJ [Many [0,11],One 11]
module tkj11m0_11 (i_0r, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  input [10:0] i_1r0;
  input [10:0] i_1r1;
  output i_1a;
  output [10:0] o_0r0;
  output [10:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [10:0] joinf_0;
  wire [10:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_1r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_1r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_1r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_1r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_1r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_1r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_1r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_1r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_1r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_1r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_1r0[10:10]);
  BUFF I11 (joint_0[0:0], i_1r1[0:0]);
  BUFF I12 (joint_0[1:1], i_1r1[1:1]);
  BUFF I13 (joint_0[2:2], i_1r1[2:2]);
  BUFF I14 (joint_0[3:3], i_1r1[3:3]);
  BUFF I15 (joint_0[4:4], i_1r1[4:4]);
  BUFF I16 (joint_0[5:5], i_1r1[5:5]);
  BUFF I17 (joint_0[6:6], i_1r1[6:6]);
  BUFF I18 (joint_0[7:7], i_1r1[7:7]);
  BUFF I19 (joint_0[8:8], i_1r1[8:8]);
  BUFF I20 (joint_0[9:9], i_1r1[9:9]);
  BUFF I21 (joint_0[10:10], i_1r1[10:10]);
  BUFF I22 (icomplete_0, i_0r);
  C2 I23 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I24 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I25 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I26 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I27 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I28 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I29 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I30 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I31 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I32 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I33 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I34 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I35 (o_0r1[1:1], joint_0[1:1]);
  BUFF I36 (o_0r1[2:2], joint_0[2:2]);
  BUFF I37 (o_0r1[3:3], joint_0[3:3]);
  BUFF I38 (o_0r1[4:4], joint_0[4:4]);
  BUFF I39 (o_0r1[5:5], joint_0[5:5]);
  BUFF I40 (o_0r1[6:6], joint_0[6:6]);
  BUFF I41 (o_0r1[7:7], joint_0[7:7]);
  BUFF I42 (o_0r1[8:8], joint_0[8:8]);
  BUFF I43 (o_0r1[9:9], joint_0[9:9]);
  BUFF I44 (o_0r1[10:10], joint_0[10:10]);
  BUFF I45 (i_0a, o_0a);
  BUFF I46 (i_1a, o_0a);
endmodule

// tks11_o0w11_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0_20o0w0_40o0w0_80o0w0_100o0w0_200o0w0_400o0w0 TeakS (0+:11
//   ) [([Imp 1 0],0),([Imp 2 0],0),([Imp 4 0],0),([Imp 8 0],0),([Imp 16 0],0),([Imp 32 0],0),([Imp 64 0]
//   ,0),([Imp 128 0],0),([Imp 256 0],0),([Imp 512 0],0),([Imp 1024 0],0)] [One 11,Many [0,0,0,0,0,0,0,0,
//   0,0,0]]
module tks11_o0w11_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0_20o0w0_40o0w0_80o0w0_100o0w0_200o0w0_400o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, o_5r, o_5a, o_6r, o_6a, o_7r, o_7a, o_8r, o_8a, o_9r, o_9a, o_10r, o_10a, reset);
  input [10:0] i_0r0;
  input [10:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  output o_7r;
  input o_7a;
  output o_8r;
  input o_8a;
  output o_9r;
  input o_9a;
  output o_10r;
  input o_10a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire sel_4;
  wire sel_5;
  wire sel_6;
  wire sel_7;
  wire sel_8;
  wire sel_9;
  wire sel_10;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire gsel_4;
  wire gsel_5;
  wire gsel_6;
  wire gsel_7;
  wire gsel_8;
  wire gsel_9;
  wire gsel_10;
  wire oack_0;
  wire match0_0;
  wire [3:0] simp261_0;
  wire [1:0] simp262_0;
  wire match1_0;
  wire [3:0] simp291_0;
  wire [1:0] simp292_0;
  wire match2_0;
  wire [3:0] simp321_0;
  wire [1:0] simp322_0;
  wire match3_0;
  wire [3:0] simp351_0;
  wire [1:0] simp352_0;
  wire match4_0;
  wire [3:0] simp381_0;
  wire [1:0] simp382_0;
  wire match5_0;
  wire [3:0] simp411_0;
  wire [1:0] simp412_0;
  wire match6_0;
  wire [3:0] simp441_0;
  wire [1:0] simp442_0;
  wire match7_0;
  wire [3:0] simp471_0;
  wire [1:0] simp472_0;
  wire match8_0;
  wire [3:0] simp501_0;
  wire [1:0] simp502_0;
  wire match9_0;
  wire [3:0] simp531_0;
  wire [1:0] simp532_0;
  wire match10_0;
  wire [3:0] simp561_0;
  wire [1:0] simp562_0;
  wire [10:0] comp_0;
  wire [3:0] simp801_0;
  wire [1:0] simp802_0;
  wire [3:0] simp921_0;
  wire [1:0] simp922_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (simp261_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I2 (simp261_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I3 (simp261_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C2 I4 (simp261_0[3:3], i_0r0[9:9], i_0r0[10:10]);
  C3 I5 (simp262_0[0:0], simp261_0[0:0], simp261_0[1:1], simp261_0[2:2]);
  BUFF I6 (simp262_0[1:1], simp261_0[3:3]);
  C2 I7 (match0_0, simp262_0[0:0], simp262_0[1:1]);
  BUFF I8 (sel_1, match1_0);
  C3 I9 (simp291_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I10 (simp291_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I11 (simp291_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C2 I12 (simp291_0[3:3], i_0r0[9:9], i_0r0[10:10]);
  C3 I13 (simp292_0[0:0], simp291_0[0:0], simp291_0[1:1], simp291_0[2:2]);
  BUFF I14 (simp292_0[1:1], simp291_0[3:3]);
  C2 I15 (match1_0, simp292_0[0:0], simp292_0[1:1]);
  BUFF I16 (sel_2, match2_0);
  C3 I17 (simp321_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I18 (simp321_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I19 (simp321_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C2 I20 (simp321_0[3:3], i_0r0[9:9], i_0r0[10:10]);
  C3 I21 (simp322_0[0:0], simp321_0[0:0], simp321_0[1:1], simp321_0[2:2]);
  BUFF I22 (simp322_0[1:1], simp321_0[3:3]);
  C2 I23 (match2_0, simp322_0[0:0], simp322_0[1:1]);
  BUFF I24 (sel_3, match3_0);
  C3 I25 (simp351_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I26 (simp351_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I27 (simp351_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C2 I28 (simp351_0[3:3], i_0r0[9:9], i_0r0[10:10]);
  C3 I29 (simp352_0[0:0], simp351_0[0:0], simp351_0[1:1], simp351_0[2:2]);
  BUFF I30 (simp352_0[1:1], simp351_0[3:3]);
  C2 I31 (match3_0, simp352_0[0:0], simp352_0[1:1]);
  BUFF I32 (sel_4, match4_0);
  C3 I33 (simp381_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I34 (simp381_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C3 I35 (simp381_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C2 I36 (simp381_0[3:3], i_0r0[9:9], i_0r0[10:10]);
  C3 I37 (simp382_0[0:0], simp381_0[0:0], simp381_0[1:1], simp381_0[2:2]);
  BUFF I38 (simp382_0[1:1], simp381_0[3:3]);
  C2 I39 (match4_0, simp382_0[0:0], simp382_0[1:1]);
  BUFF I40 (sel_5, match5_0);
  C3 I41 (simp411_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I42 (simp411_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C3 I43 (simp411_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C2 I44 (simp411_0[3:3], i_0r0[9:9], i_0r0[10:10]);
  C3 I45 (simp412_0[0:0], simp411_0[0:0], simp411_0[1:1], simp411_0[2:2]);
  BUFF I46 (simp412_0[1:1], simp411_0[3:3]);
  C2 I47 (match5_0, simp412_0[0:0], simp412_0[1:1]);
  BUFF I48 (sel_6, match6_0);
  C3 I49 (simp441_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I50 (simp441_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I51 (simp441_0[2:2], i_0r1[6:6], i_0r0[7:7], i_0r0[8:8]);
  C2 I52 (simp441_0[3:3], i_0r0[9:9], i_0r0[10:10]);
  C3 I53 (simp442_0[0:0], simp441_0[0:0], simp441_0[1:1], simp441_0[2:2]);
  BUFF I54 (simp442_0[1:1], simp441_0[3:3]);
  C2 I55 (match6_0, simp442_0[0:0], simp442_0[1:1]);
  BUFF I56 (sel_7, match7_0);
  C3 I57 (simp471_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I58 (simp471_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I59 (simp471_0[2:2], i_0r0[6:6], i_0r1[7:7], i_0r0[8:8]);
  C2 I60 (simp471_0[3:3], i_0r0[9:9], i_0r0[10:10]);
  C3 I61 (simp472_0[0:0], simp471_0[0:0], simp471_0[1:1], simp471_0[2:2]);
  BUFF I62 (simp472_0[1:1], simp471_0[3:3]);
  C2 I63 (match7_0, simp472_0[0:0], simp472_0[1:1]);
  BUFF I64 (sel_8, match8_0);
  C3 I65 (simp501_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I66 (simp501_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I67 (simp501_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r1[8:8]);
  C2 I68 (simp501_0[3:3], i_0r0[9:9], i_0r0[10:10]);
  C3 I69 (simp502_0[0:0], simp501_0[0:0], simp501_0[1:1], simp501_0[2:2]);
  BUFF I70 (simp502_0[1:1], simp501_0[3:3]);
  C2 I71 (match8_0, simp502_0[0:0], simp502_0[1:1]);
  BUFF I72 (sel_9, match9_0);
  C3 I73 (simp531_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I74 (simp531_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I75 (simp531_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C2 I76 (simp531_0[3:3], i_0r1[9:9], i_0r0[10:10]);
  C3 I77 (simp532_0[0:0], simp531_0[0:0], simp531_0[1:1], simp531_0[2:2]);
  BUFF I78 (simp532_0[1:1], simp531_0[3:3]);
  C2 I79 (match9_0, simp532_0[0:0], simp532_0[1:1]);
  BUFF I80 (sel_10, match10_0);
  C3 I81 (simp561_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I82 (simp561_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C3 I83 (simp561_0[2:2], i_0r0[6:6], i_0r0[7:7], i_0r0[8:8]);
  C2 I84 (simp561_0[3:3], i_0r0[9:9], i_0r1[10:10]);
  C3 I85 (simp562_0[0:0], simp561_0[0:0], simp561_0[1:1], simp561_0[2:2]);
  BUFF I86 (simp562_0[1:1], simp561_0[3:3]);
  C2 I87 (match10_0, simp562_0[0:0], simp562_0[1:1]);
  C2 I88 (gsel_0, sel_0, icomplete_0);
  C2 I89 (gsel_1, sel_1, icomplete_0);
  C2 I90 (gsel_2, sel_2, icomplete_0);
  C2 I91 (gsel_3, sel_3, icomplete_0);
  C2 I92 (gsel_4, sel_4, icomplete_0);
  C2 I93 (gsel_5, sel_5, icomplete_0);
  C2 I94 (gsel_6, sel_6, icomplete_0);
  C2 I95 (gsel_7, sel_7, icomplete_0);
  C2 I96 (gsel_8, sel_8, icomplete_0);
  C2 I97 (gsel_9, sel_9, icomplete_0);
  C2 I98 (gsel_10, sel_10, icomplete_0);
  OR2 I99 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I100 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I101 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I102 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I103 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I104 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I105 (comp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I106 (comp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I107 (comp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I108 (comp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I109 (comp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  C3 I110 (simp801_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I111 (simp801_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C3 I112 (simp801_0[2:2], comp_0[6:6], comp_0[7:7], comp_0[8:8]);
  C2 I113 (simp801_0[3:3], comp_0[9:9], comp_0[10:10]);
  C3 I114 (simp802_0[0:0], simp801_0[0:0], simp801_0[1:1], simp801_0[2:2]);
  BUFF I115 (simp802_0[1:1], simp801_0[3:3]);
  C2 I116 (icomplete_0, simp802_0[0:0], simp802_0[1:1]);
  BUFF I117 (o_0r, gsel_0);
  BUFF I118 (o_1r, gsel_1);
  BUFF I119 (o_2r, gsel_2);
  BUFF I120 (o_3r, gsel_3);
  BUFF I121 (o_4r, gsel_4);
  BUFF I122 (o_5r, gsel_5);
  BUFF I123 (o_6r, gsel_6);
  BUFF I124 (o_7r, gsel_7);
  BUFF I125 (o_8r, gsel_8);
  BUFF I126 (o_9r, gsel_9);
  BUFF I127 (o_10r, gsel_10);
  NOR3 I128 (simp921_0[0:0], o_0a, o_1a, o_2a);
  NOR3 I129 (simp921_0[1:1], o_3a, o_4a, o_5a);
  NOR3 I130 (simp921_0[2:2], o_6a, o_7a, o_8a);
  NOR2 I131 (simp921_0[3:3], o_9a, o_10a);
  NAND3 I132 (simp922_0[0:0], simp921_0[0:0], simp921_0[1:1], simp921_0[2:2]);
  INV I133 (simp922_0[1:1], simp921_0[3:3]);
  OR2 I134 (oack_0, simp922_0[0:0], simp922_0[1:1]);
  C2 I135 (i_0a, oack_0, icomplete_0);
endmodule

// tkj3m3_0 TeakJ [Many [3,0],One 3]
module tkj3m3_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [2:0] joinf_0;
  wire [2:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joint_0[0:0], i_0r1[0:0]);
  BUFF I4 (joint_0[1:1], i_0r1[1:1]);
  BUFF I5 (joint_0[2:2], i_0r1[2:2]);
  BUFF I6 (icomplete_0, i_1r);
  C2 I7 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I8 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I9 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I10 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I11 (o_0r1[1:1], joint_0[1:1]);
  BUFF I12 (o_0r1[2:2], joint_0[2:2]);
  BUFF I13 (i_0a, o_0a);
  BUFF I14 (i_1a, o_0a);
endmodule

// tkf4mo0w0_o0w4 TeakF [0,0] [One 4,Many [0,4]]
module tkf4mo0w0_o0w4 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [3:0] o_1r0;
  output [3:0] o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_1r0[0:0], i_0r0[0:0]);
  BUFF I3 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I4 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I5 (o_1r0[3:3], i_0r0[3:3]);
  BUFF I6 (o_1r1[0:0], i_0r1[0:0]);
  BUFF I7 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I8 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I9 (o_1r1[3:3], i_0r1[3:3]);
  BUFF I10 (o_0r, icomplete_0);
  C3 I11 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tkm11x4b TeakM [Many [4,4,4,4,4,4,4,4,4,4,4],One 4]
module tkm11x4b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, i_4r0, i_4r1, i_4a, i_5r0, i_5r1, i_5a, i_6r0, i_6r1, i_6a, i_7r0, i_7r1, i_7a, i_8r0, i_8r1, i_8a, i_9r0, i_9r1, i_9a, i_10r0, i_10r1, i_10a, o_0r0, o_0r1, o_0a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  input [3:0] i_1r0;
  input [3:0] i_1r1;
  output i_1a;
  input [3:0] i_2r0;
  input [3:0] i_2r1;
  output i_2a;
  input [3:0] i_3r0;
  input [3:0] i_3r1;
  output i_3a;
  input [3:0] i_4r0;
  input [3:0] i_4r1;
  output i_4a;
  input [3:0] i_5r0;
  input [3:0] i_5r1;
  output i_5a;
  input [3:0] i_6r0;
  input [3:0] i_6r1;
  output i_6a;
  input [3:0] i_7r0;
  input [3:0] i_7r1;
  output i_7a;
  input [3:0] i_8r0;
  input [3:0] i_8r1;
  output i_8a;
  input [3:0] i_9r0;
  input [3:0] i_9r1;
  output i_9a;
  input [3:0] i_10r0;
  input [3:0] i_10r1;
  output i_10a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  wire [3:0] gfint_0;
  wire [3:0] gfint_1;
  wire [3:0] gfint_2;
  wire [3:0] gfint_3;
  wire [3:0] gfint_4;
  wire [3:0] gfint_5;
  wire [3:0] gfint_6;
  wire [3:0] gfint_7;
  wire [3:0] gfint_8;
  wire [3:0] gfint_9;
  wire [3:0] gfint_10;
  wire [3:0] gtint_0;
  wire [3:0] gtint_1;
  wire [3:0] gtint_2;
  wire [3:0] gtint_3;
  wire [3:0] gtint_4;
  wire [3:0] gtint_5;
  wire [3:0] gtint_6;
  wire [3:0] gtint_7;
  wire [3:0] gtint_8;
  wire [3:0] gtint_9;
  wire [3:0] gtint_10;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire choice_4;
  wire choice_5;
  wire choice_6;
  wire choice_7;
  wire choice_8;
  wire choice_9;
  wire choice_10;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire icomp_3;
  wire icomp_4;
  wire icomp_5;
  wire icomp_6;
  wire icomp_7;
  wire icomp_8;
  wire icomp_9;
  wire icomp_10;
  wire nchosen_0;
  wire [3:0] simp461_0;
  wire [1:0] simp462_0;
  wire [3:0] simp471_0;
  wire [1:0] simp472_0;
  wire [3:0] simp481_0;
  wire [1:0] simp482_0;
  wire [3:0] simp491_0;
  wire [1:0] simp492_0;
  wire [3:0] simp501_0;
  wire [1:0] simp502_0;
  wire [3:0] simp511_0;
  wire [1:0] simp512_0;
  wire [3:0] simp521_0;
  wire [1:0] simp522_0;
  wire [3:0] simp531_0;
  wire [1:0] simp532_0;
  wire [3:0] comp0_0;
  wire [1:0] simp1471_0;
  wire [3:0] comp1_0;
  wire [1:0] simp1531_0;
  wire [3:0] comp2_0;
  wire [1:0] simp1591_0;
  wire [3:0] comp3_0;
  wire [1:0] simp1651_0;
  wire [3:0] comp4_0;
  wire [1:0] simp1711_0;
  wire [3:0] comp5_0;
  wire [1:0] simp1771_0;
  wire [3:0] comp6_0;
  wire [1:0] simp1831_0;
  wire [3:0] comp7_0;
  wire [1:0] simp1891_0;
  wire [3:0] comp8_0;
  wire [1:0] simp1951_0;
  wire [3:0] comp9_0;
  wire [1:0] simp2011_0;
  wire [3:0] comp10_0;
  wire [1:0] simp2071_0;
  wire [3:0] simp2191_0;
  wire [1:0] simp2192_0;
  NOR3 I0 (simp461_0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  NOR3 I1 (simp461_0[1:1], gfint_3[0:0], gfint_4[0:0], gfint_5[0:0]);
  NOR3 I2 (simp461_0[2:2], gfint_6[0:0], gfint_7[0:0], gfint_8[0:0]);
  NOR2 I3 (simp461_0[3:3], gfint_9[0:0], gfint_10[0:0]);
  NAND3 I4 (simp462_0[0:0], simp461_0[0:0], simp461_0[1:1], simp461_0[2:2]);
  INV I5 (simp462_0[1:1], simp461_0[3:3]);
  OR2 I6 (o_0r0[0:0], simp462_0[0:0], simp462_0[1:1]);
  NOR3 I7 (simp471_0[0:0], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  NOR3 I8 (simp471_0[1:1], gfint_3[1:1], gfint_4[1:1], gfint_5[1:1]);
  NOR3 I9 (simp471_0[2:2], gfint_6[1:1], gfint_7[1:1], gfint_8[1:1]);
  NOR2 I10 (simp471_0[3:3], gfint_9[1:1], gfint_10[1:1]);
  NAND3 I11 (simp472_0[0:0], simp471_0[0:0], simp471_0[1:1], simp471_0[2:2]);
  INV I12 (simp472_0[1:1], simp471_0[3:3]);
  OR2 I13 (o_0r0[1:1], simp472_0[0:0], simp472_0[1:1]);
  NOR3 I14 (simp481_0[0:0], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  NOR3 I15 (simp481_0[1:1], gfint_3[2:2], gfint_4[2:2], gfint_5[2:2]);
  NOR3 I16 (simp481_0[2:2], gfint_6[2:2], gfint_7[2:2], gfint_8[2:2]);
  NOR2 I17 (simp481_0[3:3], gfint_9[2:2], gfint_10[2:2]);
  NAND3 I18 (simp482_0[0:0], simp481_0[0:0], simp481_0[1:1], simp481_0[2:2]);
  INV I19 (simp482_0[1:1], simp481_0[3:3]);
  OR2 I20 (o_0r0[2:2], simp482_0[0:0], simp482_0[1:1]);
  NOR3 I21 (simp491_0[0:0], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  NOR3 I22 (simp491_0[1:1], gfint_3[3:3], gfint_4[3:3], gfint_5[3:3]);
  NOR3 I23 (simp491_0[2:2], gfint_6[3:3], gfint_7[3:3], gfint_8[3:3]);
  NOR2 I24 (simp491_0[3:3], gfint_9[3:3], gfint_10[3:3]);
  NAND3 I25 (simp492_0[0:0], simp491_0[0:0], simp491_0[1:1], simp491_0[2:2]);
  INV I26 (simp492_0[1:1], simp491_0[3:3]);
  OR2 I27 (o_0r0[3:3], simp492_0[0:0], simp492_0[1:1]);
  NOR3 I28 (simp501_0[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  NOR3 I29 (simp501_0[1:1], gtint_3[0:0], gtint_4[0:0], gtint_5[0:0]);
  NOR3 I30 (simp501_0[2:2], gtint_6[0:0], gtint_7[0:0], gtint_8[0:0]);
  NOR2 I31 (simp501_0[3:3], gtint_9[0:0], gtint_10[0:0]);
  NAND3 I32 (simp502_0[0:0], simp501_0[0:0], simp501_0[1:1], simp501_0[2:2]);
  INV I33 (simp502_0[1:1], simp501_0[3:3]);
  OR2 I34 (o_0r1[0:0], simp502_0[0:0], simp502_0[1:1]);
  NOR3 I35 (simp511_0[0:0], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  NOR3 I36 (simp511_0[1:1], gtint_3[1:1], gtint_4[1:1], gtint_5[1:1]);
  NOR3 I37 (simp511_0[2:2], gtint_6[1:1], gtint_7[1:1], gtint_8[1:1]);
  NOR2 I38 (simp511_0[3:3], gtint_9[1:1], gtint_10[1:1]);
  NAND3 I39 (simp512_0[0:0], simp511_0[0:0], simp511_0[1:1], simp511_0[2:2]);
  INV I40 (simp512_0[1:1], simp511_0[3:3]);
  OR2 I41 (o_0r1[1:1], simp512_0[0:0], simp512_0[1:1]);
  NOR3 I42 (simp521_0[0:0], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  NOR3 I43 (simp521_0[1:1], gtint_3[2:2], gtint_4[2:2], gtint_5[2:2]);
  NOR3 I44 (simp521_0[2:2], gtint_6[2:2], gtint_7[2:2], gtint_8[2:2]);
  NOR2 I45 (simp521_0[3:3], gtint_9[2:2], gtint_10[2:2]);
  NAND3 I46 (simp522_0[0:0], simp521_0[0:0], simp521_0[1:1], simp521_0[2:2]);
  INV I47 (simp522_0[1:1], simp521_0[3:3]);
  OR2 I48 (o_0r1[2:2], simp522_0[0:0], simp522_0[1:1]);
  NOR3 I49 (simp531_0[0:0], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  NOR3 I50 (simp531_0[1:1], gtint_3[3:3], gtint_4[3:3], gtint_5[3:3]);
  NOR3 I51 (simp531_0[2:2], gtint_6[3:3], gtint_7[3:3], gtint_8[3:3]);
  NOR2 I52 (simp531_0[3:3], gtint_9[3:3], gtint_10[3:3]);
  NAND3 I53 (simp532_0[0:0], simp531_0[0:0], simp531_0[1:1], simp531_0[2:2]);
  INV I54 (simp532_0[1:1], simp531_0[3:3]);
  OR2 I55 (o_0r1[3:3], simp532_0[0:0], simp532_0[1:1]);
  AND2 I56 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I57 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I58 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I59 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I60 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I61 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I62 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I63 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I64 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I65 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I66 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I67 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AND2 I68 (gtint_3[0:0], choice_3, i_3r1[0:0]);
  AND2 I69 (gtint_3[1:1], choice_3, i_3r1[1:1]);
  AND2 I70 (gtint_3[2:2], choice_3, i_3r1[2:2]);
  AND2 I71 (gtint_3[3:3], choice_3, i_3r1[3:3]);
  AND2 I72 (gtint_4[0:0], choice_4, i_4r1[0:0]);
  AND2 I73 (gtint_4[1:1], choice_4, i_4r1[1:1]);
  AND2 I74 (gtint_4[2:2], choice_4, i_4r1[2:2]);
  AND2 I75 (gtint_4[3:3], choice_4, i_4r1[3:3]);
  AND2 I76 (gtint_5[0:0], choice_5, i_5r1[0:0]);
  AND2 I77 (gtint_5[1:1], choice_5, i_5r1[1:1]);
  AND2 I78 (gtint_5[2:2], choice_5, i_5r1[2:2]);
  AND2 I79 (gtint_5[3:3], choice_5, i_5r1[3:3]);
  AND2 I80 (gtint_6[0:0], choice_6, i_6r1[0:0]);
  AND2 I81 (gtint_6[1:1], choice_6, i_6r1[1:1]);
  AND2 I82 (gtint_6[2:2], choice_6, i_6r1[2:2]);
  AND2 I83 (gtint_6[3:3], choice_6, i_6r1[3:3]);
  AND2 I84 (gtint_7[0:0], choice_7, i_7r1[0:0]);
  AND2 I85 (gtint_7[1:1], choice_7, i_7r1[1:1]);
  AND2 I86 (gtint_7[2:2], choice_7, i_7r1[2:2]);
  AND2 I87 (gtint_7[3:3], choice_7, i_7r1[3:3]);
  AND2 I88 (gtint_8[0:0], choice_8, i_8r1[0:0]);
  AND2 I89 (gtint_8[1:1], choice_8, i_8r1[1:1]);
  AND2 I90 (gtint_8[2:2], choice_8, i_8r1[2:2]);
  AND2 I91 (gtint_8[3:3], choice_8, i_8r1[3:3]);
  AND2 I92 (gtint_9[0:0], choice_9, i_9r1[0:0]);
  AND2 I93 (gtint_9[1:1], choice_9, i_9r1[1:1]);
  AND2 I94 (gtint_9[2:2], choice_9, i_9r1[2:2]);
  AND2 I95 (gtint_9[3:3], choice_9, i_9r1[3:3]);
  AND2 I96 (gtint_10[0:0], choice_10, i_10r1[0:0]);
  AND2 I97 (gtint_10[1:1], choice_10, i_10r1[1:1]);
  AND2 I98 (gtint_10[2:2], choice_10, i_10r1[2:2]);
  AND2 I99 (gtint_10[3:3], choice_10, i_10r1[3:3]);
  AND2 I100 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I101 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I102 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I103 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I104 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I105 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I106 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I107 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I108 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I109 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I110 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I111 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AND2 I112 (gfint_3[0:0], choice_3, i_3r0[0:0]);
  AND2 I113 (gfint_3[1:1], choice_3, i_3r0[1:1]);
  AND2 I114 (gfint_3[2:2], choice_3, i_3r0[2:2]);
  AND2 I115 (gfint_3[3:3], choice_3, i_3r0[3:3]);
  AND2 I116 (gfint_4[0:0], choice_4, i_4r0[0:0]);
  AND2 I117 (gfint_4[1:1], choice_4, i_4r0[1:1]);
  AND2 I118 (gfint_4[2:2], choice_4, i_4r0[2:2]);
  AND2 I119 (gfint_4[3:3], choice_4, i_4r0[3:3]);
  AND2 I120 (gfint_5[0:0], choice_5, i_5r0[0:0]);
  AND2 I121 (gfint_5[1:1], choice_5, i_5r0[1:1]);
  AND2 I122 (gfint_5[2:2], choice_5, i_5r0[2:2]);
  AND2 I123 (gfint_5[3:3], choice_5, i_5r0[3:3]);
  AND2 I124 (gfint_6[0:0], choice_6, i_6r0[0:0]);
  AND2 I125 (gfint_6[1:1], choice_6, i_6r0[1:1]);
  AND2 I126 (gfint_6[2:2], choice_6, i_6r0[2:2]);
  AND2 I127 (gfint_6[3:3], choice_6, i_6r0[3:3]);
  AND2 I128 (gfint_7[0:0], choice_7, i_7r0[0:0]);
  AND2 I129 (gfint_7[1:1], choice_7, i_7r0[1:1]);
  AND2 I130 (gfint_7[2:2], choice_7, i_7r0[2:2]);
  AND2 I131 (gfint_7[3:3], choice_7, i_7r0[3:3]);
  AND2 I132 (gfint_8[0:0], choice_8, i_8r0[0:0]);
  AND2 I133 (gfint_8[1:1], choice_8, i_8r0[1:1]);
  AND2 I134 (gfint_8[2:2], choice_8, i_8r0[2:2]);
  AND2 I135 (gfint_8[3:3], choice_8, i_8r0[3:3]);
  AND2 I136 (gfint_9[0:0], choice_9, i_9r0[0:0]);
  AND2 I137 (gfint_9[1:1], choice_9, i_9r0[1:1]);
  AND2 I138 (gfint_9[2:2], choice_9, i_9r0[2:2]);
  AND2 I139 (gfint_9[3:3], choice_9, i_9r0[3:3]);
  AND2 I140 (gfint_10[0:0], choice_10, i_10r0[0:0]);
  AND2 I141 (gfint_10[1:1], choice_10, i_10r0[1:1]);
  AND2 I142 (gfint_10[2:2], choice_10, i_10r0[2:2]);
  AND2 I143 (gfint_10[3:3], choice_10, i_10r0[3:3]);
  OR2 I144 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I145 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I146 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I147 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  C3 I148 (simp1471_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  BUFF I149 (simp1471_0[1:1], comp0_0[3:3]);
  C2 I150 (icomp_0, simp1471_0[0:0], simp1471_0[1:1]);
  OR2 I151 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I152 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I153 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I154 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  C3 I155 (simp1531_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  BUFF I156 (simp1531_0[1:1], comp1_0[3:3]);
  C2 I157 (icomp_1, simp1531_0[0:0], simp1531_0[1:1]);
  OR2 I158 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I159 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I160 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2 I161 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  C3 I162 (simp1591_0[0:0], comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  BUFF I163 (simp1591_0[1:1], comp2_0[3:3]);
  C2 I164 (icomp_2, simp1591_0[0:0], simp1591_0[1:1]);
  OR2 I165 (comp3_0[0:0], i_3r0[0:0], i_3r1[0:0]);
  OR2 I166 (comp3_0[1:1], i_3r0[1:1], i_3r1[1:1]);
  OR2 I167 (comp3_0[2:2], i_3r0[2:2], i_3r1[2:2]);
  OR2 I168 (comp3_0[3:3], i_3r0[3:3], i_3r1[3:3]);
  C3 I169 (simp1651_0[0:0], comp3_0[0:0], comp3_0[1:1], comp3_0[2:2]);
  BUFF I170 (simp1651_0[1:1], comp3_0[3:3]);
  C2 I171 (icomp_3, simp1651_0[0:0], simp1651_0[1:1]);
  OR2 I172 (comp4_0[0:0], i_4r0[0:0], i_4r1[0:0]);
  OR2 I173 (comp4_0[1:1], i_4r0[1:1], i_4r1[1:1]);
  OR2 I174 (comp4_0[2:2], i_4r0[2:2], i_4r1[2:2]);
  OR2 I175 (comp4_0[3:3], i_4r0[3:3], i_4r1[3:3]);
  C3 I176 (simp1711_0[0:0], comp4_0[0:0], comp4_0[1:1], comp4_0[2:2]);
  BUFF I177 (simp1711_0[1:1], comp4_0[3:3]);
  C2 I178 (icomp_4, simp1711_0[0:0], simp1711_0[1:1]);
  OR2 I179 (comp5_0[0:0], i_5r0[0:0], i_5r1[0:0]);
  OR2 I180 (comp5_0[1:1], i_5r0[1:1], i_5r1[1:1]);
  OR2 I181 (comp5_0[2:2], i_5r0[2:2], i_5r1[2:2]);
  OR2 I182 (comp5_0[3:3], i_5r0[3:3], i_5r1[3:3]);
  C3 I183 (simp1771_0[0:0], comp5_0[0:0], comp5_0[1:1], comp5_0[2:2]);
  BUFF I184 (simp1771_0[1:1], comp5_0[3:3]);
  C2 I185 (icomp_5, simp1771_0[0:0], simp1771_0[1:1]);
  OR2 I186 (comp6_0[0:0], i_6r0[0:0], i_6r1[0:0]);
  OR2 I187 (comp6_0[1:1], i_6r0[1:1], i_6r1[1:1]);
  OR2 I188 (comp6_0[2:2], i_6r0[2:2], i_6r1[2:2]);
  OR2 I189 (comp6_0[3:3], i_6r0[3:3], i_6r1[3:3]);
  C3 I190 (simp1831_0[0:0], comp6_0[0:0], comp6_0[1:1], comp6_0[2:2]);
  BUFF I191 (simp1831_0[1:1], comp6_0[3:3]);
  C2 I192 (icomp_6, simp1831_0[0:0], simp1831_0[1:1]);
  OR2 I193 (comp7_0[0:0], i_7r0[0:0], i_7r1[0:0]);
  OR2 I194 (comp7_0[1:1], i_7r0[1:1], i_7r1[1:1]);
  OR2 I195 (comp7_0[2:2], i_7r0[2:2], i_7r1[2:2]);
  OR2 I196 (comp7_0[3:3], i_7r0[3:3], i_7r1[3:3]);
  C3 I197 (simp1891_0[0:0], comp7_0[0:0], comp7_0[1:1], comp7_0[2:2]);
  BUFF I198 (simp1891_0[1:1], comp7_0[3:3]);
  C2 I199 (icomp_7, simp1891_0[0:0], simp1891_0[1:1]);
  OR2 I200 (comp8_0[0:0], i_8r0[0:0], i_8r1[0:0]);
  OR2 I201 (comp8_0[1:1], i_8r0[1:1], i_8r1[1:1]);
  OR2 I202 (comp8_0[2:2], i_8r0[2:2], i_8r1[2:2]);
  OR2 I203 (comp8_0[3:3], i_8r0[3:3], i_8r1[3:3]);
  C3 I204 (simp1951_0[0:0], comp8_0[0:0], comp8_0[1:1], comp8_0[2:2]);
  BUFF I205 (simp1951_0[1:1], comp8_0[3:3]);
  C2 I206 (icomp_8, simp1951_0[0:0], simp1951_0[1:1]);
  OR2 I207 (comp9_0[0:0], i_9r0[0:0], i_9r1[0:0]);
  OR2 I208 (comp9_0[1:1], i_9r0[1:1], i_9r1[1:1]);
  OR2 I209 (comp9_0[2:2], i_9r0[2:2], i_9r1[2:2]);
  OR2 I210 (comp9_0[3:3], i_9r0[3:3], i_9r1[3:3]);
  C3 I211 (simp2011_0[0:0], comp9_0[0:0], comp9_0[1:1], comp9_0[2:2]);
  BUFF I212 (simp2011_0[1:1], comp9_0[3:3]);
  C2 I213 (icomp_9, simp2011_0[0:0], simp2011_0[1:1]);
  OR2 I214 (comp10_0[0:0], i_10r0[0:0], i_10r1[0:0]);
  OR2 I215 (comp10_0[1:1], i_10r0[1:1], i_10r1[1:1]);
  OR2 I216 (comp10_0[2:2], i_10r0[2:2], i_10r1[2:2]);
  OR2 I217 (comp10_0[3:3], i_10r0[3:3], i_10r1[3:3]);
  C3 I218 (simp2071_0[0:0], comp10_0[0:0], comp10_0[1:1], comp10_0[2:2]);
  BUFF I219 (simp2071_0[1:1], comp10_0[3:3]);
  C2 I220 (icomp_10, simp2071_0[0:0], simp2071_0[1:1]);
  C2R I221 (choice_0, icomp_0, nchosen_0, reset);
  C2R I222 (choice_1, icomp_1, nchosen_0, reset);
  C2R I223 (choice_2, icomp_2, nchosen_0, reset);
  C2R I224 (choice_3, icomp_3, nchosen_0, reset);
  C2R I225 (choice_4, icomp_4, nchosen_0, reset);
  C2R I226 (choice_5, icomp_5, nchosen_0, reset);
  C2R I227 (choice_6, icomp_6, nchosen_0, reset);
  C2R I228 (choice_7, icomp_7, nchosen_0, reset);
  C2R I229 (choice_8, icomp_8, nchosen_0, reset);
  C2R I230 (choice_9, icomp_9, nchosen_0, reset);
  C2R I231 (choice_10, icomp_10, nchosen_0, reset);
  NOR3 I232 (simp2191_0[0:0], choice_0, choice_1, choice_2);
  NOR3 I233 (simp2191_0[1:1], choice_3, choice_4, choice_5);
  NOR3 I234 (simp2191_0[2:2], choice_6, choice_7, choice_8);
  NOR2 I235 (simp2191_0[3:3], choice_9, choice_10);
  NAND3 I236 (simp2192_0[0:0], simp2191_0[0:0], simp2191_0[1:1], simp2191_0[2:2]);
  INV I237 (simp2192_0[1:1], simp2191_0[3:3]);
  OR2 I238 (anychoice_0, simp2192_0[0:0], simp2192_0[1:1]);
  NOR2 I239 (nchosen_0, anychoice_0, o_0a);
  C2R I240 (i_0a, choice_0, o_0a, reset);
  C2R I241 (i_1a, choice_1, o_0a, reset);
  C2R I242 (i_2a, choice_2, o_0a, reset);
  C2R I243 (i_3a, choice_3, o_0a, reset);
  C2R I244 (i_4a, choice_4, o_0a, reset);
  C2R I245 (i_5a, choice_5, o_0a, reset);
  C2R I246 (i_6a, choice_6, o_0a, reset);
  C2R I247 (i_7a, choice_7, o_0a, reset);
  C2R I248 (i_8a, choice_8, o_0a, reset);
  C2R I249 (i_9a, choice_9, o_0a, reset);
  C2R I250 (i_10a, choice_10, o_0a, reset);
endmodule

// tkj4m4_0 TeakJ [Many [4,0],One 4]
module tkj4m4_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [3:0] joinf_0;
  wire [3:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joint_0[0:0], i_0r1[0:0]);
  BUFF I5 (joint_0[1:1], i_0r1[1:1]);
  BUFF I6 (joint_0[2:2], i_0r1[2:2]);
  BUFF I7 (joint_0[3:3], i_0r1[3:3]);
  BUFF I8 (icomplete_0, i_1r);
  C2 I9 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I10 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I11 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I12 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I13 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I14 (o_0r1[1:1], joint_0[1:1]);
  BUFF I15 (o_0r1[2:2], joint_0[2:2]);
  BUFF I16 (o_0r1[3:3], joint_0[3:3]);
  BUFF I17 (i_0a, o_0a);
  BUFF I18 (i_1a, o_0a);
endmodule

// tko0m15_1nm15b0 TeakO [
//     (1,TeakOConstant 15 0)] [One 0,One 15]
module tko0m15_1nm15b0 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [14:0] o_0r0;
  output [14:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r);
  BUFF I1 (o_0r0[1:1], i_0r);
  BUFF I2 (o_0r0[2:2], i_0r);
  BUFF I3 (o_0r0[3:3], i_0r);
  BUFF I4 (o_0r0[4:4], i_0r);
  BUFF I5 (o_0r0[5:5], i_0r);
  BUFF I6 (o_0r0[6:6], i_0r);
  BUFF I7 (o_0r0[7:7], i_0r);
  BUFF I8 (o_0r0[8:8], i_0r);
  BUFF I9 (o_0r0[9:9], i_0r);
  BUFF I10 (o_0r0[10:10], i_0r);
  BUFF I11 (o_0r0[11:11], i_0r);
  BUFF I12 (o_0r0[12:12], i_0r);
  BUFF I13 (o_0r0[13:13], i_0r);
  BUFF I14 (o_0r0[14:14], i_0r);
  GND I15 (o_0r1[0:0]);
  GND I16 (o_0r1[1:1]);
  GND I17 (o_0r1[2:2]);
  GND I18 (o_0r1[3:3]);
  GND I19 (o_0r1[4:4]);
  GND I20 (o_0r1[5:5]);
  GND I21 (o_0r1[6:6]);
  GND I22 (o_0r1[7:7]);
  GND I23 (o_0r1[8:8]);
  GND I24 (o_0r1[9:9]);
  GND I25 (o_0r1[10:10]);
  GND I26 (o_0r1[11:11]);
  GND I27 (o_0r1[12:12]);
  GND I28 (o_0r1[13:13]);
  GND I29 (o_0r1[14:14]);
  BUFF I30 (i_0a, o_0a);
endmodule

// tko0m6_1nm6b0 TeakO [
//     (1,TeakOConstant 6 0)] [One 0,One 6]
module tko0m6_1nm6b0 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [5:0] o_0r0;
  output [5:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r);
  BUFF I1 (o_0r0[1:1], i_0r);
  BUFF I2 (o_0r0[2:2], i_0r);
  BUFF I3 (o_0r0[3:3], i_0r);
  BUFF I4 (o_0r0[4:4], i_0r);
  BUFF I5 (o_0r0[5:5], i_0r);
  GND I6 (o_0r1[0:0]);
  GND I7 (o_0r1[1:1]);
  GND I8 (o_0r1[2:2]);
  GND I9 (o_0r1[3:3]);
  GND I10 (o_0r1[4:4]);
  GND I11 (o_0r1[5:5]);
  BUFF I12 (i_0a, o_0a);
endmodule

// tko0m2_1nm2b0 TeakO [
//     (1,TeakOConstant 2 0)] [One 0,One 2]
module tko0m2_1nm2b0 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r);
  BUFF I1 (o_0r0[1:1], i_0r);
  GND I2 (o_0r1[0:0]);
  GND I3 (o_0r1[1:1]);
  BUFF I4 (i_0a, o_0a);
endmodule

// tkj24m2_22 TeakJ [Many [2,22],One 24]
module tkj24m2_22 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  input [21:0] i_1r0;
  input [21:0] i_1r1;
  output i_1a;
  output [23:0] o_0r0;
  output [23:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [23:0] joinf_0;
  wire [23:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_1r0[0:0]);
  BUFF I3 (joinf_0[3:3], i_1r0[1:1]);
  BUFF I4 (joinf_0[4:4], i_1r0[2:2]);
  BUFF I5 (joinf_0[5:5], i_1r0[3:3]);
  BUFF I6 (joinf_0[6:6], i_1r0[4:4]);
  BUFF I7 (joinf_0[7:7], i_1r0[5:5]);
  BUFF I8 (joinf_0[8:8], i_1r0[6:6]);
  BUFF I9 (joinf_0[9:9], i_1r0[7:7]);
  BUFF I10 (joinf_0[10:10], i_1r0[8:8]);
  BUFF I11 (joinf_0[11:11], i_1r0[9:9]);
  BUFF I12 (joinf_0[12:12], i_1r0[10:10]);
  BUFF I13 (joinf_0[13:13], i_1r0[11:11]);
  BUFF I14 (joinf_0[14:14], i_1r0[12:12]);
  BUFF I15 (joinf_0[15:15], i_1r0[13:13]);
  BUFF I16 (joinf_0[16:16], i_1r0[14:14]);
  BUFF I17 (joinf_0[17:17], i_1r0[15:15]);
  BUFF I18 (joinf_0[18:18], i_1r0[16:16]);
  BUFF I19 (joinf_0[19:19], i_1r0[17:17]);
  BUFF I20 (joinf_0[20:20], i_1r0[18:18]);
  BUFF I21 (joinf_0[21:21], i_1r0[19:19]);
  BUFF I22 (joinf_0[22:22], i_1r0[20:20]);
  BUFF I23 (joinf_0[23:23], i_1r0[21:21]);
  BUFF I24 (joint_0[0:0], i_0r1[0:0]);
  BUFF I25 (joint_0[1:1], i_0r1[1:1]);
  BUFF I26 (joint_0[2:2], i_1r1[0:0]);
  BUFF I27 (joint_0[3:3], i_1r1[1:1]);
  BUFF I28 (joint_0[4:4], i_1r1[2:2]);
  BUFF I29 (joint_0[5:5], i_1r1[3:3]);
  BUFF I30 (joint_0[6:6], i_1r1[4:4]);
  BUFF I31 (joint_0[7:7], i_1r1[5:5]);
  BUFF I32 (joint_0[8:8], i_1r1[6:6]);
  BUFF I33 (joint_0[9:9], i_1r1[7:7]);
  BUFF I34 (joint_0[10:10], i_1r1[8:8]);
  BUFF I35 (joint_0[11:11], i_1r1[9:9]);
  BUFF I36 (joint_0[12:12], i_1r1[10:10]);
  BUFF I37 (joint_0[13:13], i_1r1[11:11]);
  BUFF I38 (joint_0[14:14], i_1r1[12:12]);
  BUFF I39 (joint_0[15:15], i_1r1[13:13]);
  BUFF I40 (joint_0[16:16], i_1r1[14:14]);
  BUFF I41 (joint_0[17:17], i_1r1[15:15]);
  BUFF I42 (joint_0[18:18], i_1r1[16:16]);
  BUFF I43 (joint_0[19:19], i_1r1[17:17]);
  BUFF I44 (joint_0[20:20], i_1r1[18:18]);
  BUFF I45 (joint_0[21:21], i_1r1[19:19]);
  BUFF I46 (joint_0[22:22], i_1r1[20:20]);
  BUFF I47 (joint_0[23:23], i_1r1[21:21]);
  OR2 I48 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I49 (icomplete_0, dcomplete_0);
  C2 I50 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I51 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I52 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I53 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I54 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I55 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I56 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I57 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I58 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I59 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I60 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I61 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I62 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I63 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I64 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I65 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I66 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I67 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I68 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I69 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I70 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I71 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I72 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I73 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I74 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I75 (o_0r1[1:1], joint_0[1:1]);
  BUFF I76 (o_0r1[2:2], joint_0[2:2]);
  BUFF I77 (o_0r1[3:3], joint_0[3:3]);
  BUFF I78 (o_0r1[4:4], joint_0[4:4]);
  BUFF I79 (o_0r1[5:5], joint_0[5:5]);
  BUFF I80 (o_0r1[6:6], joint_0[6:6]);
  BUFF I81 (o_0r1[7:7], joint_0[7:7]);
  BUFF I82 (o_0r1[8:8], joint_0[8:8]);
  BUFF I83 (o_0r1[9:9], joint_0[9:9]);
  BUFF I84 (o_0r1[10:10], joint_0[10:10]);
  BUFF I85 (o_0r1[11:11], joint_0[11:11]);
  BUFF I86 (o_0r1[12:12], joint_0[12:12]);
  BUFF I87 (o_0r1[13:13], joint_0[13:13]);
  BUFF I88 (o_0r1[14:14], joint_0[14:14]);
  BUFF I89 (o_0r1[15:15], joint_0[15:15]);
  BUFF I90 (o_0r1[16:16], joint_0[16:16]);
  BUFF I91 (o_0r1[17:17], joint_0[17:17]);
  BUFF I92 (o_0r1[18:18], joint_0[18:18]);
  BUFF I93 (o_0r1[19:19], joint_0[19:19]);
  BUFF I94 (o_0r1[20:20], joint_0[20:20]);
  BUFF I95 (o_0r1[21:21], joint_0[21:21]);
  BUFF I96 (o_0r1[22:22], joint_0[22:22]);
  BUFF I97 (o_0r1[23:23], joint_0[23:23]);
  BUFF I98 (i_0a, o_0a);
  BUFF I99 (i_1a, o_0a);
endmodule

// tko24m32_1ap8xi23w1b_2api0w24bt1o0w8b TeakO [
//     (1,TeakOAppend 8 [(0,23+:1)]),
//     (2,TeakOAppend 1 [(0,0+:24),(1,0+:8)])] [One 24,One 32]
module tko24m32_1ap8xi23w1b_2api0w24bt1o0w8b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [23:0] i_0r0;
  input [23:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire [7:0] termf_1;
  wire [7:0] termt_1;
  BUFF I0 (termf_1[0:0], i_0r0[23:23]);
  BUFF I1 (termt_1[0:0], i_0r1[23:23]);
  BUFF I2 (termf_1[1:1], i_0r0[23:23]);
  BUFF I3 (termt_1[1:1], i_0r1[23:23]);
  BUFF I4 (termf_1[2:2], i_0r0[23:23]);
  BUFF I5 (termt_1[2:2], i_0r1[23:23]);
  BUFF I6 (termf_1[3:3], i_0r0[23:23]);
  BUFF I7 (termt_1[3:3], i_0r1[23:23]);
  BUFF I8 (termf_1[4:4], i_0r0[23:23]);
  BUFF I9 (termt_1[4:4], i_0r1[23:23]);
  BUFF I10 (termf_1[5:5], i_0r0[23:23]);
  BUFF I11 (termt_1[5:5], i_0r1[23:23]);
  BUFF I12 (termf_1[6:6], i_0r0[23:23]);
  BUFF I13 (termt_1[6:6], i_0r1[23:23]);
  BUFF I14 (termf_1[7:7], i_0r0[23:23]);
  BUFF I15 (termt_1[7:7], i_0r1[23:23]);
  BUFF I16 (o_0r0[0:0], i_0r0[0:0]);
  BUFF I17 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I18 (o_0r0[2:2], i_0r0[2:2]);
  BUFF I19 (o_0r0[3:3], i_0r0[3:3]);
  BUFF I20 (o_0r0[4:4], i_0r0[4:4]);
  BUFF I21 (o_0r0[5:5], i_0r0[5:5]);
  BUFF I22 (o_0r0[6:6], i_0r0[6:6]);
  BUFF I23 (o_0r0[7:7], i_0r0[7:7]);
  BUFF I24 (o_0r0[8:8], i_0r0[8:8]);
  BUFF I25 (o_0r0[9:9], i_0r0[9:9]);
  BUFF I26 (o_0r0[10:10], i_0r0[10:10]);
  BUFF I27 (o_0r0[11:11], i_0r0[11:11]);
  BUFF I28 (o_0r0[12:12], i_0r0[12:12]);
  BUFF I29 (o_0r0[13:13], i_0r0[13:13]);
  BUFF I30 (o_0r0[14:14], i_0r0[14:14]);
  BUFF I31 (o_0r0[15:15], i_0r0[15:15]);
  BUFF I32 (o_0r0[16:16], i_0r0[16:16]);
  BUFF I33 (o_0r0[17:17], i_0r0[17:17]);
  BUFF I34 (o_0r0[18:18], i_0r0[18:18]);
  BUFF I35 (o_0r0[19:19], i_0r0[19:19]);
  BUFF I36 (o_0r0[20:20], i_0r0[20:20]);
  BUFF I37 (o_0r0[21:21], i_0r0[21:21]);
  BUFF I38 (o_0r0[22:22], i_0r0[22:22]);
  BUFF I39 (o_0r0[23:23], i_0r0[23:23]);
  BUFF I40 (o_0r0[24:24], termf_1[0:0]);
  BUFF I41 (o_0r0[25:25], termf_1[1:1]);
  BUFF I42 (o_0r0[26:26], termf_1[2:2]);
  BUFF I43 (o_0r0[27:27], termf_1[3:3]);
  BUFF I44 (o_0r0[28:28], termf_1[4:4]);
  BUFF I45 (o_0r0[29:29], termf_1[5:5]);
  BUFF I46 (o_0r0[30:30], termf_1[6:6]);
  BUFF I47 (o_0r0[31:31], termf_1[7:7]);
  BUFF I48 (o_0r1[0:0], i_0r1[0:0]);
  BUFF I49 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I50 (o_0r1[2:2], i_0r1[2:2]);
  BUFF I51 (o_0r1[3:3], i_0r1[3:3]);
  BUFF I52 (o_0r1[4:4], i_0r1[4:4]);
  BUFF I53 (o_0r1[5:5], i_0r1[5:5]);
  BUFF I54 (o_0r1[6:6], i_0r1[6:6]);
  BUFF I55 (o_0r1[7:7], i_0r1[7:7]);
  BUFF I56 (o_0r1[8:8], i_0r1[8:8]);
  BUFF I57 (o_0r1[9:9], i_0r1[9:9]);
  BUFF I58 (o_0r1[10:10], i_0r1[10:10]);
  BUFF I59 (o_0r1[11:11], i_0r1[11:11]);
  BUFF I60 (o_0r1[12:12], i_0r1[12:12]);
  BUFF I61 (o_0r1[13:13], i_0r1[13:13]);
  BUFF I62 (o_0r1[14:14], i_0r1[14:14]);
  BUFF I63 (o_0r1[15:15], i_0r1[15:15]);
  BUFF I64 (o_0r1[16:16], i_0r1[16:16]);
  BUFF I65 (o_0r1[17:17], i_0r1[17:17]);
  BUFF I66 (o_0r1[18:18], i_0r1[18:18]);
  BUFF I67 (o_0r1[19:19], i_0r1[19:19]);
  BUFF I68 (o_0r1[20:20], i_0r1[20:20]);
  BUFF I69 (o_0r1[21:21], i_0r1[21:21]);
  BUFF I70 (o_0r1[22:22], i_0r1[22:22]);
  BUFF I71 (o_0r1[23:23], i_0r1[23:23]);
  BUFF I72 (o_0r1[24:24], termt_1[0:0]);
  BUFF I73 (o_0r1[25:25], termt_1[1:1]);
  BUFF I74 (o_0r1[26:26], termt_1[2:2]);
  BUFF I75 (o_0r1[27:27], termt_1[3:3]);
  BUFF I76 (o_0r1[28:28], termt_1[4:4]);
  BUFF I77 (o_0r1[29:29], termt_1[5:5]);
  BUFF I78 (o_0r1[30:30], termt_1[6:6]);
  BUFF I79 (o_0r1[31:31], termt_1[7:7]);
  BUFF I80 (i_0a, o_0a);
endmodule

// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 TeakF [0,0,0,0,0,0,0,0,0,0,0] [One 0,Man
//   y [0,0,0,0,0,0,0,0,0,0,0]]
module tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, o_5r, o_5a, o_6r, o_6a, o_7r, o_7a, o_8r, o_8a, o_9r, o_9a, o_10r, o_10a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  output o_7r;
  input o_7a;
  output o_8r;
  input o_8a;
  output o_9r;
  input o_9a;
  output o_10r;
  input o_10a;
  input reset;
  wire [3:0] simp11_0;
  wire [1:0] simp12_0;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  BUFF I2 (o_2r, i_0r);
  BUFF I3 (o_3r, i_0r);
  BUFF I4 (o_4r, i_0r);
  BUFF I5 (o_5r, i_0r);
  BUFF I6 (o_6r, i_0r);
  BUFF I7 (o_7r, i_0r);
  BUFF I8 (o_8r, i_0r);
  BUFF I9 (o_9r, i_0r);
  BUFF I10 (o_10r, i_0r);
  C3 I11 (simp11_0[0:0], o_0a, o_1a, o_2a);
  C3 I12 (simp11_0[1:1], o_3a, o_4a, o_5a);
  C3 I13 (simp11_0[2:2], o_6a, o_7a, o_8a);
  C2 I14 (simp11_0[3:3], o_9a, o_10a);
  C3 I15 (simp12_0[0:0], simp11_0[0:0], simp11_0[1:1], simp11_0[2:2]);
  BUFF I16 (simp12_0[1:1], simp11_0[3:3]);
  C2 I17 (i_0a, simp12_0[0:0], simp12_0[1:1]);
endmodule

// tko0m10_1nm10b0 TeakO [
//     (1,TeakOConstant 10 0)] [One 0,One 10]
module tko0m10_1nm10b0 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [9:0] o_0r0;
  output [9:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r);
  BUFF I1 (o_0r0[1:1], i_0r);
  BUFF I2 (o_0r0[2:2], i_0r);
  BUFF I3 (o_0r0[3:3], i_0r);
  BUFF I4 (o_0r0[4:4], i_0r);
  BUFF I5 (o_0r0[5:5], i_0r);
  BUFF I6 (o_0r0[6:6], i_0r);
  BUFF I7 (o_0r0[7:7], i_0r);
  BUFF I8 (o_0r0[8:8], i_0r);
  BUFF I9 (o_0r0[9:9], i_0r);
  GND I10 (o_0r1[0:0]);
  GND I11 (o_0r1[1:1]);
  GND I12 (o_0r1[2:2]);
  GND I13 (o_0r1[3:3]);
  GND I14 (o_0r1[4:4]);
  GND I15 (o_0r1[5:5]);
  GND I16 (o_0r1[6:6]);
  GND I17 (o_0r1[7:7]);
  GND I18 (o_0r1[8:8]);
  GND I19 (o_0r1[9:9]);
  BUFF I20 (i_0a, o_0a);
endmodule

// tkj32m10_22 TeakJ [Many [10,22],One 32]
module tkj32m10_22 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [9:0] i_0r0;
  input [9:0] i_0r1;
  output i_0a;
  input [21:0] i_1r0;
  input [21:0] i_1r1;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [31:0] joinf_0;
  wire [31:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_1r0[0:0]);
  BUFF I11 (joinf_0[11:11], i_1r0[1:1]);
  BUFF I12 (joinf_0[12:12], i_1r0[2:2]);
  BUFF I13 (joinf_0[13:13], i_1r0[3:3]);
  BUFF I14 (joinf_0[14:14], i_1r0[4:4]);
  BUFF I15 (joinf_0[15:15], i_1r0[5:5]);
  BUFF I16 (joinf_0[16:16], i_1r0[6:6]);
  BUFF I17 (joinf_0[17:17], i_1r0[7:7]);
  BUFF I18 (joinf_0[18:18], i_1r0[8:8]);
  BUFF I19 (joinf_0[19:19], i_1r0[9:9]);
  BUFF I20 (joinf_0[20:20], i_1r0[10:10]);
  BUFF I21 (joinf_0[21:21], i_1r0[11:11]);
  BUFF I22 (joinf_0[22:22], i_1r0[12:12]);
  BUFF I23 (joinf_0[23:23], i_1r0[13:13]);
  BUFF I24 (joinf_0[24:24], i_1r0[14:14]);
  BUFF I25 (joinf_0[25:25], i_1r0[15:15]);
  BUFF I26 (joinf_0[26:26], i_1r0[16:16]);
  BUFF I27 (joinf_0[27:27], i_1r0[17:17]);
  BUFF I28 (joinf_0[28:28], i_1r0[18:18]);
  BUFF I29 (joinf_0[29:29], i_1r0[19:19]);
  BUFF I30 (joinf_0[30:30], i_1r0[20:20]);
  BUFF I31 (joinf_0[31:31], i_1r0[21:21]);
  BUFF I32 (joint_0[0:0], i_0r1[0:0]);
  BUFF I33 (joint_0[1:1], i_0r1[1:1]);
  BUFF I34 (joint_0[2:2], i_0r1[2:2]);
  BUFF I35 (joint_0[3:3], i_0r1[3:3]);
  BUFF I36 (joint_0[4:4], i_0r1[4:4]);
  BUFF I37 (joint_0[5:5], i_0r1[5:5]);
  BUFF I38 (joint_0[6:6], i_0r1[6:6]);
  BUFF I39 (joint_0[7:7], i_0r1[7:7]);
  BUFF I40 (joint_0[8:8], i_0r1[8:8]);
  BUFF I41 (joint_0[9:9], i_0r1[9:9]);
  BUFF I42 (joint_0[10:10], i_1r1[0:0]);
  BUFF I43 (joint_0[11:11], i_1r1[1:1]);
  BUFF I44 (joint_0[12:12], i_1r1[2:2]);
  BUFF I45 (joint_0[13:13], i_1r1[3:3]);
  BUFF I46 (joint_0[14:14], i_1r1[4:4]);
  BUFF I47 (joint_0[15:15], i_1r1[5:5]);
  BUFF I48 (joint_0[16:16], i_1r1[6:6]);
  BUFF I49 (joint_0[17:17], i_1r1[7:7]);
  BUFF I50 (joint_0[18:18], i_1r1[8:8]);
  BUFF I51 (joint_0[19:19], i_1r1[9:9]);
  BUFF I52 (joint_0[20:20], i_1r1[10:10]);
  BUFF I53 (joint_0[21:21], i_1r1[11:11]);
  BUFF I54 (joint_0[22:22], i_1r1[12:12]);
  BUFF I55 (joint_0[23:23], i_1r1[13:13]);
  BUFF I56 (joint_0[24:24], i_1r1[14:14]);
  BUFF I57 (joint_0[25:25], i_1r1[15:15]);
  BUFF I58 (joint_0[26:26], i_1r1[16:16]);
  BUFF I59 (joint_0[27:27], i_1r1[17:17]);
  BUFF I60 (joint_0[28:28], i_1r1[18:18]);
  BUFF I61 (joint_0[29:29], i_1r1[19:19]);
  BUFF I62 (joint_0[30:30], i_1r1[20:20]);
  BUFF I63 (joint_0[31:31], i_1r1[21:21]);
  OR2 I64 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I65 (icomplete_0, dcomplete_0);
  C2 I66 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I67 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I68 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I69 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I70 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I71 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I72 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I73 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I74 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I75 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I76 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I77 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I78 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I79 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I80 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I81 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I82 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I83 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I84 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I85 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I86 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I87 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I88 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I89 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I90 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I91 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I92 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I93 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I94 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I95 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I96 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I97 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I98 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I99 (o_0r1[1:1], joint_0[1:1]);
  BUFF I100 (o_0r1[2:2], joint_0[2:2]);
  BUFF I101 (o_0r1[3:3], joint_0[3:3]);
  BUFF I102 (o_0r1[4:4], joint_0[4:4]);
  BUFF I103 (o_0r1[5:5], joint_0[5:5]);
  BUFF I104 (o_0r1[6:6], joint_0[6:6]);
  BUFF I105 (o_0r1[7:7], joint_0[7:7]);
  BUFF I106 (o_0r1[8:8], joint_0[8:8]);
  BUFF I107 (o_0r1[9:9], joint_0[9:9]);
  BUFF I108 (o_0r1[10:10], joint_0[10:10]);
  BUFF I109 (o_0r1[11:11], joint_0[11:11]);
  BUFF I110 (o_0r1[12:12], joint_0[12:12]);
  BUFF I111 (o_0r1[13:13], joint_0[13:13]);
  BUFF I112 (o_0r1[14:14], joint_0[14:14]);
  BUFF I113 (o_0r1[15:15], joint_0[15:15]);
  BUFF I114 (o_0r1[16:16], joint_0[16:16]);
  BUFF I115 (o_0r1[17:17], joint_0[17:17]);
  BUFF I116 (o_0r1[18:18], joint_0[18:18]);
  BUFF I117 (o_0r1[19:19], joint_0[19:19]);
  BUFF I118 (o_0r1[20:20], joint_0[20:20]);
  BUFF I119 (o_0r1[21:21], joint_0[21:21]);
  BUFF I120 (o_0r1[22:22], joint_0[22:22]);
  BUFF I121 (o_0r1[23:23], joint_0[23:23]);
  BUFF I122 (o_0r1[24:24], joint_0[24:24]);
  BUFF I123 (o_0r1[25:25], joint_0[25:25]);
  BUFF I124 (o_0r1[26:26], joint_0[26:26]);
  BUFF I125 (o_0r1[27:27], joint_0[27:27]);
  BUFF I126 (o_0r1[28:28], joint_0[28:28]);
  BUFF I127 (o_0r1[29:29], joint_0[29:29]);
  BUFF I128 (o_0r1[30:30], joint_0[30:30]);
  BUFF I129 (o_0r1[31:31], joint_0[31:31]);
  BUFF I130 (i_0a, o_0a);
  BUFF I131 (i_1a, o_0a);
endmodule

// tks3_o0w3_0m1c6m6o0w0_2o0w0_4o0w0 TeakS (0+:3) [([Imp 0 0,Imp 1 6,Imp 6 0],0),([Imp 2 0],0),([Imp 4 
//   0],0)] [One 3,Many [0,0,0]]
module tks3_o0w3_0m1c6m6o0w0_2o0w0_4o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire oack_0;
  wire [2:0] match0_0;
  wire match1_0;
  wire match2_0;
  wire [2:0] comp_0;
  OR3 I0 (sel_0, match0_0[0:0], match0_0[1:1], match0_0[2:2]);
  C3 I1 (match0_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I2 (match0_0[1:1], i_0r1[0:0]);
  C3 I3 (match0_0[2:2], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I4 (sel_1, match1_0);
  C3 I5 (match1_0, i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I6 (sel_2, match2_0);
  C3 I7 (match2_0, i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C2 I8 (gsel_0, sel_0, icomplete_0);
  C2 I9 (gsel_1, sel_1, icomplete_0);
  C2 I10 (gsel_2, sel_2, icomplete_0);
  OR2 I11 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I12 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I13 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I14 (icomplete_0, comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  BUFF I15 (o_0r, gsel_0);
  BUFF I16 (o_1r, gsel_1);
  BUFF I17 (o_2r, gsel_2);
  OR3 I18 (oack_0, o_0a, o_1a, o_2a);
  C2 I19 (i_0a, oack_0, icomplete_0);
endmodule

// tkm3x0b TeakM [Many [0,0,0],One 0]
module tkm3x0b (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  output o_0r;
  input o_0a;
  input reset;
  wire nchosen_0;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  C2R I0 (choice_0, i_0r, nchosen_0, reset);
  C2R I1 (choice_1, i_1r, nchosen_0, reset);
  C2R I2 (choice_2, i_2r, nchosen_0, reset);
  NOR2 I3 (nchosen_0, o_0r, o_0a);
  OR3 I4 (o_0r, choice_0, choice_1, choice_2);
  C2R I5 (i_0a, choice_0, o_0a, reset);
  C2R I6 (i_1a, choice_1, o_0a, reset);
  C2R I7 (i_2a, choice_2, o_0a, reset);
endmodule

// tks2_o0w2_1o0w0_2o0w0_3o0w0_0o0w0 TeakS (0+:2) [([Imp 1 0],0),([Imp 2 0],0),([Imp 3 0],0),([Imp 0 0]
//   ,0)] [One 2,Many [0,0,0,0]]
module tks2_o0w2_1o0w0_2o0w0_3o0w0_0o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire match2_0;
  wire match3_0;
  wire [1:0] comp_0;
  wire [1:0] simp341_0;
  BUFF I0 (sel_0, match0_0);
  C2 I1 (match0_0, i_0r1[0:0], i_0r0[1:1]);
  BUFF I2 (sel_1, match1_0);
  C2 I3 (match1_0, i_0r0[0:0], i_0r1[1:1]);
  BUFF I4 (sel_2, match2_0);
  C2 I5 (match2_0, i_0r1[0:0], i_0r1[1:1]);
  BUFF I6 (sel_3, match3_0);
  C2 I7 (match3_0, i_0r0[0:0], i_0r0[1:1]);
  C2 I8 (gsel_0, sel_0, icomplete_0);
  C2 I9 (gsel_1, sel_1, icomplete_0);
  C2 I10 (gsel_2, sel_2, icomplete_0);
  C2 I11 (gsel_3, sel_3, icomplete_0);
  OR2 I12 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I13 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  C2 I14 (icomplete_0, comp_0[0:0], comp_0[1:1]);
  BUFF I15 (o_0r, gsel_0);
  BUFF I16 (o_1r, gsel_1);
  BUFF I17 (o_2r, gsel_2);
  BUFF I18 (o_3r, gsel_3);
  NOR3 I19 (simp341_0[0:0], o_0a, o_1a, o_2a);
  INV I20 (simp341_0[1:1], o_3a);
  NAND2 I21 (oack_0, simp341_0[0:0], simp341_0[1:1]);
  C2 I22 (i_0a, oack_0, icomplete_0);
endmodule

// tkm4x0b TeakM [Many [0,0,0,0],One 0]
module tkm4x0b (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, i_3r, i_3a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  output o_0r;
  input o_0a;
  input reset;
  wire nchosen_0;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire [1:0] simp101_0;
  C2R I0 (choice_0, i_0r, nchosen_0, reset);
  C2R I1 (choice_1, i_1r, nchosen_0, reset);
  C2R I2 (choice_2, i_2r, nchosen_0, reset);
  C2R I3 (choice_3, i_3r, nchosen_0, reset);
  NOR2 I4 (nchosen_0, o_0r, o_0a);
  NOR3 I5 (simp101_0[0:0], choice_0, choice_1, choice_2);
  INV I6 (simp101_0[1:1], choice_3);
  NAND2 I7 (o_0r, simp101_0[0:0], simp101_0[1:1]);
  C2R I8 (i_0a, choice_0, o_0a, reset);
  C2R I9 (i_1a, choice_1, o_0a, reset);
  C2R I10 (i_2a, choice_2, o_0a, reset);
  C2R I11 (i_3a, choice_3, o_0a, reset);
endmodule

// tko0m74_1nm74b1c00000000000000040 TeakO [
//     (1,TeakOConstant 74 8264141345021879124032)] [One 0,One 74]
module tko0m74_1nm74b1c00000000000000040 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [73:0] o_0r0;
  output [73:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[6:6], i_0r);
  BUFF I1 (o_0r1[70:70], i_0r);
  BUFF I2 (o_0r1[71:71], i_0r);
  BUFF I3 (o_0r1[72:72], i_0r);
  GND I4 (o_0r0[6:6]);
  GND I5 (o_0r0[70:70]);
  GND I6 (o_0r0[71:71]);
  GND I7 (o_0r0[72:72]);
  BUFF I8 (o_0r0[0:0], i_0r);
  BUFF I9 (o_0r0[1:1], i_0r);
  BUFF I10 (o_0r0[2:2], i_0r);
  BUFF I11 (o_0r0[3:3], i_0r);
  BUFF I12 (o_0r0[4:4], i_0r);
  BUFF I13 (o_0r0[5:5], i_0r);
  BUFF I14 (o_0r0[7:7], i_0r);
  BUFF I15 (o_0r0[8:8], i_0r);
  BUFF I16 (o_0r0[9:9], i_0r);
  BUFF I17 (o_0r0[10:10], i_0r);
  BUFF I18 (o_0r0[11:11], i_0r);
  BUFF I19 (o_0r0[12:12], i_0r);
  BUFF I20 (o_0r0[13:13], i_0r);
  BUFF I21 (o_0r0[14:14], i_0r);
  BUFF I22 (o_0r0[15:15], i_0r);
  BUFF I23 (o_0r0[16:16], i_0r);
  BUFF I24 (o_0r0[17:17], i_0r);
  BUFF I25 (o_0r0[18:18], i_0r);
  BUFF I26 (o_0r0[19:19], i_0r);
  BUFF I27 (o_0r0[20:20], i_0r);
  BUFF I28 (o_0r0[21:21], i_0r);
  BUFF I29 (o_0r0[22:22], i_0r);
  BUFF I30 (o_0r0[23:23], i_0r);
  BUFF I31 (o_0r0[24:24], i_0r);
  BUFF I32 (o_0r0[25:25], i_0r);
  BUFF I33 (o_0r0[26:26], i_0r);
  BUFF I34 (o_0r0[27:27], i_0r);
  BUFF I35 (o_0r0[28:28], i_0r);
  BUFF I36 (o_0r0[29:29], i_0r);
  BUFF I37 (o_0r0[30:30], i_0r);
  BUFF I38 (o_0r0[31:31], i_0r);
  BUFF I39 (o_0r0[32:32], i_0r);
  BUFF I40 (o_0r0[33:33], i_0r);
  BUFF I41 (o_0r0[34:34], i_0r);
  BUFF I42 (o_0r0[35:35], i_0r);
  BUFF I43 (o_0r0[36:36], i_0r);
  BUFF I44 (o_0r0[37:37], i_0r);
  BUFF I45 (o_0r0[38:38], i_0r);
  BUFF I46 (o_0r0[39:39], i_0r);
  BUFF I47 (o_0r0[40:40], i_0r);
  BUFF I48 (o_0r0[41:41], i_0r);
  BUFF I49 (o_0r0[42:42], i_0r);
  BUFF I50 (o_0r0[43:43], i_0r);
  BUFF I51 (o_0r0[44:44], i_0r);
  BUFF I52 (o_0r0[45:45], i_0r);
  BUFF I53 (o_0r0[46:46], i_0r);
  BUFF I54 (o_0r0[47:47], i_0r);
  BUFF I55 (o_0r0[48:48], i_0r);
  BUFF I56 (o_0r0[49:49], i_0r);
  BUFF I57 (o_0r0[50:50], i_0r);
  BUFF I58 (o_0r0[51:51], i_0r);
  BUFF I59 (o_0r0[52:52], i_0r);
  BUFF I60 (o_0r0[53:53], i_0r);
  BUFF I61 (o_0r0[54:54], i_0r);
  BUFF I62 (o_0r0[55:55], i_0r);
  BUFF I63 (o_0r0[56:56], i_0r);
  BUFF I64 (o_0r0[57:57], i_0r);
  BUFF I65 (o_0r0[58:58], i_0r);
  BUFF I66 (o_0r0[59:59], i_0r);
  BUFF I67 (o_0r0[60:60], i_0r);
  BUFF I68 (o_0r0[61:61], i_0r);
  BUFF I69 (o_0r0[62:62], i_0r);
  BUFF I70 (o_0r0[63:63], i_0r);
  BUFF I71 (o_0r0[64:64], i_0r);
  BUFF I72 (o_0r0[65:65], i_0r);
  BUFF I73 (o_0r0[66:66], i_0r);
  BUFF I74 (o_0r0[67:67], i_0r);
  BUFF I75 (o_0r0[68:68], i_0r);
  BUFF I76 (o_0r0[69:69], i_0r);
  BUFF I77 (o_0r0[73:73], i_0r);
  GND I78 (o_0r1[0:0]);
  GND I79 (o_0r1[1:1]);
  GND I80 (o_0r1[2:2]);
  GND I81 (o_0r1[3:3]);
  GND I82 (o_0r1[4:4]);
  GND I83 (o_0r1[5:5]);
  GND I84 (o_0r1[7:7]);
  GND I85 (o_0r1[8:8]);
  GND I86 (o_0r1[9:9]);
  GND I87 (o_0r1[10:10]);
  GND I88 (o_0r1[11:11]);
  GND I89 (o_0r1[12:12]);
  GND I90 (o_0r1[13:13]);
  GND I91 (o_0r1[14:14]);
  GND I92 (o_0r1[15:15]);
  GND I93 (o_0r1[16:16]);
  GND I94 (o_0r1[17:17]);
  GND I95 (o_0r1[18:18]);
  GND I96 (o_0r1[19:19]);
  GND I97 (o_0r1[20:20]);
  GND I98 (o_0r1[21:21]);
  GND I99 (o_0r1[22:22]);
  GND I100 (o_0r1[23:23]);
  GND I101 (o_0r1[24:24]);
  GND I102 (o_0r1[25:25]);
  GND I103 (o_0r1[26:26]);
  GND I104 (o_0r1[27:27]);
  GND I105 (o_0r1[28:28]);
  GND I106 (o_0r1[29:29]);
  GND I107 (o_0r1[30:30]);
  GND I108 (o_0r1[31:31]);
  GND I109 (o_0r1[32:32]);
  GND I110 (o_0r1[33:33]);
  GND I111 (o_0r1[34:34]);
  GND I112 (o_0r1[35:35]);
  GND I113 (o_0r1[36:36]);
  GND I114 (o_0r1[37:37]);
  GND I115 (o_0r1[38:38]);
  GND I116 (o_0r1[39:39]);
  GND I117 (o_0r1[40:40]);
  GND I118 (o_0r1[41:41]);
  GND I119 (o_0r1[42:42]);
  GND I120 (o_0r1[43:43]);
  GND I121 (o_0r1[44:44]);
  GND I122 (o_0r1[45:45]);
  GND I123 (o_0r1[46:46]);
  GND I124 (o_0r1[47:47]);
  GND I125 (o_0r1[48:48]);
  GND I126 (o_0r1[49:49]);
  GND I127 (o_0r1[50:50]);
  GND I128 (o_0r1[51:51]);
  GND I129 (o_0r1[52:52]);
  GND I130 (o_0r1[53:53]);
  GND I131 (o_0r1[54:54]);
  GND I132 (o_0r1[55:55]);
  GND I133 (o_0r1[56:56]);
  GND I134 (o_0r1[57:57]);
  GND I135 (o_0r1[58:58]);
  GND I136 (o_0r1[59:59]);
  GND I137 (o_0r1[60:60]);
  GND I138 (o_0r1[61:61]);
  GND I139 (o_0r1[62:62]);
  GND I140 (o_0r1[63:63]);
  GND I141 (o_0r1[64:64]);
  GND I142 (o_0r1[65:65]);
  GND I143 (o_0r1[66:66]);
  GND I144 (o_0r1[67:67]);
  GND I145 (o_0r1[68:68]);
  GND I146 (o_0r1[69:69]);
  GND I147 (o_0r1[73:73]);
  BUFF I148 (i_0a, o_0a);
endmodule

// tko0m4_1nm4b1 TeakO [
//     (1,TeakOConstant 4 1)] [One 0,One 4]
module tko0m4_1nm4b1 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  GND I1 (o_0r0[0:0]);
  BUFF I2 (o_0r0[1:1], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  GND I5 (o_0r1[1:1]);
  GND I6 (o_0r1[2:2]);
  GND I7 (o_0r1[3:3]);
  BUFF I8 (i_0a, o_0a);
endmodule

// tkm4x4b TeakM [Many [4,4,4,4],One 4]
module tkm4x4b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, o_0r0, o_0r1, o_0a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  input [3:0] i_1r0;
  input [3:0] i_1r1;
  output i_1a;
  input [3:0] i_2r0;
  input [3:0] i_2r1;
  output i_2a;
  input [3:0] i_3r0;
  input [3:0] i_3r1;
  output i_3a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  wire [3:0] gfint_0;
  wire [3:0] gfint_1;
  wire [3:0] gfint_2;
  wire [3:0] gfint_3;
  wire [3:0] gtint_0;
  wire [3:0] gtint_1;
  wire [3:0] gtint_2;
  wire [3:0] gtint_3;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire icomp_3;
  wire nchosen_0;
  wire [1:0] simp181_0;
  wire [1:0] simp191_0;
  wire [1:0] simp201_0;
  wire [1:0] simp211_0;
  wire [1:0] simp221_0;
  wire [1:0] simp231_0;
  wire [1:0] simp241_0;
  wire [1:0] simp251_0;
  wire [3:0] comp0_0;
  wire [1:0] simp631_0;
  wire [3:0] comp1_0;
  wire [1:0] simp691_0;
  wire [3:0] comp2_0;
  wire [1:0] simp751_0;
  wire [3:0] comp3_0;
  wire [1:0] simp811_0;
  wire [1:0] simp861_0;
  NOR3 I0 (simp181_0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  INV I1 (simp181_0[1:1], gfint_3[0:0]);
  NAND2 I2 (o_0r0[0:0], simp181_0[0:0], simp181_0[1:1]);
  NOR3 I3 (simp191_0[0:0], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  INV I4 (simp191_0[1:1], gfint_3[1:1]);
  NAND2 I5 (o_0r0[1:1], simp191_0[0:0], simp191_0[1:1]);
  NOR3 I6 (simp201_0[0:0], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  INV I7 (simp201_0[1:1], gfint_3[2:2]);
  NAND2 I8 (o_0r0[2:2], simp201_0[0:0], simp201_0[1:1]);
  NOR3 I9 (simp211_0[0:0], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  INV I10 (simp211_0[1:1], gfint_3[3:3]);
  NAND2 I11 (o_0r0[3:3], simp211_0[0:0], simp211_0[1:1]);
  NOR3 I12 (simp221_0[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  INV I13 (simp221_0[1:1], gtint_3[0:0]);
  NAND2 I14 (o_0r1[0:0], simp221_0[0:0], simp221_0[1:1]);
  NOR3 I15 (simp231_0[0:0], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  INV I16 (simp231_0[1:1], gtint_3[1:1]);
  NAND2 I17 (o_0r1[1:1], simp231_0[0:0], simp231_0[1:1]);
  NOR3 I18 (simp241_0[0:0], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  INV I19 (simp241_0[1:1], gtint_3[2:2]);
  NAND2 I20 (o_0r1[2:2], simp241_0[0:0], simp241_0[1:1]);
  NOR3 I21 (simp251_0[0:0], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  INV I22 (simp251_0[1:1], gtint_3[3:3]);
  NAND2 I23 (o_0r1[3:3], simp251_0[0:0], simp251_0[1:1]);
  AND2 I24 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I25 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I26 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I27 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I28 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I29 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I30 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I31 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I32 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I33 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I34 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I35 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AND2 I36 (gtint_3[0:0], choice_3, i_3r1[0:0]);
  AND2 I37 (gtint_3[1:1], choice_3, i_3r1[1:1]);
  AND2 I38 (gtint_3[2:2], choice_3, i_3r1[2:2]);
  AND2 I39 (gtint_3[3:3], choice_3, i_3r1[3:3]);
  AND2 I40 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I41 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I42 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I43 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I44 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I45 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I46 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I47 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I48 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I49 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I50 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I51 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AND2 I52 (gfint_3[0:0], choice_3, i_3r0[0:0]);
  AND2 I53 (gfint_3[1:1], choice_3, i_3r0[1:1]);
  AND2 I54 (gfint_3[2:2], choice_3, i_3r0[2:2]);
  AND2 I55 (gfint_3[3:3], choice_3, i_3r0[3:3]);
  OR2 I56 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I57 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I58 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I59 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  C3 I60 (simp631_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  BUFF I61 (simp631_0[1:1], comp0_0[3:3]);
  C2 I62 (icomp_0, simp631_0[0:0], simp631_0[1:1]);
  OR2 I63 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I64 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I65 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I66 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  C3 I67 (simp691_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  BUFF I68 (simp691_0[1:1], comp1_0[3:3]);
  C2 I69 (icomp_1, simp691_0[0:0], simp691_0[1:1]);
  OR2 I70 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I71 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I72 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2 I73 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  C3 I74 (simp751_0[0:0], comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  BUFF I75 (simp751_0[1:1], comp2_0[3:3]);
  C2 I76 (icomp_2, simp751_0[0:0], simp751_0[1:1]);
  OR2 I77 (comp3_0[0:0], i_3r0[0:0], i_3r1[0:0]);
  OR2 I78 (comp3_0[1:1], i_3r0[1:1], i_3r1[1:1]);
  OR2 I79 (comp3_0[2:2], i_3r0[2:2], i_3r1[2:2]);
  OR2 I80 (comp3_0[3:3], i_3r0[3:3], i_3r1[3:3]);
  C3 I81 (simp811_0[0:0], comp3_0[0:0], comp3_0[1:1], comp3_0[2:2]);
  BUFF I82 (simp811_0[1:1], comp3_0[3:3]);
  C2 I83 (icomp_3, simp811_0[0:0], simp811_0[1:1]);
  C2R I84 (choice_0, icomp_0, nchosen_0, reset);
  C2R I85 (choice_1, icomp_1, nchosen_0, reset);
  C2R I86 (choice_2, icomp_2, nchosen_0, reset);
  C2R I87 (choice_3, icomp_3, nchosen_0, reset);
  NOR3 I88 (simp861_0[0:0], choice_0, choice_1, choice_2);
  INV I89 (simp861_0[1:1], choice_3);
  NAND2 I90 (anychoice_0, simp861_0[0:0], simp861_0[1:1]);
  NOR2 I91 (nchosen_0, anychoice_0, o_0a);
  C2R I92 (i_0a, choice_0, o_0a, reset);
  C2R I93 (i_1a, choice_1, o_0a, reset);
  C2R I94 (i_2a, choice_2, o_0a, reset);
  C2R I95 (i_3a, choice_3, o_0a, reset);
endmodule

// tkj4m0_4 TeakJ [Many [0,4],One 4]
module tkj4m0_4 (i_0r, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  input [3:0] i_1r0;
  input [3:0] i_1r1;
  output i_1a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [3:0] joinf_0;
  wire [3:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_1r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_1r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_1r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_1r0[3:3]);
  BUFF I4 (joint_0[0:0], i_1r1[0:0]);
  BUFF I5 (joint_0[1:1], i_1r1[1:1]);
  BUFF I6 (joint_0[2:2], i_1r1[2:2]);
  BUFF I7 (joint_0[3:3], i_1r1[3:3]);
  BUFF I8 (icomplete_0, i_0r);
  C2 I9 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I10 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I11 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I12 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I13 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I14 (o_0r1[1:1], joint_0[1:1]);
  BUFF I15 (o_0r1[2:2], joint_0[2:2]);
  BUFF I16 (o_0r1[3:3], joint_0[3:3]);
  BUFF I17 (i_0a, o_0a);
  BUFF I18 (i_1a, o_0a);
endmodule

// tks4_o0w4_1o0w0_2o0w0_4o0w0_8o0w0 TeakS (0+:4) [([Imp 1 0],0),([Imp 2 0],0),([Imp 4 0],0),([Imp 8 0]
//   ,0)] [One 4,Many [0,0,0,0]]
module tks4_o0w4_1o0w0_2o0w0_4o0w0_8o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire oack_0;
  wire match0_0;
  wire [1:0] simp121_0;
  wire match1_0;
  wire [1:0] simp151_0;
  wire match2_0;
  wire [1:0] simp181_0;
  wire match3_0;
  wire [1:0] simp211_0;
  wire [3:0] comp_0;
  wire [1:0] simp311_0;
  wire [1:0] simp361_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (simp121_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I2 (simp121_0[1:1], i_0r0[3:3]);
  C2 I3 (match0_0, simp121_0[0:0], simp121_0[1:1]);
  BUFF I4 (sel_1, match1_0);
  C3 I5 (simp151_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I6 (simp151_0[1:1], i_0r0[3:3]);
  C2 I7 (match1_0, simp151_0[0:0], simp151_0[1:1]);
  BUFF I8 (sel_2, match2_0);
  C3 I9 (simp181_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I10 (simp181_0[1:1], i_0r0[3:3]);
  C2 I11 (match2_0, simp181_0[0:0], simp181_0[1:1]);
  BUFF I12 (sel_3, match3_0);
  C3 I13 (simp211_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I14 (simp211_0[1:1], i_0r1[3:3]);
  C2 I15 (match3_0, simp211_0[0:0], simp211_0[1:1]);
  C2 I16 (gsel_0, sel_0, icomplete_0);
  C2 I17 (gsel_1, sel_1, icomplete_0);
  C2 I18 (gsel_2, sel_2, icomplete_0);
  C2 I19 (gsel_3, sel_3, icomplete_0);
  OR2 I20 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I21 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I22 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I23 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  C3 I24 (simp311_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  BUFF I25 (simp311_0[1:1], comp_0[3:3]);
  C2 I26 (icomplete_0, simp311_0[0:0], simp311_0[1:1]);
  BUFF I27 (o_0r, gsel_0);
  BUFF I28 (o_1r, gsel_1);
  BUFF I29 (o_2r, gsel_2);
  BUFF I30 (o_3r, gsel_3);
  NOR3 I31 (simp361_0[0:0], o_0a, o_1a, o_2a);
  INV I32 (simp361_0[1:1], o_3a);
  NAND2 I33 (oack_0, simp361_0[0:0], simp361_0[1:1]);
  C2 I34 (i_0a, oack_0, icomplete_0);
endmodule

// tkvir65_wo0w65_ro0w22o25w5o0w22o25w4o22w3o19w6o13w1o0w13o19w6o25w5o25w5o0w5o14w5o13w1o13w1o0w13o19w6
//   o25w5o0w5o14w5o13w1o19w6o30w2o32w33 TeakV "ir" 65 [] [0] [0,25,0,25,22,19,13,0,19,25,25,0,14,13,13,0
//   ,19,25,0,14,13,19,30,32] [Many [65],Many [0],Many [0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0],
//   Many [22,5,22,4,3,6,1,13,6,5,5,5,5,1,1,13,6,5,5,5,1,6,2,33]]
module tkvir65_wo0w65_ro0w22o25w5o0w22o25w4o22w3o19w6o13w1o0w13o19w6o25w5o25w5o0w5o14w5o13w1o13w1o0w13o19w6o25w5o0w5o14w5o13w1o19w6o30w2o32w33 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rg_5r, rg_5a, rg_6r, rg_6a, rg_7r, rg_7a, rg_8r, rg_8a, rg_9r, rg_9a, rg_10r, rg_10a, rg_11r, rg_11a, rg_12r, rg_12a, rg_13r, rg_13a, rg_14r, rg_14a, rg_15r, rg_15a, rg_16r, rg_16a, rg_17r, rg_17a, rg_18r, rg_18a, rg_19r, rg_19a, rg_20r, rg_20a, rg_21r, rg_21a, rg_22r, rg_22a, rg_23r, rg_23a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, rd_5r0, rd_5r1, rd_5a, rd_6r0, rd_6r1, rd_6a, rd_7r0, rd_7r1, rd_7a, rd_8r0, rd_8r1, rd_8a, rd_9r0, rd_9r1, rd_9a, rd_10r0, rd_10r1, rd_10a, rd_11r0, rd_11r1, rd_11a, rd_12r0, rd_12r1, rd_12a, rd_13r0, rd_13r1, rd_13a, rd_14r0, rd_14r1, rd_14a, rd_15r0, rd_15r1, rd_15a, rd_16r0, rd_16r1, rd_16a, rd_17r0, rd_17r1, rd_17a, rd_18r0, rd_18r1, rd_18a, rd_19r0, rd_19r1, rd_19a, rd_20r0, rd_20r1, rd_20a, rd_21r0, rd_21r1, rd_21a, rd_22r0, rd_22r1, rd_22a, rd_23r0, rd_23r1, rd_23a, reset);
  input [64:0] wg_0r0;
  input [64:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  input rg_5r;
  output rg_5a;
  input rg_6r;
  output rg_6a;
  input rg_7r;
  output rg_7a;
  input rg_8r;
  output rg_8a;
  input rg_9r;
  output rg_9a;
  input rg_10r;
  output rg_10a;
  input rg_11r;
  output rg_11a;
  input rg_12r;
  output rg_12a;
  input rg_13r;
  output rg_13a;
  input rg_14r;
  output rg_14a;
  input rg_15r;
  output rg_15a;
  input rg_16r;
  output rg_16a;
  input rg_17r;
  output rg_17a;
  input rg_18r;
  output rg_18a;
  input rg_19r;
  output rg_19a;
  input rg_20r;
  output rg_20a;
  input rg_21r;
  output rg_21a;
  input rg_22r;
  output rg_22a;
  input rg_23r;
  output rg_23a;
  output [21:0] rd_0r0;
  output [21:0] rd_0r1;
  input rd_0a;
  output [4:0] rd_1r0;
  output [4:0] rd_1r1;
  input rd_1a;
  output [21:0] rd_2r0;
  output [21:0] rd_2r1;
  input rd_2a;
  output [3:0] rd_3r0;
  output [3:0] rd_3r1;
  input rd_3a;
  output [2:0] rd_4r0;
  output [2:0] rd_4r1;
  input rd_4a;
  output [5:0] rd_5r0;
  output [5:0] rd_5r1;
  input rd_5a;
  output rd_6r0;
  output rd_6r1;
  input rd_6a;
  output [12:0] rd_7r0;
  output [12:0] rd_7r1;
  input rd_7a;
  output [5:0] rd_8r0;
  output [5:0] rd_8r1;
  input rd_8a;
  output [4:0] rd_9r0;
  output [4:0] rd_9r1;
  input rd_9a;
  output [4:0] rd_10r0;
  output [4:0] rd_10r1;
  input rd_10a;
  output [4:0] rd_11r0;
  output [4:0] rd_11r1;
  input rd_11a;
  output [4:0] rd_12r0;
  output [4:0] rd_12r1;
  input rd_12a;
  output rd_13r0;
  output rd_13r1;
  input rd_13a;
  output rd_14r0;
  output rd_14r1;
  input rd_14a;
  output [12:0] rd_15r0;
  output [12:0] rd_15r1;
  input rd_15a;
  output [5:0] rd_16r0;
  output [5:0] rd_16r1;
  input rd_16a;
  output [4:0] rd_17r0;
  output [4:0] rd_17r1;
  input rd_17a;
  output [4:0] rd_18r0;
  output [4:0] rd_18r1;
  input rd_18a;
  output [4:0] rd_19r0;
  output [4:0] rd_19r1;
  input rd_19a;
  output rd_20r0;
  output rd_20r1;
  input rd_20a;
  output [5:0] rd_21r0;
  output [5:0] rd_21r1;
  input rd_21a;
  output [1:0] rd_22r0;
  output [1:0] rd_22r1;
  input rd_22a;
  output [32:0] rd_23r0;
  output [32:0] rd_23r1;
  input rd_23a;
  input reset;
  wire [64:0] wf_0;
  wire [64:0] wt_0;
  wire [64:0] df_0;
  wire [64:0] dt_0;
  wire wc_0;
  wire [64:0] wacks_0;
  wire [64:0] wenr_0;
  wire [64:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [64:0] drlgf_0;
  wire [64:0] drlgt_0;
  wire [64:0] comp0_0;
  wire [21:0] simp4691_0;
  wire [7:0] simp4692_0;
  wire [2:0] simp4693_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [64:0] conwgit_0;
  wire [64:0] conwgif_0;
  wire conwig_0;
  wire [21:0] simp8031_0;
  wire [7:0] simp8032_0;
  wire [2:0] simp8033_0;
  wire [15:0] simp11641_0;
  wire [5:0] simp11642_0;
  wire [1:0] simp11643_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (wen_0[32:32], wenr_0[32:32], nreset_0);
  AND2 I34 (wen_0[33:33], wenr_0[33:33], nreset_0);
  AND2 I35 (wen_0[34:34], wenr_0[34:34], nreset_0);
  AND2 I36 (wen_0[35:35], wenr_0[35:35], nreset_0);
  AND2 I37 (wen_0[36:36], wenr_0[36:36], nreset_0);
  AND2 I38 (wen_0[37:37], wenr_0[37:37], nreset_0);
  AND2 I39 (wen_0[38:38], wenr_0[38:38], nreset_0);
  AND2 I40 (wen_0[39:39], wenr_0[39:39], nreset_0);
  AND2 I41 (wen_0[40:40], wenr_0[40:40], nreset_0);
  AND2 I42 (wen_0[41:41], wenr_0[41:41], nreset_0);
  AND2 I43 (wen_0[42:42], wenr_0[42:42], nreset_0);
  AND2 I44 (wen_0[43:43], wenr_0[43:43], nreset_0);
  AND2 I45 (wen_0[44:44], wenr_0[44:44], nreset_0);
  AND2 I46 (wen_0[45:45], wenr_0[45:45], nreset_0);
  AND2 I47 (wen_0[46:46], wenr_0[46:46], nreset_0);
  AND2 I48 (wen_0[47:47], wenr_0[47:47], nreset_0);
  AND2 I49 (wen_0[48:48], wenr_0[48:48], nreset_0);
  AND2 I50 (wen_0[49:49], wenr_0[49:49], nreset_0);
  AND2 I51 (wen_0[50:50], wenr_0[50:50], nreset_0);
  AND2 I52 (wen_0[51:51], wenr_0[51:51], nreset_0);
  AND2 I53 (wen_0[52:52], wenr_0[52:52], nreset_0);
  AND2 I54 (wen_0[53:53], wenr_0[53:53], nreset_0);
  AND2 I55 (wen_0[54:54], wenr_0[54:54], nreset_0);
  AND2 I56 (wen_0[55:55], wenr_0[55:55], nreset_0);
  AND2 I57 (wen_0[56:56], wenr_0[56:56], nreset_0);
  AND2 I58 (wen_0[57:57], wenr_0[57:57], nreset_0);
  AND2 I59 (wen_0[58:58], wenr_0[58:58], nreset_0);
  AND2 I60 (wen_0[59:59], wenr_0[59:59], nreset_0);
  AND2 I61 (wen_0[60:60], wenr_0[60:60], nreset_0);
  AND2 I62 (wen_0[61:61], wenr_0[61:61], nreset_0);
  AND2 I63 (wen_0[62:62], wenr_0[62:62], nreset_0);
  AND2 I64 (wen_0[63:63], wenr_0[63:63], nreset_0);
  AND2 I65 (wen_0[64:64], wenr_0[64:64], nreset_0);
  AND2 I66 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I67 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I68 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I69 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I70 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I71 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I72 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I73 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I74 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I75 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I76 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I77 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I78 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I79 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I80 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I81 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I82 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I83 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I84 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I85 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I86 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I87 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I88 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I89 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I90 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I91 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I92 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I93 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I94 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I95 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I96 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I97 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I98 (drlgf_0[32:32], wf_0[32:32], wen_0[32:32]);
  AND2 I99 (drlgf_0[33:33], wf_0[33:33], wen_0[33:33]);
  AND2 I100 (drlgf_0[34:34], wf_0[34:34], wen_0[34:34]);
  AND2 I101 (drlgf_0[35:35], wf_0[35:35], wen_0[35:35]);
  AND2 I102 (drlgf_0[36:36], wf_0[36:36], wen_0[36:36]);
  AND2 I103 (drlgf_0[37:37], wf_0[37:37], wen_0[37:37]);
  AND2 I104 (drlgf_0[38:38], wf_0[38:38], wen_0[38:38]);
  AND2 I105 (drlgf_0[39:39], wf_0[39:39], wen_0[39:39]);
  AND2 I106 (drlgf_0[40:40], wf_0[40:40], wen_0[40:40]);
  AND2 I107 (drlgf_0[41:41], wf_0[41:41], wen_0[41:41]);
  AND2 I108 (drlgf_0[42:42], wf_0[42:42], wen_0[42:42]);
  AND2 I109 (drlgf_0[43:43], wf_0[43:43], wen_0[43:43]);
  AND2 I110 (drlgf_0[44:44], wf_0[44:44], wen_0[44:44]);
  AND2 I111 (drlgf_0[45:45], wf_0[45:45], wen_0[45:45]);
  AND2 I112 (drlgf_0[46:46], wf_0[46:46], wen_0[46:46]);
  AND2 I113 (drlgf_0[47:47], wf_0[47:47], wen_0[47:47]);
  AND2 I114 (drlgf_0[48:48], wf_0[48:48], wen_0[48:48]);
  AND2 I115 (drlgf_0[49:49], wf_0[49:49], wen_0[49:49]);
  AND2 I116 (drlgf_0[50:50], wf_0[50:50], wen_0[50:50]);
  AND2 I117 (drlgf_0[51:51], wf_0[51:51], wen_0[51:51]);
  AND2 I118 (drlgf_0[52:52], wf_0[52:52], wen_0[52:52]);
  AND2 I119 (drlgf_0[53:53], wf_0[53:53], wen_0[53:53]);
  AND2 I120 (drlgf_0[54:54], wf_0[54:54], wen_0[54:54]);
  AND2 I121 (drlgf_0[55:55], wf_0[55:55], wen_0[55:55]);
  AND2 I122 (drlgf_0[56:56], wf_0[56:56], wen_0[56:56]);
  AND2 I123 (drlgf_0[57:57], wf_0[57:57], wen_0[57:57]);
  AND2 I124 (drlgf_0[58:58], wf_0[58:58], wen_0[58:58]);
  AND2 I125 (drlgf_0[59:59], wf_0[59:59], wen_0[59:59]);
  AND2 I126 (drlgf_0[60:60], wf_0[60:60], wen_0[60:60]);
  AND2 I127 (drlgf_0[61:61], wf_0[61:61], wen_0[61:61]);
  AND2 I128 (drlgf_0[62:62], wf_0[62:62], wen_0[62:62]);
  AND2 I129 (drlgf_0[63:63], wf_0[63:63], wen_0[63:63]);
  AND2 I130 (drlgf_0[64:64], wf_0[64:64], wen_0[64:64]);
  AND2 I131 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I132 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I133 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I134 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I135 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I136 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I137 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I138 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I139 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I140 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I141 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I142 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I143 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I144 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I145 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I146 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I147 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I148 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I149 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I150 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I151 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I152 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I153 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I154 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I155 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I156 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I157 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I158 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I159 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I160 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I161 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I162 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  AND2 I163 (drlgt_0[32:32], wt_0[32:32], wen_0[32:32]);
  AND2 I164 (drlgt_0[33:33], wt_0[33:33], wen_0[33:33]);
  AND2 I165 (drlgt_0[34:34], wt_0[34:34], wen_0[34:34]);
  AND2 I166 (drlgt_0[35:35], wt_0[35:35], wen_0[35:35]);
  AND2 I167 (drlgt_0[36:36], wt_0[36:36], wen_0[36:36]);
  AND2 I168 (drlgt_0[37:37], wt_0[37:37], wen_0[37:37]);
  AND2 I169 (drlgt_0[38:38], wt_0[38:38], wen_0[38:38]);
  AND2 I170 (drlgt_0[39:39], wt_0[39:39], wen_0[39:39]);
  AND2 I171 (drlgt_0[40:40], wt_0[40:40], wen_0[40:40]);
  AND2 I172 (drlgt_0[41:41], wt_0[41:41], wen_0[41:41]);
  AND2 I173 (drlgt_0[42:42], wt_0[42:42], wen_0[42:42]);
  AND2 I174 (drlgt_0[43:43], wt_0[43:43], wen_0[43:43]);
  AND2 I175 (drlgt_0[44:44], wt_0[44:44], wen_0[44:44]);
  AND2 I176 (drlgt_0[45:45], wt_0[45:45], wen_0[45:45]);
  AND2 I177 (drlgt_0[46:46], wt_0[46:46], wen_0[46:46]);
  AND2 I178 (drlgt_0[47:47], wt_0[47:47], wen_0[47:47]);
  AND2 I179 (drlgt_0[48:48], wt_0[48:48], wen_0[48:48]);
  AND2 I180 (drlgt_0[49:49], wt_0[49:49], wen_0[49:49]);
  AND2 I181 (drlgt_0[50:50], wt_0[50:50], wen_0[50:50]);
  AND2 I182 (drlgt_0[51:51], wt_0[51:51], wen_0[51:51]);
  AND2 I183 (drlgt_0[52:52], wt_0[52:52], wen_0[52:52]);
  AND2 I184 (drlgt_0[53:53], wt_0[53:53], wen_0[53:53]);
  AND2 I185 (drlgt_0[54:54], wt_0[54:54], wen_0[54:54]);
  AND2 I186 (drlgt_0[55:55], wt_0[55:55], wen_0[55:55]);
  AND2 I187 (drlgt_0[56:56], wt_0[56:56], wen_0[56:56]);
  AND2 I188 (drlgt_0[57:57], wt_0[57:57], wen_0[57:57]);
  AND2 I189 (drlgt_0[58:58], wt_0[58:58], wen_0[58:58]);
  AND2 I190 (drlgt_0[59:59], wt_0[59:59], wen_0[59:59]);
  AND2 I191 (drlgt_0[60:60], wt_0[60:60], wen_0[60:60]);
  AND2 I192 (drlgt_0[61:61], wt_0[61:61], wen_0[61:61]);
  AND2 I193 (drlgt_0[62:62], wt_0[62:62], wen_0[62:62]);
  AND2 I194 (drlgt_0[63:63], wt_0[63:63], wen_0[63:63]);
  AND2 I195 (drlgt_0[64:64], wt_0[64:64], wen_0[64:64]);
  NOR2 I196 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I197 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I198 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I199 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I200 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I201 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I202 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I203 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I204 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I205 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I206 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I207 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I208 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I209 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I210 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I211 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I212 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I213 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I214 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I215 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I216 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I217 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I218 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I219 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I220 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I221 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I222 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I223 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I224 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I225 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I226 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I227 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR2 I228 (df_0[32:32], dt_0[32:32], drlgt_0[32:32]);
  NOR2 I229 (df_0[33:33], dt_0[33:33], drlgt_0[33:33]);
  NOR2 I230 (df_0[34:34], dt_0[34:34], drlgt_0[34:34]);
  NOR2 I231 (df_0[35:35], dt_0[35:35], drlgt_0[35:35]);
  NOR2 I232 (df_0[36:36], dt_0[36:36], drlgt_0[36:36]);
  NOR2 I233 (df_0[37:37], dt_0[37:37], drlgt_0[37:37]);
  NOR2 I234 (df_0[38:38], dt_0[38:38], drlgt_0[38:38]);
  NOR2 I235 (df_0[39:39], dt_0[39:39], drlgt_0[39:39]);
  NOR2 I236 (df_0[40:40], dt_0[40:40], drlgt_0[40:40]);
  NOR2 I237 (df_0[41:41], dt_0[41:41], drlgt_0[41:41]);
  NOR2 I238 (df_0[42:42], dt_0[42:42], drlgt_0[42:42]);
  NOR2 I239 (df_0[43:43], dt_0[43:43], drlgt_0[43:43]);
  NOR2 I240 (df_0[44:44], dt_0[44:44], drlgt_0[44:44]);
  NOR2 I241 (df_0[45:45], dt_0[45:45], drlgt_0[45:45]);
  NOR2 I242 (df_0[46:46], dt_0[46:46], drlgt_0[46:46]);
  NOR2 I243 (df_0[47:47], dt_0[47:47], drlgt_0[47:47]);
  NOR2 I244 (df_0[48:48], dt_0[48:48], drlgt_0[48:48]);
  NOR2 I245 (df_0[49:49], dt_0[49:49], drlgt_0[49:49]);
  NOR2 I246 (df_0[50:50], dt_0[50:50], drlgt_0[50:50]);
  NOR2 I247 (df_0[51:51], dt_0[51:51], drlgt_0[51:51]);
  NOR2 I248 (df_0[52:52], dt_0[52:52], drlgt_0[52:52]);
  NOR2 I249 (df_0[53:53], dt_0[53:53], drlgt_0[53:53]);
  NOR2 I250 (df_0[54:54], dt_0[54:54], drlgt_0[54:54]);
  NOR2 I251 (df_0[55:55], dt_0[55:55], drlgt_0[55:55]);
  NOR2 I252 (df_0[56:56], dt_0[56:56], drlgt_0[56:56]);
  NOR2 I253 (df_0[57:57], dt_0[57:57], drlgt_0[57:57]);
  NOR2 I254 (df_0[58:58], dt_0[58:58], drlgt_0[58:58]);
  NOR2 I255 (df_0[59:59], dt_0[59:59], drlgt_0[59:59]);
  NOR2 I256 (df_0[60:60], dt_0[60:60], drlgt_0[60:60]);
  NOR2 I257 (df_0[61:61], dt_0[61:61], drlgt_0[61:61]);
  NOR2 I258 (df_0[62:62], dt_0[62:62], drlgt_0[62:62]);
  NOR2 I259 (df_0[63:63], dt_0[63:63], drlgt_0[63:63]);
  NOR2 I260 (df_0[64:64], dt_0[64:64], drlgt_0[64:64]);
  NOR3 I261 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I262 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I263 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I264 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I265 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I266 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I267 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I268 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I269 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I270 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I271 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I272 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I273 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I274 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I275 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I276 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I277 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I278 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I279 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I280 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I281 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I282 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I283 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I284 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I285 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I286 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I287 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I288 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I289 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I290 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I291 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I292 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  NOR3 I293 (dt_0[32:32], df_0[32:32], drlgf_0[32:32], reset);
  NOR3 I294 (dt_0[33:33], df_0[33:33], drlgf_0[33:33], reset);
  NOR3 I295 (dt_0[34:34], df_0[34:34], drlgf_0[34:34], reset);
  NOR3 I296 (dt_0[35:35], df_0[35:35], drlgf_0[35:35], reset);
  NOR3 I297 (dt_0[36:36], df_0[36:36], drlgf_0[36:36], reset);
  NOR3 I298 (dt_0[37:37], df_0[37:37], drlgf_0[37:37], reset);
  NOR3 I299 (dt_0[38:38], df_0[38:38], drlgf_0[38:38], reset);
  NOR3 I300 (dt_0[39:39], df_0[39:39], drlgf_0[39:39], reset);
  NOR3 I301 (dt_0[40:40], df_0[40:40], drlgf_0[40:40], reset);
  NOR3 I302 (dt_0[41:41], df_0[41:41], drlgf_0[41:41], reset);
  NOR3 I303 (dt_0[42:42], df_0[42:42], drlgf_0[42:42], reset);
  NOR3 I304 (dt_0[43:43], df_0[43:43], drlgf_0[43:43], reset);
  NOR3 I305 (dt_0[44:44], df_0[44:44], drlgf_0[44:44], reset);
  NOR3 I306 (dt_0[45:45], df_0[45:45], drlgf_0[45:45], reset);
  NOR3 I307 (dt_0[46:46], df_0[46:46], drlgf_0[46:46], reset);
  NOR3 I308 (dt_0[47:47], df_0[47:47], drlgf_0[47:47], reset);
  NOR3 I309 (dt_0[48:48], df_0[48:48], drlgf_0[48:48], reset);
  NOR3 I310 (dt_0[49:49], df_0[49:49], drlgf_0[49:49], reset);
  NOR3 I311 (dt_0[50:50], df_0[50:50], drlgf_0[50:50], reset);
  NOR3 I312 (dt_0[51:51], df_0[51:51], drlgf_0[51:51], reset);
  NOR3 I313 (dt_0[52:52], df_0[52:52], drlgf_0[52:52], reset);
  NOR3 I314 (dt_0[53:53], df_0[53:53], drlgf_0[53:53], reset);
  NOR3 I315 (dt_0[54:54], df_0[54:54], drlgf_0[54:54], reset);
  NOR3 I316 (dt_0[55:55], df_0[55:55], drlgf_0[55:55], reset);
  NOR3 I317 (dt_0[56:56], df_0[56:56], drlgf_0[56:56], reset);
  NOR3 I318 (dt_0[57:57], df_0[57:57], drlgf_0[57:57], reset);
  NOR3 I319 (dt_0[58:58], df_0[58:58], drlgf_0[58:58], reset);
  NOR3 I320 (dt_0[59:59], df_0[59:59], drlgf_0[59:59], reset);
  NOR3 I321 (dt_0[60:60], df_0[60:60], drlgf_0[60:60], reset);
  NOR3 I322 (dt_0[61:61], df_0[61:61], drlgf_0[61:61], reset);
  NOR3 I323 (dt_0[62:62], df_0[62:62], drlgf_0[62:62], reset);
  NOR3 I324 (dt_0[63:63], df_0[63:63], drlgf_0[63:63], reset);
  NOR3 I325 (dt_0[64:64], df_0[64:64], drlgf_0[64:64], reset);
  AO22 I326 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I327 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I328 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I329 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I330 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I331 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I332 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I333 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I334 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I335 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I336 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I337 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I338 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I339 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I340 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I341 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I342 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I343 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I344 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I345 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I346 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I347 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I348 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I349 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I350 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I351 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I352 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I353 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I354 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I355 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I356 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I357 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  AO22 I358 (wacks_0[32:32], drlgf_0[32:32], df_0[32:32], drlgt_0[32:32], dt_0[32:32]);
  AO22 I359 (wacks_0[33:33], drlgf_0[33:33], df_0[33:33], drlgt_0[33:33], dt_0[33:33]);
  AO22 I360 (wacks_0[34:34], drlgf_0[34:34], df_0[34:34], drlgt_0[34:34], dt_0[34:34]);
  AO22 I361 (wacks_0[35:35], drlgf_0[35:35], df_0[35:35], drlgt_0[35:35], dt_0[35:35]);
  AO22 I362 (wacks_0[36:36], drlgf_0[36:36], df_0[36:36], drlgt_0[36:36], dt_0[36:36]);
  AO22 I363 (wacks_0[37:37], drlgf_0[37:37], df_0[37:37], drlgt_0[37:37], dt_0[37:37]);
  AO22 I364 (wacks_0[38:38], drlgf_0[38:38], df_0[38:38], drlgt_0[38:38], dt_0[38:38]);
  AO22 I365 (wacks_0[39:39], drlgf_0[39:39], df_0[39:39], drlgt_0[39:39], dt_0[39:39]);
  AO22 I366 (wacks_0[40:40], drlgf_0[40:40], df_0[40:40], drlgt_0[40:40], dt_0[40:40]);
  AO22 I367 (wacks_0[41:41], drlgf_0[41:41], df_0[41:41], drlgt_0[41:41], dt_0[41:41]);
  AO22 I368 (wacks_0[42:42], drlgf_0[42:42], df_0[42:42], drlgt_0[42:42], dt_0[42:42]);
  AO22 I369 (wacks_0[43:43], drlgf_0[43:43], df_0[43:43], drlgt_0[43:43], dt_0[43:43]);
  AO22 I370 (wacks_0[44:44], drlgf_0[44:44], df_0[44:44], drlgt_0[44:44], dt_0[44:44]);
  AO22 I371 (wacks_0[45:45], drlgf_0[45:45], df_0[45:45], drlgt_0[45:45], dt_0[45:45]);
  AO22 I372 (wacks_0[46:46], drlgf_0[46:46], df_0[46:46], drlgt_0[46:46], dt_0[46:46]);
  AO22 I373 (wacks_0[47:47], drlgf_0[47:47], df_0[47:47], drlgt_0[47:47], dt_0[47:47]);
  AO22 I374 (wacks_0[48:48], drlgf_0[48:48], df_0[48:48], drlgt_0[48:48], dt_0[48:48]);
  AO22 I375 (wacks_0[49:49], drlgf_0[49:49], df_0[49:49], drlgt_0[49:49], dt_0[49:49]);
  AO22 I376 (wacks_0[50:50], drlgf_0[50:50], df_0[50:50], drlgt_0[50:50], dt_0[50:50]);
  AO22 I377 (wacks_0[51:51], drlgf_0[51:51], df_0[51:51], drlgt_0[51:51], dt_0[51:51]);
  AO22 I378 (wacks_0[52:52], drlgf_0[52:52], df_0[52:52], drlgt_0[52:52], dt_0[52:52]);
  AO22 I379 (wacks_0[53:53], drlgf_0[53:53], df_0[53:53], drlgt_0[53:53], dt_0[53:53]);
  AO22 I380 (wacks_0[54:54], drlgf_0[54:54], df_0[54:54], drlgt_0[54:54], dt_0[54:54]);
  AO22 I381 (wacks_0[55:55], drlgf_0[55:55], df_0[55:55], drlgt_0[55:55], dt_0[55:55]);
  AO22 I382 (wacks_0[56:56], drlgf_0[56:56], df_0[56:56], drlgt_0[56:56], dt_0[56:56]);
  AO22 I383 (wacks_0[57:57], drlgf_0[57:57], df_0[57:57], drlgt_0[57:57], dt_0[57:57]);
  AO22 I384 (wacks_0[58:58], drlgf_0[58:58], df_0[58:58], drlgt_0[58:58], dt_0[58:58]);
  AO22 I385 (wacks_0[59:59], drlgf_0[59:59], df_0[59:59], drlgt_0[59:59], dt_0[59:59]);
  AO22 I386 (wacks_0[60:60], drlgf_0[60:60], df_0[60:60], drlgt_0[60:60], dt_0[60:60]);
  AO22 I387 (wacks_0[61:61], drlgf_0[61:61], df_0[61:61], drlgt_0[61:61], dt_0[61:61]);
  AO22 I388 (wacks_0[62:62], drlgf_0[62:62], df_0[62:62], drlgt_0[62:62], dt_0[62:62]);
  AO22 I389 (wacks_0[63:63], drlgf_0[63:63], df_0[63:63], drlgt_0[63:63], dt_0[63:63]);
  AO22 I390 (wacks_0[64:64], drlgf_0[64:64], df_0[64:64], drlgt_0[64:64], dt_0[64:64]);
  OR2 I391 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I392 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I393 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I394 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I395 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I396 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I397 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I398 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I399 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I400 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I401 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I402 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I403 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I404 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I405 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I406 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I407 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I408 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I409 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I410 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I411 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I412 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I413 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I414 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I415 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I416 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I417 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I418 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I419 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I420 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I421 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I422 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  OR2 I423 (comp0_0[32:32], wg_0r0[32:32], wg_0r1[32:32]);
  OR2 I424 (comp0_0[33:33], wg_0r0[33:33], wg_0r1[33:33]);
  OR2 I425 (comp0_0[34:34], wg_0r0[34:34], wg_0r1[34:34]);
  OR2 I426 (comp0_0[35:35], wg_0r0[35:35], wg_0r1[35:35]);
  OR2 I427 (comp0_0[36:36], wg_0r0[36:36], wg_0r1[36:36]);
  OR2 I428 (comp0_0[37:37], wg_0r0[37:37], wg_0r1[37:37]);
  OR2 I429 (comp0_0[38:38], wg_0r0[38:38], wg_0r1[38:38]);
  OR2 I430 (comp0_0[39:39], wg_0r0[39:39], wg_0r1[39:39]);
  OR2 I431 (comp0_0[40:40], wg_0r0[40:40], wg_0r1[40:40]);
  OR2 I432 (comp0_0[41:41], wg_0r0[41:41], wg_0r1[41:41]);
  OR2 I433 (comp0_0[42:42], wg_0r0[42:42], wg_0r1[42:42]);
  OR2 I434 (comp0_0[43:43], wg_0r0[43:43], wg_0r1[43:43]);
  OR2 I435 (comp0_0[44:44], wg_0r0[44:44], wg_0r1[44:44]);
  OR2 I436 (comp0_0[45:45], wg_0r0[45:45], wg_0r1[45:45]);
  OR2 I437 (comp0_0[46:46], wg_0r0[46:46], wg_0r1[46:46]);
  OR2 I438 (comp0_0[47:47], wg_0r0[47:47], wg_0r1[47:47]);
  OR2 I439 (comp0_0[48:48], wg_0r0[48:48], wg_0r1[48:48]);
  OR2 I440 (comp0_0[49:49], wg_0r0[49:49], wg_0r1[49:49]);
  OR2 I441 (comp0_0[50:50], wg_0r0[50:50], wg_0r1[50:50]);
  OR2 I442 (comp0_0[51:51], wg_0r0[51:51], wg_0r1[51:51]);
  OR2 I443 (comp0_0[52:52], wg_0r0[52:52], wg_0r1[52:52]);
  OR2 I444 (comp0_0[53:53], wg_0r0[53:53], wg_0r1[53:53]);
  OR2 I445 (comp0_0[54:54], wg_0r0[54:54], wg_0r1[54:54]);
  OR2 I446 (comp0_0[55:55], wg_0r0[55:55], wg_0r1[55:55]);
  OR2 I447 (comp0_0[56:56], wg_0r0[56:56], wg_0r1[56:56]);
  OR2 I448 (comp0_0[57:57], wg_0r0[57:57], wg_0r1[57:57]);
  OR2 I449 (comp0_0[58:58], wg_0r0[58:58], wg_0r1[58:58]);
  OR2 I450 (comp0_0[59:59], wg_0r0[59:59], wg_0r1[59:59]);
  OR2 I451 (comp0_0[60:60], wg_0r0[60:60], wg_0r1[60:60]);
  OR2 I452 (comp0_0[61:61], wg_0r0[61:61], wg_0r1[61:61]);
  OR2 I453 (comp0_0[62:62], wg_0r0[62:62], wg_0r1[62:62]);
  OR2 I454 (comp0_0[63:63], wg_0r0[63:63], wg_0r1[63:63]);
  OR2 I455 (comp0_0[64:64], wg_0r0[64:64], wg_0r1[64:64]);
  C3 I456 (simp4691_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I457 (simp4691_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I458 (simp4691_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I459 (simp4691_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I460 (simp4691_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I461 (simp4691_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I462 (simp4691_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I463 (simp4691_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I464 (simp4691_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I465 (simp4691_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C3 I466 (simp4691_0[10:10], comp0_0[30:30], comp0_0[31:31], comp0_0[32:32]);
  C3 I467 (simp4691_0[11:11], comp0_0[33:33], comp0_0[34:34], comp0_0[35:35]);
  C3 I468 (simp4691_0[12:12], comp0_0[36:36], comp0_0[37:37], comp0_0[38:38]);
  C3 I469 (simp4691_0[13:13], comp0_0[39:39], comp0_0[40:40], comp0_0[41:41]);
  C3 I470 (simp4691_0[14:14], comp0_0[42:42], comp0_0[43:43], comp0_0[44:44]);
  C3 I471 (simp4691_0[15:15], comp0_0[45:45], comp0_0[46:46], comp0_0[47:47]);
  C3 I472 (simp4691_0[16:16], comp0_0[48:48], comp0_0[49:49], comp0_0[50:50]);
  C3 I473 (simp4691_0[17:17], comp0_0[51:51], comp0_0[52:52], comp0_0[53:53]);
  C3 I474 (simp4691_0[18:18], comp0_0[54:54], comp0_0[55:55], comp0_0[56:56]);
  C3 I475 (simp4691_0[19:19], comp0_0[57:57], comp0_0[58:58], comp0_0[59:59]);
  C3 I476 (simp4691_0[20:20], comp0_0[60:60], comp0_0[61:61], comp0_0[62:62]);
  C2 I477 (simp4691_0[21:21], comp0_0[63:63], comp0_0[64:64]);
  C3 I478 (simp4692_0[0:0], simp4691_0[0:0], simp4691_0[1:1], simp4691_0[2:2]);
  C3 I479 (simp4692_0[1:1], simp4691_0[3:3], simp4691_0[4:4], simp4691_0[5:5]);
  C3 I480 (simp4692_0[2:2], simp4691_0[6:6], simp4691_0[7:7], simp4691_0[8:8]);
  C3 I481 (simp4692_0[3:3], simp4691_0[9:9], simp4691_0[10:10], simp4691_0[11:11]);
  C3 I482 (simp4692_0[4:4], simp4691_0[12:12], simp4691_0[13:13], simp4691_0[14:14]);
  C3 I483 (simp4692_0[5:5], simp4691_0[15:15], simp4691_0[16:16], simp4691_0[17:17]);
  C3 I484 (simp4692_0[6:6], simp4691_0[18:18], simp4691_0[19:19], simp4691_0[20:20]);
  BUFF I485 (simp4692_0[7:7], simp4691_0[21:21]);
  C3 I486 (simp4693_0[0:0], simp4692_0[0:0], simp4692_0[1:1], simp4692_0[2:2]);
  C3 I487 (simp4693_0[1:1], simp4692_0[3:3], simp4692_0[4:4], simp4692_0[5:5]);
  C2 I488 (simp4693_0[2:2], simp4692_0[6:6], simp4692_0[7:7]);
  C3 I489 (wc_0, simp4693_0[0:0], simp4693_0[1:1], simp4693_0[2:2]);
  AND2 I490 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I491 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I492 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I493 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I494 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I495 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I496 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I497 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I498 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I499 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I500 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I501 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I502 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I503 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I504 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I505 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I506 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I507 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I508 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I509 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I510 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I511 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I512 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I513 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I514 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I515 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I516 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I517 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I518 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I519 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I520 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I521 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I522 (conwgif_0[32:32], wg_0r0[32:32], conwig_0);
  AND2 I523 (conwgif_0[33:33], wg_0r0[33:33], conwig_0);
  AND2 I524 (conwgif_0[34:34], wg_0r0[34:34], conwig_0);
  AND2 I525 (conwgif_0[35:35], wg_0r0[35:35], conwig_0);
  AND2 I526 (conwgif_0[36:36], wg_0r0[36:36], conwig_0);
  AND2 I527 (conwgif_0[37:37], wg_0r0[37:37], conwig_0);
  AND2 I528 (conwgif_0[38:38], wg_0r0[38:38], conwig_0);
  AND2 I529 (conwgif_0[39:39], wg_0r0[39:39], conwig_0);
  AND2 I530 (conwgif_0[40:40], wg_0r0[40:40], conwig_0);
  AND2 I531 (conwgif_0[41:41], wg_0r0[41:41], conwig_0);
  AND2 I532 (conwgif_0[42:42], wg_0r0[42:42], conwig_0);
  AND2 I533 (conwgif_0[43:43], wg_0r0[43:43], conwig_0);
  AND2 I534 (conwgif_0[44:44], wg_0r0[44:44], conwig_0);
  AND2 I535 (conwgif_0[45:45], wg_0r0[45:45], conwig_0);
  AND2 I536 (conwgif_0[46:46], wg_0r0[46:46], conwig_0);
  AND2 I537 (conwgif_0[47:47], wg_0r0[47:47], conwig_0);
  AND2 I538 (conwgif_0[48:48], wg_0r0[48:48], conwig_0);
  AND2 I539 (conwgif_0[49:49], wg_0r0[49:49], conwig_0);
  AND2 I540 (conwgif_0[50:50], wg_0r0[50:50], conwig_0);
  AND2 I541 (conwgif_0[51:51], wg_0r0[51:51], conwig_0);
  AND2 I542 (conwgif_0[52:52], wg_0r0[52:52], conwig_0);
  AND2 I543 (conwgif_0[53:53], wg_0r0[53:53], conwig_0);
  AND2 I544 (conwgif_0[54:54], wg_0r0[54:54], conwig_0);
  AND2 I545 (conwgif_0[55:55], wg_0r0[55:55], conwig_0);
  AND2 I546 (conwgif_0[56:56], wg_0r0[56:56], conwig_0);
  AND2 I547 (conwgif_0[57:57], wg_0r0[57:57], conwig_0);
  AND2 I548 (conwgif_0[58:58], wg_0r0[58:58], conwig_0);
  AND2 I549 (conwgif_0[59:59], wg_0r0[59:59], conwig_0);
  AND2 I550 (conwgif_0[60:60], wg_0r0[60:60], conwig_0);
  AND2 I551 (conwgif_0[61:61], wg_0r0[61:61], conwig_0);
  AND2 I552 (conwgif_0[62:62], wg_0r0[62:62], conwig_0);
  AND2 I553 (conwgif_0[63:63], wg_0r0[63:63], conwig_0);
  AND2 I554 (conwgif_0[64:64], wg_0r0[64:64], conwig_0);
  AND2 I555 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I556 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I557 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I558 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I559 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I560 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I561 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I562 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I563 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I564 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I565 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I566 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I567 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I568 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I569 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I570 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I571 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I572 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I573 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I574 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I575 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I576 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I577 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I578 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I579 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I580 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I581 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I582 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I583 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I584 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I585 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I586 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  AND2 I587 (conwgit_0[32:32], wg_0r1[32:32], conwig_0);
  AND2 I588 (conwgit_0[33:33], wg_0r1[33:33], conwig_0);
  AND2 I589 (conwgit_0[34:34], wg_0r1[34:34], conwig_0);
  AND2 I590 (conwgit_0[35:35], wg_0r1[35:35], conwig_0);
  AND2 I591 (conwgit_0[36:36], wg_0r1[36:36], conwig_0);
  AND2 I592 (conwgit_0[37:37], wg_0r1[37:37], conwig_0);
  AND2 I593 (conwgit_0[38:38], wg_0r1[38:38], conwig_0);
  AND2 I594 (conwgit_0[39:39], wg_0r1[39:39], conwig_0);
  AND2 I595 (conwgit_0[40:40], wg_0r1[40:40], conwig_0);
  AND2 I596 (conwgit_0[41:41], wg_0r1[41:41], conwig_0);
  AND2 I597 (conwgit_0[42:42], wg_0r1[42:42], conwig_0);
  AND2 I598 (conwgit_0[43:43], wg_0r1[43:43], conwig_0);
  AND2 I599 (conwgit_0[44:44], wg_0r1[44:44], conwig_0);
  AND2 I600 (conwgit_0[45:45], wg_0r1[45:45], conwig_0);
  AND2 I601 (conwgit_0[46:46], wg_0r1[46:46], conwig_0);
  AND2 I602 (conwgit_0[47:47], wg_0r1[47:47], conwig_0);
  AND2 I603 (conwgit_0[48:48], wg_0r1[48:48], conwig_0);
  AND2 I604 (conwgit_0[49:49], wg_0r1[49:49], conwig_0);
  AND2 I605 (conwgit_0[50:50], wg_0r1[50:50], conwig_0);
  AND2 I606 (conwgit_0[51:51], wg_0r1[51:51], conwig_0);
  AND2 I607 (conwgit_0[52:52], wg_0r1[52:52], conwig_0);
  AND2 I608 (conwgit_0[53:53], wg_0r1[53:53], conwig_0);
  AND2 I609 (conwgit_0[54:54], wg_0r1[54:54], conwig_0);
  AND2 I610 (conwgit_0[55:55], wg_0r1[55:55], conwig_0);
  AND2 I611 (conwgit_0[56:56], wg_0r1[56:56], conwig_0);
  AND2 I612 (conwgit_0[57:57], wg_0r1[57:57], conwig_0);
  AND2 I613 (conwgit_0[58:58], wg_0r1[58:58], conwig_0);
  AND2 I614 (conwgit_0[59:59], wg_0r1[59:59], conwig_0);
  AND2 I615 (conwgit_0[60:60], wg_0r1[60:60], conwig_0);
  AND2 I616 (conwgit_0[61:61], wg_0r1[61:61], conwig_0);
  AND2 I617 (conwgit_0[62:62], wg_0r1[62:62], conwig_0);
  AND2 I618 (conwgit_0[63:63], wg_0r1[63:63], conwig_0);
  AND2 I619 (conwgit_0[64:64], wg_0r1[64:64], conwig_0);
  BUFF I620 (conwigc_0, wc_0);
  AO22 I621 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I622 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I623 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I624 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I625 (wenr_0[0:0], wc_0);
  BUFF I626 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I627 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I628 (wenr_0[1:1], wc_0);
  BUFF I629 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I630 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I631 (wenr_0[2:2], wc_0);
  BUFF I632 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I633 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I634 (wenr_0[3:3], wc_0);
  BUFF I635 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I636 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I637 (wenr_0[4:4], wc_0);
  BUFF I638 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I639 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I640 (wenr_0[5:5], wc_0);
  BUFF I641 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I642 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I643 (wenr_0[6:6], wc_0);
  BUFF I644 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I645 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I646 (wenr_0[7:7], wc_0);
  BUFF I647 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I648 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I649 (wenr_0[8:8], wc_0);
  BUFF I650 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I651 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I652 (wenr_0[9:9], wc_0);
  BUFF I653 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I654 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I655 (wenr_0[10:10], wc_0);
  BUFF I656 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I657 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I658 (wenr_0[11:11], wc_0);
  BUFF I659 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I660 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I661 (wenr_0[12:12], wc_0);
  BUFF I662 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I663 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I664 (wenr_0[13:13], wc_0);
  BUFF I665 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I666 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I667 (wenr_0[14:14], wc_0);
  BUFF I668 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I669 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I670 (wenr_0[15:15], wc_0);
  BUFF I671 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I672 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I673 (wenr_0[16:16], wc_0);
  BUFF I674 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I675 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I676 (wenr_0[17:17], wc_0);
  BUFF I677 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I678 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I679 (wenr_0[18:18], wc_0);
  BUFF I680 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I681 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I682 (wenr_0[19:19], wc_0);
  BUFF I683 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I684 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I685 (wenr_0[20:20], wc_0);
  BUFF I686 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I687 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I688 (wenr_0[21:21], wc_0);
  BUFF I689 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I690 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I691 (wenr_0[22:22], wc_0);
  BUFF I692 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I693 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I694 (wenr_0[23:23], wc_0);
  BUFF I695 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I696 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I697 (wenr_0[24:24], wc_0);
  BUFF I698 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I699 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I700 (wenr_0[25:25], wc_0);
  BUFF I701 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I702 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I703 (wenr_0[26:26], wc_0);
  BUFF I704 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I705 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I706 (wenr_0[27:27], wc_0);
  BUFF I707 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I708 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I709 (wenr_0[28:28], wc_0);
  BUFF I710 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I711 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I712 (wenr_0[29:29], wc_0);
  BUFF I713 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I714 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I715 (wenr_0[30:30], wc_0);
  BUFF I716 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I717 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I718 (wenr_0[31:31], wc_0);
  BUFF I719 (wf_0[32:32], conwgif_0[32:32]);
  BUFF I720 (wt_0[32:32], conwgit_0[32:32]);
  BUFF I721 (wenr_0[32:32], wc_0);
  BUFF I722 (wf_0[33:33], conwgif_0[33:33]);
  BUFF I723 (wt_0[33:33], conwgit_0[33:33]);
  BUFF I724 (wenr_0[33:33], wc_0);
  BUFF I725 (wf_0[34:34], conwgif_0[34:34]);
  BUFF I726 (wt_0[34:34], conwgit_0[34:34]);
  BUFF I727 (wenr_0[34:34], wc_0);
  BUFF I728 (wf_0[35:35], conwgif_0[35:35]);
  BUFF I729 (wt_0[35:35], conwgit_0[35:35]);
  BUFF I730 (wenr_0[35:35], wc_0);
  BUFF I731 (wf_0[36:36], conwgif_0[36:36]);
  BUFF I732 (wt_0[36:36], conwgit_0[36:36]);
  BUFF I733 (wenr_0[36:36], wc_0);
  BUFF I734 (wf_0[37:37], conwgif_0[37:37]);
  BUFF I735 (wt_0[37:37], conwgit_0[37:37]);
  BUFF I736 (wenr_0[37:37], wc_0);
  BUFF I737 (wf_0[38:38], conwgif_0[38:38]);
  BUFF I738 (wt_0[38:38], conwgit_0[38:38]);
  BUFF I739 (wenr_0[38:38], wc_0);
  BUFF I740 (wf_0[39:39], conwgif_0[39:39]);
  BUFF I741 (wt_0[39:39], conwgit_0[39:39]);
  BUFF I742 (wenr_0[39:39], wc_0);
  BUFF I743 (wf_0[40:40], conwgif_0[40:40]);
  BUFF I744 (wt_0[40:40], conwgit_0[40:40]);
  BUFF I745 (wenr_0[40:40], wc_0);
  BUFF I746 (wf_0[41:41], conwgif_0[41:41]);
  BUFF I747 (wt_0[41:41], conwgit_0[41:41]);
  BUFF I748 (wenr_0[41:41], wc_0);
  BUFF I749 (wf_0[42:42], conwgif_0[42:42]);
  BUFF I750 (wt_0[42:42], conwgit_0[42:42]);
  BUFF I751 (wenr_0[42:42], wc_0);
  BUFF I752 (wf_0[43:43], conwgif_0[43:43]);
  BUFF I753 (wt_0[43:43], conwgit_0[43:43]);
  BUFF I754 (wenr_0[43:43], wc_0);
  BUFF I755 (wf_0[44:44], conwgif_0[44:44]);
  BUFF I756 (wt_0[44:44], conwgit_0[44:44]);
  BUFF I757 (wenr_0[44:44], wc_0);
  BUFF I758 (wf_0[45:45], conwgif_0[45:45]);
  BUFF I759 (wt_0[45:45], conwgit_0[45:45]);
  BUFF I760 (wenr_0[45:45], wc_0);
  BUFF I761 (wf_0[46:46], conwgif_0[46:46]);
  BUFF I762 (wt_0[46:46], conwgit_0[46:46]);
  BUFF I763 (wenr_0[46:46], wc_0);
  BUFF I764 (wf_0[47:47], conwgif_0[47:47]);
  BUFF I765 (wt_0[47:47], conwgit_0[47:47]);
  BUFF I766 (wenr_0[47:47], wc_0);
  BUFF I767 (wf_0[48:48], conwgif_0[48:48]);
  BUFF I768 (wt_0[48:48], conwgit_0[48:48]);
  BUFF I769 (wenr_0[48:48], wc_0);
  BUFF I770 (wf_0[49:49], conwgif_0[49:49]);
  BUFF I771 (wt_0[49:49], conwgit_0[49:49]);
  BUFF I772 (wenr_0[49:49], wc_0);
  BUFF I773 (wf_0[50:50], conwgif_0[50:50]);
  BUFF I774 (wt_0[50:50], conwgit_0[50:50]);
  BUFF I775 (wenr_0[50:50], wc_0);
  BUFF I776 (wf_0[51:51], conwgif_0[51:51]);
  BUFF I777 (wt_0[51:51], conwgit_0[51:51]);
  BUFF I778 (wenr_0[51:51], wc_0);
  BUFF I779 (wf_0[52:52], conwgif_0[52:52]);
  BUFF I780 (wt_0[52:52], conwgit_0[52:52]);
  BUFF I781 (wenr_0[52:52], wc_0);
  BUFF I782 (wf_0[53:53], conwgif_0[53:53]);
  BUFF I783 (wt_0[53:53], conwgit_0[53:53]);
  BUFF I784 (wenr_0[53:53], wc_0);
  BUFF I785 (wf_0[54:54], conwgif_0[54:54]);
  BUFF I786 (wt_0[54:54], conwgit_0[54:54]);
  BUFF I787 (wenr_0[54:54], wc_0);
  BUFF I788 (wf_0[55:55], conwgif_0[55:55]);
  BUFF I789 (wt_0[55:55], conwgit_0[55:55]);
  BUFF I790 (wenr_0[55:55], wc_0);
  BUFF I791 (wf_0[56:56], conwgif_0[56:56]);
  BUFF I792 (wt_0[56:56], conwgit_0[56:56]);
  BUFF I793 (wenr_0[56:56], wc_0);
  BUFF I794 (wf_0[57:57], conwgif_0[57:57]);
  BUFF I795 (wt_0[57:57], conwgit_0[57:57]);
  BUFF I796 (wenr_0[57:57], wc_0);
  BUFF I797 (wf_0[58:58], conwgif_0[58:58]);
  BUFF I798 (wt_0[58:58], conwgit_0[58:58]);
  BUFF I799 (wenr_0[58:58], wc_0);
  BUFF I800 (wf_0[59:59], conwgif_0[59:59]);
  BUFF I801 (wt_0[59:59], conwgit_0[59:59]);
  BUFF I802 (wenr_0[59:59], wc_0);
  BUFF I803 (wf_0[60:60], conwgif_0[60:60]);
  BUFF I804 (wt_0[60:60], conwgit_0[60:60]);
  BUFF I805 (wenr_0[60:60], wc_0);
  BUFF I806 (wf_0[61:61], conwgif_0[61:61]);
  BUFF I807 (wt_0[61:61], conwgit_0[61:61]);
  BUFF I808 (wenr_0[61:61], wc_0);
  BUFF I809 (wf_0[62:62], conwgif_0[62:62]);
  BUFF I810 (wt_0[62:62], conwgit_0[62:62]);
  BUFF I811 (wenr_0[62:62], wc_0);
  BUFF I812 (wf_0[63:63], conwgif_0[63:63]);
  BUFF I813 (wt_0[63:63], conwgit_0[63:63]);
  BUFF I814 (wenr_0[63:63], wc_0);
  BUFF I815 (wf_0[64:64], conwgif_0[64:64]);
  BUFF I816 (wt_0[64:64], conwgit_0[64:64]);
  BUFF I817 (wenr_0[64:64], wc_0);
  C3 I818 (simp8031_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I819 (simp8031_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I820 (simp8031_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I821 (simp8031_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I822 (simp8031_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I823 (simp8031_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I824 (simp8031_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I825 (simp8031_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I826 (simp8031_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I827 (simp8031_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I828 (simp8031_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I829 (simp8031_0[11:11], wacks_0[32:32], wacks_0[33:33], wacks_0[34:34]);
  C3 I830 (simp8031_0[12:12], wacks_0[35:35], wacks_0[36:36], wacks_0[37:37]);
  C3 I831 (simp8031_0[13:13], wacks_0[38:38], wacks_0[39:39], wacks_0[40:40]);
  C3 I832 (simp8031_0[14:14], wacks_0[41:41], wacks_0[42:42], wacks_0[43:43]);
  C3 I833 (simp8031_0[15:15], wacks_0[44:44], wacks_0[45:45], wacks_0[46:46]);
  C3 I834 (simp8031_0[16:16], wacks_0[47:47], wacks_0[48:48], wacks_0[49:49]);
  C3 I835 (simp8031_0[17:17], wacks_0[50:50], wacks_0[51:51], wacks_0[52:52]);
  C3 I836 (simp8031_0[18:18], wacks_0[53:53], wacks_0[54:54], wacks_0[55:55]);
  C3 I837 (simp8031_0[19:19], wacks_0[56:56], wacks_0[57:57], wacks_0[58:58]);
  C3 I838 (simp8031_0[20:20], wacks_0[59:59], wacks_0[60:60], wacks_0[61:61]);
  C3 I839 (simp8031_0[21:21], wacks_0[62:62], wacks_0[63:63], wacks_0[64:64]);
  C3 I840 (simp8032_0[0:0], simp8031_0[0:0], simp8031_0[1:1], simp8031_0[2:2]);
  C3 I841 (simp8032_0[1:1], simp8031_0[3:3], simp8031_0[4:4], simp8031_0[5:5]);
  C3 I842 (simp8032_0[2:2], simp8031_0[6:6], simp8031_0[7:7], simp8031_0[8:8]);
  C3 I843 (simp8032_0[3:3], simp8031_0[9:9], simp8031_0[10:10], simp8031_0[11:11]);
  C3 I844 (simp8032_0[4:4], simp8031_0[12:12], simp8031_0[13:13], simp8031_0[14:14]);
  C3 I845 (simp8032_0[5:5], simp8031_0[15:15], simp8031_0[16:16], simp8031_0[17:17]);
  C3 I846 (simp8032_0[6:6], simp8031_0[18:18], simp8031_0[19:19], simp8031_0[20:20]);
  BUFF I847 (simp8032_0[7:7], simp8031_0[21:21]);
  C3 I848 (simp8033_0[0:0], simp8032_0[0:0], simp8032_0[1:1], simp8032_0[2:2]);
  C3 I849 (simp8033_0[1:1], simp8032_0[3:3], simp8032_0[4:4], simp8032_0[5:5]);
  C2 I850 (simp8033_0[2:2], simp8032_0[6:6], simp8032_0[7:7]);
  C3 I851 (wd_0r, simp8033_0[0:0], simp8033_0[1:1], simp8033_0[2:2]);
  AND2 I852 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I853 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I854 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I855 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I856 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I857 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I858 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I859 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I860 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I861 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I862 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I863 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I864 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I865 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I866 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I867 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I868 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I869 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I870 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I871 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I872 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I873 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I874 (rd_1r0[0:0], df_0[25:25], rg_1r);
  AND2 I875 (rd_1r0[1:1], df_0[26:26], rg_1r);
  AND2 I876 (rd_1r0[2:2], df_0[27:27], rg_1r);
  AND2 I877 (rd_1r0[3:3], df_0[28:28], rg_1r);
  AND2 I878 (rd_1r0[4:4], df_0[29:29], rg_1r);
  AND2 I879 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I880 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I881 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I882 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I883 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I884 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I885 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I886 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I887 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I888 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I889 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I890 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I891 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I892 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I893 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I894 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I895 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I896 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I897 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I898 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I899 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I900 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I901 (rd_3r0[0:0], df_0[25:25], rg_3r);
  AND2 I902 (rd_3r0[1:1], df_0[26:26], rg_3r);
  AND2 I903 (rd_3r0[2:2], df_0[27:27], rg_3r);
  AND2 I904 (rd_3r0[3:3], df_0[28:28], rg_3r);
  AND2 I905 (rd_4r0[0:0], df_0[22:22], rg_4r);
  AND2 I906 (rd_4r0[1:1], df_0[23:23], rg_4r);
  AND2 I907 (rd_4r0[2:2], df_0[24:24], rg_4r);
  AND2 I908 (rd_5r0[0:0], df_0[19:19], rg_5r);
  AND2 I909 (rd_5r0[1:1], df_0[20:20], rg_5r);
  AND2 I910 (rd_5r0[2:2], df_0[21:21], rg_5r);
  AND2 I911 (rd_5r0[3:3], df_0[22:22], rg_5r);
  AND2 I912 (rd_5r0[4:4], df_0[23:23], rg_5r);
  AND2 I913 (rd_5r0[5:5], df_0[24:24], rg_5r);
  AND2 I914 (rd_6r0, df_0[13:13], rg_6r);
  AND2 I915 (rd_7r0[0:0], df_0[0:0], rg_7r);
  AND2 I916 (rd_7r0[1:1], df_0[1:1], rg_7r);
  AND2 I917 (rd_7r0[2:2], df_0[2:2], rg_7r);
  AND2 I918 (rd_7r0[3:3], df_0[3:3], rg_7r);
  AND2 I919 (rd_7r0[4:4], df_0[4:4], rg_7r);
  AND2 I920 (rd_7r0[5:5], df_0[5:5], rg_7r);
  AND2 I921 (rd_7r0[6:6], df_0[6:6], rg_7r);
  AND2 I922 (rd_7r0[7:7], df_0[7:7], rg_7r);
  AND2 I923 (rd_7r0[8:8], df_0[8:8], rg_7r);
  AND2 I924 (rd_7r0[9:9], df_0[9:9], rg_7r);
  AND2 I925 (rd_7r0[10:10], df_0[10:10], rg_7r);
  AND2 I926 (rd_7r0[11:11], df_0[11:11], rg_7r);
  AND2 I927 (rd_7r0[12:12], df_0[12:12], rg_7r);
  AND2 I928 (rd_8r0[0:0], df_0[19:19], rg_8r);
  AND2 I929 (rd_8r0[1:1], df_0[20:20], rg_8r);
  AND2 I930 (rd_8r0[2:2], df_0[21:21], rg_8r);
  AND2 I931 (rd_8r0[3:3], df_0[22:22], rg_8r);
  AND2 I932 (rd_8r0[4:4], df_0[23:23], rg_8r);
  AND2 I933 (rd_8r0[5:5], df_0[24:24], rg_8r);
  AND2 I934 (rd_9r0[0:0], df_0[25:25], rg_9r);
  AND2 I935 (rd_9r0[1:1], df_0[26:26], rg_9r);
  AND2 I936 (rd_9r0[2:2], df_0[27:27], rg_9r);
  AND2 I937 (rd_9r0[3:3], df_0[28:28], rg_9r);
  AND2 I938 (rd_9r0[4:4], df_0[29:29], rg_9r);
  AND2 I939 (rd_10r0[0:0], df_0[25:25], rg_10r);
  AND2 I940 (rd_10r0[1:1], df_0[26:26], rg_10r);
  AND2 I941 (rd_10r0[2:2], df_0[27:27], rg_10r);
  AND2 I942 (rd_10r0[3:3], df_0[28:28], rg_10r);
  AND2 I943 (rd_10r0[4:4], df_0[29:29], rg_10r);
  AND2 I944 (rd_11r0[0:0], df_0[0:0], rg_11r);
  AND2 I945 (rd_11r0[1:1], df_0[1:1], rg_11r);
  AND2 I946 (rd_11r0[2:2], df_0[2:2], rg_11r);
  AND2 I947 (rd_11r0[3:3], df_0[3:3], rg_11r);
  AND2 I948 (rd_11r0[4:4], df_0[4:4], rg_11r);
  AND2 I949 (rd_12r0[0:0], df_0[14:14], rg_12r);
  AND2 I950 (rd_12r0[1:1], df_0[15:15], rg_12r);
  AND2 I951 (rd_12r0[2:2], df_0[16:16], rg_12r);
  AND2 I952 (rd_12r0[3:3], df_0[17:17], rg_12r);
  AND2 I953 (rd_12r0[4:4], df_0[18:18], rg_12r);
  AND2 I954 (rd_13r0, df_0[13:13], rg_13r);
  AND2 I955 (rd_14r0, df_0[13:13], rg_14r);
  AND2 I956 (rd_15r0[0:0], df_0[0:0], rg_15r);
  AND2 I957 (rd_15r0[1:1], df_0[1:1], rg_15r);
  AND2 I958 (rd_15r0[2:2], df_0[2:2], rg_15r);
  AND2 I959 (rd_15r0[3:3], df_0[3:3], rg_15r);
  AND2 I960 (rd_15r0[4:4], df_0[4:4], rg_15r);
  AND2 I961 (rd_15r0[5:5], df_0[5:5], rg_15r);
  AND2 I962 (rd_15r0[6:6], df_0[6:6], rg_15r);
  AND2 I963 (rd_15r0[7:7], df_0[7:7], rg_15r);
  AND2 I964 (rd_15r0[8:8], df_0[8:8], rg_15r);
  AND2 I965 (rd_15r0[9:9], df_0[9:9], rg_15r);
  AND2 I966 (rd_15r0[10:10], df_0[10:10], rg_15r);
  AND2 I967 (rd_15r0[11:11], df_0[11:11], rg_15r);
  AND2 I968 (rd_15r0[12:12], df_0[12:12], rg_15r);
  AND2 I969 (rd_16r0[0:0], df_0[19:19], rg_16r);
  AND2 I970 (rd_16r0[1:1], df_0[20:20], rg_16r);
  AND2 I971 (rd_16r0[2:2], df_0[21:21], rg_16r);
  AND2 I972 (rd_16r0[3:3], df_0[22:22], rg_16r);
  AND2 I973 (rd_16r0[4:4], df_0[23:23], rg_16r);
  AND2 I974 (rd_16r0[5:5], df_0[24:24], rg_16r);
  AND2 I975 (rd_17r0[0:0], df_0[25:25], rg_17r);
  AND2 I976 (rd_17r0[1:1], df_0[26:26], rg_17r);
  AND2 I977 (rd_17r0[2:2], df_0[27:27], rg_17r);
  AND2 I978 (rd_17r0[3:3], df_0[28:28], rg_17r);
  AND2 I979 (rd_17r0[4:4], df_0[29:29], rg_17r);
  AND2 I980 (rd_18r0[0:0], df_0[0:0], rg_18r);
  AND2 I981 (rd_18r0[1:1], df_0[1:1], rg_18r);
  AND2 I982 (rd_18r0[2:2], df_0[2:2], rg_18r);
  AND2 I983 (rd_18r0[3:3], df_0[3:3], rg_18r);
  AND2 I984 (rd_18r0[4:4], df_0[4:4], rg_18r);
  AND2 I985 (rd_19r0[0:0], df_0[14:14], rg_19r);
  AND2 I986 (rd_19r0[1:1], df_0[15:15], rg_19r);
  AND2 I987 (rd_19r0[2:2], df_0[16:16], rg_19r);
  AND2 I988 (rd_19r0[3:3], df_0[17:17], rg_19r);
  AND2 I989 (rd_19r0[4:4], df_0[18:18], rg_19r);
  AND2 I990 (rd_20r0, df_0[13:13], rg_20r);
  AND2 I991 (rd_21r0[0:0], df_0[19:19], rg_21r);
  AND2 I992 (rd_21r0[1:1], df_0[20:20], rg_21r);
  AND2 I993 (rd_21r0[2:2], df_0[21:21], rg_21r);
  AND2 I994 (rd_21r0[3:3], df_0[22:22], rg_21r);
  AND2 I995 (rd_21r0[4:4], df_0[23:23], rg_21r);
  AND2 I996 (rd_21r0[5:5], df_0[24:24], rg_21r);
  AND2 I997 (rd_22r0[0:0], df_0[30:30], rg_22r);
  AND2 I998 (rd_22r0[1:1], df_0[31:31], rg_22r);
  AND2 I999 (rd_23r0[0:0], df_0[32:32], rg_23r);
  AND2 I1000 (rd_23r0[1:1], df_0[33:33], rg_23r);
  AND2 I1001 (rd_23r0[2:2], df_0[34:34], rg_23r);
  AND2 I1002 (rd_23r0[3:3], df_0[35:35], rg_23r);
  AND2 I1003 (rd_23r0[4:4], df_0[36:36], rg_23r);
  AND2 I1004 (rd_23r0[5:5], df_0[37:37], rg_23r);
  AND2 I1005 (rd_23r0[6:6], df_0[38:38], rg_23r);
  AND2 I1006 (rd_23r0[7:7], df_0[39:39], rg_23r);
  AND2 I1007 (rd_23r0[8:8], df_0[40:40], rg_23r);
  AND2 I1008 (rd_23r0[9:9], df_0[41:41], rg_23r);
  AND2 I1009 (rd_23r0[10:10], df_0[42:42], rg_23r);
  AND2 I1010 (rd_23r0[11:11], df_0[43:43], rg_23r);
  AND2 I1011 (rd_23r0[12:12], df_0[44:44], rg_23r);
  AND2 I1012 (rd_23r0[13:13], df_0[45:45], rg_23r);
  AND2 I1013 (rd_23r0[14:14], df_0[46:46], rg_23r);
  AND2 I1014 (rd_23r0[15:15], df_0[47:47], rg_23r);
  AND2 I1015 (rd_23r0[16:16], df_0[48:48], rg_23r);
  AND2 I1016 (rd_23r0[17:17], df_0[49:49], rg_23r);
  AND2 I1017 (rd_23r0[18:18], df_0[50:50], rg_23r);
  AND2 I1018 (rd_23r0[19:19], df_0[51:51], rg_23r);
  AND2 I1019 (rd_23r0[20:20], df_0[52:52], rg_23r);
  AND2 I1020 (rd_23r0[21:21], df_0[53:53], rg_23r);
  AND2 I1021 (rd_23r0[22:22], df_0[54:54], rg_23r);
  AND2 I1022 (rd_23r0[23:23], df_0[55:55], rg_23r);
  AND2 I1023 (rd_23r0[24:24], df_0[56:56], rg_23r);
  AND2 I1024 (rd_23r0[25:25], df_0[57:57], rg_23r);
  AND2 I1025 (rd_23r0[26:26], df_0[58:58], rg_23r);
  AND2 I1026 (rd_23r0[27:27], df_0[59:59], rg_23r);
  AND2 I1027 (rd_23r0[28:28], df_0[60:60], rg_23r);
  AND2 I1028 (rd_23r0[29:29], df_0[61:61], rg_23r);
  AND2 I1029 (rd_23r0[30:30], df_0[62:62], rg_23r);
  AND2 I1030 (rd_23r0[31:31], df_0[63:63], rg_23r);
  AND2 I1031 (rd_23r0[32:32], df_0[64:64], rg_23r);
  AND2 I1032 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I1033 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I1034 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I1035 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I1036 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I1037 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I1038 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I1039 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I1040 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I1041 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I1042 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I1043 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I1044 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I1045 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I1046 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I1047 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I1048 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I1049 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I1050 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I1051 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I1052 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I1053 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I1054 (rd_1r1[0:0], dt_0[25:25], rg_1r);
  AND2 I1055 (rd_1r1[1:1], dt_0[26:26], rg_1r);
  AND2 I1056 (rd_1r1[2:2], dt_0[27:27], rg_1r);
  AND2 I1057 (rd_1r1[3:3], dt_0[28:28], rg_1r);
  AND2 I1058 (rd_1r1[4:4], dt_0[29:29], rg_1r);
  AND2 I1059 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I1060 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I1061 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I1062 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I1063 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I1064 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I1065 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I1066 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I1067 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I1068 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I1069 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I1070 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I1071 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I1072 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I1073 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I1074 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I1075 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I1076 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I1077 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I1078 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I1079 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I1080 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I1081 (rd_3r1[0:0], dt_0[25:25], rg_3r);
  AND2 I1082 (rd_3r1[1:1], dt_0[26:26], rg_3r);
  AND2 I1083 (rd_3r1[2:2], dt_0[27:27], rg_3r);
  AND2 I1084 (rd_3r1[3:3], dt_0[28:28], rg_3r);
  AND2 I1085 (rd_4r1[0:0], dt_0[22:22], rg_4r);
  AND2 I1086 (rd_4r1[1:1], dt_0[23:23], rg_4r);
  AND2 I1087 (rd_4r1[2:2], dt_0[24:24], rg_4r);
  AND2 I1088 (rd_5r1[0:0], dt_0[19:19], rg_5r);
  AND2 I1089 (rd_5r1[1:1], dt_0[20:20], rg_5r);
  AND2 I1090 (rd_5r1[2:2], dt_0[21:21], rg_5r);
  AND2 I1091 (rd_5r1[3:3], dt_0[22:22], rg_5r);
  AND2 I1092 (rd_5r1[4:4], dt_0[23:23], rg_5r);
  AND2 I1093 (rd_5r1[5:5], dt_0[24:24], rg_5r);
  AND2 I1094 (rd_6r1, dt_0[13:13], rg_6r);
  AND2 I1095 (rd_7r1[0:0], dt_0[0:0], rg_7r);
  AND2 I1096 (rd_7r1[1:1], dt_0[1:1], rg_7r);
  AND2 I1097 (rd_7r1[2:2], dt_0[2:2], rg_7r);
  AND2 I1098 (rd_7r1[3:3], dt_0[3:3], rg_7r);
  AND2 I1099 (rd_7r1[4:4], dt_0[4:4], rg_7r);
  AND2 I1100 (rd_7r1[5:5], dt_0[5:5], rg_7r);
  AND2 I1101 (rd_7r1[6:6], dt_0[6:6], rg_7r);
  AND2 I1102 (rd_7r1[7:7], dt_0[7:7], rg_7r);
  AND2 I1103 (rd_7r1[8:8], dt_0[8:8], rg_7r);
  AND2 I1104 (rd_7r1[9:9], dt_0[9:9], rg_7r);
  AND2 I1105 (rd_7r1[10:10], dt_0[10:10], rg_7r);
  AND2 I1106 (rd_7r1[11:11], dt_0[11:11], rg_7r);
  AND2 I1107 (rd_7r1[12:12], dt_0[12:12], rg_7r);
  AND2 I1108 (rd_8r1[0:0], dt_0[19:19], rg_8r);
  AND2 I1109 (rd_8r1[1:1], dt_0[20:20], rg_8r);
  AND2 I1110 (rd_8r1[2:2], dt_0[21:21], rg_8r);
  AND2 I1111 (rd_8r1[3:3], dt_0[22:22], rg_8r);
  AND2 I1112 (rd_8r1[4:4], dt_0[23:23], rg_8r);
  AND2 I1113 (rd_8r1[5:5], dt_0[24:24], rg_8r);
  AND2 I1114 (rd_9r1[0:0], dt_0[25:25], rg_9r);
  AND2 I1115 (rd_9r1[1:1], dt_0[26:26], rg_9r);
  AND2 I1116 (rd_9r1[2:2], dt_0[27:27], rg_9r);
  AND2 I1117 (rd_9r1[3:3], dt_0[28:28], rg_9r);
  AND2 I1118 (rd_9r1[4:4], dt_0[29:29], rg_9r);
  AND2 I1119 (rd_10r1[0:0], dt_0[25:25], rg_10r);
  AND2 I1120 (rd_10r1[1:1], dt_0[26:26], rg_10r);
  AND2 I1121 (rd_10r1[2:2], dt_0[27:27], rg_10r);
  AND2 I1122 (rd_10r1[3:3], dt_0[28:28], rg_10r);
  AND2 I1123 (rd_10r1[4:4], dt_0[29:29], rg_10r);
  AND2 I1124 (rd_11r1[0:0], dt_0[0:0], rg_11r);
  AND2 I1125 (rd_11r1[1:1], dt_0[1:1], rg_11r);
  AND2 I1126 (rd_11r1[2:2], dt_0[2:2], rg_11r);
  AND2 I1127 (rd_11r1[3:3], dt_0[3:3], rg_11r);
  AND2 I1128 (rd_11r1[4:4], dt_0[4:4], rg_11r);
  AND2 I1129 (rd_12r1[0:0], dt_0[14:14], rg_12r);
  AND2 I1130 (rd_12r1[1:1], dt_0[15:15], rg_12r);
  AND2 I1131 (rd_12r1[2:2], dt_0[16:16], rg_12r);
  AND2 I1132 (rd_12r1[3:3], dt_0[17:17], rg_12r);
  AND2 I1133 (rd_12r1[4:4], dt_0[18:18], rg_12r);
  AND2 I1134 (rd_13r1, dt_0[13:13], rg_13r);
  AND2 I1135 (rd_14r1, dt_0[13:13], rg_14r);
  AND2 I1136 (rd_15r1[0:0], dt_0[0:0], rg_15r);
  AND2 I1137 (rd_15r1[1:1], dt_0[1:1], rg_15r);
  AND2 I1138 (rd_15r1[2:2], dt_0[2:2], rg_15r);
  AND2 I1139 (rd_15r1[3:3], dt_0[3:3], rg_15r);
  AND2 I1140 (rd_15r1[4:4], dt_0[4:4], rg_15r);
  AND2 I1141 (rd_15r1[5:5], dt_0[5:5], rg_15r);
  AND2 I1142 (rd_15r1[6:6], dt_0[6:6], rg_15r);
  AND2 I1143 (rd_15r1[7:7], dt_0[7:7], rg_15r);
  AND2 I1144 (rd_15r1[8:8], dt_0[8:8], rg_15r);
  AND2 I1145 (rd_15r1[9:9], dt_0[9:9], rg_15r);
  AND2 I1146 (rd_15r1[10:10], dt_0[10:10], rg_15r);
  AND2 I1147 (rd_15r1[11:11], dt_0[11:11], rg_15r);
  AND2 I1148 (rd_15r1[12:12], dt_0[12:12], rg_15r);
  AND2 I1149 (rd_16r1[0:0], dt_0[19:19], rg_16r);
  AND2 I1150 (rd_16r1[1:1], dt_0[20:20], rg_16r);
  AND2 I1151 (rd_16r1[2:2], dt_0[21:21], rg_16r);
  AND2 I1152 (rd_16r1[3:3], dt_0[22:22], rg_16r);
  AND2 I1153 (rd_16r1[4:4], dt_0[23:23], rg_16r);
  AND2 I1154 (rd_16r1[5:5], dt_0[24:24], rg_16r);
  AND2 I1155 (rd_17r1[0:0], dt_0[25:25], rg_17r);
  AND2 I1156 (rd_17r1[1:1], dt_0[26:26], rg_17r);
  AND2 I1157 (rd_17r1[2:2], dt_0[27:27], rg_17r);
  AND2 I1158 (rd_17r1[3:3], dt_0[28:28], rg_17r);
  AND2 I1159 (rd_17r1[4:4], dt_0[29:29], rg_17r);
  AND2 I1160 (rd_18r1[0:0], dt_0[0:0], rg_18r);
  AND2 I1161 (rd_18r1[1:1], dt_0[1:1], rg_18r);
  AND2 I1162 (rd_18r1[2:2], dt_0[2:2], rg_18r);
  AND2 I1163 (rd_18r1[3:3], dt_0[3:3], rg_18r);
  AND2 I1164 (rd_18r1[4:4], dt_0[4:4], rg_18r);
  AND2 I1165 (rd_19r1[0:0], dt_0[14:14], rg_19r);
  AND2 I1166 (rd_19r1[1:1], dt_0[15:15], rg_19r);
  AND2 I1167 (rd_19r1[2:2], dt_0[16:16], rg_19r);
  AND2 I1168 (rd_19r1[3:3], dt_0[17:17], rg_19r);
  AND2 I1169 (rd_19r1[4:4], dt_0[18:18], rg_19r);
  AND2 I1170 (rd_20r1, dt_0[13:13], rg_20r);
  AND2 I1171 (rd_21r1[0:0], dt_0[19:19], rg_21r);
  AND2 I1172 (rd_21r1[1:1], dt_0[20:20], rg_21r);
  AND2 I1173 (rd_21r1[2:2], dt_0[21:21], rg_21r);
  AND2 I1174 (rd_21r1[3:3], dt_0[22:22], rg_21r);
  AND2 I1175 (rd_21r1[4:4], dt_0[23:23], rg_21r);
  AND2 I1176 (rd_21r1[5:5], dt_0[24:24], rg_21r);
  AND2 I1177 (rd_22r1[0:0], dt_0[30:30], rg_22r);
  AND2 I1178 (rd_22r1[1:1], dt_0[31:31], rg_22r);
  AND2 I1179 (rd_23r1[0:0], dt_0[32:32], rg_23r);
  AND2 I1180 (rd_23r1[1:1], dt_0[33:33], rg_23r);
  AND2 I1181 (rd_23r1[2:2], dt_0[34:34], rg_23r);
  AND2 I1182 (rd_23r1[3:3], dt_0[35:35], rg_23r);
  AND2 I1183 (rd_23r1[4:4], dt_0[36:36], rg_23r);
  AND2 I1184 (rd_23r1[5:5], dt_0[37:37], rg_23r);
  AND2 I1185 (rd_23r1[6:6], dt_0[38:38], rg_23r);
  AND2 I1186 (rd_23r1[7:7], dt_0[39:39], rg_23r);
  AND2 I1187 (rd_23r1[8:8], dt_0[40:40], rg_23r);
  AND2 I1188 (rd_23r1[9:9], dt_0[41:41], rg_23r);
  AND2 I1189 (rd_23r1[10:10], dt_0[42:42], rg_23r);
  AND2 I1190 (rd_23r1[11:11], dt_0[43:43], rg_23r);
  AND2 I1191 (rd_23r1[12:12], dt_0[44:44], rg_23r);
  AND2 I1192 (rd_23r1[13:13], dt_0[45:45], rg_23r);
  AND2 I1193 (rd_23r1[14:14], dt_0[46:46], rg_23r);
  AND2 I1194 (rd_23r1[15:15], dt_0[47:47], rg_23r);
  AND2 I1195 (rd_23r1[16:16], dt_0[48:48], rg_23r);
  AND2 I1196 (rd_23r1[17:17], dt_0[49:49], rg_23r);
  AND2 I1197 (rd_23r1[18:18], dt_0[50:50], rg_23r);
  AND2 I1198 (rd_23r1[19:19], dt_0[51:51], rg_23r);
  AND2 I1199 (rd_23r1[20:20], dt_0[52:52], rg_23r);
  AND2 I1200 (rd_23r1[21:21], dt_0[53:53], rg_23r);
  AND2 I1201 (rd_23r1[22:22], dt_0[54:54], rg_23r);
  AND2 I1202 (rd_23r1[23:23], dt_0[55:55], rg_23r);
  AND2 I1203 (rd_23r1[24:24], dt_0[56:56], rg_23r);
  AND2 I1204 (rd_23r1[25:25], dt_0[57:57], rg_23r);
  AND2 I1205 (rd_23r1[26:26], dt_0[58:58], rg_23r);
  AND2 I1206 (rd_23r1[27:27], dt_0[59:59], rg_23r);
  AND2 I1207 (rd_23r1[28:28], dt_0[60:60], rg_23r);
  AND2 I1208 (rd_23r1[29:29], dt_0[61:61], rg_23r);
  AND2 I1209 (rd_23r1[30:30], dt_0[62:62], rg_23r);
  AND2 I1210 (rd_23r1[31:31], dt_0[63:63], rg_23r);
  AND2 I1211 (rd_23r1[32:32], dt_0[64:64], rg_23r);
  NOR3 I1212 (simp11641_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I1213 (simp11641_0[1:1], rg_3r, rg_4r, rg_5r);
  NOR3 I1214 (simp11641_0[2:2], rg_6r, rg_7r, rg_8r);
  NOR3 I1215 (simp11641_0[3:3], rg_9r, rg_10r, rg_11r);
  NOR3 I1216 (simp11641_0[4:4], rg_12r, rg_13r, rg_14r);
  NOR3 I1217 (simp11641_0[5:5], rg_15r, rg_16r, rg_17r);
  NOR3 I1218 (simp11641_0[6:6], rg_18r, rg_19r, rg_20r);
  NOR3 I1219 (simp11641_0[7:7], rg_21r, rg_22r, rg_23r);
  NOR3 I1220 (simp11641_0[8:8], rg_0a, rg_1a, rg_2a);
  NOR3 I1221 (simp11641_0[9:9], rg_3a, rg_4a, rg_5a);
  NOR3 I1222 (simp11641_0[10:10], rg_6a, rg_7a, rg_8a);
  NOR3 I1223 (simp11641_0[11:11], rg_9a, rg_10a, rg_11a);
  NOR3 I1224 (simp11641_0[12:12], rg_12a, rg_13a, rg_14a);
  NOR3 I1225 (simp11641_0[13:13], rg_15a, rg_16a, rg_17a);
  NOR3 I1226 (simp11641_0[14:14], rg_18a, rg_19a, rg_20a);
  NOR3 I1227 (simp11641_0[15:15], rg_21a, rg_22a, rg_23a);
  NAND3 I1228 (simp11642_0[0:0], simp11641_0[0:0], simp11641_0[1:1], simp11641_0[2:2]);
  NAND3 I1229 (simp11642_0[1:1], simp11641_0[3:3], simp11641_0[4:4], simp11641_0[5:5]);
  NAND3 I1230 (simp11642_0[2:2], simp11641_0[6:6], simp11641_0[7:7], simp11641_0[8:8]);
  NAND3 I1231 (simp11642_0[3:3], simp11641_0[9:9], simp11641_0[10:10], simp11641_0[11:11]);
  NAND3 I1232 (simp11642_0[4:4], simp11641_0[12:12], simp11641_0[13:13], simp11641_0[14:14]);
  INV I1233 (simp11642_0[5:5], simp11641_0[15:15]);
  NOR3 I1234 (simp11643_0[0:0], simp11642_0[0:0], simp11642_0[1:1], simp11642_0[2:2]);
  NOR3 I1235 (simp11643_0[1:1], simp11642_0[3:3], simp11642_0[4:4], simp11642_0[5:5]);
  NAND2 I1236 (anyread_0, simp11643_0[0:0], simp11643_0[1:1]);
  BUFF I1237 (wg_0a, wd_0a);
  BUFF I1238 (rg_0a, rd_0a);
  BUFF I1239 (rg_1a, rd_1a);
  BUFF I1240 (rg_2a, rd_2a);
  BUFF I1241 (rg_3a, rd_3a);
  BUFF I1242 (rg_4a, rd_4a);
  BUFF I1243 (rg_5a, rd_5a);
  BUFF I1244 (rg_6a, rd_6a);
  BUFF I1245 (rg_7a, rd_7a);
  BUFF I1246 (rg_8a, rd_8a);
  BUFF I1247 (rg_9a, rd_9a);
  BUFF I1248 (rg_10a, rd_10a);
  BUFF I1249 (rg_11a, rd_11a);
  BUFF I1250 (rg_12a, rd_12a);
  BUFF I1251 (rg_13a, rd_13a);
  BUFF I1252 (rg_14a, rd_14a);
  BUFF I1253 (rg_15a, rd_15a);
  BUFF I1254 (rg_16a, rd_16a);
  BUFF I1255 (rg_17a, rd_17a);
  BUFF I1256 (rg_18a, rd_18a);
  BUFF I1257 (rg_19a, rd_19a);
  BUFF I1258 (rg_20a, rd_20a);
  BUFF I1259 (rg_21a, rd_21a);
  BUFF I1260 (rg_22a, rd_22a);
  BUFF I1261 (rg_23a, rd_23a);
endmodule

// tkj65m65_0 TeakJ [Many [65,0],One 65]
module tkj65m65_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [64:0] i_0r0;
  input [64:0] i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  output [64:0] o_0r0;
  output [64:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [64:0] joinf_0;
  wire [64:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joinf_0[32:32], i_0r0[32:32]);
  BUFF I33 (joinf_0[33:33], i_0r0[33:33]);
  BUFF I34 (joinf_0[34:34], i_0r0[34:34]);
  BUFF I35 (joinf_0[35:35], i_0r0[35:35]);
  BUFF I36 (joinf_0[36:36], i_0r0[36:36]);
  BUFF I37 (joinf_0[37:37], i_0r0[37:37]);
  BUFF I38 (joinf_0[38:38], i_0r0[38:38]);
  BUFF I39 (joinf_0[39:39], i_0r0[39:39]);
  BUFF I40 (joinf_0[40:40], i_0r0[40:40]);
  BUFF I41 (joinf_0[41:41], i_0r0[41:41]);
  BUFF I42 (joinf_0[42:42], i_0r0[42:42]);
  BUFF I43 (joinf_0[43:43], i_0r0[43:43]);
  BUFF I44 (joinf_0[44:44], i_0r0[44:44]);
  BUFF I45 (joinf_0[45:45], i_0r0[45:45]);
  BUFF I46 (joinf_0[46:46], i_0r0[46:46]);
  BUFF I47 (joinf_0[47:47], i_0r0[47:47]);
  BUFF I48 (joinf_0[48:48], i_0r0[48:48]);
  BUFF I49 (joinf_0[49:49], i_0r0[49:49]);
  BUFF I50 (joinf_0[50:50], i_0r0[50:50]);
  BUFF I51 (joinf_0[51:51], i_0r0[51:51]);
  BUFF I52 (joinf_0[52:52], i_0r0[52:52]);
  BUFF I53 (joinf_0[53:53], i_0r0[53:53]);
  BUFF I54 (joinf_0[54:54], i_0r0[54:54]);
  BUFF I55 (joinf_0[55:55], i_0r0[55:55]);
  BUFF I56 (joinf_0[56:56], i_0r0[56:56]);
  BUFF I57 (joinf_0[57:57], i_0r0[57:57]);
  BUFF I58 (joinf_0[58:58], i_0r0[58:58]);
  BUFF I59 (joinf_0[59:59], i_0r0[59:59]);
  BUFF I60 (joinf_0[60:60], i_0r0[60:60]);
  BUFF I61 (joinf_0[61:61], i_0r0[61:61]);
  BUFF I62 (joinf_0[62:62], i_0r0[62:62]);
  BUFF I63 (joinf_0[63:63], i_0r0[63:63]);
  BUFF I64 (joinf_0[64:64], i_0r0[64:64]);
  BUFF I65 (joint_0[0:0], i_0r1[0:0]);
  BUFF I66 (joint_0[1:1], i_0r1[1:1]);
  BUFF I67 (joint_0[2:2], i_0r1[2:2]);
  BUFF I68 (joint_0[3:3], i_0r1[3:3]);
  BUFF I69 (joint_0[4:4], i_0r1[4:4]);
  BUFF I70 (joint_0[5:5], i_0r1[5:5]);
  BUFF I71 (joint_0[6:6], i_0r1[6:6]);
  BUFF I72 (joint_0[7:7], i_0r1[7:7]);
  BUFF I73 (joint_0[8:8], i_0r1[8:8]);
  BUFF I74 (joint_0[9:9], i_0r1[9:9]);
  BUFF I75 (joint_0[10:10], i_0r1[10:10]);
  BUFF I76 (joint_0[11:11], i_0r1[11:11]);
  BUFF I77 (joint_0[12:12], i_0r1[12:12]);
  BUFF I78 (joint_0[13:13], i_0r1[13:13]);
  BUFF I79 (joint_0[14:14], i_0r1[14:14]);
  BUFF I80 (joint_0[15:15], i_0r1[15:15]);
  BUFF I81 (joint_0[16:16], i_0r1[16:16]);
  BUFF I82 (joint_0[17:17], i_0r1[17:17]);
  BUFF I83 (joint_0[18:18], i_0r1[18:18]);
  BUFF I84 (joint_0[19:19], i_0r1[19:19]);
  BUFF I85 (joint_0[20:20], i_0r1[20:20]);
  BUFF I86 (joint_0[21:21], i_0r1[21:21]);
  BUFF I87 (joint_0[22:22], i_0r1[22:22]);
  BUFF I88 (joint_0[23:23], i_0r1[23:23]);
  BUFF I89 (joint_0[24:24], i_0r1[24:24]);
  BUFF I90 (joint_0[25:25], i_0r1[25:25]);
  BUFF I91 (joint_0[26:26], i_0r1[26:26]);
  BUFF I92 (joint_0[27:27], i_0r1[27:27]);
  BUFF I93 (joint_0[28:28], i_0r1[28:28]);
  BUFF I94 (joint_0[29:29], i_0r1[29:29]);
  BUFF I95 (joint_0[30:30], i_0r1[30:30]);
  BUFF I96 (joint_0[31:31], i_0r1[31:31]);
  BUFF I97 (joint_0[32:32], i_0r1[32:32]);
  BUFF I98 (joint_0[33:33], i_0r1[33:33]);
  BUFF I99 (joint_0[34:34], i_0r1[34:34]);
  BUFF I100 (joint_0[35:35], i_0r1[35:35]);
  BUFF I101 (joint_0[36:36], i_0r1[36:36]);
  BUFF I102 (joint_0[37:37], i_0r1[37:37]);
  BUFF I103 (joint_0[38:38], i_0r1[38:38]);
  BUFF I104 (joint_0[39:39], i_0r1[39:39]);
  BUFF I105 (joint_0[40:40], i_0r1[40:40]);
  BUFF I106 (joint_0[41:41], i_0r1[41:41]);
  BUFF I107 (joint_0[42:42], i_0r1[42:42]);
  BUFF I108 (joint_0[43:43], i_0r1[43:43]);
  BUFF I109 (joint_0[44:44], i_0r1[44:44]);
  BUFF I110 (joint_0[45:45], i_0r1[45:45]);
  BUFF I111 (joint_0[46:46], i_0r1[46:46]);
  BUFF I112 (joint_0[47:47], i_0r1[47:47]);
  BUFF I113 (joint_0[48:48], i_0r1[48:48]);
  BUFF I114 (joint_0[49:49], i_0r1[49:49]);
  BUFF I115 (joint_0[50:50], i_0r1[50:50]);
  BUFF I116 (joint_0[51:51], i_0r1[51:51]);
  BUFF I117 (joint_0[52:52], i_0r1[52:52]);
  BUFF I118 (joint_0[53:53], i_0r1[53:53]);
  BUFF I119 (joint_0[54:54], i_0r1[54:54]);
  BUFF I120 (joint_0[55:55], i_0r1[55:55]);
  BUFF I121 (joint_0[56:56], i_0r1[56:56]);
  BUFF I122 (joint_0[57:57], i_0r1[57:57]);
  BUFF I123 (joint_0[58:58], i_0r1[58:58]);
  BUFF I124 (joint_0[59:59], i_0r1[59:59]);
  BUFF I125 (joint_0[60:60], i_0r1[60:60]);
  BUFF I126 (joint_0[61:61], i_0r1[61:61]);
  BUFF I127 (joint_0[62:62], i_0r1[62:62]);
  BUFF I128 (joint_0[63:63], i_0r1[63:63]);
  BUFF I129 (joint_0[64:64], i_0r1[64:64]);
  BUFF I130 (icomplete_0, i_1r);
  C2 I131 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I132 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I133 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I134 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I135 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I136 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I137 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I138 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I139 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I140 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I141 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I142 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I143 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I144 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I145 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I146 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I147 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I148 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I149 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I150 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I151 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I152 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I153 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I154 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I155 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I156 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I157 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I158 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I159 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I160 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I161 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I162 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I163 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I164 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I165 (o_0r0[33:33], joinf_0[33:33]);
  BUFF I166 (o_0r0[34:34], joinf_0[34:34]);
  BUFF I167 (o_0r0[35:35], joinf_0[35:35]);
  BUFF I168 (o_0r0[36:36], joinf_0[36:36]);
  BUFF I169 (o_0r0[37:37], joinf_0[37:37]);
  BUFF I170 (o_0r0[38:38], joinf_0[38:38]);
  BUFF I171 (o_0r0[39:39], joinf_0[39:39]);
  BUFF I172 (o_0r0[40:40], joinf_0[40:40]);
  BUFF I173 (o_0r0[41:41], joinf_0[41:41]);
  BUFF I174 (o_0r0[42:42], joinf_0[42:42]);
  BUFF I175 (o_0r0[43:43], joinf_0[43:43]);
  BUFF I176 (o_0r0[44:44], joinf_0[44:44]);
  BUFF I177 (o_0r0[45:45], joinf_0[45:45]);
  BUFF I178 (o_0r0[46:46], joinf_0[46:46]);
  BUFF I179 (o_0r0[47:47], joinf_0[47:47]);
  BUFF I180 (o_0r0[48:48], joinf_0[48:48]);
  BUFF I181 (o_0r0[49:49], joinf_0[49:49]);
  BUFF I182 (o_0r0[50:50], joinf_0[50:50]);
  BUFF I183 (o_0r0[51:51], joinf_0[51:51]);
  BUFF I184 (o_0r0[52:52], joinf_0[52:52]);
  BUFF I185 (o_0r0[53:53], joinf_0[53:53]);
  BUFF I186 (o_0r0[54:54], joinf_0[54:54]);
  BUFF I187 (o_0r0[55:55], joinf_0[55:55]);
  BUFF I188 (o_0r0[56:56], joinf_0[56:56]);
  BUFF I189 (o_0r0[57:57], joinf_0[57:57]);
  BUFF I190 (o_0r0[58:58], joinf_0[58:58]);
  BUFF I191 (o_0r0[59:59], joinf_0[59:59]);
  BUFF I192 (o_0r0[60:60], joinf_0[60:60]);
  BUFF I193 (o_0r0[61:61], joinf_0[61:61]);
  BUFF I194 (o_0r0[62:62], joinf_0[62:62]);
  BUFF I195 (o_0r0[63:63], joinf_0[63:63]);
  BUFF I196 (o_0r0[64:64], joinf_0[64:64]);
  BUFF I197 (o_0r1[1:1], joint_0[1:1]);
  BUFF I198 (o_0r1[2:2], joint_0[2:2]);
  BUFF I199 (o_0r1[3:3], joint_0[3:3]);
  BUFF I200 (o_0r1[4:4], joint_0[4:4]);
  BUFF I201 (o_0r1[5:5], joint_0[5:5]);
  BUFF I202 (o_0r1[6:6], joint_0[6:6]);
  BUFF I203 (o_0r1[7:7], joint_0[7:7]);
  BUFF I204 (o_0r1[8:8], joint_0[8:8]);
  BUFF I205 (o_0r1[9:9], joint_0[9:9]);
  BUFF I206 (o_0r1[10:10], joint_0[10:10]);
  BUFF I207 (o_0r1[11:11], joint_0[11:11]);
  BUFF I208 (o_0r1[12:12], joint_0[12:12]);
  BUFF I209 (o_0r1[13:13], joint_0[13:13]);
  BUFF I210 (o_0r1[14:14], joint_0[14:14]);
  BUFF I211 (o_0r1[15:15], joint_0[15:15]);
  BUFF I212 (o_0r1[16:16], joint_0[16:16]);
  BUFF I213 (o_0r1[17:17], joint_0[17:17]);
  BUFF I214 (o_0r1[18:18], joint_0[18:18]);
  BUFF I215 (o_0r1[19:19], joint_0[19:19]);
  BUFF I216 (o_0r1[20:20], joint_0[20:20]);
  BUFF I217 (o_0r1[21:21], joint_0[21:21]);
  BUFF I218 (o_0r1[22:22], joint_0[22:22]);
  BUFF I219 (o_0r1[23:23], joint_0[23:23]);
  BUFF I220 (o_0r1[24:24], joint_0[24:24]);
  BUFF I221 (o_0r1[25:25], joint_0[25:25]);
  BUFF I222 (o_0r1[26:26], joint_0[26:26]);
  BUFF I223 (o_0r1[27:27], joint_0[27:27]);
  BUFF I224 (o_0r1[28:28], joint_0[28:28]);
  BUFF I225 (o_0r1[29:29], joint_0[29:29]);
  BUFF I226 (o_0r1[30:30], joint_0[30:30]);
  BUFF I227 (o_0r1[31:31], joint_0[31:31]);
  BUFF I228 (o_0r1[32:32], joint_0[32:32]);
  BUFF I229 (o_0r1[33:33], joint_0[33:33]);
  BUFF I230 (o_0r1[34:34], joint_0[34:34]);
  BUFF I231 (o_0r1[35:35], joint_0[35:35]);
  BUFF I232 (o_0r1[36:36], joint_0[36:36]);
  BUFF I233 (o_0r1[37:37], joint_0[37:37]);
  BUFF I234 (o_0r1[38:38], joint_0[38:38]);
  BUFF I235 (o_0r1[39:39], joint_0[39:39]);
  BUFF I236 (o_0r1[40:40], joint_0[40:40]);
  BUFF I237 (o_0r1[41:41], joint_0[41:41]);
  BUFF I238 (o_0r1[42:42], joint_0[42:42]);
  BUFF I239 (o_0r1[43:43], joint_0[43:43]);
  BUFF I240 (o_0r1[44:44], joint_0[44:44]);
  BUFF I241 (o_0r1[45:45], joint_0[45:45]);
  BUFF I242 (o_0r1[46:46], joint_0[46:46]);
  BUFF I243 (o_0r1[47:47], joint_0[47:47]);
  BUFF I244 (o_0r1[48:48], joint_0[48:48]);
  BUFF I245 (o_0r1[49:49], joint_0[49:49]);
  BUFF I246 (o_0r1[50:50], joint_0[50:50]);
  BUFF I247 (o_0r1[51:51], joint_0[51:51]);
  BUFF I248 (o_0r1[52:52], joint_0[52:52]);
  BUFF I249 (o_0r1[53:53], joint_0[53:53]);
  BUFF I250 (o_0r1[54:54], joint_0[54:54]);
  BUFF I251 (o_0r1[55:55], joint_0[55:55]);
  BUFF I252 (o_0r1[56:56], joint_0[56:56]);
  BUFF I253 (o_0r1[57:57], joint_0[57:57]);
  BUFF I254 (o_0r1[58:58], joint_0[58:58]);
  BUFF I255 (o_0r1[59:59], joint_0[59:59]);
  BUFF I256 (o_0r1[60:60], joint_0[60:60]);
  BUFF I257 (o_0r1[61:61], joint_0[61:61]);
  BUFF I258 (o_0r1[62:62], joint_0[62:62]);
  BUFF I259 (o_0r1[63:63], joint_0[63:63]);
  BUFF I260 (o_0r1[64:64], joint_0[64:64]);
  BUFF I261 (i_0a, o_0a);
  BUFF I262 (i_1a, o_0a);
endmodule

// tkf74mo0w0_o0w74 TeakF [0,0] [One 74,Many [0,74]]
module tkf74mo0w0_o0w74 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [73:0] i_0r0;
  input [73:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [73:0] o_1r0;
  output [73:0] o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_1r0[0:0], i_0r0[0:0]);
  BUFF I3 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I4 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I5 (o_1r0[3:3], i_0r0[3:3]);
  BUFF I6 (o_1r0[4:4], i_0r0[4:4]);
  BUFF I7 (o_1r0[5:5], i_0r0[5:5]);
  BUFF I8 (o_1r0[6:6], i_0r0[6:6]);
  BUFF I9 (o_1r0[7:7], i_0r0[7:7]);
  BUFF I10 (o_1r0[8:8], i_0r0[8:8]);
  BUFF I11 (o_1r0[9:9], i_0r0[9:9]);
  BUFF I12 (o_1r0[10:10], i_0r0[10:10]);
  BUFF I13 (o_1r0[11:11], i_0r0[11:11]);
  BUFF I14 (o_1r0[12:12], i_0r0[12:12]);
  BUFF I15 (o_1r0[13:13], i_0r0[13:13]);
  BUFF I16 (o_1r0[14:14], i_0r0[14:14]);
  BUFF I17 (o_1r0[15:15], i_0r0[15:15]);
  BUFF I18 (o_1r0[16:16], i_0r0[16:16]);
  BUFF I19 (o_1r0[17:17], i_0r0[17:17]);
  BUFF I20 (o_1r0[18:18], i_0r0[18:18]);
  BUFF I21 (o_1r0[19:19], i_0r0[19:19]);
  BUFF I22 (o_1r0[20:20], i_0r0[20:20]);
  BUFF I23 (o_1r0[21:21], i_0r0[21:21]);
  BUFF I24 (o_1r0[22:22], i_0r0[22:22]);
  BUFF I25 (o_1r0[23:23], i_0r0[23:23]);
  BUFF I26 (o_1r0[24:24], i_0r0[24:24]);
  BUFF I27 (o_1r0[25:25], i_0r0[25:25]);
  BUFF I28 (o_1r0[26:26], i_0r0[26:26]);
  BUFF I29 (o_1r0[27:27], i_0r0[27:27]);
  BUFF I30 (o_1r0[28:28], i_0r0[28:28]);
  BUFF I31 (o_1r0[29:29], i_0r0[29:29]);
  BUFF I32 (o_1r0[30:30], i_0r0[30:30]);
  BUFF I33 (o_1r0[31:31], i_0r0[31:31]);
  BUFF I34 (o_1r0[32:32], i_0r0[32:32]);
  BUFF I35 (o_1r0[33:33], i_0r0[33:33]);
  BUFF I36 (o_1r0[34:34], i_0r0[34:34]);
  BUFF I37 (o_1r0[35:35], i_0r0[35:35]);
  BUFF I38 (o_1r0[36:36], i_0r0[36:36]);
  BUFF I39 (o_1r0[37:37], i_0r0[37:37]);
  BUFF I40 (o_1r0[38:38], i_0r0[38:38]);
  BUFF I41 (o_1r0[39:39], i_0r0[39:39]);
  BUFF I42 (o_1r0[40:40], i_0r0[40:40]);
  BUFF I43 (o_1r0[41:41], i_0r0[41:41]);
  BUFF I44 (o_1r0[42:42], i_0r0[42:42]);
  BUFF I45 (o_1r0[43:43], i_0r0[43:43]);
  BUFF I46 (o_1r0[44:44], i_0r0[44:44]);
  BUFF I47 (o_1r0[45:45], i_0r0[45:45]);
  BUFF I48 (o_1r0[46:46], i_0r0[46:46]);
  BUFF I49 (o_1r0[47:47], i_0r0[47:47]);
  BUFF I50 (o_1r0[48:48], i_0r0[48:48]);
  BUFF I51 (o_1r0[49:49], i_0r0[49:49]);
  BUFF I52 (o_1r0[50:50], i_0r0[50:50]);
  BUFF I53 (o_1r0[51:51], i_0r0[51:51]);
  BUFF I54 (o_1r0[52:52], i_0r0[52:52]);
  BUFF I55 (o_1r0[53:53], i_0r0[53:53]);
  BUFF I56 (o_1r0[54:54], i_0r0[54:54]);
  BUFF I57 (o_1r0[55:55], i_0r0[55:55]);
  BUFF I58 (o_1r0[56:56], i_0r0[56:56]);
  BUFF I59 (o_1r0[57:57], i_0r0[57:57]);
  BUFF I60 (o_1r0[58:58], i_0r0[58:58]);
  BUFF I61 (o_1r0[59:59], i_0r0[59:59]);
  BUFF I62 (o_1r0[60:60], i_0r0[60:60]);
  BUFF I63 (o_1r0[61:61], i_0r0[61:61]);
  BUFF I64 (o_1r0[62:62], i_0r0[62:62]);
  BUFF I65 (o_1r0[63:63], i_0r0[63:63]);
  BUFF I66 (o_1r0[64:64], i_0r0[64:64]);
  BUFF I67 (o_1r0[65:65], i_0r0[65:65]);
  BUFF I68 (o_1r0[66:66], i_0r0[66:66]);
  BUFF I69 (o_1r0[67:67], i_0r0[67:67]);
  BUFF I70 (o_1r0[68:68], i_0r0[68:68]);
  BUFF I71 (o_1r0[69:69], i_0r0[69:69]);
  BUFF I72 (o_1r0[70:70], i_0r0[70:70]);
  BUFF I73 (o_1r0[71:71], i_0r0[71:71]);
  BUFF I74 (o_1r0[72:72], i_0r0[72:72]);
  BUFF I75 (o_1r0[73:73], i_0r0[73:73]);
  BUFF I76 (o_1r1[0:0], i_0r1[0:0]);
  BUFF I77 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I78 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I79 (o_1r1[3:3], i_0r1[3:3]);
  BUFF I80 (o_1r1[4:4], i_0r1[4:4]);
  BUFF I81 (o_1r1[5:5], i_0r1[5:5]);
  BUFF I82 (o_1r1[6:6], i_0r1[6:6]);
  BUFF I83 (o_1r1[7:7], i_0r1[7:7]);
  BUFF I84 (o_1r1[8:8], i_0r1[8:8]);
  BUFF I85 (o_1r1[9:9], i_0r1[9:9]);
  BUFF I86 (o_1r1[10:10], i_0r1[10:10]);
  BUFF I87 (o_1r1[11:11], i_0r1[11:11]);
  BUFF I88 (o_1r1[12:12], i_0r1[12:12]);
  BUFF I89 (o_1r1[13:13], i_0r1[13:13]);
  BUFF I90 (o_1r1[14:14], i_0r1[14:14]);
  BUFF I91 (o_1r1[15:15], i_0r1[15:15]);
  BUFF I92 (o_1r1[16:16], i_0r1[16:16]);
  BUFF I93 (o_1r1[17:17], i_0r1[17:17]);
  BUFF I94 (o_1r1[18:18], i_0r1[18:18]);
  BUFF I95 (o_1r1[19:19], i_0r1[19:19]);
  BUFF I96 (o_1r1[20:20], i_0r1[20:20]);
  BUFF I97 (o_1r1[21:21], i_0r1[21:21]);
  BUFF I98 (o_1r1[22:22], i_0r1[22:22]);
  BUFF I99 (o_1r1[23:23], i_0r1[23:23]);
  BUFF I100 (o_1r1[24:24], i_0r1[24:24]);
  BUFF I101 (o_1r1[25:25], i_0r1[25:25]);
  BUFF I102 (o_1r1[26:26], i_0r1[26:26]);
  BUFF I103 (o_1r1[27:27], i_0r1[27:27]);
  BUFF I104 (o_1r1[28:28], i_0r1[28:28]);
  BUFF I105 (o_1r1[29:29], i_0r1[29:29]);
  BUFF I106 (o_1r1[30:30], i_0r1[30:30]);
  BUFF I107 (o_1r1[31:31], i_0r1[31:31]);
  BUFF I108 (o_1r1[32:32], i_0r1[32:32]);
  BUFF I109 (o_1r1[33:33], i_0r1[33:33]);
  BUFF I110 (o_1r1[34:34], i_0r1[34:34]);
  BUFF I111 (o_1r1[35:35], i_0r1[35:35]);
  BUFF I112 (o_1r1[36:36], i_0r1[36:36]);
  BUFF I113 (o_1r1[37:37], i_0r1[37:37]);
  BUFF I114 (o_1r1[38:38], i_0r1[38:38]);
  BUFF I115 (o_1r1[39:39], i_0r1[39:39]);
  BUFF I116 (o_1r1[40:40], i_0r1[40:40]);
  BUFF I117 (o_1r1[41:41], i_0r1[41:41]);
  BUFF I118 (o_1r1[42:42], i_0r1[42:42]);
  BUFF I119 (o_1r1[43:43], i_0r1[43:43]);
  BUFF I120 (o_1r1[44:44], i_0r1[44:44]);
  BUFF I121 (o_1r1[45:45], i_0r1[45:45]);
  BUFF I122 (o_1r1[46:46], i_0r1[46:46]);
  BUFF I123 (o_1r1[47:47], i_0r1[47:47]);
  BUFF I124 (o_1r1[48:48], i_0r1[48:48]);
  BUFF I125 (o_1r1[49:49], i_0r1[49:49]);
  BUFF I126 (o_1r1[50:50], i_0r1[50:50]);
  BUFF I127 (o_1r1[51:51], i_0r1[51:51]);
  BUFF I128 (o_1r1[52:52], i_0r1[52:52]);
  BUFF I129 (o_1r1[53:53], i_0r1[53:53]);
  BUFF I130 (o_1r1[54:54], i_0r1[54:54]);
  BUFF I131 (o_1r1[55:55], i_0r1[55:55]);
  BUFF I132 (o_1r1[56:56], i_0r1[56:56]);
  BUFF I133 (o_1r1[57:57], i_0r1[57:57]);
  BUFF I134 (o_1r1[58:58], i_0r1[58:58]);
  BUFF I135 (o_1r1[59:59], i_0r1[59:59]);
  BUFF I136 (o_1r1[60:60], i_0r1[60:60]);
  BUFF I137 (o_1r1[61:61], i_0r1[61:61]);
  BUFF I138 (o_1r1[62:62], i_0r1[62:62]);
  BUFF I139 (o_1r1[63:63], i_0r1[63:63]);
  BUFF I140 (o_1r1[64:64], i_0r1[64:64]);
  BUFF I141 (o_1r1[65:65], i_0r1[65:65]);
  BUFF I142 (o_1r1[66:66], i_0r1[66:66]);
  BUFF I143 (o_1r1[67:67], i_0r1[67:67]);
  BUFF I144 (o_1r1[68:68], i_0r1[68:68]);
  BUFF I145 (o_1r1[69:69], i_0r1[69:69]);
  BUFF I146 (o_1r1[70:70], i_0r1[70:70]);
  BUFF I147 (o_1r1[71:71], i_0r1[71:71]);
  BUFF I148 (o_1r1[72:72], i_0r1[72:72]);
  BUFF I149 (o_1r1[73:73], i_0r1[73:73]);
  BUFF I150 (o_0r, icomplete_0);
  C3 I151 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tkm5x74b TeakM [Many [74,74,74,74,74],One 74]
module tkm5x74b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, i_4r0, i_4r1, i_4a, o_0r0, o_0r1, o_0a, reset);
  input [73:0] i_0r0;
  input [73:0] i_0r1;
  output i_0a;
  input [73:0] i_1r0;
  input [73:0] i_1r1;
  output i_1a;
  input [73:0] i_2r0;
  input [73:0] i_2r1;
  output i_2a;
  input [73:0] i_3r0;
  input [73:0] i_3r1;
  output i_3a;
  input [73:0] i_4r0;
  input [73:0] i_4r1;
  output i_4a;
  output [73:0] o_0r0;
  output [73:0] o_0r1;
  input o_0a;
  input reset;
  wire [73:0] gfint_0;
  wire [73:0] gfint_1;
  wire [73:0] gfint_2;
  wire [73:0] gfint_3;
  wire [73:0] gfint_4;
  wire [73:0] gtint_0;
  wire [73:0] gtint_1;
  wire [73:0] gtint_2;
  wire [73:0] gtint_3;
  wire [73:0] gtint_4;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire choice_4;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire icomp_3;
  wire icomp_4;
  wire nchosen_0;
  wire [1:0] simp221_0;
  wire [1:0] simp231_0;
  wire [1:0] simp241_0;
  wire [1:0] simp251_0;
  wire [1:0] simp261_0;
  wire [1:0] simp271_0;
  wire [1:0] simp281_0;
  wire [1:0] simp291_0;
  wire [1:0] simp301_0;
  wire [1:0] simp311_0;
  wire [1:0] simp321_0;
  wire [1:0] simp331_0;
  wire [1:0] simp341_0;
  wire [1:0] simp351_0;
  wire [1:0] simp361_0;
  wire [1:0] simp371_0;
  wire [1:0] simp381_0;
  wire [1:0] simp391_0;
  wire [1:0] simp401_0;
  wire [1:0] simp411_0;
  wire [1:0] simp421_0;
  wire [1:0] simp431_0;
  wire [1:0] simp441_0;
  wire [1:0] simp451_0;
  wire [1:0] simp461_0;
  wire [1:0] simp471_0;
  wire [1:0] simp481_0;
  wire [1:0] simp491_0;
  wire [1:0] simp501_0;
  wire [1:0] simp511_0;
  wire [1:0] simp521_0;
  wire [1:0] simp531_0;
  wire [1:0] simp541_0;
  wire [1:0] simp551_0;
  wire [1:0] simp561_0;
  wire [1:0] simp571_0;
  wire [1:0] simp581_0;
  wire [1:0] simp591_0;
  wire [1:0] simp601_0;
  wire [1:0] simp611_0;
  wire [1:0] simp621_0;
  wire [1:0] simp631_0;
  wire [1:0] simp641_0;
  wire [1:0] simp651_0;
  wire [1:0] simp661_0;
  wire [1:0] simp671_0;
  wire [1:0] simp681_0;
  wire [1:0] simp691_0;
  wire [1:0] simp701_0;
  wire [1:0] simp711_0;
  wire [1:0] simp721_0;
  wire [1:0] simp731_0;
  wire [1:0] simp741_0;
  wire [1:0] simp751_0;
  wire [1:0] simp761_0;
  wire [1:0] simp771_0;
  wire [1:0] simp781_0;
  wire [1:0] simp791_0;
  wire [1:0] simp801_0;
  wire [1:0] simp811_0;
  wire [1:0] simp821_0;
  wire [1:0] simp831_0;
  wire [1:0] simp841_0;
  wire [1:0] simp851_0;
  wire [1:0] simp861_0;
  wire [1:0] simp871_0;
  wire [1:0] simp881_0;
  wire [1:0] simp891_0;
  wire [1:0] simp901_0;
  wire [1:0] simp911_0;
  wire [1:0] simp921_0;
  wire [1:0] simp931_0;
  wire [1:0] simp941_0;
  wire [1:0] simp951_0;
  wire [1:0] simp961_0;
  wire [1:0] simp971_0;
  wire [1:0] simp981_0;
  wire [1:0] simp991_0;
  wire [1:0] simp1001_0;
  wire [1:0] simp1011_0;
  wire [1:0] simp1021_0;
  wire [1:0] simp1031_0;
  wire [1:0] simp1041_0;
  wire [1:0] simp1051_0;
  wire [1:0] simp1061_0;
  wire [1:0] simp1071_0;
  wire [1:0] simp1081_0;
  wire [1:0] simp1091_0;
  wire [1:0] simp1101_0;
  wire [1:0] simp1111_0;
  wire [1:0] simp1121_0;
  wire [1:0] simp1131_0;
  wire [1:0] simp1141_0;
  wire [1:0] simp1151_0;
  wire [1:0] simp1161_0;
  wire [1:0] simp1171_0;
  wire [1:0] simp1181_0;
  wire [1:0] simp1191_0;
  wire [1:0] simp1201_0;
  wire [1:0] simp1211_0;
  wire [1:0] simp1221_0;
  wire [1:0] simp1231_0;
  wire [1:0] simp1241_0;
  wire [1:0] simp1251_0;
  wire [1:0] simp1261_0;
  wire [1:0] simp1271_0;
  wire [1:0] simp1281_0;
  wire [1:0] simp1291_0;
  wire [1:0] simp1301_0;
  wire [1:0] simp1311_0;
  wire [1:0] simp1321_0;
  wire [1:0] simp1331_0;
  wire [1:0] simp1341_0;
  wire [1:0] simp1351_0;
  wire [1:0] simp1361_0;
  wire [1:0] simp1371_0;
  wire [1:0] simp1381_0;
  wire [1:0] simp1391_0;
  wire [1:0] simp1401_0;
  wire [1:0] simp1411_0;
  wire [1:0] simp1421_0;
  wire [1:0] simp1431_0;
  wire [1:0] simp1441_0;
  wire [1:0] simp1451_0;
  wire [1:0] simp1461_0;
  wire [1:0] simp1471_0;
  wire [1:0] simp1481_0;
  wire [1:0] simp1491_0;
  wire [1:0] simp1501_0;
  wire [1:0] simp1511_0;
  wire [1:0] simp1521_0;
  wire [1:0] simp1531_0;
  wire [1:0] simp1541_0;
  wire [1:0] simp1551_0;
  wire [1:0] simp1561_0;
  wire [1:0] simp1571_0;
  wire [1:0] simp1581_0;
  wire [1:0] simp1591_0;
  wire [1:0] simp1601_0;
  wire [1:0] simp1611_0;
  wire [1:0] simp1621_0;
  wire [1:0] simp1631_0;
  wire [1:0] simp1641_0;
  wire [1:0] simp1651_0;
  wire [1:0] simp1661_0;
  wire [1:0] simp1671_0;
  wire [1:0] simp1681_0;
  wire [1:0] simp1691_0;
  wire [73:0] comp0_0;
  wire [24:0] simp9851_0;
  wire [8:0] simp9852_0;
  wire [2:0] simp9853_0;
  wire [73:0] comp1_0;
  wire [24:0] simp10611_0;
  wire [8:0] simp10612_0;
  wire [2:0] simp10613_0;
  wire [73:0] comp2_0;
  wire [24:0] simp11371_0;
  wire [8:0] simp11372_0;
  wire [2:0] simp11373_0;
  wire [73:0] comp3_0;
  wire [24:0] simp12131_0;
  wire [8:0] simp12132_0;
  wire [2:0] simp12133_0;
  wire [73:0] comp4_0;
  wire [24:0] simp12891_0;
  wire [8:0] simp12892_0;
  wire [2:0] simp12893_0;
  wire [1:0] simp12951_0;
  NOR3 I0 (simp221_0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  NOR2 I1 (simp221_0[1:1], gfint_3[0:0], gfint_4[0:0]);
  NAND2 I2 (o_0r0[0:0], simp221_0[0:0], simp221_0[1:1]);
  NOR3 I3 (simp231_0[0:0], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  NOR2 I4 (simp231_0[1:1], gfint_3[1:1], gfint_4[1:1]);
  NAND2 I5 (o_0r0[1:1], simp231_0[0:0], simp231_0[1:1]);
  NOR3 I6 (simp241_0[0:0], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  NOR2 I7 (simp241_0[1:1], gfint_3[2:2], gfint_4[2:2]);
  NAND2 I8 (o_0r0[2:2], simp241_0[0:0], simp241_0[1:1]);
  NOR3 I9 (simp251_0[0:0], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  NOR2 I10 (simp251_0[1:1], gfint_3[3:3], gfint_4[3:3]);
  NAND2 I11 (o_0r0[3:3], simp251_0[0:0], simp251_0[1:1]);
  NOR3 I12 (simp261_0[0:0], gfint_0[4:4], gfint_1[4:4], gfint_2[4:4]);
  NOR2 I13 (simp261_0[1:1], gfint_3[4:4], gfint_4[4:4]);
  NAND2 I14 (o_0r0[4:4], simp261_0[0:0], simp261_0[1:1]);
  NOR3 I15 (simp271_0[0:0], gfint_0[5:5], gfint_1[5:5], gfint_2[5:5]);
  NOR2 I16 (simp271_0[1:1], gfint_3[5:5], gfint_4[5:5]);
  NAND2 I17 (o_0r0[5:5], simp271_0[0:0], simp271_0[1:1]);
  NOR3 I18 (simp281_0[0:0], gfint_0[6:6], gfint_1[6:6], gfint_2[6:6]);
  NOR2 I19 (simp281_0[1:1], gfint_3[6:6], gfint_4[6:6]);
  NAND2 I20 (o_0r0[6:6], simp281_0[0:0], simp281_0[1:1]);
  NOR3 I21 (simp291_0[0:0], gfint_0[7:7], gfint_1[7:7], gfint_2[7:7]);
  NOR2 I22 (simp291_0[1:1], gfint_3[7:7], gfint_4[7:7]);
  NAND2 I23 (o_0r0[7:7], simp291_0[0:0], simp291_0[1:1]);
  NOR3 I24 (simp301_0[0:0], gfint_0[8:8], gfint_1[8:8], gfint_2[8:8]);
  NOR2 I25 (simp301_0[1:1], gfint_3[8:8], gfint_4[8:8]);
  NAND2 I26 (o_0r0[8:8], simp301_0[0:0], simp301_0[1:1]);
  NOR3 I27 (simp311_0[0:0], gfint_0[9:9], gfint_1[9:9], gfint_2[9:9]);
  NOR2 I28 (simp311_0[1:1], gfint_3[9:9], gfint_4[9:9]);
  NAND2 I29 (o_0r0[9:9], simp311_0[0:0], simp311_0[1:1]);
  NOR3 I30 (simp321_0[0:0], gfint_0[10:10], gfint_1[10:10], gfint_2[10:10]);
  NOR2 I31 (simp321_0[1:1], gfint_3[10:10], gfint_4[10:10]);
  NAND2 I32 (o_0r0[10:10], simp321_0[0:0], simp321_0[1:1]);
  NOR3 I33 (simp331_0[0:0], gfint_0[11:11], gfint_1[11:11], gfint_2[11:11]);
  NOR2 I34 (simp331_0[1:1], gfint_3[11:11], gfint_4[11:11]);
  NAND2 I35 (o_0r0[11:11], simp331_0[0:0], simp331_0[1:1]);
  NOR3 I36 (simp341_0[0:0], gfint_0[12:12], gfint_1[12:12], gfint_2[12:12]);
  NOR2 I37 (simp341_0[1:1], gfint_3[12:12], gfint_4[12:12]);
  NAND2 I38 (o_0r0[12:12], simp341_0[0:0], simp341_0[1:1]);
  NOR3 I39 (simp351_0[0:0], gfint_0[13:13], gfint_1[13:13], gfint_2[13:13]);
  NOR2 I40 (simp351_0[1:1], gfint_3[13:13], gfint_4[13:13]);
  NAND2 I41 (o_0r0[13:13], simp351_0[0:0], simp351_0[1:1]);
  NOR3 I42 (simp361_0[0:0], gfint_0[14:14], gfint_1[14:14], gfint_2[14:14]);
  NOR2 I43 (simp361_0[1:1], gfint_3[14:14], gfint_4[14:14]);
  NAND2 I44 (o_0r0[14:14], simp361_0[0:0], simp361_0[1:1]);
  NOR3 I45 (simp371_0[0:0], gfint_0[15:15], gfint_1[15:15], gfint_2[15:15]);
  NOR2 I46 (simp371_0[1:1], gfint_3[15:15], gfint_4[15:15]);
  NAND2 I47 (o_0r0[15:15], simp371_0[0:0], simp371_0[1:1]);
  NOR3 I48 (simp381_0[0:0], gfint_0[16:16], gfint_1[16:16], gfint_2[16:16]);
  NOR2 I49 (simp381_0[1:1], gfint_3[16:16], gfint_4[16:16]);
  NAND2 I50 (o_0r0[16:16], simp381_0[0:0], simp381_0[1:1]);
  NOR3 I51 (simp391_0[0:0], gfint_0[17:17], gfint_1[17:17], gfint_2[17:17]);
  NOR2 I52 (simp391_0[1:1], gfint_3[17:17], gfint_4[17:17]);
  NAND2 I53 (o_0r0[17:17], simp391_0[0:0], simp391_0[1:1]);
  NOR3 I54 (simp401_0[0:0], gfint_0[18:18], gfint_1[18:18], gfint_2[18:18]);
  NOR2 I55 (simp401_0[1:1], gfint_3[18:18], gfint_4[18:18]);
  NAND2 I56 (o_0r0[18:18], simp401_0[0:0], simp401_0[1:1]);
  NOR3 I57 (simp411_0[0:0], gfint_0[19:19], gfint_1[19:19], gfint_2[19:19]);
  NOR2 I58 (simp411_0[1:1], gfint_3[19:19], gfint_4[19:19]);
  NAND2 I59 (o_0r0[19:19], simp411_0[0:0], simp411_0[1:1]);
  NOR3 I60 (simp421_0[0:0], gfint_0[20:20], gfint_1[20:20], gfint_2[20:20]);
  NOR2 I61 (simp421_0[1:1], gfint_3[20:20], gfint_4[20:20]);
  NAND2 I62 (o_0r0[20:20], simp421_0[0:0], simp421_0[1:1]);
  NOR3 I63 (simp431_0[0:0], gfint_0[21:21], gfint_1[21:21], gfint_2[21:21]);
  NOR2 I64 (simp431_0[1:1], gfint_3[21:21], gfint_4[21:21]);
  NAND2 I65 (o_0r0[21:21], simp431_0[0:0], simp431_0[1:1]);
  NOR3 I66 (simp441_0[0:0], gfint_0[22:22], gfint_1[22:22], gfint_2[22:22]);
  NOR2 I67 (simp441_0[1:1], gfint_3[22:22], gfint_4[22:22]);
  NAND2 I68 (o_0r0[22:22], simp441_0[0:0], simp441_0[1:1]);
  NOR3 I69 (simp451_0[0:0], gfint_0[23:23], gfint_1[23:23], gfint_2[23:23]);
  NOR2 I70 (simp451_0[1:1], gfint_3[23:23], gfint_4[23:23]);
  NAND2 I71 (o_0r0[23:23], simp451_0[0:0], simp451_0[1:1]);
  NOR3 I72 (simp461_0[0:0], gfint_0[24:24], gfint_1[24:24], gfint_2[24:24]);
  NOR2 I73 (simp461_0[1:1], gfint_3[24:24], gfint_4[24:24]);
  NAND2 I74 (o_0r0[24:24], simp461_0[0:0], simp461_0[1:1]);
  NOR3 I75 (simp471_0[0:0], gfint_0[25:25], gfint_1[25:25], gfint_2[25:25]);
  NOR2 I76 (simp471_0[1:1], gfint_3[25:25], gfint_4[25:25]);
  NAND2 I77 (o_0r0[25:25], simp471_0[0:0], simp471_0[1:1]);
  NOR3 I78 (simp481_0[0:0], gfint_0[26:26], gfint_1[26:26], gfint_2[26:26]);
  NOR2 I79 (simp481_0[1:1], gfint_3[26:26], gfint_4[26:26]);
  NAND2 I80 (o_0r0[26:26], simp481_0[0:0], simp481_0[1:1]);
  NOR3 I81 (simp491_0[0:0], gfint_0[27:27], gfint_1[27:27], gfint_2[27:27]);
  NOR2 I82 (simp491_0[1:1], gfint_3[27:27], gfint_4[27:27]);
  NAND2 I83 (o_0r0[27:27], simp491_0[0:0], simp491_0[1:1]);
  NOR3 I84 (simp501_0[0:0], gfint_0[28:28], gfint_1[28:28], gfint_2[28:28]);
  NOR2 I85 (simp501_0[1:1], gfint_3[28:28], gfint_4[28:28]);
  NAND2 I86 (o_0r0[28:28], simp501_0[0:0], simp501_0[1:1]);
  NOR3 I87 (simp511_0[0:0], gfint_0[29:29], gfint_1[29:29], gfint_2[29:29]);
  NOR2 I88 (simp511_0[1:1], gfint_3[29:29], gfint_4[29:29]);
  NAND2 I89 (o_0r0[29:29], simp511_0[0:0], simp511_0[1:1]);
  NOR3 I90 (simp521_0[0:0], gfint_0[30:30], gfint_1[30:30], gfint_2[30:30]);
  NOR2 I91 (simp521_0[1:1], gfint_3[30:30], gfint_4[30:30]);
  NAND2 I92 (o_0r0[30:30], simp521_0[0:0], simp521_0[1:1]);
  NOR3 I93 (simp531_0[0:0], gfint_0[31:31], gfint_1[31:31], gfint_2[31:31]);
  NOR2 I94 (simp531_0[1:1], gfint_3[31:31], gfint_4[31:31]);
  NAND2 I95 (o_0r0[31:31], simp531_0[0:0], simp531_0[1:1]);
  NOR3 I96 (simp541_0[0:0], gfint_0[32:32], gfint_1[32:32], gfint_2[32:32]);
  NOR2 I97 (simp541_0[1:1], gfint_3[32:32], gfint_4[32:32]);
  NAND2 I98 (o_0r0[32:32], simp541_0[0:0], simp541_0[1:1]);
  NOR3 I99 (simp551_0[0:0], gfint_0[33:33], gfint_1[33:33], gfint_2[33:33]);
  NOR2 I100 (simp551_0[1:1], gfint_3[33:33], gfint_4[33:33]);
  NAND2 I101 (o_0r0[33:33], simp551_0[0:0], simp551_0[1:1]);
  NOR3 I102 (simp561_0[0:0], gfint_0[34:34], gfint_1[34:34], gfint_2[34:34]);
  NOR2 I103 (simp561_0[1:1], gfint_3[34:34], gfint_4[34:34]);
  NAND2 I104 (o_0r0[34:34], simp561_0[0:0], simp561_0[1:1]);
  NOR3 I105 (simp571_0[0:0], gfint_0[35:35], gfint_1[35:35], gfint_2[35:35]);
  NOR2 I106 (simp571_0[1:1], gfint_3[35:35], gfint_4[35:35]);
  NAND2 I107 (o_0r0[35:35], simp571_0[0:0], simp571_0[1:1]);
  NOR3 I108 (simp581_0[0:0], gfint_0[36:36], gfint_1[36:36], gfint_2[36:36]);
  NOR2 I109 (simp581_0[1:1], gfint_3[36:36], gfint_4[36:36]);
  NAND2 I110 (o_0r0[36:36], simp581_0[0:0], simp581_0[1:1]);
  NOR3 I111 (simp591_0[0:0], gfint_0[37:37], gfint_1[37:37], gfint_2[37:37]);
  NOR2 I112 (simp591_0[1:1], gfint_3[37:37], gfint_4[37:37]);
  NAND2 I113 (o_0r0[37:37], simp591_0[0:0], simp591_0[1:1]);
  NOR3 I114 (simp601_0[0:0], gfint_0[38:38], gfint_1[38:38], gfint_2[38:38]);
  NOR2 I115 (simp601_0[1:1], gfint_3[38:38], gfint_4[38:38]);
  NAND2 I116 (o_0r0[38:38], simp601_0[0:0], simp601_0[1:1]);
  NOR3 I117 (simp611_0[0:0], gfint_0[39:39], gfint_1[39:39], gfint_2[39:39]);
  NOR2 I118 (simp611_0[1:1], gfint_3[39:39], gfint_4[39:39]);
  NAND2 I119 (o_0r0[39:39], simp611_0[0:0], simp611_0[1:1]);
  NOR3 I120 (simp621_0[0:0], gfint_0[40:40], gfint_1[40:40], gfint_2[40:40]);
  NOR2 I121 (simp621_0[1:1], gfint_3[40:40], gfint_4[40:40]);
  NAND2 I122 (o_0r0[40:40], simp621_0[0:0], simp621_0[1:1]);
  NOR3 I123 (simp631_0[0:0], gfint_0[41:41], gfint_1[41:41], gfint_2[41:41]);
  NOR2 I124 (simp631_0[1:1], gfint_3[41:41], gfint_4[41:41]);
  NAND2 I125 (o_0r0[41:41], simp631_0[0:0], simp631_0[1:1]);
  NOR3 I126 (simp641_0[0:0], gfint_0[42:42], gfint_1[42:42], gfint_2[42:42]);
  NOR2 I127 (simp641_0[1:1], gfint_3[42:42], gfint_4[42:42]);
  NAND2 I128 (o_0r0[42:42], simp641_0[0:0], simp641_0[1:1]);
  NOR3 I129 (simp651_0[0:0], gfint_0[43:43], gfint_1[43:43], gfint_2[43:43]);
  NOR2 I130 (simp651_0[1:1], gfint_3[43:43], gfint_4[43:43]);
  NAND2 I131 (o_0r0[43:43], simp651_0[0:0], simp651_0[1:1]);
  NOR3 I132 (simp661_0[0:0], gfint_0[44:44], gfint_1[44:44], gfint_2[44:44]);
  NOR2 I133 (simp661_0[1:1], gfint_3[44:44], gfint_4[44:44]);
  NAND2 I134 (o_0r0[44:44], simp661_0[0:0], simp661_0[1:1]);
  NOR3 I135 (simp671_0[0:0], gfint_0[45:45], gfint_1[45:45], gfint_2[45:45]);
  NOR2 I136 (simp671_0[1:1], gfint_3[45:45], gfint_4[45:45]);
  NAND2 I137 (o_0r0[45:45], simp671_0[0:0], simp671_0[1:1]);
  NOR3 I138 (simp681_0[0:0], gfint_0[46:46], gfint_1[46:46], gfint_2[46:46]);
  NOR2 I139 (simp681_0[1:1], gfint_3[46:46], gfint_4[46:46]);
  NAND2 I140 (o_0r0[46:46], simp681_0[0:0], simp681_0[1:1]);
  NOR3 I141 (simp691_0[0:0], gfint_0[47:47], gfint_1[47:47], gfint_2[47:47]);
  NOR2 I142 (simp691_0[1:1], gfint_3[47:47], gfint_4[47:47]);
  NAND2 I143 (o_0r0[47:47], simp691_0[0:0], simp691_0[1:1]);
  NOR3 I144 (simp701_0[0:0], gfint_0[48:48], gfint_1[48:48], gfint_2[48:48]);
  NOR2 I145 (simp701_0[1:1], gfint_3[48:48], gfint_4[48:48]);
  NAND2 I146 (o_0r0[48:48], simp701_0[0:0], simp701_0[1:1]);
  NOR3 I147 (simp711_0[0:0], gfint_0[49:49], gfint_1[49:49], gfint_2[49:49]);
  NOR2 I148 (simp711_0[1:1], gfint_3[49:49], gfint_4[49:49]);
  NAND2 I149 (o_0r0[49:49], simp711_0[0:0], simp711_0[1:1]);
  NOR3 I150 (simp721_0[0:0], gfint_0[50:50], gfint_1[50:50], gfint_2[50:50]);
  NOR2 I151 (simp721_0[1:1], gfint_3[50:50], gfint_4[50:50]);
  NAND2 I152 (o_0r0[50:50], simp721_0[0:0], simp721_0[1:1]);
  NOR3 I153 (simp731_0[0:0], gfint_0[51:51], gfint_1[51:51], gfint_2[51:51]);
  NOR2 I154 (simp731_0[1:1], gfint_3[51:51], gfint_4[51:51]);
  NAND2 I155 (o_0r0[51:51], simp731_0[0:0], simp731_0[1:1]);
  NOR3 I156 (simp741_0[0:0], gfint_0[52:52], gfint_1[52:52], gfint_2[52:52]);
  NOR2 I157 (simp741_0[1:1], gfint_3[52:52], gfint_4[52:52]);
  NAND2 I158 (o_0r0[52:52], simp741_0[0:0], simp741_0[1:1]);
  NOR3 I159 (simp751_0[0:0], gfint_0[53:53], gfint_1[53:53], gfint_2[53:53]);
  NOR2 I160 (simp751_0[1:1], gfint_3[53:53], gfint_4[53:53]);
  NAND2 I161 (o_0r0[53:53], simp751_0[0:0], simp751_0[1:1]);
  NOR3 I162 (simp761_0[0:0], gfint_0[54:54], gfint_1[54:54], gfint_2[54:54]);
  NOR2 I163 (simp761_0[1:1], gfint_3[54:54], gfint_4[54:54]);
  NAND2 I164 (o_0r0[54:54], simp761_0[0:0], simp761_0[1:1]);
  NOR3 I165 (simp771_0[0:0], gfint_0[55:55], gfint_1[55:55], gfint_2[55:55]);
  NOR2 I166 (simp771_0[1:1], gfint_3[55:55], gfint_4[55:55]);
  NAND2 I167 (o_0r0[55:55], simp771_0[0:0], simp771_0[1:1]);
  NOR3 I168 (simp781_0[0:0], gfint_0[56:56], gfint_1[56:56], gfint_2[56:56]);
  NOR2 I169 (simp781_0[1:1], gfint_3[56:56], gfint_4[56:56]);
  NAND2 I170 (o_0r0[56:56], simp781_0[0:0], simp781_0[1:1]);
  NOR3 I171 (simp791_0[0:0], gfint_0[57:57], gfint_1[57:57], gfint_2[57:57]);
  NOR2 I172 (simp791_0[1:1], gfint_3[57:57], gfint_4[57:57]);
  NAND2 I173 (o_0r0[57:57], simp791_0[0:0], simp791_0[1:1]);
  NOR3 I174 (simp801_0[0:0], gfint_0[58:58], gfint_1[58:58], gfint_2[58:58]);
  NOR2 I175 (simp801_0[1:1], gfint_3[58:58], gfint_4[58:58]);
  NAND2 I176 (o_0r0[58:58], simp801_0[0:0], simp801_0[1:1]);
  NOR3 I177 (simp811_0[0:0], gfint_0[59:59], gfint_1[59:59], gfint_2[59:59]);
  NOR2 I178 (simp811_0[1:1], gfint_3[59:59], gfint_4[59:59]);
  NAND2 I179 (o_0r0[59:59], simp811_0[0:0], simp811_0[1:1]);
  NOR3 I180 (simp821_0[0:0], gfint_0[60:60], gfint_1[60:60], gfint_2[60:60]);
  NOR2 I181 (simp821_0[1:1], gfint_3[60:60], gfint_4[60:60]);
  NAND2 I182 (o_0r0[60:60], simp821_0[0:0], simp821_0[1:1]);
  NOR3 I183 (simp831_0[0:0], gfint_0[61:61], gfint_1[61:61], gfint_2[61:61]);
  NOR2 I184 (simp831_0[1:1], gfint_3[61:61], gfint_4[61:61]);
  NAND2 I185 (o_0r0[61:61], simp831_0[0:0], simp831_0[1:1]);
  NOR3 I186 (simp841_0[0:0], gfint_0[62:62], gfint_1[62:62], gfint_2[62:62]);
  NOR2 I187 (simp841_0[1:1], gfint_3[62:62], gfint_4[62:62]);
  NAND2 I188 (o_0r0[62:62], simp841_0[0:0], simp841_0[1:1]);
  NOR3 I189 (simp851_0[0:0], gfint_0[63:63], gfint_1[63:63], gfint_2[63:63]);
  NOR2 I190 (simp851_0[1:1], gfint_3[63:63], gfint_4[63:63]);
  NAND2 I191 (o_0r0[63:63], simp851_0[0:0], simp851_0[1:1]);
  NOR3 I192 (simp861_0[0:0], gfint_0[64:64], gfint_1[64:64], gfint_2[64:64]);
  NOR2 I193 (simp861_0[1:1], gfint_3[64:64], gfint_4[64:64]);
  NAND2 I194 (o_0r0[64:64], simp861_0[0:0], simp861_0[1:1]);
  NOR3 I195 (simp871_0[0:0], gfint_0[65:65], gfint_1[65:65], gfint_2[65:65]);
  NOR2 I196 (simp871_0[1:1], gfint_3[65:65], gfint_4[65:65]);
  NAND2 I197 (o_0r0[65:65], simp871_0[0:0], simp871_0[1:1]);
  NOR3 I198 (simp881_0[0:0], gfint_0[66:66], gfint_1[66:66], gfint_2[66:66]);
  NOR2 I199 (simp881_0[1:1], gfint_3[66:66], gfint_4[66:66]);
  NAND2 I200 (o_0r0[66:66], simp881_0[0:0], simp881_0[1:1]);
  NOR3 I201 (simp891_0[0:0], gfint_0[67:67], gfint_1[67:67], gfint_2[67:67]);
  NOR2 I202 (simp891_0[1:1], gfint_3[67:67], gfint_4[67:67]);
  NAND2 I203 (o_0r0[67:67], simp891_0[0:0], simp891_0[1:1]);
  NOR3 I204 (simp901_0[0:0], gfint_0[68:68], gfint_1[68:68], gfint_2[68:68]);
  NOR2 I205 (simp901_0[1:1], gfint_3[68:68], gfint_4[68:68]);
  NAND2 I206 (o_0r0[68:68], simp901_0[0:0], simp901_0[1:1]);
  NOR3 I207 (simp911_0[0:0], gfint_0[69:69], gfint_1[69:69], gfint_2[69:69]);
  NOR2 I208 (simp911_0[1:1], gfint_3[69:69], gfint_4[69:69]);
  NAND2 I209 (o_0r0[69:69], simp911_0[0:0], simp911_0[1:1]);
  NOR3 I210 (simp921_0[0:0], gfint_0[70:70], gfint_1[70:70], gfint_2[70:70]);
  NOR2 I211 (simp921_0[1:1], gfint_3[70:70], gfint_4[70:70]);
  NAND2 I212 (o_0r0[70:70], simp921_0[0:0], simp921_0[1:1]);
  NOR3 I213 (simp931_0[0:0], gfint_0[71:71], gfint_1[71:71], gfint_2[71:71]);
  NOR2 I214 (simp931_0[1:1], gfint_3[71:71], gfint_4[71:71]);
  NAND2 I215 (o_0r0[71:71], simp931_0[0:0], simp931_0[1:1]);
  NOR3 I216 (simp941_0[0:0], gfint_0[72:72], gfint_1[72:72], gfint_2[72:72]);
  NOR2 I217 (simp941_0[1:1], gfint_3[72:72], gfint_4[72:72]);
  NAND2 I218 (o_0r0[72:72], simp941_0[0:0], simp941_0[1:1]);
  NOR3 I219 (simp951_0[0:0], gfint_0[73:73], gfint_1[73:73], gfint_2[73:73]);
  NOR2 I220 (simp951_0[1:1], gfint_3[73:73], gfint_4[73:73]);
  NAND2 I221 (o_0r0[73:73], simp951_0[0:0], simp951_0[1:1]);
  NOR3 I222 (simp961_0[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  NOR2 I223 (simp961_0[1:1], gtint_3[0:0], gtint_4[0:0]);
  NAND2 I224 (o_0r1[0:0], simp961_0[0:0], simp961_0[1:1]);
  NOR3 I225 (simp971_0[0:0], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  NOR2 I226 (simp971_0[1:1], gtint_3[1:1], gtint_4[1:1]);
  NAND2 I227 (o_0r1[1:1], simp971_0[0:0], simp971_0[1:1]);
  NOR3 I228 (simp981_0[0:0], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  NOR2 I229 (simp981_0[1:1], gtint_3[2:2], gtint_4[2:2]);
  NAND2 I230 (o_0r1[2:2], simp981_0[0:0], simp981_0[1:1]);
  NOR3 I231 (simp991_0[0:0], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  NOR2 I232 (simp991_0[1:1], gtint_3[3:3], gtint_4[3:3]);
  NAND2 I233 (o_0r1[3:3], simp991_0[0:0], simp991_0[1:1]);
  NOR3 I234 (simp1001_0[0:0], gtint_0[4:4], gtint_1[4:4], gtint_2[4:4]);
  NOR2 I235 (simp1001_0[1:1], gtint_3[4:4], gtint_4[4:4]);
  NAND2 I236 (o_0r1[4:4], simp1001_0[0:0], simp1001_0[1:1]);
  NOR3 I237 (simp1011_0[0:0], gtint_0[5:5], gtint_1[5:5], gtint_2[5:5]);
  NOR2 I238 (simp1011_0[1:1], gtint_3[5:5], gtint_4[5:5]);
  NAND2 I239 (o_0r1[5:5], simp1011_0[0:0], simp1011_0[1:1]);
  NOR3 I240 (simp1021_0[0:0], gtint_0[6:6], gtint_1[6:6], gtint_2[6:6]);
  NOR2 I241 (simp1021_0[1:1], gtint_3[6:6], gtint_4[6:6]);
  NAND2 I242 (o_0r1[6:6], simp1021_0[0:0], simp1021_0[1:1]);
  NOR3 I243 (simp1031_0[0:0], gtint_0[7:7], gtint_1[7:7], gtint_2[7:7]);
  NOR2 I244 (simp1031_0[1:1], gtint_3[7:7], gtint_4[7:7]);
  NAND2 I245 (o_0r1[7:7], simp1031_0[0:0], simp1031_0[1:1]);
  NOR3 I246 (simp1041_0[0:0], gtint_0[8:8], gtint_1[8:8], gtint_2[8:8]);
  NOR2 I247 (simp1041_0[1:1], gtint_3[8:8], gtint_4[8:8]);
  NAND2 I248 (o_0r1[8:8], simp1041_0[0:0], simp1041_0[1:1]);
  NOR3 I249 (simp1051_0[0:0], gtint_0[9:9], gtint_1[9:9], gtint_2[9:9]);
  NOR2 I250 (simp1051_0[1:1], gtint_3[9:9], gtint_4[9:9]);
  NAND2 I251 (o_0r1[9:9], simp1051_0[0:0], simp1051_0[1:1]);
  NOR3 I252 (simp1061_0[0:0], gtint_0[10:10], gtint_1[10:10], gtint_2[10:10]);
  NOR2 I253 (simp1061_0[1:1], gtint_3[10:10], gtint_4[10:10]);
  NAND2 I254 (o_0r1[10:10], simp1061_0[0:0], simp1061_0[1:1]);
  NOR3 I255 (simp1071_0[0:0], gtint_0[11:11], gtint_1[11:11], gtint_2[11:11]);
  NOR2 I256 (simp1071_0[1:1], gtint_3[11:11], gtint_4[11:11]);
  NAND2 I257 (o_0r1[11:11], simp1071_0[0:0], simp1071_0[1:1]);
  NOR3 I258 (simp1081_0[0:0], gtint_0[12:12], gtint_1[12:12], gtint_2[12:12]);
  NOR2 I259 (simp1081_0[1:1], gtint_3[12:12], gtint_4[12:12]);
  NAND2 I260 (o_0r1[12:12], simp1081_0[0:0], simp1081_0[1:1]);
  NOR3 I261 (simp1091_0[0:0], gtint_0[13:13], gtint_1[13:13], gtint_2[13:13]);
  NOR2 I262 (simp1091_0[1:1], gtint_3[13:13], gtint_4[13:13]);
  NAND2 I263 (o_0r1[13:13], simp1091_0[0:0], simp1091_0[1:1]);
  NOR3 I264 (simp1101_0[0:0], gtint_0[14:14], gtint_1[14:14], gtint_2[14:14]);
  NOR2 I265 (simp1101_0[1:1], gtint_3[14:14], gtint_4[14:14]);
  NAND2 I266 (o_0r1[14:14], simp1101_0[0:0], simp1101_0[1:1]);
  NOR3 I267 (simp1111_0[0:0], gtint_0[15:15], gtint_1[15:15], gtint_2[15:15]);
  NOR2 I268 (simp1111_0[1:1], gtint_3[15:15], gtint_4[15:15]);
  NAND2 I269 (o_0r1[15:15], simp1111_0[0:0], simp1111_0[1:1]);
  NOR3 I270 (simp1121_0[0:0], gtint_0[16:16], gtint_1[16:16], gtint_2[16:16]);
  NOR2 I271 (simp1121_0[1:1], gtint_3[16:16], gtint_4[16:16]);
  NAND2 I272 (o_0r1[16:16], simp1121_0[0:0], simp1121_0[1:1]);
  NOR3 I273 (simp1131_0[0:0], gtint_0[17:17], gtint_1[17:17], gtint_2[17:17]);
  NOR2 I274 (simp1131_0[1:1], gtint_3[17:17], gtint_4[17:17]);
  NAND2 I275 (o_0r1[17:17], simp1131_0[0:0], simp1131_0[1:1]);
  NOR3 I276 (simp1141_0[0:0], gtint_0[18:18], gtint_1[18:18], gtint_2[18:18]);
  NOR2 I277 (simp1141_0[1:1], gtint_3[18:18], gtint_4[18:18]);
  NAND2 I278 (o_0r1[18:18], simp1141_0[0:0], simp1141_0[1:1]);
  NOR3 I279 (simp1151_0[0:0], gtint_0[19:19], gtint_1[19:19], gtint_2[19:19]);
  NOR2 I280 (simp1151_0[1:1], gtint_3[19:19], gtint_4[19:19]);
  NAND2 I281 (o_0r1[19:19], simp1151_0[0:0], simp1151_0[1:1]);
  NOR3 I282 (simp1161_0[0:0], gtint_0[20:20], gtint_1[20:20], gtint_2[20:20]);
  NOR2 I283 (simp1161_0[1:1], gtint_3[20:20], gtint_4[20:20]);
  NAND2 I284 (o_0r1[20:20], simp1161_0[0:0], simp1161_0[1:1]);
  NOR3 I285 (simp1171_0[0:0], gtint_0[21:21], gtint_1[21:21], gtint_2[21:21]);
  NOR2 I286 (simp1171_0[1:1], gtint_3[21:21], gtint_4[21:21]);
  NAND2 I287 (o_0r1[21:21], simp1171_0[0:0], simp1171_0[1:1]);
  NOR3 I288 (simp1181_0[0:0], gtint_0[22:22], gtint_1[22:22], gtint_2[22:22]);
  NOR2 I289 (simp1181_0[1:1], gtint_3[22:22], gtint_4[22:22]);
  NAND2 I290 (o_0r1[22:22], simp1181_0[0:0], simp1181_0[1:1]);
  NOR3 I291 (simp1191_0[0:0], gtint_0[23:23], gtint_1[23:23], gtint_2[23:23]);
  NOR2 I292 (simp1191_0[1:1], gtint_3[23:23], gtint_4[23:23]);
  NAND2 I293 (o_0r1[23:23], simp1191_0[0:0], simp1191_0[1:1]);
  NOR3 I294 (simp1201_0[0:0], gtint_0[24:24], gtint_1[24:24], gtint_2[24:24]);
  NOR2 I295 (simp1201_0[1:1], gtint_3[24:24], gtint_4[24:24]);
  NAND2 I296 (o_0r1[24:24], simp1201_0[0:0], simp1201_0[1:1]);
  NOR3 I297 (simp1211_0[0:0], gtint_0[25:25], gtint_1[25:25], gtint_2[25:25]);
  NOR2 I298 (simp1211_0[1:1], gtint_3[25:25], gtint_4[25:25]);
  NAND2 I299 (o_0r1[25:25], simp1211_0[0:0], simp1211_0[1:1]);
  NOR3 I300 (simp1221_0[0:0], gtint_0[26:26], gtint_1[26:26], gtint_2[26:26]);
  NOR2 I301 (simp1221_0[1:1], gtint_3[26:26], gtint_4[26:26]);
  NAND2 I302 (o_0r1[26:26], simp1221_0[0:0], simp1221_0[1:1]);
  NOR3 I303 (simp1231_0[0:0], gtint_0[27:27], gtint_1[27:27], gtint_2[27:27]);
  NOR2 I304 (simp1231_0[1:1], gtint_3[27:27], gtint_4[27:27]);
  NAND2 I305 (o_0r1[27:27], simp1231_0[0:0], simp1231_0[1:1]);
  NOR3 I306 (simp1241_0[0:0], gtint_0[28:28], gtint_1[28:28], gtint_2[28:28]);
  NOR2 I307 (simp1241_0[1:1], gtint_3[28:28], gtint_4[28:28]);
  NAND2 I308 (o_0r1[28:28], simp1241_0[0:0], simp1241_0[1:1]);
  NOR3 I309 (simp1251_0[0:0], gtint_0[29:29], gtint_1[29:29], gtint_2[29:29]);
  NOR2 I310 (simp1251_0[1:1], gtint_3[29:29], gtint_4[29:29]);
  NAND2 I311 (o_0r1[29:29], simp1251_0[0:0], simp1251_0[1:1]);
  NOR3 I312 (simp1261_0[0:0], gtint_0[30:30], gtint_1[30:30], gtint_2[30:30]);
  NOR2 I313 (simp1261_0[1:1], gtint_3[30:30], gtint_4[30:30]);
  NAND2 I314 (o_0r1[30:30], simp1261_0[0:0], simp1261_0[1:1]);
  NOR3 I315 (simp1271_0[0:0], gtint_0[31:31], gtint_1[31:31], gtint_2[31:31]);
  NOR2 I316 (simp1271_0[1:1], gtint_3[31:31], gtint_4[31:31]);
  NAND2 I317 (o_0r1[31:31], simp1271_0[0:0], simp1271_0[1:1]);
  NOR3 I318 (simp1281_0[0:0], gtint_0[32:32], gtint_1[32:32], gtint_2[32:32]);
  NOR2 I319 (simp1281_0[1:1], gtint_3[32:32], gtint_4[32:32]);
  NAND2 I320 (o_0r1[32:32], simp1281_0[0:0], simp1281_0[1:1]);
  NOR3 I321 (simp1291_0[0:0], gtint_0[33:33], gtint_1[33:33], gtint_2[33:33]);
  NOR2 I322 (simp1291_0[1:1], gtint_3[33:33], gtint_4[33:33]);
  NAND2 I323 (o_0r1[33:33], simp1291_0[0:0], simp1291_0[1:1]);
  NOR3 I324 (simp1301_0[0:0], gtint_0[34:34], gtint_1[34:34], gtint_2[34:34]);
  NOR2 I325 (simp1301_0[1:1], gtint_3[34:34], gtint_4[34:34]);
  NAND2 I326 (o_0r1[34:34], simp1301_0[0:0], simp1301_0[1:1]);
  NOR3 I327 (simp1311_0[0:0], gtint_0[35:35], gtint_1[35:35], gtint_2[35:35]);
  NOR2 I328 (simp1311_0[1:1], gtint_3[35:35], gtint_4[35:35]);
  NAND2 I329 (o_0r1[35:35], simp1311_0[0:0], simp1311_0[1:1]);
  NOR3 I330 (simp1321_0[0:0], gtint_0[36:36], gtint_1[36:36], gtint_2[36:36]);
  NOR2 I331 (simp1321_0[1:1], gtint_3[36:36], gtint_4[36:36]);
  NAND2 I332 (o_0r1[36:36], simp1321_0[0:0], simp1321_0[1:1]);
  NOR3 I333 (simp1331_0[0:0], gtint_0[37:37], gtint_1[37:37], gtint_2[37:37]);
  NOR2 I334 (simp1331_0[1:1], gtint_3[37:37], gtint_4[37:37]);
  NAND2 I335 (o_0r1[37:37], simp1331_0[0:0], simp1331_0[1:1]);
  NOR3 I336 (simp1341_0[0:0], gtint_0[38:38], gtint_1[38:38], gtint_2[38:38]);
  NOR2 I337 (simp1341_0[1:1], gtint_3[38:38], gtint_4[38:38]);
  NAND2 I338 (o_0r1[38:38], simp1341_0[0:0], simp1341_0[1:1]);
  NOR3 I339 (simp1351_0[0:0], gtint_0[39:39], gtint_1[39:39], gtint_2[39:39]);
  NOR2 I340 (simp1351_0[1:1], gtint_3[39:39], gtint_4[39:39]);
  NAND2 I341 (o_0r1[39:39], simp1351_0[0:0], simp1351_0[1:1]);
  NOR3 I342 (simp1361_0[0:0], gtint_0[40:40], gtint_1[40:40], gtint_2[40:40]);
  NOR2 I343 (simp1361_0[1:1], gtint_3[40:40], gtint_4[40:40]);
  NAND2 I344 (o_0r1[40:40], simp1361_0[0:0], simp1361_0[1:1]);
  NOR3 I345 (simp1371_0[0:0], gtint_0[41:41], gtint_1[41:41], gtint_2[41:41]);
  NOR2 I346 (simp1371_0[1:1], gtint_3[41:41], gtint_4[41:41]);
  NAND2 I347 (o_0r1[41:41], simp1371_0[0:0], simp1371_0[1:1]);
  NOR3 I348 (simp1381_0[0:0], gtint_0[42:42], gtint_1[42:42], gtint_2[42:42]);
  NOR2 I349 (simp1381_0[1:1], gtint_3[42:42], gtint_4[42:42]);
  NAND2 I350 (o_0r1[42:42], simp1381_0[0:0], simp1381_0[1:1]);
  NOR3 I351 (simp1391_0[0:0], gtint_0[43:43], gtint_1[43:43], gtint_2[43:43]);
  NOR2 I352 (simp1391_0[1:1], gtint_3[43:43], gtint_4[43:43]);
  NAND2 I353 (o_0r1[43:43], simp1391_0[0:0], simp1391_0[1:1]);
  NOR3 I354 (simp1401_0[0:0], gtint_0[44:44], gtint_1[44:44], gtint_2[44:44]);
  NOR2 I355 (simp1401_0[1:1], gtint_3[44:44], gtint_4[44:44]);
  NAND2 I356 (o_0r1[44:44], simp1401_0[0:0], simp1401_0[1:1]);
  NOR3 I357 (simp1411_0[0:0], gtint_0[45:45], gtint_1[45:45], gtint_2[45:45]);
  NOR2 I358 (simp1411_0[1:1], gtint_3[45:45], gtint_4[45:45]);
  NAND2 I359 (o_0r1[45:45], simp1411_0[0:0], simp1411_0[1:1]);
  NOR3 I360 (simp1421_0[0:0], gtint_0[46:46], gtint_1[46:46], gtint_2[46:46]);
  NOR2 I361 (simp1421_0[1:1], gtint_3[46:46], gtint_4[46:46]);
  NAND2 I362 (o_0r1[46:46], simp1421_0[0:0], simp1421_0[1:1]);
  NOR3 I363 (simp1431_0[0:0], gtint_0[47:47], gtint_1[47:47], gtint_2[47:47]);
  NOR2 I364 (simp1431_0[1:1], gtint_3[47:47], gtint_4[47:47]);
  NAND2 I365 (o_0r1[47:47], simp1431_0[0:0], simp1431_0[1:1]);
  NOR3 I366 (simp1441_0[0:0], gtint_0[48:48], gtint_1[48:48], gtint_2[48:48]);
  NOR2 I367 (simp1441_0[1:1], gtint_3[48:48], gtint_4[48:48]);
  NAND2 I368 (o_0r1[48:48], simp1441_0[0:0], simp1441_0[1:1]);
  NOR3 I369 (simp1451_0[0:0], gtint_0[49:49], gtint_1[49:49], gtint_2[49:49]);
  NOR2 I370 (simp1451_0[1:1], gtint_3[49:49], gtint_4[49:49]);
  NAND2 I371 (o_0r1[49:49], simp1451_0[0:0], simp1451_0[1:1]);
  NOR3 I372 (simp1461_0[0:0], gtint_0[50:50], gtint_1[50:50], gtint_2[50:50]);
  NOR2 I373 (simp1461_0[1:1], gtint_3[50:50], gtint_4[50:50]);
  NAND2 I374 (o_0r1[50:50], simp1461_0[0:0], simp1461_0[1:1]);
  NOR3 I375 (simp1471_0[0:0], gtint_0[51:51], gtint_1[51:51], gtint_2[51:51]);
  NOR2 I376 (simp1471_0[1:1], gtint_3[51:51], gtint_4[51:51]);
  NAND2 I377 (o_0r1[51:51], simp1471_0[0:0], simp1471_0[1:1]);
  NOR3 I378 (simp1481_0[0:0], gtint_0[52:52], gtint_1[52:52], gtint_2[52:52]);
  NOR2 I379 (simp1481_0[1:1], gtint_3[52:52], gtint_4[52:52]);
  NAND2 I380 (o_0r1[52:52], simp1481_0[0:0], simp1481_0[1:1]);
  NOR3 I381 (simp1491_0[0:0], gtint_0[53:53], gtint_1[53:53], gtint_2[53:53]);
  NOR2 I382 (simp1491_0[1:1], gtint_3[53:53], gtint_4[53:53]);
  NAND2 I383 (o_0r1[53:53], simp1491_0[0:0], simp1491_0[1:1]);
  NOR3 I384 (simp1501_0[0:0], gtint_0[54:54], gtint_1[54:54], gtint_2[54:54]);
  NOR2 I385 (simp1501_0[1:1], gtint_3[54:54], gtint_4[54:54]);
  NAND2 I386 (o_0r1[54:54], simp1501_0[0:0], simp1501_0[1:1]);
  NOR3 I387 (simp1511_0[0:0], gtint_0[55:55], gtint_1[55:55], gtint_2[55:55]);
  NOR2 I388 (simp1511_0[1:1], gtint_3[55:55], gtint_4[55:55]);
  NAND2 I389 (o_0r1[55:55], simp1511_0[0:0], simp1511_0[1:1]);
  NOR3 I390 (simp1521_0[0:0], gtint_0[56:56], gtint_1[56:56], gtint_2[56:56]);
  NOR2 I391 (simp1521_0[1:1], gtint_3[56:56], gtint_4[56:56]);
  NAND2 I392 (o_0r1[56:56], simp1521_0[0:0], simp1521_0[1:1]);
  NOR3 I393 (simp1531_0[0:0], gtint_0[57:57], gtint_1[57:57], gtint_2[57:57]);
  NOR2 I394 (simp1531_0[1:1], gtint_3[57:57], gtint_4[57:57]);
  NAND2 I395 (o_0r1[57:57], simp1531_0[0:0], simp1531_0[1:1]);
  NOR3 I396 (simp1541_0[0:0], gtint_0[58:58], gtint_1[58:58], gtint_2[58:58]);
  NOR2 I397 (simp1541_0[1:1], gtint_3[58:58], gtint_4[58:58]);
  NAND2 I398 (o_0r1[58:58], simp1541_0[0:0], simp1541_0[1:1]);
  NOR3 I399 (simp1551_0[0:0], gtint_0[59:59], gtint_1[59:59], gtint_2[59:59]);
  NOR2 I400 (simp1551_0[1:1], gtint_3[59:59], gtint_4[59:59]);
  NAND2 I401 (o_0r1[59:59], simp1551_0[0:0], simp1551_0[1:1]);
  NOR3 I402 (simp1561_0[0:0], gtint_0[60:60], gtint_1[60:60], gtint_2[60:60]);
  NOR2 I403 (simp1561_0[1:1], gtint_3[60:60], gtint_4[60:60]);
  NAND2 I404 (o_0r1[60:60], simp1561_0[0:0], simp1561_0[1:1]);
  NOR3 I405 (simp1571_0[0:0], gtint_0[61:61], gtint_1[61:61], gtint_2[61:61]);
  NOR2 I406 (simp1571_0[1:1], gtint_3[61:61], gtint_4[61:61]);
  NAND2 I407 (o_0r1[61:61], simp1571_0[0:0], simp1571_0[1:1]);
  NOR3 I408 (simp1581_0[0:0], gtint_0[62:62], gtint_1[62:62], gtint_2[62:62]);
  NOR2 I409 (simp1581_0[1:1], gtint_3[62:62], gtint_4[62:62]);
  NAND2 I410 (o_0r1[62:62], simp1581_0[0:0], simp1581_0[1:1]);
  NOR3 I411 (simp1591_0[0:0], gtint_0[63:63], gtint_1[63:63], gtint_2[63:63]);
  NOR2 I412 (simp1591_0[1:1], gtint_3[63:63], gtint_4[63:63]);
  NAND2 I413 (o_0r1[63:63], simp1591_0[0:0], simp1591_0[1:1]);
  NOR3 I414 (simp1601_0[0:0], gtint_0[64:64], gtint_1[64:64], gtint_2[64:64]);
  NOR2 I415 (simp1601_0[1:1], gtint_3[64:64], gtint_4[64:64]);
  NAND2 I416 (o_0r1[64:64], simp1601_0[0:0], simp1601_0[1:1]);
  NOR3 I417 (simp1611_0[0:0], gtint_0[65:65], gtint_1[65:65], gtint_2[65:65]);
  NOR2 I418 (simp1611_0[1:1], gtint_3[65:65], gtint_4[65:65]);
  NAND2 I419 (o_0r1[65:65], simp1611_0[0:0], simp1611_0[1:1]);
  NOR3 I420 (simp1621_0[0:0], gtint_0[66:66], gtint_1[66:66], gtint_2[66:66]);
  NOR2 I421 (simp1621_0[1:1], gtint_3[66:66], gtint_4[66:66]);
  NAND2 I422 (o_0r1[66:66], simp1621_0[0:0], simp1621_0[1:1]);
  NOR3 I423 (simp1631_0[0:0], gtint_0[67:67], gtint_1[67:67], gtint_2[67:67]);
  NOR2 I424 (simp1631_0[1:1], gtint_3[67:67], gtint_4[67:67]);
  NAND2 I425 (o_0r1[67:67], simp1631_0[0:0], simp1631_0[1:1]);
  NOR3 I426 (simp1641_0[0:0], gtint_0[68:68], gtint_1[68:68], gtint_2[68:68]);
  NOR2 I427 (simp1641_0[1:1], gtint_3[68:68], gtint_4[68:68]);
  NAND2 I428 (o_0r1[68:68], simp1641_0[0:0], simp1641_0[1:1]);
  NOR3 I429 (simp1651_0[0:0], gtint_0[69:69], gtint_1[69:69], gtint_2[69:69]);
  NOR2 I430 (simp1651_0[1:1], gtint_3[69:69], gtint_4[69:69]);
  NAND2 I431 (o_0r1[69:69], simp1651_0[0:0], simp1651_0[1:1]);
  NOR3 I432 (simp1661_0[0:0], gtint_0[70:70], gtint_1[70:70], gtint_2[70:70]);
  NOR2 I433 (simp1661_0[1:1], gtint_3[70:70], gtint_4[70:70]);
  NAND2 I434 (o_0r1[70:70], simp1661_0[0:0], simp1661_0[1:1]);
  NOR3 I435 (simp1671_0[0:0], gtint_0[71:71], gtint_1[71:71], gtint_2[71:71]);
  NOR2 I436 (simp1671_0[1:1], gtint_3[71:71], gtint_4[71:71]);
  NAND2 I437 (o_0r1[71:71], simp1671_0[0:0], simp1671_0[1:1]);
  NOR3 I438 (simp1681_0[0:0], gtint_0[72:72], gtint_1[72:72], gtint_2[72:72]);
  NOR2 I439 (simp1681_0[1:1], gtint_3[72:72], gtint_4[72:72]);
  NAND2 I440 (o_0r1[72:72], simp1681_0[0:0], simp1681_0[1:1]);
  NOR3 I441 (simp1691_0[0:0], gtint_0[73:73], gtint_1[73:73], gtint_2[73:73]);
  NOR2 I442 (simp1691_0[1:1], gtint_3[73:73], gtint_4[73:73]);
  NAND2 I443 (o_0r1[73:73], simp1691_0[0:0], simp1691_0[1:1]);
  AND2 I444 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I445 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I446 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I447 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I448 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I449 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I450 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I451 (gtint_0[7:7], choice_0, i_0r1[7:7]);
  AND2 I452 (gtint_0[8:8], choice_0, i_0r1[8:8]);
  AND2 I453 (gtint_0[9:9], choice_0, i_0r1[9:9]);
  AND2 I454 (gtint_0[10:10], choice_0, i_0r1[10:10]);
  AND2 I455 (gtint_0[11:11], choice_0, i_0r1[11:11]);
  AND2 I456 (gtint_0[12:12], choice_0, i_0r1[12:12]);
  AND2 I457 (gtint_0[13:13], choice_0, i_0r1[13:13]);
  AND2 I458 (gtint_0[14:14], choice_0, i_0r1[14:14]);
  AND2 I459 (gtint_0[15:15], choice_0, i_0r1[15:15]);
  AND2 I460 (gtint_0[16:16], choice_0, i_0r1[16:16]);
  AND2 I461 (gtint_0[17:17], choice_0, i_0r1[17:17]);
  AND2 I462 (gtint_0[18:18], choice_0, i_0r1[18:18]);
  AND2 I463 (gtint_0[19:19], choice_0, i_0r1[19:19]);
  AND2 I464 (gtint_0[20:20], choice_0, i_0r1[20:20]);
  AND2 I465 (gtint_0[21:21], choice_0, i_0r1[21:21]);
  AND2 I466 (gtint_0[22:22], choice_0, i_0r1[22:22]);
  AND2 I467 (gtint_0[23:23], choice_0, i_0r1[23:23]);
  AND2 I468 (gtint_0[24:24], choice_0, i_0r1[24:24]);
  AND2 I469 (gtint_0[25:25], choice_0, i_0r1[25:25]);
  AND2 I470 (gtint_0[26:26], choice_0, i_0r1[26:26]);
  AND2 I471 (gtint_0[27:27], choice_0, i_0r1[27:27]);
  AND2 I472 (gtint_0[28:28], choice_0, i_0r1[28:28]);
  AND2 I473 (gtint_0[29:29], choice_0, i_0r1[29:29]);
  AND2 I474 (gtint_0[30:30], choice_0, i_0r1[30:30]);
  AND2 I475 (gtint_0[31:31], choice_0, i_0r1[31:31]);
  AND2 I476 (gtint_0[32:32], choice_0, i_0r1[32:32]);
  AND2 I477 (gtint_0[33:33], choice_0, i_0r1[33:33]);
  AND2 I478 (gtint_0[34:34], choice_0, i_0r1[34:34]);
  AND2 I479 (gtint_0[35:35], choice_0, i_0r1[35:35]);
  AND2 I480 (gtint_0[36:36], choice_0, i_0r1[36:36]);
  AND2 I481 (gtint_0[37:37], choice_0, i_0r1[37:37]);
  AND2 I482 (gtint_0[38:38], choice_0, i_0r1[38:38]);
  AND2 I483 (gtint_0[39:39], choice_0, i_0r1[39:39]);
  AND2 I484 (gtint_0[40:40], choice_0, i_0r1[40:40]);
  AND2 I485 (gtint_0[41:41], choice_0, i_0r1[41:41]);
  AND2 I486 (gtint_0[42:42], choice_0, i_0r1[42:42]);
  AND2 I487 (gtint_0[43:43], choice_0, i_0r1[43:43]);
  AND2 I488 (gtint_0[44:44], choice_0, i_0r1[44:44]);
  AND2 I489 (gtint_0[45:45], choice_0, i_0r1[45:45]);
  AND2 I490 (gtint_0[46:46], choice_0, i_0r1[46:46]);
  AND2 I491 (gtint_0[47:47], choice_0, i_0r1[47:47]);
  AND2 I492 (gtint_0[48:48], choice_0, i_0r1[48:48]);
  AND2 I493 (gtint_0[49:49], choice_0, i_0r1[49:49]);
  AND2 I494 (gtint_0[50:50], choice_0, i_0r1[50:50]);
  AND2 I495 (gtint_0[51:51], choice_0, i_0r1[51:51]);
  AND2 I496 (gtint_0[52:52], choice_0, i_0r1[52:52]);
  AND2 I497 (gtint_0[53:53], choice_0, i_0r1[53:53]);
  AND2 I498 (gtint_0[54:54], choice_0, i_0r1[54:54]);
  AND2 I499 (gtint_0[55:55], choice_0, i_0r1[55:55]);
  AND2 I500 (gtint_0[56:56], choice_0, i_0r1[56:56]);
  AND2 I501 (gtint_0[57:57], choice_0, i_0r1[57:57]);
  AND2 I502 (gtint_0[58:58], choice_0, i_0r1[58:58]);
  AND2 I503 (gtint_0[59:59], choice_0, i_0r1[59:59]);
  AND2 I504 (gtint_0[60:60], choice_0, i_0r1[60:60]);
  AND2 I505 (gtint_0[61:61], choice_0, i_0r1[61:61]);
  AND2 I506 (gtint_0[62:62], choice_0, i_0r1[62:62]);
  AND2 I507 (gtint_0[63:63], choice_0, i_0r1[63:63]);
  AND2 I508 (gtint_0[64:64], choice_0, i_0r1[64:64]);
  AND2 I509 (gtint_0[65:65], choice_0, i_0r1[65:65]);
  AND2 I510 (gtint_0[66:66], choice_0, i_0r1[66:66]);
  AND2 I511 (gtint_0[67:67], choice_0, i_0r1[67:67]);
  AND2 I512 (gtint_0[68:68], choice_0, i_0r1[68:68]);
  AND2 I513 (gtint_0[69:69], choice_0, i_0r1[69:69]);
  AND2 I514 (gtint_0[70:70], choice_0, i_0r1[70:70]);
  AND2 I515 (gtint_0[71:71], choice_0, i_0r1[71:71]);
  AND2 I516 (gtint_0[72:72], choice_0, i_0r1[72:72]);
  AND2 I517 (gtint_0[73:73], choice_0, i_0r1[73:73]);
  AND2 I518 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I519 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I520 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I521 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I522 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I523 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I524 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I525 (gtint_1[7:7], choice_1, i_1r1[7:7]);
  AND2 I526 (gtint_1[8:8], choice_1, i_1r1[8:8]);
  AND2 I527 (gtint_1[9:9], choice_1, i_1r1[9:9]);
  AND2 I528 (gtint_1[10:10], choice_1, i_1r1[10:10]);
  AND2 I529 (gtint_1[11:11], choice_1, i_1r1[11:11]);
  AND2 I530 (gtint_1[12:12], choice_1, i_1r1[12:12]);
  AND2 I531 (gtint_1[13:13], choice_1, i_1r1[13:13]);
  AND2 I532 (gtint_1[14:14], choice_1, i_1r1[14:14]);
  AND2 I533 (gtint_1[15:15], choice_1, i_1r1[15:15]);
  AND2 I534 (gtint_1[16:16], choice_1, i_1r1[16:16]);
  AND2 I535 (gtint_1[17:17], choice_1, i_1r1[17:17]);
  AND2 I536 (gtint_1[18:18], choice_1, i_1r1[18:18]);
  AND2 I537 (gtint_1[19:19], choice_1, i_1r1[19:19]);
  AND2 I538 (gtint_1[20:20], choice_1, i_1r1[20:20]);
  AND2 I539 (gtint_1[21:21], choice_1, i_1r1[21:21]);
  AND2 I540 (gtint_1[22:22], choice_1, i_1r1[22:22]);
  AND2 I541 (gtint_1[23:23], choice_1, i_1r1[23:23]);
  AND2 I542 (gtint_1[24:24], choice_1, i_1r1[24:24]);
  AND2 I543 (gtint_1[25:25], choice_1, i_1r1[25:25]);
  AND2 I544 (gtint_1[26:26], choice_1, i_1r1[26:26]);
  AND2 I545 (gtint_1[27:27], choice_1, i_1r1[27:27]);
  AND2 I546 (gtint_1[28:28], choice_1, i_1r1[28:28]);
  AND2 I547 (gtint_1[29:29], choice_1, i_1r1[29:29]);
  AND2 I548 (gtint_1[30:30], choice_1, i_1r1[30:30]);
  AND2 I549 (gtint_1[31:31], choice_1, i_1r1[31:31]);
  AND2 I550 (gtint_1[32:32], choice_1, i_1r1[32:32]);
  AND2 I551 (gtint_1[33:33], choice_1, i_1r1[33:33]);
  AND2 I552 (gtint_1[34:34], choice_1, i_1r1[34:34]);
  AND2 I553 (gtint_1[35:35], choice_1, i_1r1[35:35]);
  AND2 I554 (gtint_1[36:36], choice_1, i_1r1[36:36]);
  AND2 I555 (gtint_1[37:37], choice_1, i_1r1[37:37]);
  AND2 I556 (gtint_1[38:38], choice_1, i_1r1[38:38]);
  AND2 I557 (gtint_1[39:39], choice_1, i_1r1[39:39]);
  AND2 I558 (gtint_1[40:40], choice_1, i_1r1[40:40]);
  AND2 I559 (gtint_1[41:41], choice_1, i_1r1[41:41]);
  AND2 I560 (gtint_1[42:42], choice_1, i_1r1[42:42]);
  AND2 I561 (gtint_1[43:43], choice_1, i_1r1[43:43]);
  AND2 I562 (gtint_1[44:44], choice_1, i_1r1[44:44]);
  AND2 I563 (gtint_1[45:45], choice_1, i_1r1[45:45]);
  AND2 I564 (gtint_1[46:46], choice_1, i_1r1[46:46]);
  AND2 I565 (gtint_1[47:47], choice_1, i_1r1[47:47]);
  AND2 I566 (gtint_1[48:48], choice_1, i_1r1[48:48]);
  AND2 I567 (gtint_1[49:49], choice_1, i_1r1[49:49]);
  AND2 I568 (gtint_1[50:50], choice_1, i_1r1[50:50]);
  AND2 I569 (gtint_1[51:51], choice_1, i_1r1[51:51]);
  AND2 I570 (gtint_1[52:52], choice_1, i_1r1[52:52]);
  AND2 I571 (gtint_1[53:53], choice_1, i_1r1[53:53]);
  AND2 I572 (gtint_1[54:54], choice_1, i_1r1[54:54]);
  AND2 I573 (gtint_1[55:55], choice_1, i_1r1[55:55]);
  AND2 I574 (gtint_1[56:56], choice_1, i_1r1[56:56]);
  AND2 I575 (gtint_1[57:57], choice_1, i_1r1[57:57]);
  AND2 I576 (gtint_1[58:58], choice_1, i_1r1[58:58]);
  AND2 I577 (gtint_1[59:59], choice_1, i_1r1[59:59]);
  AND2 I578 (gtint_1[60:60], choice_1, i_1r1[60:60]);
  AND2 I579 (gtint_1[61:61], choice_1, i_1r1[61:61]);
  AND2 I580 (gtint_1[62:62], choice_1, i_1r1[62:62]);
  AND2 I581 (gtint_1[63:63], choice_1, i_1r1[63:63]);
  AND2 I582 (gtint_1[64:64], choice_1, i_1r1[64:64]);
  AND2 I583 (gtint_1[65:65], choice_1, i_1r1[65:65]);
  AND2 I584 (gtint_1[66:66], choice_1, i_1r1[66:66]);
  AND2 I585 (gtint_1[67:67], choice_1, i_1r1[67:67]);
  AND2 I586 (gtint_1[68:68], choice_1, i_1r1[68:68]);
  AND2 I587 (gtint_1[69:69], choice_1, i_1r1[69:69]);
  AND2 I588 (gtint_1[70:70], choice_1, i_1r1[70:70]);
  AND2 I589 (gtint_1[71:71], choice_1, i_1r1[71:71]);
  AND2 I590 (gtint_1[72:72], choice_1, i_1r1[72:72]);
  AND2 I591 (gtint_1[73:73], choice_1, i_1r1[73:73]);
  AND2 I592 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I593 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I594 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I595 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AND2 I596 (gtint_2[4:4], choice_2, i_2r1[4:4]);
  AND2 I597 (gtint_2[5:5], choice_2, i_2r1[5:5]);
  AND2 I598 (gtint_2[6:6], choice_2, i_2r1[6:6]);
  AND2 I599 (gtint_2[7:7], choice_2, i_2r1[7:7]);
  AND2 I600 (gtint_2[8:8], choice_2, i_2r1[8:8]);
  AND2 I601 (gtint_2[9:9], choice_2, i_2r1[9:9]);
  AND2 I602 (gtint_2[10:10], choice_2, i_2r1[10:10]);
  AND2 I603 (gtint_2[11:11], choice_2, i_2r1[11:11]);
  AND2 I604 (gtint_2[12:12], choice_2, i_2r1[12:12]);
  AND2 I605 (gtint_2[13:13], choice_2, i_2r1[13:13]);
  AND2 I606 (gtint_2[14:14], choice_2, i_2r1[14:14]);
  AND2 I607 (gtint_2[15:15], choice_2, i_2r1[15:15]);
  AND2 I608 (gtint_2[16:16], choice_2, i_2r1[16:16]);
  AND2 I609 (gtint_2[17:17], choice_2, i_2r1[17:17]);
  AND2 I610 (gtint_2[18:18], choice_2, i_2r1[18:18]);
  AND2 I611 (gtint_2[19:19], choice_2, i_2r1[19:19]);
  AND2 I612 (gtint_2[20:20], choice_2, i_2r1[20:20]);
  AND2 I613 (gtint_2[21:21], choice_2, i_2r1[21:21]);
  AND2 I614 (gtint_2[22:22], choice_2, i_2r1[22:22]);
  AND2 I615 (gtint_2[23:23], choice_2, i_2r1[23:23]);
  AND2 I616 (gtint_2[24:24], choice_2, i_2r1[24:24]);
  AND2 I617 (gtint_2[25:25], choice_2, i_2r1[25:25]);
  AND2 I618 (gtint_2[26:26], choice_2, i_2r1[26:26]);
  AND2 I619 (gtint_2[27:27], choice_2, i_2r1[27:27]);
  AND2 I620 (gtint_2[28:28], choice_2, i_2r1[28:28]);
  AND2 I621 (gtint_2[29:29], choice_2, i_2r1[29:29]);
  AND2 I622 (gtint_2[30:30], choice_2, i_2r1[30:30]);
  AND2 I623 (gtint_2[31:31], choice_2, i_2r1[31:31]);
  AND2 I624 (gtint_2[32:32], choice_2, i_2r1[32:32]);
  AND2 I625 (gtint_2[33:33], choice_2, i_2r1[33:33]);
  AND2 I626 (gtint_2[34:34], choice_2, i_2r1[34:34]);
  AND2 I627 (gtint_2[35:35], choice_2, i_2r1[35:35]);
  AND2 I628 (gtint_2[36:36], choice_2, i_2r1[36:36]);
  AND2 I629 (gtint_2[37:37], choice_2, i_2r1[37:37]);
  AND2 I630 (gtint_2[38:38], choice_2, i_2r1[38:38]);
  AND2 I631 (gtint_2[39:39], choice_2, i_2r1[39:39]);
  AND2 I632 (gtint_2[40:40], choice_2, i_2r1[40:40]);
  AND2 I633 (gtint_2[41:41], choice_2, i_2r1[41:41]);
  AND2 I634 (gtint_2[42:42], choice_2, i_2r1[42:42]);
  AND2 I635 (gtint_2[43:43], choice_2, i_2r1[43:43]);
  AND2 I636 (gtint_2[44:44], choice_2, i_2r1[44:44]);
  AND2 I637 (gtint_2[45:45], choice_2, i_2r1[45:45]);
  AND2 I638 (gtint_2[46:46], choice_2, i_2r1[46:46]);
  AND2 I639 (gtint_2[47:47], choice_2, i_2r1[47:47]);
  AND2 I640 (gtint_2[48:48], choice_2, i_2r1[48:48]);
  AND2 I641 (gtint_2[49:49], choice_2, i_2r1[49:49]);
  AND2 I642 (gtint_2[50:50], choice_2, i_2r1[50:50]);
  AND2 I643 (gtint_2[51:51], choice_2, i_2r1[51:51]);
  AND2 I644 (gtint_2[52:52], choice_2, i_2r1[52:52]);
  AND2 I645 (gtint_2[53:53], choice_2, i_2r1[53:53]);
  AND2 I646 (gtint_2[54:54], choice_2, i_2r1[54:54]);
  AND2 I647 (gtint_2[55:55], choice_2, i_2r1[55:55]);
  AND2 I648 (gtint_2[56:56], choice_2, i_2r1[56:56]);
  AND2 I649 (gtint_2[57:57], choice_2, i_2r1[57:57]);
  AND2 I650 (gtint_2[58:58], choice_2, i_2r1[58:58]);
  AND2 I651 (gtint_2[59:59], choice_2, i_2r1[59:59]);
  AND2 I652 (gtint_2[60:60], choice_2, i_2r1[60:60]);
  AND2 I653 (gtint_2[61:61], choice_2, i_2r1[61:61]);
  AND2 I654 (gtint_2[62:62], choice_2, i_2r1[62:62]);
  AND2 I655 (gtint_2[63:63], choice_2, i_2r1[63:63]);
  AND2 I656 (gtint_2[64:64], choice_2, i_2r1[64:64]);
  AND2 I657 (gtint_2[65:65], choice_2, i_2r1[65:65]);
  AND2 I658 (gtint_2[66:66], choice_2, i_2r1[66:66]);
  AND2 I659 (gtint_2[67:67], choice_2, i_2r1[67:67]);
  AND2 I660 (gtint_2[68:68], choice_2, i_2r1[68:68]);
  AND2 I661 (gtint_2[69:69], choice_2, i_2r1[69:69]);
  AND2 I662 (gtint_2[70:70], choice_2, i_2r1[70:70]);
  AND2 I663 (gtint_2[71:71], choice_2, i_2r1[71:71]);
  AND2 I664 (gtint_2[72:72], choice_2, i_2r1[72:72]);
  AND2 I665 (gtint_2[73:73], choice_2, i_2r1[73:73]);
  AND2 I666 (gtint_3[0:0], choice_3, i_3r1[0:0]);
  AND2 I667 (gtint_3[1:1], choice_3, i_3r1[1:1]);
  AND2 I668 (gtint_3[2:2], choice_3, i_3r1[2:2]);
  AND2 I669 (gtint_3[3:3], choice_3, i_3r1[3:3]);
  AND2 I670 (gtint_3[4:4], choice_3, i_3r1[4:4]);
  AND2 I671 (gtint_3[5:5], choice_3, i_3r1[5:5]);
  AND2 I672 (gtint_3[6:6], choice_3, i_3r1[6:6]);
  AND2 I673 (gtint_3[7:7], choice_3, i_3r1[7:7]);
  AND2 I674 (gtint_3[8:8], choice_3, i_3r1[8:8]);
  AND2 I675 (gtint_3[9:9], choice_3, i_3r1[9:9]);
  AND2 I676 (gtint_3[10:10], choice_3, i_3r1[10:10]);
  AND2 I677 (gtint_3[11:11], choice_3, i_3r1[11:11]);
  AND2 I678 (gtint_3[12:12], choice_3, i_3r1[12:12]);
  AND2 I679 (gtint_3[13:13], choice_3, i_3r1[13:13]);
  AND2 I680 (gtint_3[14:14], choice_3, i_3r1[14:14]);
  AND2 I681 (gtint_3[15:15], choice_3, i_3r1[15:15]);
  AND2 I682 (gtint_3[16:16], choice_3, i_3r1[16:16]);
  AND2 I683 (gtint_3[17:17], choice_3, i_3r1[17:17]);
  AND2 I684 (gtint_3[18:18], choice_3, i_3r1[18:18]);
  AND2 I685 (gtint_3[19:19], choice_3, i_3r1[19:19]);
  AND2 I686 (gtint_3[20:20], choice_3, i_3r1[20:20]);
  AND2 I687 (gtint_3[21:21], choice_3, i_3r1[21:21]);
  AND2 I688 (gtint_3[22:22], choice_3, i_3r1[22:22]);
  AND2 I689 (gtint_3[23:23], choice_3, i_3r1[23:23]);
  AND2 I690 (gtint_3[24:24], choice_3, i_3r1[24:24]);
  AND2 I691 (gtint_3[25:25], choice_3, i_3r1[25:25]);
  AND2 I692 (gtint_3[26:26], choice_3, i_3r1[26:26]);
  AND2 I693 (gtint_3[27:27], choice_3, i_3r1[27:27]);
  AND2 I694 (gtint_3[28:28], choice_3, i_3r1[28:28]);
  AND2 I695 (gtint_3[29:29], choice_3, i_3r1[29:29]);
  AND2 I696 (gtint_3[30:30], choice_3, i_3r1[30:30]);
  AND2 I697 (gtint_3[31:31], choice_3, i_3r1[31:31]);
  AND2 I698 (gtint_3[32:32], choice_3, i_3r1[32:32]);
  AND2 I699 (gtint_3[33:33], choice_3, i_3r1[33:33]);
  AND2 I700 (gtint_3[34:34], choice_3, i_3r1[34:34]);
  AND2 I701 (gtint_3[35:35], choice_3, i_3r1[35:35]);
  AND2 I702 (gtint_3[36:36], choice_3, i_3r1[36:36]);
  AND2 I703 (gtint_3[37:37], choice_3, i_3r1[37:37]);
  AND2 I704 (gtint_3[38:38], choice_3, i_3r1[38:38]);
  AND2 I705 (gtint_3[39:39], choice_3, i_3r1[39:39]);
  AND2 I706 (gtint_3[40:40], choice_3, i_3r1[40:40]);
  AND2 I707 (gtint_3[41:41], choice_3, i_3r1[41:41]);
  AND2 I708 (gtint_3[42:42], choice_3, i_3r1[42:42]);
  AND2 I709 (gtint_3[43:43], choice_3, i_3r1[43:43]);
  AND2 I710 (gtint_3[44:44], choice_3, i_3r1[44:44]);
  AND2 I711 (gtint_3[45:45], choice_3, i_3r1[45:45]);
  AND2 I712 (gtint_3[46:46], choice_3, i_3r1[46:46]);
  AND2 I713 (gtint_3[47:47], choice_3, i_3r1[47:47]);
  AND2 I714 (gtint_3[48:48], choice_3, i_3r1[48:48]);
  AND2 I715 (gtint_3[49:49], choice_3, i_3r1[49:49]);
  AND2 I716 (gtint_3[50:50], choice_3, i_3r1[50:50]);
  AND2 I717 (gtint_3[51:51], choice_3, i_3r1[51:51]);
  AND2 I718 (gtint_3[52:52], choice_3, i_3r1[52:52]);
  AND2 I719 (gtint_3[53:53], choice_3, i_3r1[53:53]);
  AND2 I720 (gtint_3[54:54], choice_3, i_3r1[54:54]);
  AND2 I721 (gtint_3[55:55], choice_3, i_3r1[55:55]);
  AND2 I722 (gtint_3[56:56], choice_3, i_3r1[56:56]);
  AND2 I723 (gtint_3[57:57], choice_3, i_3r1[57:57]);
  AND2 I724 (gtint_3[58:58], choice_3, i_3r1[58:58]);
  AND2 I725 (gtint_3[59:59], choice_3, i_3r1[59:59]);
  AND2 I726 (gtint_3[60:60], choice_3, i_3r1[60:60]);
  AND2 I727 (gtint_3[61:61], choice_3, i_3r1[61:61]);
  AND2 I728 (gtint_3[62:62], choice_3, i_3r1[62:62]);
  AND2 I729 (gtint_3[63:63], choice_3, i_3r1[63:63]);
  AND2 I730 (gtint_3[64:64], choice_3, i_3r1[64:64]);
  AND2 I731 (gtint_3[65:65], choice_3, i_3r1[65:65]);
  AND2 I732 (gtint_3[66:66], choice_3, i_3r1[66:66]);
  AND2 I733 (gtint_3[67:67], choice_3, i_3r1[67:67]);
  AND2 I734 (gtint_3[68:68], choice_3, i_3r1[68:68]);
  AND2 I735 (gtint_3[69:69], choice_3, i_3r1[69:69]);
  AND2 I736 (gtint_3[70:70], choice_3, i_3r1[70:70]);
  AND2 I737 (gtint_3[71:71], choice_3, i_3r1[71:71]);
  AND2 I738 (gtint_3[72:72], choice_3, i_3r1[72:72]);
  AND2 I739 (gtint_3[73:73], choice_3, i_3r1[73:73]);
  AND2 I740 (gtint_4[0:0], choice_4, i_4r1[0:0]);
  AND2 I741 (gtint_4[1:1], choice_4, i_4r1[1:1]);
  AND2 I742 (gtint_4[2:2], choice_4, i_4r1[2:2]);
  AND2 I743 (gtint_4[3:3], choice_4, i_4r1[3:3]);
  AND2 I744 (gtint_4[4:4], choice_4, i_4r1[4:4]);
  AND2 I745 (gtint_4[5:5], choice_4, i_4r1[5:5]);
  AND2 I746 (gtint_4[6:6], choice_4, i_4r1[6:6]);
  AND2 I747 (gtint_4[7:7], choice_4, i_4r1[7:7]);
  AND2 I748 (gtint_4[8:8], choice_4, i_4r1[8:8]);
  AND2 I749 (gtint_4[9:9], choice_4, i_4r1[9:9]);
  AND2 I750 (gtint_4[10:10], choice_4, i_4r1[10:10]);
  AND2 I751 (gtint_4[11:11], choice_4, i_4r1[11:11]);
  AND2 I752 (gtint_4[12:12], choice_4, i_4r1[12:12]);
  AND2 I753 (gtint_4[13:13], choice_4, i_4r1[13:13]);
  AND2 I754 (gtint_4[14:14], choice_4, i_4r1[14:14]);
  AND2 I755 (gtint_4[15:15], choice_4, i_4r1[15:15]);
  AND2 I756 (gtint_4[16:16], choice_4, i_4r1[16:16]);
  AND2 I757 (gtint_4[17:17], choice_4, i_4r1[17:17]);
  AND2 I758 (gtint_4[18:18], choice_4, i_4r1[18:18]);
  AND2 I759 (gtint_4[19:19], choice_4, i_4r1[19:19]);
  AND2 I760 (gtint_4[20:20], choice_4, i_4r1[20:20]);
  AND2 I761 (gtint_4[21:21], choice_4, i_4r1[21:21]);
  AND2 I762 (gtint_4[22:22], choice_4, i_4r1[22:22]);
  AND2 I763 (gtint_4[23:23], choice_4, i_4r1[23:23]);
  AND2 I764 (gtint_4[24:24], choice_4, i_4r1[24:24]);
  AND2 I765 (gtint_4[25:25], choice_4, i_4r1[25:25]);
  AND2 I766 (gtint_4[26:26], choice_4, i_4r1[26:26]);
  AND2 I767 (gtint_4[27:27], choice_4, i_4r1[27:27]);
  AND2 I768 (gtint_4[28:28], choice_4, i_4r1[28:28]);
  AND2 I769 (gtint_4[29:29], choice_4, i_4r1[29:29]);
  AND2 I770 (gtint_4[30:30], choice_4, i_4r1[30:30]);
  AND2 I771 (gtint_4[31:31], choice_4, i_4r1[31:31]);
  AND2 I772 (gtint_4[32:32], choice_4, i_4r1[32:32]);
  AND2 I773 (gtint_4[33:33], choice_4, i_4r1[33:33]);
  AND2 I774 (gtint_4[34:34], choice_4, i_4r1[34:34]);
  AND2 I775 (gtint_4[35:35], choice_4, i_4r1[35:35]);
  AND2 I776 (gtint_4[36:36], choice_4, i_4r1[36:36]);
  AND2 I777 (gtint_4[37:37], choice_4, i_4r1[37:37]);
  AND2 I778 (gtint_4[38:38], choice_4, i_4r1[38:38]);
  AND2 I779 (gtint_4[39:39], choice_4, i_4r1[39:39]);
  AND2 I780 (gtint_4[40:40], choice_4, i_4r1[40:40]);
  AND2 I781 (gtint_4[41:41], choice_4, i_4r1[41:41]);
  AND2 I782 (gtint_4[42:42], choice_4, i_4r1[42:42]);
  AND2 I783 (gtint_4[43:43], choice_4, i_4r1[43:43]);
  AND2 I784 (gtint_4[44:44], choice_4, i_4r1[44:44]);
  AND2 I785 (gtint_4[45:45], choice_4, i_4r1[45:45]);
  AND2 I786 (gtint_4[46:46], choice_4, i_4r1[46:46]);
  AND2 I787 (gtint_4[47:47], choice_4, i_4r1[47:47]);
  AND2 I788 (gtint_4[48:48], choice_4, i_4r1[48:48]);
  AND2 I789 (gtint_4[49:49], choice_4, i_4r1[49:49]);
  AND2 I790 (gtint_4[50:50], choice_4, i_4r1[50:50]);
  AND2 I791 (gtint_4[51:51], choice_4, i_4r1[51:51]);
  AND2 I792 (gtint_4[52:52], choice_4, i_4r1[52:52]);
  AND2 I793 (gtint_4[53:53], choice_4, i_4r1[53:53]);
  AND2 I794 (gtint_4[54:54], choice_4, i_4r1[54:54]);
  AND2 I795 (gtint_4[55:55], choice_4, i_4r1[55:55]);
  AND2 I796 (gtint_4[56:56], choice_4, i_4r1[56:56]);
  AND2 I797 (gtint_4[57:57], choice_4, i_4r1[57:57]);
  AND2 I798 (gtint_4[58:58], choice_4, i_4r1[58:58]);
  AND2 I799 (gtint_4[59:59], choice_4, i_4r1[59:59]);
  AND2 I800 (gtint_4[60:60], choice_4, i_4r1[60:60]);
  AND2 I801 (gtint_4[61:61], choice_4, i_4r1[61:61]);
  AND2 I802 (gtint_4[62:62], choice_4, i_4r1[62:62]);
  AND2 I803 (gtint_4[63:63], choice_4, i_4r1[63:63]);
  AND2 I804 (gtint_4[64:64], choice_4, i_4r1[64:64]);
  AND2 I805 (gtint_4[65:65], choice_4, i_4r1[65:65]);
  AND2 I806 (gtint_4[66:66], choice_4, i_4r1[66:66]);
  AND2 I807 (gtint_4[67:67], choice_4, i_4r1[67:67]);
  AND2 I808 (gtint_4[68:68], choice_4, i_4r1[68:68]);
  AND2 I809 (gtint_4[69:69], choice_4, i_4r1[69:69]);
  AND2 I810 (gtint_4[70:70], choice_4, i_4r1[70:70]);
  AND2 I811 (gtint_4[71:71], choice_4, i_4r1[71:71]);
  AND2 I812 (gtint_4[72:72], choice_4, i_4r1[72:72]);
  AND2 I813 (gtint_4[73:73], choice_4, i_4r1[73:73]);
  AND2 I814 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I815 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I816 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I817 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I818 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I819 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I820 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I821 (gfint_0[7:7], choice_0, i_0r0[7:7]);
  AND2 I822 (gfint_0[8:8], choice_0, i_0r0[8:8]);
  AND2 I823 (gfint_0[9:9], choice_0, i_0r0[9:9]);
  AND2 I824 (gfint_0[10:10], choice_0, i_0r0[10:10]);
  AND2 I825 (gfint_0[11:11], choice_0, i_0r0[11:11]);
  AND2 I826 (gfint_0[12:12], choice_0, i_0r0[12:12]);
  AND2 I827 (gfint_0[13:13], choice_0, i_0r0[13:13]);
  AND2 I828 (gfint_0[14:14], choice_0, i_0r0[14:14]);
  AND2 I829 (gfint_0[15:15], choice_0, i_0r0[15:15]);
  AND2 I830 (gfint_0[16:16], choice_0, i_0r0[16:16]);
  AND2 I831 (gfint_0[17:17], choice_0, i_0r0[17:17]);
  AND2 I832 (gfint_0[18:18], choice_0, i_0r0[18:18]);
  AND2 I833 (gfint_0[19:19], choice_0, i_0r0[19:19]);
  AND2 I834 (gfint_0[20:20], choice_0, i_0r0[20:20]);
  AND2 I835 (gfint_0[21:21], choice_0, i_0r0[21:21]);
  AND2 I836 (gfint_0[22:22], choice_0, i_0r0[22:22]);
  AND2 I837 (gfint_0[23:23], choice_0, i_0r0[23:23]);
  AND2 I838 (gfint_0[24:24], choice_0, i_0r0[24:24]);
  AND2 I839 (gfint_0[25:25], choice_0, i_0r0[25:25]);
  AND2 I840 (gfint_0[26:26], choice_0, i_0r0[26:26]);
  AND2 I841 (gfint_0[27:27], choice_0, i_0r0[27:27]);
  AND2 I842 (gfint_0[28:28], choice_0, i_0r0[28:28]);
  AND2 I843 (gfint_0[29:29], choice_0, i_0r0[29:29]);
  AND2 I844 (gfint_0[30:30], choice_0, i_0r0[30:30]);
  AND2 I845 (gfint_0[31:31], choice_0, i_0r0[31:31]);
  AND2 I846 (gfint_0[32:32], choice_0, i_0r0[32:32]);
  AND2 I847 (gfint_0[33:33], choice_0, i_0r0[33:33]);
  AND2 I848 (gfint_0[34:34], choice_0, i_0r0[34:34]);
  AND2 I849 (gfint_0[35:35], choice_0, i_0r0[35:35]);
  AND2 I850 (gfint_0[36:36], choice_0, i_0r0[36:36]);
  AND2 I851 (gfint_0[37:37], choice_0, i_0r0[37:37]);
  AND2 I852 (gfint_0[38:38], choice_0, i_0r0[38:38]);
  AND2 I853 (gfint_0[39:39], choice_0, i_0r0[39:39]);
  AND2 I854 (gfint_0[40:40], choice_0, i_0r0[40:40]);
  AND2 I855 (gfint_0[41:41], choice_0, i_0r0[41:41]);
  AND2 I856 (gfint_0[42:42], choice_0, i_0r0[42:42]);
  AND2 I857 (gfint_0[43:43], choice_0, i_0r0[43:43]);
  AND2 I858 (gfint_0[44:44], choice_0, i_0r0[44:44]);
  AND2 I859 (gfint_0[45:45], choice_0, i_0r0[45:45]);
  AND2 I860 (gfint_0[46:46], choice_0, i_0r0[46:46]);
  AND2 I861 (gfint_0[47:47], choice_0, i_0r0[47:47]);
  AND2 I862 (gfint_0[48:48], choice_0, i_0r0[48:48]);
  AND2 I863 (gfint_0[49:49], choice_0, i_0r0[49:49]);
  AND2 I864 (gfint_0[50:50], choice_0, i_0r0[50:50]);
  AND2 I865 (gfint_0[51:51], choice_0, i_0r0[51:51]);
  AND2 I866 (gfint_0[52:52], choice_0, i_0r0[52:52]);
  AND2 I867 (gfint_0[53:53], choice_0, i_0r0[53:53]);
  AND2 I868 (gfint_0[54:54], choice_0, i_0r0[54:54]);
  AND2 I869 (gfint_0[55:55], choice_0, i_0r0[55:55]);
  AND2 I870 (gfint_0[56:56], choice_0, i_0r0[56:56]);
  AND2 I871 (gfint_0[57:57], choice_0, i_0r0[57:57]);
  AND2 I872 (gfint_0[58:58], choice_0, i_0r0[58:58]);
  AND2 I873 (gfint_0[59:59], choice_0, i_0r0[59:59]);
  AND2 I874 (gfint_0[60:60], choice_0, i_0r0[60:60]);
  AND2 I875 (gfint_0[61:61], choice_0, i_0r0[61:61]);
  AND2 I876 (gfint_0[62:62], choice_0, i_0r0[62:62]);
  AND2 I877 (gfint_0[63:63], choice_0, i_0r0[63:63]);
  AND2 I878 (gfint_0[64:64], choice_0, i_0r0[64:64]);
  AND2 I879 (gfint_0[65:65], choice_0, i_0r0[65:65]);
  AND2 I880 (gfint_0[66:66], choice_0, i_0r0[66:66]);
  AND2 I881 (gfint_0[67:67], choice_0, i_0r0[67:67]);
  AND2 I882 (gfint_0[68:68], choice_0, i_0r0[68:68]);
  AND2 I883 (gfint_0[69:69], choice_0, i_0r0[69:69]);
  AND2 I884 (gfint_0[70:70], choice_0, i_0r0[70:70]);
  AND2 I885 (gfint_0[71:71], choice_0, i_0r0[71:71]);
  AND2 I886 (gfint_0[72:72], choice_0, i_0r0[72:72]);
  AND2 I887 (gfint_0[73:73], choice_0, i_0r0[73:73]);
  AND2 I888 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I889 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I890 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I891 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I892 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I893 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I894 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I895 (gfint_1[7:7], choice_1, i_1r0[7:7]);
  AND2 I896 (gfint_1[8:8], choice_1, i_1r0[8:8]);
  AND2 I897 (gfint_1[9:9], choice_1, i_1r0[9:9]);
  AND2 I898 (gfint_1[10:10], choice_1, i_1r0[10:10]);
  AND2 I899 (gfint_1[11:11], choice_1, i_1r0[11:11]);
  AND2 I900 (gfint_1[12:12], choice_1, i_1r0[12:12]);
  AND2 I901 (gfint_1[13:13], choice_1, i_1r0[13:13]);
  AND2 I902 (gfint_1[14:14], choice_1, i_1r0[14:14]);
  AND2 I903 (gfint_1[15:15], choice_1, i_1r0[15:15]);
  AND2 I904 (gfint_1[16:16], choice_1, i_1r0[16:16]);
  AND2 I905 (gfint_1[17:17], choice_1, i_1r0[17:17]);
  AND2 I906 (gfint_1[18:18], choice_1, i_1r0[18:18]);
  AND2 I907 (gfint_1[19:19], choice_1, i_1r0[19:19]);
  AND2 I908 (gfint_1[20:20], choice_1, i_1r0[20:20]);
  AND2 I909 (gfint_1[21:21], choice_1, i_1r0[21:21]);
  AND2 I910 (gfint_1[22:22], choice_1, i_1r0[22:22]);
  AND2 I911 (gfint_1[23:23], choice_1, i_1r0[23:23]);
  AND2 I912 (gfint_1[24:24], choice_1, i_1r0[24:24]);
  AND2 I913 (gfint_1[25:25], choice_1, i_1r0[25:25]);
  AND2 I914 (gfint_1[26:26], choice_1, i_1r0[26:26]);
  AND2 I915 (gfint_1[27:27], choice_1, i_1r0[27:27]);
  AND2 I916 (gfint_1[28:28], choice_1, i_1r0[28:28]);
  AND2 I917 (gfint_1[29:29], choice_1, i_1r0[29:29]);
  AND2 I918 (gfint_1[30:30], choice_1, i_1r0[30:30]);
  AND2 I919 (gfint_1[31:31], choice_1, i_1r0[31:31]);
  AND2 I920 (gfint_1[32:32], choice_1, i_1r0[32:32]);
  AND2 I921 (gfint_1[33:33], choice_1, i_1r0[33:33]);
  AND2 I922 (gfint_1[34:34], choice_1, i_1r0[34:34]);
  AND2 I923 (gfint_1[35:35], choice_1, i_1r0[35:35]);
  AND2 I924 (gfint_1[36:36], choice_1, i_1r0[36:36]);
  AND2 I925 (gfint_1[37:37], choice_1, i_1r0[37:37]);
  AND2 I926 (gfint_1[38:38], choice_1, i_1r0[38:38]);
  AND2 I927 (gfint_1[39:39], choice_1, i_1r0[39:39]);
  AND2 I928 (gfint_1[40:40], choice_1, i_1r0[40:40]);
  AND2 I929 (gfint_1[41:41], choice_1, i_1r0[41:41]);
  AND2 I930 (gfint_1[42:42], choice_1, i_1r0[42:42]);
  AND2 I931 (gfint_1[43:43], choice_1, i_1r0[43:43]);
  AND2 I932 (gfint_1[44:44], choice_1, i_1r0[44:44]);
  AND2 I933 (gfint_1[45:45], choice_1, i_1r0[45:45]);
  AND2 I934 (gfint_1[46:46], choice_1, i_1r0[46:46]);
  AND2 I935 (gfint_1[47:47], choice_1, i_1r0[47:47]);
  AND2 I936 (gfint_1[48:48], choice_1, i_1r0[48:48]);
  AND2 I937 (gfint_1[49:49], choice_1, i_1r0[49:49]);
  AND2 I938 (gfint_1[50:50], choice_1, i_1r0[50:50]);
  AND2 I939 (gfint_1[51:51], choice_1, i_1r0[51:51]);
  AND2 I940 (gfint_1[52:52], choice_1, i_1r0[52:52]);
  AND2 I941 (gfint_1[53:53], choice_1, i_1r0[53:53]);
  AND2 I942 (gfint_1[54:54], choice_1, i_1r0[54:54]);
  AND2 I943 (gfint_1[55:55], choice_1, i_1r0[55:55]);
  AND2 I944 (gfint_1[56:56], choice_1, i_1r0[56:56]);
  AND2 I945 (gfint_1[57:57], choice_1, i_1r0[57:57]);
  AND2 I946 (gfint_1[58:58], choice_1, i_1r0[58:58]);
  AND2 I947 (gfint_1[59:59], choice_1, i_1r0[59:59]);
  AND2 I948 (gfint_1[60:60], choice_1, i_1r0[60:60]);
  AND2 I949 (gfint_1[61:61], choice_1, i_1r0[61:61]);
  AND2 I950 (gfint_1[62:62], choice_1, i_1r0[62:62]);
  AND2 I951 (gfint_1[63:63], choice_1, i_1r0[63:63]);
  AND2 I952 (gfint_1[64:64], choice_1, i_1r0[64:64]);
  AND2 I953 (gfint_1[65:65], choice_1, i_1r0[65:65]);
  AND2 I954 (gfint_1[66:66], choice_1, i_1r0[66:66]);
  AND2 I955 (gfint_1[67:67], choice_1, i_1r0[67:67]);
  AND2 I956 (gfint_1[68:68], choice_1, i_1r0[68:68]);
  AND2 I957 (gfint_1[69:69], choice_1, i_1r0[69:69]);
  AND2 I958 (gfint_1[70:70], choice_1, i_1r0[70:70]);
  AND2 I959 (gfint_1[71:71], choice_1, i_1r0[71:71]);
  AND2 I960 (gfint_1[72:72], choice_1, i_1r0[72:72]);
  AND2 I961 (gfint_1[73:73], choice_1, i_1r0[73:73]);
  AND2 I962 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I963 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I964 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I965 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AND2 I966 (gfint_2[4:4], choice_2, i_2r0[4:4]);
  AND2 I967 (gfint_2[5:5], choice_2, i_2r0[5:5]);
  AND2 I968 (gfint_2[6:6], choice_2, i_2r0[6:6]);
  AND2 I969 (gfint_2[7:7], choice_2, i_2r0[7:7]);
  AND2 I970 (gfint_2[8:8], choice_2, i_2r0[8:8]);
  AND2 I971 (gfint_2[9:9], choice_2, i_2r0[9:9]);
  AND2 I972 (gfint_2[10:10], choice_2, i_2r0[10:10]);
  AND2 I973 (gfint_2[11:11], choice_2, i_2r0[11:11]);
  AND2 I974 (gfint_2[12:12], choice_2, i_2r0[12:12]);
  AND2 I975 (gfint_2[13:13], choice_2, i_2r0[13:13]);
  AND2 I976 (gfint_2[14:14], choice_2, i_2r0[14:14]);
  AND2 I977 (gfint_2[15:15], choice_2, i_2r0[15:15]);
  AND2 I978 (gfint_2[16:16], choice_2, i_2r0[16:16]);
  AND2 I979 (gfint_2[17:17], choice_2, i_2r0[17:17]);
  AND2 I980 (gfint_2[18:18], choice_2, i_2r0[18:18]);
  AND2 I981 (gfint_2[19:19], choice_2, i_2r0[19:19]);
  AND2 I982 (gfint_2[20:20], choice_2, i_2r0[20:20]);
  AND2 I983 (gfint_2[21:21], choice_2, i_2r0[21:21]);
  AND2 I984 (gfint_2[22:22], choice_2, i_2r0[22:22]);
  AND2 I985 (gfint_2[23:23], choice_2, i_2r0[23:23]);
  AND2 I986 (gfint_2[24:24], choice_2, i_2r0[24:24]);
  AND2 I987 (gfint_2[25:25], choice_2, i_2r0[25:25]);
  AND2 I988 (gfint_2[26:26], choice_2, i_2r0[26:26]);
  AND2 I989 (gfint_2[27:27], choice_2, i_2r0[27:27]);
  AND2 I990 (gfint_2[28:28], choice_2, i_2r0[28:28]);
  AND2 I991 (gfint_2[29:29], choice_2, i_2r0[29:29]);
  AND2 I992 (gfint_2[30:30], choice_2, i_2r0[30:30]);
  AND2 I993 (gfint_2[31:31], choice_2, i_2r0[31:31]);
  AND2 I994 (gfint_2[32:32], choice_2, i_2r0[32:32]);
  AND2 I995 (gfint_2[33:33], choice_2, i_2r0[33:33]);
  AND2 I996 (gfint_2[34:34], choice_2, i_2r0[34:34]);
  AND2 I997 (gfint_2[35:35], choice_2, i_2r0[35:35]);
  AND2 I998 (gfint_2[36:36], choice_2, i_2r0[36:36]);
  AND2 I999 (gfint_2[37:37], choice_2, i_2r0[37:37]);
  AND2 I1000 (gfint_2[38:38], choice_2, i_2r0[38:38]);
  AND2 I1001 (gfint_2[39:39], choice_2, i_2r0[39:39]);
  AND2 I1002 (gfint_2[40:40], choice_2, i_2r0[40:40]);
  AND2 I1003 (gfint_2[41:41], choice_2, i_2r0[41:41]);
  AND2 I1004 (gfint_2[42:42], choice_2, i_2r0[42:42]);
  AND2 I1005 (gfint_2[43:43], choice_2, i_2r0[43:43]);
  AND2 I1006 (gfint_2[44:44], choice_2, i_2r0[44:44]);
  AND2 I1007 (gfint_2[45:45], choice_2, i_2r0[45:45]);
  AND2 I1008 (gfint_2[46:46], choice_2, i_2r0[46:46]);
  AND2 I1009 (gfint_2[47:47], choice_2, i_2r0[47:47]);
  AND2 I1010 (gfint_2[48:48], choice_2, i_2r0[48:48]);
  AND2 I1011 (gfint_2[49:49], choice_2, i_2r0[49:49]);
  AND2 I1012 (gfint_2[50:50], choice_2, i_2r0[50:50]);
  AND2 I1013 (gfint_2[51:51], choice_2, i_2r0[51:51]);
  AND2 I1014 (gfint_2[52:52], choice_2, i_2r0[52:52]);
  AND2 I1015 (gfint_2[53:53], choice_2, i_2r0[53:53]);
  AND2 I1016 (gfint_2[54:54], choice_2, i_2r0[54:54]);
  AND2 I1017 (gfint_2[55:55], choice_2, i_2r0[55:55]);
  AND2 I1018 (gfint_2[56:56], choice_2, i_2r0[56:56]);
  AND2 I1019 (gfint_2[57:57], choice_2, i_2r0[57:57]);
  AND2 I1020 (gfint_2[58:58], choice_2, i_2r0[58:58]);
  AND2 I1021 (gfint_2[59:59], choice_2, i_2r0[59:59]);
  AND2 I1022 (gfint_2[60:60], choice_2, i_2r0[60:60]);
  AND2 I1023 (gfint_2[61:61], choice_2, i_2r0[61:61]);
  AND2 I1024 (gfint_2[62:62], choice_2, i_2r0[62:62]);
  AND2 I1025 (gfint_2[63:63], choice_2, i_2r0[63:63]);
  AND2 I1026 (gfint_2[64:64], choice_2, i_2r0[64:64]);
  AND2 I1027 (gfint_2[65:65], choice_2, i_2r0[65:65]);
  AND2 I1028 (gfint_2[66:66], choice_2, i_2r0[66:66]);
  AND2 I1029 (gfint_2[67:67], choice_2, i_2r0[67:67]);
  AND2 I1030 (gfint_2[68:68], choice_2, i_2r0[68:68]);
  AND2 I1031 (gfint_2[69:69], choice_2, i_2r0[69:69]);
  AND2 I1032 (gfint_2[70:70], choice_2, i_2r0[70:70]);
  AND2 I1033 (gfint_2[71:71], choice_2, i_2r0[71:71]);
  AND2 I1034 (gfint_2[72:72], choice_2, i_2r0[72:72]);
  AND2 I1035 (gfint_2[73:73], choice_2, i_2r0[73:73]);
  AND2 I1036 (gfint_3[0:0], choice_3, i_3r0[0:0]);
  AND2 I1037 (gfint_3[1:1], choice_3, i_3r0[1:1]);
  AND2 I1038 (gfint_3[2:2], choice_3, i_3r0[2:2]);
  AND2 I1039 (gfint_3[3:3], choice_3, i_3r0[3:3]);
  AND2 I1040 (gfint_3[4:4], choice_3, i_3r0[4:4]);
  AND2 I1041 (gfint_3[5:5], choice_3, i_3r0[5:5]);
  AND2 I1042 (gfint_3[6:6], choice_3, i_3r0[6:6]);
  AND2 I1043 (gfint_3[7:7], choice_3, i_3r0[7:7]);
  AND2 I1044 (gfint_3[8:8], choice_3, i_3r0[8:8]);
  AND2 I1045 (gfint_3[9:9], choice_3, i_3r0[9:9]);
  AND2 I1046 (gfint_3[10:10], choice_3, i_3r0[10:10]);
  AND2 I1047 (gfint_3[11:11], choice_3, i_3r0[11:11]);
  AND2 I1048 (gfint_3[12:12], choice_3, i_3r0[12:12]);
  AND2 I1049 (gfint_3[13:13], choice_3, i_3r0[13:13]);
  AND2 I1050 (gfint_3[14:14], choice_3, i_3r0[14:14]);
  AND2 I1051 (gfint_3[15:15], choice_3, i_3r0[15:15]);
  AND2 I1052 (gfint_3[16:16], choice_3, i_3r0[16:16]);
  AND2 I1053 (gfint_3[17:17], choice_3, i_3r0[17:17]);
  AND2 I1054 (gfint_3[18:18], choice_3, i_3r0[18:18]);
  AND2 I1055 (gfint_3[19:19], choice_3, i_3r0[19:19]);
  AND2 I1056 (gfint_3[20:20], choice_3, i_3r0[20:20]);
  AND2 I1057 (gfint_3[21:21], choice_3, i_3r0[21:21]);
  AND2 I1058 (gfint_3[22:22], choice_3, i_3r0[22:22]);
  AND2 I1059 (gfint_3[23:23], choice_3, i_3r0[23:23]);
  AND2 I1060 (gfint_3[24:24], choice_3, i_3r0[24:24]);
  AND2 I1061 (gfint_3[25:25], choice_3, i_3r0[25:25]);
  AND2 I1062 (gfint_3[26:26], choice_3, i_3r0[26:26]);
  AND2 I1063 (gfint_3[27:27], choice_3, i_3r0[27:27]);
  AND2 I1064 (gfint_3[28:28], choice_3, i_3r0[28:28]);
  AND2 I1065 (gfint_3[29:29], choice_3, i_3r0[29:29]);
  AND2 I1066 (gfint_3[30:30], choice_3, i_3r0[30:30]);
  AND2 I1067 (gfint_3[31:31], choice_3, i_3r0[31:31]);
  AND2 I1068 (gfint_3[32:32], choice_3, i_3r0[32:32]);
  AND2 I1069 (gfint_3[33:33], choice_3, i_3r0[33:33]);
  AND2 I1070 (gfint_3[34:34], choice_3, i_3r0[34:34]);
  AND2 I1071 (gfint_3[35:35], choice_3, i_3r0[35:35]);
  AND2 I1072 (gfint_3[36:36], choice_3, i_3r0[36:36]);
  AND2 I1073 (gfint_3[37:37], choice_3, i_3r0[37:37]);
  AND2 I1074 (gfint_3[38:38], choice_3, i_3r0[38:38]);
  AND2 I1075 (gfint_3[39:39], choice_3, i_3r0[39:39]);
  AND2 I1076 (gfint_3[40:40], choice_3, i_3r0[40:40]);
  AND2 I1077 (gfint_3[41:41], choice_3, i_3r0[41:41]);
  AND2 I1078 (gfint_3[42:42], choice_3, i_3r0[42:42]);
  AND2 I1079 (gfint_3[43:43], choice_3, i_3r0[43:43]);
  AND2 I1080 (gfint_3[44:44], choice_3, i_3r0[44:44]);
  AND2 I1081 (gfint_3[45:45], choice_3, i_3r0[45:45]);
  AND2 I1082 (gfint_3[46:46], choice_3, i_3r0[46:46]);
  AND2 I1083 (gfint_3[47:47], choice_3, i_3r0[47:47]);
  AND2 I1084 (gfint_3[48:48], choice_3, i_3r0[48:48]);
  AND2 I1085 (gfint_3[49:49], choice_3, i_3r0[49:49]);
  AND2 I1086 (gfint_3[50:50], choice_3, i_3r0[50:50]);
  AND2 I1087 (gfint_3[51:51], choice_3, i_3r0[51:51]);
  AND2 I1088 (gfint_3[52:52], choice_3, i_3r0[52:52]);
  AND2 I1089 (gfint_3[53:53], choice_3, i_3r0[53:53]);
  AND2 I1090 (gfint_3[54:54], choice_3, i_3r0[54:54]);
  AND2 I1091 (gfint_3[55:55], choice_3, i_3r0[55:55]);
  AND2 I1092 (gfint_3[56:56], choice_3, i_3r0[56:56]);
  AND2 I1093 (gfint_3[57:57], choice_3, i_3r0[57:57]);
  AND2 I1094 (gfint_3[58:58], choice_3, i_3r0[58:58]);
  AND2 I1095 (gfint_3[59:59], choice_3, i_3r0[59:59]);
  AND2 I1096 (gfint_3[60:60], choice_3, i_3r0[60:60]);
  AND2 I1097 (gfint_3[61:61], choice_3, i_3r0[61:61]);
  AND2 I1098 (gfint_3[62:62], choice_3, i_3r0[62:62]);
  AND2 I1099 (gfint_3[63:63], choice_3, i_3r0[63:63]);
  AND2 I1100 (gfint_3[64:64], choice_3, i_3r0[64:64]);
  AND2 I1101 (gfint_3[65:65], choice_3, i_3r0[65:65]);
  AND2 I1102 (gfint_3[66:66], choice_3, i_3r0[66:66]);
  AND2 I1103 (gfint_3[67:67], choice_3, i_3r0[67:67]);
  AND2 I1104 (gfint_3[68:68], choice_3, i_3r0[68:68]);
  AND2 I1105 (gfint_3[69:69], choice_3, i_3r0[69:69]);
  AND2 I1106 (gfint_3[70:70], choice_3, i_3r0[70:70]);
  AND2 I1107 (gfint_3[71:71], choice_3, i_3r0[71:71]);
  AND2 I1108 (gfint_3[72:72], choice_3, i_3r0[72:72]);
  AND2 I1109 (gfint_3[73:73], choice_3, i_3r0[73:73]);
  AND2 I1110 (gfint_4[0:0], choice_4, i_4r0[0:0]);
  AND2 I1111 (gfint_4[1:1], choice_4, i_4r0[1:1]);
  AND2 I1112 (gfint_4[2:2], choice_4, i_4r0[2:2]);
  AND2 I1113 (gfint_4[3:3], choice_4, i_4r0[3:3]);
  AND2 I1114 (gfint_4[4:4], choice_4, i_4r0[4:4]);
  AND2 I1115 (gfint_4[5:5], choice_4, i_4r0[5:5]);
  AND2 I1116 (gfint_4[6:6], choice_4, i_4r0[6:6]);
  AND2 I1117 (gfint_4[7:7], choice_4, i_4r0[7:7]);
  AND2 I1118 (gfint_4[8:8], choice_4, i_4r0[8:8]);
  AND2 I1119 (gfint_4[9:9], choice_4, i_4r0[9:9]);
  AND2 I1120 (gfint_4[10:10], choice_4, i_4r0[10:10]);
  AND2 I1121 (gfint_4[11:11], choice_4, i_4r0[11:11]);
  AND2 I1122 (gfint_4[12:12], choice_4, i_4r0[12:12]);
  AND2 I1123 (gfint_4[13:13], choice_4, i_4r0[13:13]);
  AND2 I1124 (gfint_4[14:14], choice_4, i_4r0[14:14]);
  AND2 I1125 (gfint_4[15:15], choice_4, i_4r0[15:15]);
  AND2 I1126 (gfint_4[16:16], choice_4, i_4r0[16:16]);
  AND2 I1127 (gfint_4[17:17], choice_4, i_4r0[17:17]);
  AND2 I1128 (gfint_4[18:18], choice_4, i_4r0[18:18]);
  AND2 I1129 (gfint_4[19:19], choice_4, i_4r0[19:19]);
  AND2 I1130 (gfint_4[20:20], choice_4, i_4r0[20:20]);
  AND2 I1131 (gfint_4[21:21], choice_4, i_4r0[21:21]);
  AND2 I1132 (gfint_4[22:22], choice_4, i_4r0[22:22]);
  AND2 I1133 (gfint_4[23:23], choice_4, i_4r0[23:23]);
  AND2 I1134 (gfint_4[24:24], choice_4, i_4r0[24:24]);
  AND2 I1135 (gfint_4[25:25], choice_4, i_4r0[25:25]);
  AND2 I1136 (gfint_4[26:26], choice_4, i_4r0[26:26]);
  AND2 I1137 (gfint_4[27:27], choice_4, i_4r0[27:27]);
  AND2 I1138 (gfint_4[28:28], choice_4, i_4r0[28:28]);
  AND2 I1139 (gfint_4[29:29], choice_4, i_4r0[29:29]);
  AND2 I1140 (gfint_4[30:30], choice_4, i_4r0[30:30]);
  AND2 I1141 (gfint_4[31:31], choice_4, i_4r0[31:31]);
  AND2 I1142 (gfint_4[32:32], choice_4, i_4r0[32:32]);
  AND2 I1143 (gfint_4[33:33], choice_4, i_4r0[33:33]);
  AND2 I1144 (gfint_4[34:34], choice_4, i_4r0[34:34]);
  AND2 I1145 (gfint_4[35:35], choice_4, i_4r0[35:35]);
  AND2 I1146 (gfint_4[36:36], choice_4, i_4r0[36:36]);
  AND2 I1147 (gfint_4[37:37], choice_4, i_4r0[37:37]);
  AND2 I1148 (gfint_4[38:38], choice_4, i_4r0[38:38]);
  AND2 I1149 (gfint_4[39:39], choice_4, i_4r0[39:39]);
  AND2 I1150 (gfint_4[40:40], choice_4, i_4r0[40:40]);
  AND2 I1151 (gfint_4[41:41], choice_4, i_4r0[41:41]);
  AND2 I1152 (gfint_4[42:42], choice_4, i_4r0[42:42]);
  AND2 I1153 (gfint_4[43:43], choice_4, i_4r0[43:43]);
  AND2 I1154 (gfint_4[44:44], choice_4, i_4r0[44:44]);
  AND2 I1155 (gfint_4[45:45], choice_4, i_4r0[45:45]);
  AND2 I1156 (gfint_4[46:46], choice_4, i_4r0[46:46]);
  AND2 I1157 (gfint_4[47:47], choice_4, i_4r0[47:47]);
  AND2 I1158 (gfint_4[48:48], choice_4, i_4r0[48:48]);
  AND2 I1159 (gfint_4[49:49], choice_4, i_4r0[49:49]);
  AND2 I1160 (gfint_4[50:50], choice_4, i_4r0[50:50]);
  AND2 I1161 (gfint_4[51:51], choice_4, i_4r0[51:51]);
  AND2 I1162 (gfint_4[52:52], choice_4, i_4r0[52:52]);
  AND2 I1163 (gfint_4[53:53], choice_4, i_4r0[53:53]);
  AND2 I1164 (gfint_4[54:54], choice_4, i_4r0[54:54]);
  AND2 I1165 (gfint_4[55:55], choice_4, i_4r0[55:55]);
  AND2 I1166 (gfint_4[56:56], choice_4, i_4r0[56:56]);
  AND2 I1167 (gfint_4[57:57], choice_4, i_4r0[57:57]);
  AND2 I1168 (gfint_4[58:58], choice_4, i_4r0[58:58]);
  AND2 I1169 (gfint_4[59:59], choice_4, i_4r0[59:59]);
  AND2 I1170 (gfint_4[60:60], choice_4, i_4r0[60:60]);
  AND2 I1171 (gfint_4[61:61], choice_4, i_4r0[61:61]);
  AND2 I1172 (gfint_4[62:62], choice_4, i_4r0[62:62]);
  AND2 I1173 (gfint_4[63:63], choice_4, i_4r0[63:63]);
  AND2 I1174 (gfint_4[64:64], choice_4, i_4r0[64:64]);
  AND2 I1175 (gfint_4[65:65], choice_4, i_4r0[65:65]);
  AND2 I1176 (gfint_4[66:66], choice_4, i_4r0[66:66]);
  AND2 I1177 (gfint_4[67:67], choice_4, i_4r0[67:67]);
  AND2 I1178 (gfint_4[68:68], choice_4, i_4r0[68:68]);
  AND2 I1179 (gfint_4[69:69], choice_4, i_4r0[69:69]);
  AND2 I1180 (gfint_4[70:70], choice_4, i_4r0[70:70]);
  AND2 I1181 (gfint_4[71:71], choice_4, i_4r0[71:71]);
  AND2 I1182 (gfint_4[72:72], choice_4, i_4r0[72:72]);
  AND2 I1183 (gfint_4[73:73], choice_4, i_4r0[73:73]);
  OR2 I1184 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1185 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I1186 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I1187 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I1188 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I1189 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I1190 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I1191 (comp0_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I1192 (comp0_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I1193 (comp0_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I1194 (comp0_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I1195 (comp0_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I1196 (comp0_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I1197 (comp0_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I1198 (comp0_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I1199 (comp0_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I1200 (comp0_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I1201 (comp0_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I1202 (comp0_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I1203 (comp0_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I1204 (comp0_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I1205 (comp0_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I1206 (comp0_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I1207 (comp0_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I1208 (comp0_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I1209 (comp0_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I1210 (comp0_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I1211 (comp0_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I1212 (comp0_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I1213 (comp0_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I1214 (comp0_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I1215 (comp0_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I1216 (comp0_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  OR2 I1217 (comp0_0[33:33], i_0r0[33:33], i_0r1[33:33]);
  OR2 I1218 (comp0_0[34:34], i_0r0[34:34], i_0r1[34:34]);
  OR2 I1219 (comp0_0[35:35], i_0r0[35:35], i_0r1[35:35]);
  OR2 I1220 (comp0_0[36:36], i_0r0[36:36], i_0r1[36:36]);
  OR2 I1221 (comp0_0[37:37], i_0r0[37:37], i_0r1[37:37]);
  OR2 I1222 (comp0_0[38:38], i_0r0[38:38], i_0r1[38:38]);
  OR2 I1223 (comp0_0[39:39], i_0r0[39:39], i_0r1[39:39]);
  OR2 I1224 (comp0_0[40:40], i_0r0[40:40], i_0r1[40:40]);
  OR2 I1225 (comp0_0[41:41], i_0r0[41:41], i_0r1[41:41]);
  OR2 I1226 (comp0_0[42:42], i_0r0[42:42], i_0r1[42:42]);
  OR2 I1227 (comp0_0[43:43], i_0r0[43:43], i_0r1[43:43]);
  OR2 I1228 (comp0_0[44:44], i_0r0[44:44], i_0r1[44:44]);
  OR2 I1229 (comp0_0[45:45], i_0r0[45:45], i_0r1[45:45]);
  OR2 I1230 (comp0_0[46:46], i_0r0[46:46], i_0r1[46:46]);
  OR2 I1231 (comp0_0[47:47], i_0r0[47:47], i_0r1[47:47]);
  OR2 I1232 (comp0_0[48:48], i_0r0[48:48], i_0r1[48:48]);
  OR2 I1233 (comp0_0[49:49], i_0r0[49:49], i_0r1[49:49]);
  OR2 I1234 (comp0_0[50:50], i_0r0[50:50], i_0r1[50:50]);
  OR2 I1235 (comp0_0[51:51], i_0r0[51:51], i_0r1[51:51]);
  OR2 I1236 (comp0_0[52:52], i_0r0[52:52], i_0r1[52:52]);
  OR2 I1237 (comp0_0[53:53], i_0r0[53:53], i_0r1[53:53]);
  OR2 I1238 (comp0_0[54:54], i_0r0[54:54], i_0r1[54:54]);
  OR2 I1239 (comp0_0[55:55], i_0r0[55:55], i_0r1[55:55]);
  OR2 I1240 (comp0_0[56:56], i_0r0[56:56], i_0r1[56:56]);
  OR2 I1241 (comp0_0[57:57], i_0r0[57:57], i_0r1[57:57]);
  OR2 I1242 (comp0_0[58:58], i_0r0[58:58], i_0r1[58:58]);
  OR2 I1243 (comp0_0[59:59], i_0r0[59:59], i_0r1[59:59]);
  OR2 I1244 (comp0_0[60:60], i_0r0[60:60], i_0r1[60:60]);
  OR2 I1245 (comp0_0[61:61], i_0r0[61:61], i_0r1[61:61]);
  OR2 I1246 (comp0_0[62:62], i_0r0[62:62], i_0r1[62:62]);
  OR2 I1247 (comp0_0[63:63], i_0r0[63:63], i_0r1[63:63]);
  OR2 I1248 (comp0_0[64:64], i_0r0[64:64], i_0r1[64:64]);
  OR2 I1249 (comp0_0[65:65], i_0r0[65:65], i_0r1[65:65]);
  OR2 I1250 (comp0_0[66:66], i_0r0[66:66], i_0r1[66:66]);
  OR2 I1251 (comp0_0[67:67], i_0r0[67:67], i_0r1[67:67]);
  OR2 I1252 (comp0_0[68:68], i_0r0[68:68], i_0r1[68:68]);
  OR2 I1253 (comp0_0[69:69], i_0r0[69:69], i_0r1[69:69]);
  OR2 I1254 (comp0_0[70:70], i_0r0[70:70], i_0r1[70:70]);
  OR2 I1255 (comp0_0[71:71], i_0r0[71:71], i_0r1[71:71]);
  OR2 I1256 (comp0_0[72:72], i_0r0[72:72], i_0r1[72:72]);
  OR2 I1257 (comp0_0[73:73], i_0r0[73:73], i_0r1[73:73]);
  C3 I1258 (simp9851_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I1259 (simp9851_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I1260 (simp9851_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I1261 (simp9851_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I1262 (simp9851_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I1263 (simp9851_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I1264 (simp9851_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I1265 (simp9851_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I1266 (simp9851_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I1267 (simp9851_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C3 I1268 (simp9851_0[10:10], comp0_0[30:30], comp0_0[31:31], comp0_0[32:32]);
  C3 I1269 (simp9851_0[11:11], comp0_0[33:33], comp0_0[34:34], comp0_0[35:35]);
  C3 I1270 (simp9851_0[12:12], comp0_0[36:36], comp0_0[37:37], comp0_0[38:38]);
  C3 I1271 (simp9851_0[13:13], comp0_0[39:39], comp0_0[40:40], comp0_0[41:41]);
  C3 I1272 (simp9851_0[14:14], comp0_0[42:42], comp0_0[43:43], comp0_0[44:44]);
  C3 I1273 (simp9851_0[15:15], comp0_0[45:45], comp0_0[46:46], comp0_0[47:47]);
  C3 I1274 (simp9851_0[16:16], comp0_0[48:48], comp0_0[49:49], comp0_0[50:50]);
  C3 I1275 (simp9851_0[17:17], comp0_0[51:51], comp0_0[52:52], comp0_0[53:53]);
  C3 I1276 (simp9851_0[18:18], comp0_0[54:54], comp0_0[55:55], comp0_0[56:56]);
  C3 I1277 (simp9851_0[19:19], comp0_0[57:57], comp0_0[58:58], comp0_0[59:59]);
  C3 I1278 (simp9851_0[20:20], comp0_0[60:60], comp0_0[61:61], comp0_0[62:62]);
  C3 I1279 (simp9851_0[21:21], comp0_0[63:63], comp0_0[64:64], comp0_0[65:65]);
  C3 I1280 (simp9851_0[22:22], comp0_0[66:66], comp0_0[67:67], comp0_0[68:68]);
  C3 I1281 (simp9851_0[23:23], comp0_0[69:69], comp0_0[70:70], comp0_0[71:71]);
  C2 I1282 (simp9851_0[24:24], comp0_0[72:72], comp0_0[73:73]);
  C3 I1283 (simp9852_0[0:0], simp9851_0[0:0], simp9851_0[1:1], simp9851_0[2:2]);
  C3 I1284 (simp9852_0[1:1], simp9851_0[3:3], simp9851_0[4:4], simp9851_0[5:5]);
  C3 I1285 (simp9852_0[2:2], simp9851_0[6:6], simp9851_0[7:7], simp9851_0[8:8]);
  C3 I1286 (simp9852_0[3:3], simp9851_0[9:9], simp9851_0[10:10], simp9851_0[11:11]);
  C3 I1287 (simp9852_0[4:4], simp9851_0[12:12], simp9851_0[13:13], simp9851_0[14:14]);
  C3 I1288 (simp9852_0[5:5], simp9851_0[15:15], simp9851_0[16:16], simp9851_0[17:17]);
  C3 I1289 (simp9852_0[6:6], simp9851_0[18:18], simp9851_0[19:19], simp9851_0[20:20]);
  C3 I1290 (simp9852_0[7:7], simp9851_0[21:21], simp9851_0[22:22], simp9851_0[23:23]);
  BUFF I1291 (simp9852_0[8:8], simp9851_0[24:24]);
  C3 I1292 (simp9853_0[0:0], simp9852_0[0:0], simp9852_0[1:1], simp9852_0[2:2]);
  C3 I1293 (simp9853_0[1:1], simp9852_0[3:3], simp9852_0[4:4], simp9852_0[5:5]);
  C3 I1294 (simp9853_0[2:2], simp9852_0[6:6], simp9852_0[7:7], simp9852_0[8:8]);
  C3 I1295 (icomp_0, simp9853_0[0:0], simp9853_0[1:1], simp9853_0[2:2]);
  OR2 I1296 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I1297 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I1298 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I1299 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I1300 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I1301 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I1302 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  OR2 I1303 (comp1_0[7:7], i_1r0[7:7], i_1r1[7:7]);
  OR2 I1304 (comp1_0[8:8], i_1r0[8:8], i_1r1[8:8]);
  OR2 I1305 (comp1_0[9:9], i_1r0[9:9], i_1r1[9:9]);
  OR2 I1306 (comp1_0[10:10], i_1r0[10:10], i_1r1[10:10]);
  OR2 I1307 (comp1_0[11:11], i_1r0[11:11], i_1r1[11:11]);
  OR2 I1308 (comp1_0[12:12], i_1r0[12:12], i_1r1[12:12]);
  OR2 I1309 (comp1_0[13:13], i_1r0[13:13], i_1r1[13:13]);
  OR2 I1310 (comp1_0[14:14], i_1r0[14:14], i_1r1[14:14]);
  OR2 I1311 (comp1_0[15:15], i_1r0[15:15], i_1r1[15:15]);
  OR2 I1312 (comp1_0[16:16], i_1r0[16:16], i_1r1[16:16]);
  OR2 I1313 (comp1_0[17:17], i_1r0[17:17], i_1r1[17:17]);
  OR2 I1314 (comp1_0[18:18], i_1r0[18:18], i_1r1[18:18]);
  OR2 I1315 (comp1_0[19:19], i_1r0[19:19], i_1r1[19:19]);
  OR2 I1316 (comp1_0[20:20], i_1r0[20:20], i_1r1[20:20]);
  OR2 I1317 (comp1_0[21:21], i_1r0[21:21], i_1r1[21:21]);
  OR2 I1318 (comp1_0[22:22], i_1r0[22:22], i_1r1[22:22]);
  OR2 I1319 (comp1_0[23:23], i_1r0[23:23], i_1r1[23:23]);
  OR2 I1320 (comp1_0[24:24], i_1r0[24:24], i_1r1[24:24]);
  OR2 I1321 (comp1_0[25:25], i_1r0[25:25], i_1r1[25:25]);
  OR2 I1322 (comp1_0[26:26], i_1r0[26:26], i_1r1[26:26]);
  OR2 I1323 (comp1_0[27:27], i_1r0[27:27], i_1r1[27:27]);
  OR2 I1324 (comp1_0[28:28], i_1r0[28:28], i_1r1[28:28]);
  OR2 I1325 (comp1_0[29:29], i_1r0[29:29], i_1r1[29:29]);
  OR2 I1326 (comp1_0[30:30], i_1r0[30:30], i_1r1[30:30]);
  OR2 I1327 (comp1_0[31:31], i_1r0[31:31], i_1r1[31:31]);
  OR2 I1328 (comp1_0[32:32], i_1r0[32:32], i_1r1[32:32]);
  OR2 I1329 (comp1_0[33:33], i_1r0[33:33], i_1r1[33:33]);
  OR2 I1330 (comp1_0[34:34], i_1r0[34:34], i_1r1[34:34]);
  OR2 I1331 (comp1_0[35:35], i_1r0[35:35], i_1r1[35:35]);
  OR2 I1332 (comp1_0[36:36], i_1r0[36:36], i_1r1[36:36]);
  OR2 I1333 (comp1_0[37:37], i_1r0[37:37], i_1r1[37:37]);
  OR2 I1334 (comp1_0[38:38], i_1r0[38:38], i_1r1[38:38]);
  OR2 I1335 (comp1_0[39:39], i_1r0[39:39], i_1r1[39:39]);
  OR2 I1336 (comp1_0[40:40], i_1r0[40:40], i_1r1[40:40]);
  OR2 I1337 (comp1_0[41:41], i_1r0[41:41], i_1r1[41:41]);
  OR2 I1338 (comp1_0[42:42], i_1r0[42:42], i_1r1[42:42]);
  OR2 I1339 (comp1_0[43:43], i_1r0[43:43], i_1r1[43:43]);
  OR2 I1340 (comp1_0[44:44], i_1r0[44:44], i_1r1[44:44]);
  OR2 I1341 (comp1_0[45:45], i_1r0[45:45], i_1r1[45:45]);
  OR2 I1342 (comp1_0[46:46], i_1r0[46:46], i_1r1[46:46]);
  OR2 I1343 (comp1_0[47:47], i_1r0[47:47], i_1r1[47:47]);
  OR2 I1344 (comp1_0[48:48], i_1r0[48:48], i_1r1[48:48]);
  OR2 I1345 (comp1_0[49:49], i_1r0[49:49], i_1r1[49:49]);
  OR2 I1346 (comp1_0[50:50], i_1r0[50:50], i_1r1[50:50]);
  OR2 I1347 (comp1_0[51:51], i_1r0[51:51], i_1r1[51:51]);
  OR2 I1348 (comp1_0[52:52], i_1r0[52:52], i_1r1[52:52]);
  OR2 I1349 (comp1_0[53:53], i_1r0[53:53], i_1r1[53:53]);
  OR2 I1350 (comp1_0[54:54], i_1r0[54:54], i_1r1[54:54]);
  OR2 I1351 (comp1_0[55:55], i_1r0[55:55], i_1r1[55:55]);
  OR2 I1352 (comp1_0[56:56], i_1r0[56:56], i_1r1[56:56]);
  OR2 I1353 (comp1_0[57:57], i_1r0[57:57], i_1r1[57:57]);
  OR2 I1354 (comp1_0[58:58], i_1r0[58:58], i_1r1[58:58]);
  OR2 I1355 (comp1_0[59:59], i_1r0[59:59], i_1r1[59:59]);
  OR2 I1356 (comp1_0[60:60], i_1r0[60:60], i_1r1[60:60]);
  OR2 I1357 (comp1_0[61:61], i_1r0[61:61], i_1r1[61:61]);
  OR2 I1358 (comp1_0[62:62], i_1r0[62:62], i_1r1[62:62]);
  OR2 I1359 (comp1_0[63:63], i_1r0[63:63], i_1r1[63:63]);
  OR2 I1360 (comp1_0[64:64], i_1r0[64:64], i_1r1[64:64]);
  OR2 I1361 (comp1_0[65:65], i_1r0[65:65], i_1r1[65:65]);
  OR2 I1362 (comp1_0[66:66], i_1r0[66:66], i_1r1[66:66]);
  OR2 I1363 (comp1_0[67:67], i_1r0[67:67], i_1r1[67:67]);
  OR2 I1364 (comp1_0[68:68], i_1r0[68:68], i_1r1[68:68]);
  OR2 I1365 (comp1_0[69:69], i_1r0[69:69], i_1r1[69:69]);
  OR2 I1366 (comp1_0[70:70], i_1r0[70:70], i_1r1[70:70]);
  OR2 I1367 (comp1_0[71:71], i_1r0[71:71], i_1r1[71:71]);
  OR2 I1368 (comp1_0[72:72], i_1r0[72:72], i_1r1[72:72]);
  OR2 I1369 (comp1_0[73:73], i_1r0[73:73], i_1r1[73:73]);
  C3 I1370 (simp10611_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I1371 (simp10611_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  C3 I1372 (simp10611_0[2:2], comp1_0[6:6], comp1_0[7:7], comp1_0[8:8]);
  C3 I1373 (simp10611_0[3:3], comp1_0[9:9], comp1_0[10:10], comp1_0[11:11]);
  C3 I1374 (simp10611_0[4:4], comp1_0[12:12], comp1_0[13:13], comp1_0[14:14]);
  C3 I1375 (simp10611_0[5:5], comp1_0[15:15], comp1_0[16:16], comp1_0[17:17]);
  C3 I1376 (simp10611_0[6:6], comp1_0[18:18], comp1_0[19:19], comp1_0[20:20]);
  C3 I1377 (simp10611_0[7:7], comp1_0[21:21], comp1_0[22:22], comp1_0[23:23]);
  C3 I1378 (simp10611_0[8:8], comp1_0[24:24], comp1_0[25:25], comp1_0[26:26]);
  C3 I1379 (simp10611_0[9:9], comp1_0[27:27], comp1_0[28:28], comp1_0[29:29]);
  C3 I1380 (simp10611_0[10:10], comp1_0[30:30], comp1_0[31:31], comp1_0[32:32]);
  C3 I1381 (simp10611_0[11:11], comp1_0[33:33], comp1_0[34:34], comp1_0[35:35]);
  C3 I1382 (simp10611_0[12:12], comp1_0[36:36], comp1_0[37:37], comp1_0[38:38]);
  C3 I1383 (simp10611_0[13:13], comp1_0[39:39], comp1_0[40:40], comp1_0[41:41]);
  C3 I1384 (simp10611_0[14:14], comp1_0[42:42], comp1_0[43:43], comp1_0[44:44]);
  C3 I1385 (simp10611_0[15:15], comp1_0[45:45], comp1_0[46:46], comp1_0[47:47]);
  C3 I1386 (simp10611_0[16:16], comp1_0[48:48], comp1_0[49:49], comp1_0[50:50]);
  C3 I1387 (simp10611_0[17:17], comp1_0[51:51], comp1_0[52:52], comp1_0[53:53]);
  C3 I1388 (simp10611_0[18:18], comp1_0[54:54], comp1_0[55:55], comp1_0[56:56]);
  C3 I1389 (simp10611_0[19:19], comp1_0[57:57], comp1_0[58:58], comp1_0[59:59]);
  C3 I1390 (simp10611_0[20:20], comp1_0[60:60], comp1_0[61:61], comp1_0[62:62]);
  C3 I1391 (simp10611_0[21:21], comp1_0[63:63], comp1_0[64:64], comp1_0[65:65]);
  C3 I1392 (simp10611_0[22:22], comp1_0[66:66], comp1_0[67:67], comp1_0[68:68]);
  C3 I1393 (simp10611_0[23:23], comp1_0[69:69], comp1_0[70:70], comp1_0[71:71]);
  C2 I1394 (simp10611_0[24:24], comp1_0[72:72], comp1_0[73:73]);
  C3 I1395 (simp10612_0[0:0], simp10611_0[0:0], simp10611_0[1:1], simp10611_0[2:2]);
  C3 I1396 (simp10612_0[1:1], simp10611_0[3:3], simp10611_0[4:4], simp10611_0[5:5]);
  C3 I1397 (simp10612_0[2:2], simp10611_0[6:6], simp10611_0[7:7], simp10611_0[8:8]);
  C3 I1398 (simp10612_0[3:3], simp10611_0[9:9], simp10611_0[10:10], simp10611_0[11:11]);
  C3 I1399 (simp10612_0[4:4], simp10611_0[12:12], simp10611_0[13:13], simp10611_0[14:14]);
  C3 I1400 (simp10612_0[5:5], simp10611_0[15:15], simp10611_0[16:16], simp10611_0[17:17]);
  C3 I1401 (simp10612_0[6:6], simp10611_0[18:18], simp10611_0[19:19], simp10611_0[20:20]);
  C3 I1402 (simp10612_0[7:7], simp10611_0[21:21], simp10611_0[22:22], simp10611_0[23:23]);
  BUFF I1403 (simp10612_0[8:8], simp10611_0[24:24]);
  C3 I1404 (simp10613_0[0:0], simp10612_0[0:0], simp10612_0[1:1], simp10612_0[2:2]);
  C3 I1405 (simp10613_0[1:1], simp10612_0[3:3], simp10612_0[4:4], simp10612_0[5:5]);
  C3 I1406 (simp10613_0[2:2], simp10612_0[6:6], simp10612_0[7:7], simp10612_0[8:8]);
  C3 I1407 (icomp_1, simp10613_0[0:0], simp10613_0[1:1], simp10613_0[2:2]);
  OR2 I1408 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I1409 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I1410 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2 I1411 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  OR2 I1412 (comp2_0[4:4], i_2r0[4:4], i_2r1[4:4]);
  OR2 I1413 (comp2_0[5:5], i_2r0[5:5], i_2r1[5:5]);
  OR2 I1414 (comp2_0[6:6], i_2r0[6:6], i_2r1[6:6]);
  OR2 I1415 (comp2_0[7:7], i_2r0[7:7], i_2r1[7:7]);
  OR2 I1416 (comp2_0[8:8], i_2r0[8:8], i_2r1[8:8]);
  OR2 I1417 (comp2_0[9:9], i_2r0[9:9], i_2r1[9:9]);
  OR2 I1418 (comp2_0[10:10], i_2r0[10:10], i_2r1[10:10]);
  OR2 I1419 (comp2_0[11:11], i_2r0[11:11], i_2r1[11:11]);
  OR2 I1420 (comp2_0[12:12], i_2r0[12:12], i_2r1[12:12]);
  OR2 I1421 (comp2_0[13:13], i_2r0[13:13], i_2r1[13:13]);
  OR2 I1422 (comp2_0[14:14], i_2r0[14:14], i_2r1[14:14]);
  OR2 I1423 (comp2_0[15:15], i_2r0[15:15], i_2r1[15:15]);
  OR2 I1424 (comp2_0[16:16], i_2r0[16:16], i_2r1[16:16]);
  OR2 I1425 (comp2_0[17:17], i_2r0[17:17], i_2r1[17:17]);
  OR2 I1426 (comp2_0[18:18], i_2r0[18:18], i_2r1[18:18]);
  OR2 I1427 (comp2_0[19:19], i_2r0[19:19], i_2r1[19:19]);
  OR2 I1428 (comp2_0[20:20], i_2r0[20:20], i_2r1[20:20]);
  OR2 I1429 (comp2_0[21:21], i_2r0[21:21], i_2r1[21:21]);
  OR2 I1430 (comp2_0[22:22], i_2r0[22:22], i_2r1[22:22]);
  OR2 I1431 (comp2_0[23:23], i_2r0[23:23], i_2r1[23:23]);
  OR2 I1432 (comp2_0[24:24], i_2r0[24:24], i_2r1[24:24]);
  OR2 I1433 (comp2_0[25:25], i_2r0[25:25], i_2r1[25:25]);
  OR2 I1434 (comp2_0[26:26], i_2r0[26:26], i_2r1[26:26]);
  OR2 I1435 (comp2_0[27:27], i_2r0[27:27], i_2r1[27:27]);
  OR2 I1436 (comp2_0[28:28], i_2r0[28:28], i_2r1[28:28]);
  OR2 I1437 (comp2_0[29:29], i_2r0[29:29], i_2r1[29:29]);
  OR2 I1438 (comp2_0[30:30], i_2r0[30:30], i_2r1[30:30]);
  OR2 I1439 (comp2_0[31:31], i_2r0[31:31], i_2r1[31:31]);
  OR2 I1440 (comp2_0[32:32], i_2r0[32:32], i_2r1[32:32]);
  OR2 I1441 (comp2_0[33:33], i_2r0[33:33], i_2r1[33:33]);
  OR2 I1442 (comp2_0[34:34], i_2r0[34:34], i_2r1[34:34]);
  OR2 I1443 (comp2_0[35:35], i_2r0[35:35], i_2r1[35:35]);
  OR2 I1444 (comp2_0[36:36], i_2r0[36:36], i_2r1[36:36]);
  OR2 I1445 (comp2_0[37:37], i_2r0[37:37], i_2r1[37:37]);
  OR2 I1446 (comp2_0[38:38], i_2r0[38:38], i_2r1[38:38]);
  OR2 I1447 (comp2_0[39:39], i_2r0[39:39], i_2r1[39:39]);
  OR2 I1448 (comp2_0[40:40], i_2r0[40:40], i_2r1[40:40]);
  OR2 I1449 (comp2_0[41:41], i_2r0[41:41], i_2r1[41:41]);
  OR2 I1450 (comp2_0[42:42], i_2r0[42:42], i_2r1[42:42]);
  OR2 I1451 (comp2_0[43:43], i_2r0[43:43], i_2r1[43:43]);
  OR2 I1452 (comp2_0[44:44], i_2r0[44:44], i_2r1[44:44]);
  OR2 I1453 (comp2_0[45:45], i_2r0[45:45], i_2r1[45:45]);
  OR2 I1454 (comp2_0[46:46], i_2r0[46:46], i_2r1[46:46]);
  OR2 I1455 (comp2_0[47:47], i_2r0[47:47], i_2r1[47:47]);
  OR2 I1456 (comp2_0[48:48], i_2r0[48:48], i_2r1[48:48]);
  OR2 I1457 (comp2_0[49:49], i_2r0[49:49], i_2r1[49:49]);
  OR2 I1458 (comp2_0[50:50], i_2r0[50:50], i_2r1[50:50]);
  OR2 I1459 (comp2_0[51:51], i_2r0[51:51], i_2r1[51:51]);
  OR2 I1460 (comp2_0[52:52], i_2r0[52:52], i_2r1[52:52]);
  OR2 I1461 (comp2_0[53:53], i_2r0[53:53], i_2r1[53:53]);
  OR2 I1462 (comp2_0[54:54], i_2r0[54:54], i_2r1[54:54]);
  OR2 I1463 (comp2_0[55:55], i_2r0[55:55], i_2r1[55:55]);
  OR2 I1464 (comp2_0[56:56], i_2r0[56:56], i_2r1[56:56]);
  OR2 I1465 (comp2_0[57:57], i_2r0[57:57], i_2r1[57:57]);
  OR2 I1466 (comp2_0[58:58], i_2r0[58:58], i_2r1[58:58]);
  OR2 I1467 (comp2_0[59:59], i_2r0[59:59], i_2r1[59:59]);
  OR2 I1468 (comp2_0[60:60], i_2r0[60:60], i_2r1[60:60]);
  OR2 I1469 (comp2_0[61:61], i_2r0[61:61], i_2r1[61:61]);
  OR2 I1470 (comp2_0[62:62], i_2r0[62:62], i_2r1[62:62]);
  OR2 I1471 (comp2_0[63:63], i_2r0[63:63], i_2r1[63:63]);
  OR2 I1472 (comp2_0[64:64], i_2r0[64:64], i_2r1[64:64]);
  OR2 I1473 (comp2_0[65:65], i_2r0[65:65], i_2r1[65:65]);
  OR2 I1474 (comp2_0[66:66], i_2r0[66:66], i_2r1[66:66]);
  OR2 I1475 (comp2_0[67:67], i_2r0[67:67], i_2r1[67:67]);
  OR2 I1476 (comp2_0[68:68], i_2r0[68:68], i_2r1[68:68]);
  OR2 I1477 (comp2_0[69:69], i_2r0[69:69], i_2r1[69:69]);
  OR2 I1478 (comp2_0[70:70], i_2r0[70:70], i_2r1[70:70]);
  OR2 I1479 (comp2_0[71:71], i_2r0[71:71], i_2r1[71:71]);
  OR2 I1480 (comp2_0[72:72], i_2r0[72:72], i_2r1[72:72]);
  OR2 I1481 (comp2_0[73:73], i_2r0[73:73], i_2r1[73:73]);
  C3 I1482 (simp11371_0[0:0], comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C3 I1483 (simp11371_0[1:1], comp2_0[3:3], comp2_0[4:4], comp2_0[5:5]);
  C3 I1484 (simp11371_0[2:2], comp2_0[6:6], comp2_0[7:7], comp2_0[8:8]);
  C3 I1485 (simp11371_0[3:3], comp2_0[9:9], comp2_0[10:10], comp2_0[11:11]);
  C3 I1486 (simp11371_0[4:4], comp2_0[12:12], comp2_0[13:13], comp2_0[14:14]);
  C3 I1487 (simp11371_0[5:5], comp2_0[15:15], comp2_0[16:16], comp2_0[17:17]);
  C3 I1488 (simp11371_0[6:6], comp2_0[18:18], comp2_0[19:19], comp2_0[20:20]);
  C3 I1489 (simp11371_0[7:7], comp2_0[21:21], comp2_0[22:22], comp2_0[23:23]);
  C3 I1490 (simp11371_0[8:8], comp2_0[24:24], comp2_0[25:25], comp2_0[26:26]);
  C3 I1491 (simp11371_0[9:9], comp2_0[27:27], comp2_0[28:28], comp2_0[29:29]);
  C3 I1492 (simp11371_0[10:10], comp2_0[30:30], comp2_0[31:31], comp2_0[32:32]);
  C3 I1493 (simp11371_0[11:11], comp2_0[33:33], comp2_0[34:34], comp2_0[35:35]);
  C3 I1494 (simp11371_0[12:12], comp2_0[36:36], comp2_0[37:37], comp2_0[38:38]);
  C3 I1495 (simp11371_0[13:13], comp2_0[39:39], comp2_0[40:40], comp2_0[41:41]);
  C3 I1496 (simp11371_0[14:14], comp2_0[42:42], comp2_0[43:43], comp2_0[44:44]);
  C3 I1497 (simp11371_0[15:15], comp2_0[45:45], comp2_0[46:46], comp2_0[47:47]);
  C3 I1498 (simp11371_0[16:16], comp2_0[48:48], comp2_0[49:49], comp2_0[50:50]);
  C3 I1499 (simp11371_0[17:17], comp2_0[51:51], comp2_0[52:52], comp2_0[53:53]);
  C3 I1500 (simp11371_0[18:18], comp2_0[54:54], comp2_0[55:55], comp2_0[56:56]);
  C3 I1501 (simp11371_0[19:19], comp2_0[57:57], comp2_0[58:58], comp2_0[59:59]);
  C3 I1502 (simp11371_0[20:20], comp2_0[60:60], comp2_0[61:61], comp2_0[62:62]);
  C3 I1503 (simp11371_0[21:21], comp2_0[63:63], comp2_0[64:64], comp2_0[65:65]);
  C3 I1504 (simp11371_0[22:22], comp2_0[66:66], comp2_0[67:67], comp2_0[68:68]);
  C3 I1505 (simp11371_0[23:23], comp2_0[69:69], comp2_0[70:70], comp2_0[71:71]);
  C2 I1506 (simp11371_0[24:24], comp2_0[72:72], comp2_0[73:73]);
  C3 I1507 (simp11372_0[0:0], simp11371_0[0:0], simp11371_0[1:1], simp11371_0[2:2]);
  C3 I1508 (simp11372_0[1:1], simp11371_0[3:3], simp11371_0[4:4], simp11371_0[5:5]);
  C3 I1509 (simp11372_0[2:2], simp11371_0[6:6], simp11371_0[7:7], simp11371_0[8:8]);
  C3 I1510 (simp11372_0[3:3], simp11371_0[9:9], simp11371_0[10:10], simp11371_0[11:11]);
  C3 I1511 (simp11372_0[4:4], simp11371_0[12:12], simp11371_0[13:13], simp11371_0[14:14]);
  C3 I1512 (simp11372_0[5:5], simp11371_0[15:15], simp11371_0[16:16], simp11371_0[17:17]);
  C3 I1513 (simp11372_0[6:6], simp11371_0[18:18], simp11371_0[19:19], simp11371_0[20:20]);
  C3 I1514 (simp11372_0[7:7], simp11371_0[21:21], simp11371_0[22:22], simp11371_0[23:23]);
  BUFF I1515 (simp11372_0[8:8], simp11371_0[24:24]);
  C3 I1516 (simp11373_0[0:0], simp11372_0[0:0], simp11372_0[1:1], simp11372_0[2:2]);
  C3 I1517 (simp11373_0[1:1], simp11372_0[3:3], simp11372_0[4:4], simp11372_0[5:5]);
  C3 I1518 (simp11373_0[2:2], simp11372_0[6:6], simp11372_0[7:7], simp11372_0[8:8]);
  C3 I1519 (icomp_2, simp11373_0[0:0], simp11373_0[1:1], simp11373_0[2:2]);
  OR2 I1520 (comp3_0[0:0], i_3r0[0:0], i_3r1[0:0]);
  OR2 I1521 (comp3_0[1:1], i_3r0[1:1], i_3r1[1:1]);
  OR2 I1522 (comp3_0[2:2], i_3r0[2:2], i_3r1[2:2]);
  OR2 I1523 (comp3_0[3:3], i_3r0[3:3], i_3r1[3:3]);
  OR2 I1524 (comp3_0[4:4], i_3r0[4:4], i_3r1[4:4]);
  OR2 I1525 (comp3_0[5:5], i_3r0[5:5], i_3r1[5:5]);
  OR2 I1526 (comp3_0[6:6], i_3r0[6:6], i_3r1[6:6]);
  OR2 I1527 (comp3_0[7:7], i_3r0[7:7], i_3r1[7:7]);
  OR2 I1528 (comp3_0[8:8], i_3r0[8:8], i_3r1[8:8]);
  OR2 I1529 (comp3_0[9:9], i_3r0[9:9], i_3r1[9:9]);
  OR2 I1530 (comp3_0[10:10], i_3r0[10:10], i_3r1[10:10]);
  OR2 I1531 (comp3_0[11:11], i_3r0[11:11], i_3r1[11:11]);
  OR2 I1532 (comp3_0[12:12], i_3r0[12:12], i_3r1[12:12]);
  OR2 I1533 (comp3_0[13:13], i_3r0[13:13], i_3r1[13:13]);
  OR2 I1534 (comp3_0[14:14], i_3r0[14:14], i_3r1[14:14]);
  OR2 I1535 (comp3_0[15:15], i_3r0[15:15], i_3r1[15:15]);
  OR2 I1536 (comp3_0[16:16], i_3r0[16:16], i_3r1[16:16]);
  OR2 I1537 (comp3_0[17:17], i_3r0[17:17], i_3r1[17:17]);
  OR2 I1538 (comp3_0[18:18], i_3r0[18:18], i_3r1[18:18]);
  OR2 I1539 (comp3_0[19:19], i_3r0[19:19], i_3r1[19:19]);
  OR2 I1540 (comp3_0[20:20], i_3r0[20:20], i_3r1[20:20]);
  OR2 I1541 (comp3_0[21:21], i_3r0[21:21], i_3r1[21:21]);
  OR2 I1542 (comp3_0[22:22], i_3r0[22:22], i_3r1[22:22]);
  OR2 I1543 (comp3_0[23:23], i_3r0[23:23], i_3r1[23:23]);
  OR2 I1544 (comp3_0[24:24], i_3r0[24:24], i_3r1[24:24]);
  OR2 I1545 (comp3_0[25:25], i_3r0[25:25], i_3r1[25:25]);
  OR2 I1546 (comp3_0[26:26], i_3r0[26:26], i_3r1[26:26]);
  OR2 I1547 (comp3_0[27:27], i_3r0[27:27], i_3r1[27:27]);
  OR2 I1548 (comp3_0[28:28], i_3r0[28:28], i_3r1[28:28]);
  OR2 I1549 (comp3_0[29:29], i_3r0[29:29], i_3r1[29:29]);
  OR2 I1550 (comp3_0[30:30], i_3r0[30:30], i_3r1[30:30]);
  OR2 I1551 (comp3_0[31:31], i_3r0[31:31], i_3r1[31:31]);
  OR2 I1552 (comp3_0[32:32], i_3r0[32:32], i_3r1[32:32]);
  OR2 I1553 (comp3_0[33:33], i_3r0[33:33], i_3r1[33:33]);
  OR2 I1554 (comp3_0[34:34], i_3r0[34:34], i_3r1[34:34]);
  OR2 I1555 (comp3_0[35:35], i_3r0[35:35], i_3r1[35:35]);
  OR2 I1556 (comp3_0[36:36], i_3r0[36:36], i_3r1[36:36]);
  OR2 I1557 (comp3_0[37:37], i_3r0[37:37], i_3r1[37:37]);
  OR2 I1558 (comp3_0[38:38], i_3r0[38:38], i_3r1[38:38]);
  OR2 I1559 (comp3_0[39:39], i_3r0[39:39], i_3r1[39:39]);
  OR2 I1560 (comp3_0[40:40], i_3r0[40:40], i_3r1[40:40]);
  OR2 I1561 (comp3_0[41:41], i_3r0[41:41], i_3r1[41:41]);
  OR2 I1562 (comp3_0[42:42], i_3r0[42:42], i_3r1[42:42]);
  OR2 I1563 (comp3_0[43:43], i_3r0[43:43], i_3r1[43:43]);
  OR2 I1564 (comp3_0[44:44], i_3r0[44:44], i_3r1[44:44]);
  OR2 I1565 (comp3_0[45:45], i_3r0[45:45], i_3r1[45:45]);
  OR2 I1566 (comp3_0[46:46], i_3r0[46:46], i_3r1[46:46]);
  OR2 I1567 (comp3_0[47:47], i_3r0[47:47], i_3r1[47:47]);
  OR2 I1568 (comp3_0[48:48], i_3r0[48:48], i_3r1[48:48]);
  OR2 I1569 (comp3_0[49:49], i_3r0[49:49], i_3r1[49:49]);
  OR2 I1570 (comp3_0[50:50], i_3r0[50:50], i_3r1[50:50]);
  OR2 I1571 (comp3_0[51:51], i_3r0[51:51], i_3r1[51:51]);
  OR2 I1572 (comp3_0[52:52], i_3r0[52:52], i_3r1[52:52]);
  OR2 I1573 (comp3_0[53:53], i_3r0[53:53], i_3r1[53:53]);
  OR2 I1574 (comp3_0[54:54], i_3r0[54:54], i_3r1[54:54]);
  OR2 I1575 (comp3_0[55:55], i_3r0[55:55], i_3r1[55:55]);
  OR2 I1576 (comp3_0[56:56], i_3r0[56:56], i_3r1[56:56]);
  OR2 I1577 (comp3_0[57:57], i_3r0[57:57], i_3r1[57:57]);
  OR2 I1578 (comp3_0[58:58], i_3r0[58:58], i_3r1[58:58]);
  OR2 I1579 (comp3_0[59:59], i_3r0[59:59], i_3r1[59:59]);
  OR2 I1580 (comp3_0[60:60], i_3r0[60:60], i_3r1[60:60]);
  OR2 I1581 (comp3_0[61:61], i_3r0[61:61], i_3r1[61:61]);
  OR2 I1582 (comp3_0[62:62], i_3r0[62:62], i_3r1[62:62]);
  OR2 I1583 (comp3_0[63:63], i_3r0[63:63], i_3r1[63:63]);
  OR2 I1584 (comp3_0[64:64], i_3r0[64:64], i_3r1[64:64]);
  OR2 I1585 (comp3_0[65:65], i_3r0[65:65], i_3r1[65:65]);
  OR2 I1586 (comp3_0[66:66], i_3r0[66:66], i_3r1[66:66]);
  OR2 I1587 (comp3_0[67:67], i_3r0[67:67], i_3r1[67:67]);
  OR2 I1588 (comp3_0[68:68], i_3r0[68:68], i_3r1[68:68]);
  OR2 I1589 (comp3_0[69:69], i_3r0[69:69], i_3r1[69:69]);
  OR2 I1590 (comp3_0[70:70], i_3r0[70:70], i_3r1[70:70]);
  OR2 I1591 (comp3_0[71:71], i_3r0[71:71], i_3r1[71:71]);
  OR2 I1592 (comp3_0[72:72], i_3r0[72:72], i_3r1[72:72]);
  OR2 I1593 (comp3_0[73:73], i_3r0[73:73], i_3r1[73:73]);
  C3 I1594 (simp12131_0[0:0], comp3_0[0:0], comp3_0[1:1], comp3_0[2:2]);
  C3 I1595 (simp12131_0[1:1], comp3_0[3:3], comp3_0[4:4], comp3_0[5:5]);
  C3 I1596 (simp12131_0[2:2], comp3_0[6:6], comp3_0[7:7], comp3_0[8:8]);
  C3 I1597 (simp12131_0[3:3], comp3_0[9:9], comp3_0[10:10], comp3_0[11:11]);
  C3 I1598 (simp12131_0[4:4], comp3_0[12:12], comp3_0[13:13], comp3_0[14:14]);
  C3 I1599 (simp12131_0[5:5], comp3_0[15:15], comp3_0[16:16], comp3_0[17:17]);
  C3 I1600 (simp12131_0[6:6], comp3_0[18:18], comp3_0[19:19], comp3_0[20:20]);
  C3 I1601 (simp12131_0[7:7], comp3_0[21:21], comp3_0[22:22], comp3_0[23:23]);
  C3 I1602 (simp12131_0[8:8], comp3_0[24:24], comp3_0[25:25], comp3_0[26:26]);
  C3 I1603 (simp12131_0[9:9], comp3_0[27:27], comp3_0[28:28], comp3_0[29:29]);
  C3 I1604 (simp12131_0[10:10], comp3_0[30:30], comp3_0[31:31], comp3_0[32:32]);
  C3 I1605 (simp12131_0[11:11], comp3_0[33:33], comp3_0[34:34], comp3_0[35:35]);
  C3 I1606 (simp12131_0[12:12], comp3_0[36:36], comp3_0[37:37], comp3_0[38:38]);
  C3 I1607 (simp12131_0[13:13], comp3_0[39:39], comp3_0[40:40], comp3_0[41:41]);
  C3 I1608 (simp12131_0[14:14], comp3_0[42:42], comp3_0[43:43], comp3_0[44:44]);
  C3 I1609 (simp12131_0[15:15], comp3_0[45:45], comp3_0[46:46], comp3_0[47:47]);
  C3 I1610 (simp12131_0[16:16], comp3_0[48:48], comp3_0[49:49], comp3_0[50:50]);
  C3 I1611 (simp12131_0[17:17], comp3_0[51:51], comp3_0[52:52], comp3_0[53:53]);
  C3 I1612 (simp12131_0[18:18], comp3_0[54:54], comp3_0[55:55], comp3_0[56:56]);
  C3 I1613 (simp12131_0[19:19], comp3_0[57:57], comp3_0[58:58], comp3_0[59:59]);
  C3 I1614 (simp12131_0[20:20], comp3_0[60:60], comp3_0[61:61], comp3_0[62:62]);
  C3 I1615 (simp12131_0[21:21], comp3_0[63:63], comp3_0[64:64], comp3_0[65:65]);
  C3 I1616 (simp12131_0[22:22], comp3_0[66:66], comp3_0[67:67], comp3_0[68:68]);
  C3 I1617 (simp12131_0[23:23], comp3_0[69:69], comp3_0[70:70], comp3_0[71:71]);
  C2 I1618 (simp12131_0[24:24], comp3_0[72:72], comp3_0[73:73]);
  C3 I1619 (simp12132_0[0:0], simp12131_0[0:0], simp12131_0[1:1], simp12131_0[2:2]);
  C3 I1620 (simp12132_0[1:1], simp12131_0[3:3], simp12131_0[4:4], simp12131_0[5:5]);
  C3 I1621 (simp12132_0[2:2], simp12131_0[6:6], simp12131_0[7:7], simp12131_0[8:8]);
  C3 I1622 (simp12132_0[3:3], simp12131_0[9:9], simp12131_0[10:10], simp12131_0[11:11]);
  C3 I1623 (simp12132_0[4:4], simp12131_0[12:12], simp12131_0[13:13], simp12131_0[14:14]);
  C3 I1624 (simp12132_0[5:5], simp12131_0[15:15], simp12131_0[16:16], simp12131_0[17:17]);
  C3 I1625 (simp12132_0[6:6], simp12131_0[18:18], simp12131_0[19:19], simp12131_0[20:20]);
  C3 I1626 (simp12132_0[7:7], simp12131_0[21:21], simp12131_0[22:22], simp12131_0[23:23]);
  BUFF I1627 (simp12132_0[8:8], simp12131_0[24:24]);
  C3 I1628 (simp12133_0[0:0], simp12132_0[0:0], simp12132_0[1:1], simp12132_0[2:2]);
  C3 I1629 (simp12133_0[1:1], simp12132_0[3:3], simp12132_0[4:4], simp12132_0[5:5]);
  C3 I1630 (simp12133_0[2:2], simp12132_0[6:6], simp12132_0[7:7], simp12132_0[8:8]);
  C3 I1631 (icomp_3, simp12133_0[0:0], simp12133_0[1:1], simp12133_0[2:2]);
  OR2 I1632 (comp4_0[0:0], i_4r0[0:0], i_4r1[0:0]);
  OR2 I1633 (comp4_0[1:1], i_4r0[1:1], i_4r1[1:1]);
  OR2 I1634 (comp4_0[2:2], i_4r0[2:2], i_4r1[2:2]);
  OR2 I1635 (comp4_0[3:3], i_4r0[3:3], i_4r1[3:3]);
  OR2 I1636 (comp4_0[4:4], i_4r0[4:4], i_4r1[4:4]);
  OR2 I1637 (comp4_0[5:5], i_4r0[5:5], i_4r1[5:5]);
  OR2 I1638 (comp4_0[6:6], i_4r0[6:6], i_4r1[6:6]);
  OR2 I1639 (comp4_0[7:7], i_4r0[7:7], i_4r1[7:7]);
  OR2 I1640 (comp4_0[8:8], i_4r0[8:8], i_4r1[8:8]);
  OR2 I1641 (comp4_0[9:9], i_4r0[9:9], i_4r1[9:9]);
  OR2 I1642 (comp4_0[10:10], i_4r0[10:10], i_4r1[10:10]);
  OR2 I1643 (comp4_0[11:11], i_4r0[11:11], i_4r1[11:11]);
  OR2 I1644 (comp4_0[12:12], i_4r0[12:12], i_4r1[12:12]);
  OR2 I1645 (comp4_0[13:13], i_4r0[13:13], i_4r1[13:13]);
  OR2 I1646 (comp4_0[14:14], i_4r0[14:14], i_4r1[14:14]);
  OR2 I1647 (comp4_0[15:15], i_4r0[15:15], i_4r1[15:15]);
  OR2 I1648 (comp4_0[16:16], i_4r0[16:16], i_4r1[16:16]);
  OR2 I1649 (comp4_0[17:17], i_4r0[17:17], i_4r1[17:17]);
  OR2 I1650 (comp4_0[18:18], i_4r0[18:18], i_4r1[18:18]);
  OR2 I1651 (comp4_0[19:19], i_4r0[19:19], i_4r1[19:19]);
  OR2 I1652 (comp4_0[20:20], i_4r0[20:20], i_4r1[20:20]);
  OR2 I1653 (comp4_0[21:21], i_4r0[21:21], i_4r1[21:21]);
  OR2 I1654 (comp4_0[22:22], i_4r0[22:22], i_4r1[22:22]);
  OR2 I1655 (comp4_0[23:23], i_4r0[23:23], i_4r1[23:23]);
  OR2 I1656 (comp4_0[24:24], i_4r0[24:24], i_4r1[24:24]);
  OR2 I1657 (comp4_0[25:25], i_4r0[25:25], i_4r1[25:25]);
  OR2 I1658 (comp4_0[26:26], i_4r0[26:26], i_4r1[26:26]);
  OR2 I1659 (comp4_0[27:27], i_4r0[27:27], i_4r1[27:27]);
  OR2 I1660 (comp4_0[28:28], i_4r0[28:28], i_4r1[28:28]);
  OR2 I1661 (comp4_0[29:29], i_4r0[29:29], i_4r1[29:29]);
  OR2 I1662 (comp4_0[30:30], i_4r0[30:30], i_4r1[30:30]);
  OR2 I1663 (comp4_0[31:31], i_4r0[31:31], i_4r1[31:31]);
  OR2 I1664 (comp4_0[32:32], i_4r0[32:32], i_4r1[32:32]);
  OR2 I1665 (comp4_0[33:33], i_4r0[33:33], i_4r1[33:33]);
  OR2 I1666 (comp4_0[34:34], i_4r0[34:34], i_4r1[34:34]);
  OR2 I1667 (comp4_0[35:35], i_4r0[35:35], i_4r1[35:35]);
  OR2 I1668 (comp4_0[36:36], i_4r0[36:36], i_4r1[36:36]);
  OR2 I1669 (comp4_0[37:37], i_4r0[37:37], i_4r1[37:37]);
  OR2 I1670 (comp4_0[38:38], i_4r0[38:38], i_4r1[38:38]);
  OR2 I1671 (comp4_0[39:39], i_4r0[39:39], i_4r1[39:39]);
  OR2 I1672 (comp4_0[40:40], i_4r0[40:40], i_4r1[40:40]);
  OR2 I1673 (comp4_0[41:41], i_4r0[41:41], i_4r1[41:41]);
  OR2 I1674 (comp4_0[42:42], i_4r0[42:42], i_4r1[42:42]);
  OR2 I1675 (comp4_0[43:43], i_4r0[43:43], i_4r1[43:43]);
  OR2 I1676 (comp4_0[44:44], i_4r0[44:44], i_4r1[44:44]);
  OR2 I1677 (comp4_0[45:45], i_4r0[45:45], i_4r1[45:45]);
  OR2 I1678 (comp4_0[46:46], i_4r0[46:46], i_4r1[46:46]);
  OR2 I1679 (comp4_0[47:47], i_4r0[47:47], i_4r1[47:47]);
  OR2 I1680 (comp4_0[48:48], i_4r0[48:48], i_4r1[48:48]);
  OR2 I1681 (comp4_0[49:49], i_4r0[49:49], i_4r1[49:49]);
  OR2 I1682 (comp4_0[50:50], i_4r0[50:50], i_4r1[50:50]);
  OR2 I1683 (comp4_0[51:51], i_4r0[51:51], i_4r1[51:51]);
  OR2 I1684 (comp4_0[52:52], i_4r0[52:52], i_4r1[52:52]);
  OR2 I1685 (comp4_0[53:53], i_4r0[53:53], i_4r1[53:53]);
  OR2 I1686 (comp4_0[54:54], i_4r0[54:54], i_4r1[54:54]);
  OR2 I1687 (comp4_0[55:55], i_4r0[55:55], i_4r1[55:55]);
  OR2 I1688 (comp4_0[56:56], i_4r0[56:56], i_4r1[56:56]);
  OR2 I1689 (comp4_0[57:57], i_4r0[57:57], i_4r1[57:57]);
  OR2 I1690 (comp4_0[58:58], i_4r0[58:58], i_4r1[58:58]);
  OR2 I1691 (comp4_0[59:59], i_4r0[59:59], i_4r1[59:59]);
  OR2 I1692 (comp4_0[60:60], i_4r0[60:60], i_4r1[60:60]);
  OR2 I1693 (comp4_0[61:61], i_4r0[61:61], i_4r1[61:61]);
  OR2 I1694 (comp4_0[62:62], i_4r0[62:62], i_4r1[62:62]);
  OR2 I1695 (comp4_0[63:63], i_4r0[63:63], i_4r1[63:63]);
  OR2 I1696 (comp4_0[64:64], i_4r0[64:64], i_4r1[64:64]);
  OR2 I1697 (comp4_0[65:65], i_4r0[65:65], i_4r1[65:65]);
  OR2 I1698 (comp4_0[66:66], i_4r0[66:66], i_4r1[66:66]);
  OR2 I1699 (comp4_0[67:67], i_4r0[67:67], i_4r1[67:67]);
  OR2 I1700 (comp4_0[68:68], i_4r0[68:68], i_4r1[68:68]);
  OR2 I1701 (comp4_0[69:69], i_4r0[69:69], i_4r1[69:69]);
  OR2 I1702 (comp4_0[70:70], i_4r0[70:70], i_4r1[70:70]);
  OR2 I1703 (comp4_0[71:71], i_4r0[71:71], i_4r1[71:71]);
  OR2 I1704 (comp4_0[72:72], i_4r0[72:72], i_4r1[72:72]);
  OR2 I1705 (comp4_0[73:73], i_4r0[73:73], i_4r1[73:73]);
  C3 I1706 (simp12891_0[0:0], comp4_0[0:0], comp4_0[1:1], comp4_0[2:2]);
  C3 I1707 (simp12891_0[1:1], comp4_0[3:3], comp4_0[4:4], comp4_0[5:5]);
  C3 I1708 (simp12891_0[2:2], comp4_0[6:6], comp4_0[7:7], comp4_0[8:8]);
  C3 I1709 (simp12891_0[3:3], comp4_0[9:9], comp4_0[10:10], comp4_0[11:11]);
  C3 I1710 (simp12891_0[4:4], comp4_0[12:12], comp4_0[13:13], comp4_0[14:14]);
  C3 I1711 (simp12891_0[5:5], comp4_0[15:15], comp4_0[16:16], comp4_0[17:17]);
  C3 I1712 (simp12891_0[6:6], comp4_0[18:18], comp4_0[19:19], comp4_0[20:20]);
  C3 I1713 (simp12891_0[7:7], comp4_0[21:21], comp4_0[22:22], comp4_0[23:23]);
  C3 I1714 (simp12891_0[8:8], comp4_0[24:24], comp4_0[25:25], comp4_0[26:26]);
  C3 I1715 (simp12891_0[9:9], comp4_0[27:27], comp4_0[28:28], comp4_0[29:29]);
  C3 I1716 (simp12891_0[10:10], comp4_0[30:30], comp4_0[31:31], comp4_0[32:32]);
  C3 I1717 (simp12891_0[11:11], comp4_0[33:33], comp4_0[34:34], comp4_0[35:35]);
  C3 I1718 (simp12891_0[12:12], comp4_0[36:36], comp4_0[37:37], comp4_0[38:38]);
  C3 I1719 (simp12891_0[13:13], comp4_0[39:39], comp4_0[40:40], comp4_0[41:41]);
  C3 I1720 (simp12891_0[14:14], comp4_0[42:42], comp4_0[43:43], comp4_0[44:44]);
  C3 I1721 (simp12891_0[15:15], comp4_0[45:45], comp4_0[46:46], comp4_0[47:47]);
  C3 I1722 (simp12891_0[16:16], comp4_0[48:48], comp4_0[49:49], comp4_0[50:50]);
  C3 I1723 (simp12891_0[17:17], comp4_0[51:51], comp4_0[52:52], comp4_0[53:53]);
  C3 I1724 (simp12891_0[18:18], comp4_0[54:54], comp4_0[55:55], comp4_0[56:56]);
  C3 I1725 (simp12891_0[19:19], comp4_0[57:57], comp4_0[58:58], comp4_0[59:59]);
  C3 I1726 (simp12891_0[20:20], comp4_0[60:60], comp4_0[61:61], comp4_0[62:62]);
  C3 I1727 (simp12891_0[21:21], comp4_0[63:63], comp4_0[64:64], comp4_0[65:65]);
  C3 I1728 (simp12891_0[22:22], comp4_0[66:66], comp4_0[67:67], comp4_0[68:68]);
  C3 I1729 (simp12891_0[23:23], comp4_0[69:69], comp4_0[70:70], comp4_0[71:71]);
  C2 I1730 (simp12891_0[24:24], comp4_0[72:72], comp4_0[73:73]);
  C3 I1731 (simp12892_0[0:0], simp12891_0[0:0], simp12891_0[1:1], simp12891_0[2:2]);
  C3 I1732 (simp12892_0[1:1], simp12891_0[3:3], simp12891_0[4:4], simp12891_0[5:5]);
  C3 I1733 (simp12892_0[2:2], simp12891_0[6:6], simp12891_0[7:7], simp12891_0[8:8]);
  C3 I1734 (simp12892_0[3:3], simp12891_0[9:9], simp12891_0[10:10], simp12891_0[11:11]);
  C3 I1735 (simp12892_0[4:4], simp12891_0[12:12], simp12891_0[13:13], simp12891_0[14:14]);
  C3 I1736 (simp12892_0[5:5], simp12891_0[15:15], simp12891_0[16:16], simp12891_0[17:17]);
  C3 I1737 (simp12892_0[6:6], simp12891_0[18:18], simp12891_0[19:19], simp12891_0[20:20]);
  C3 I1738 (simp12892_0[7:7], simp12891_0[21:21], simp12891_0[22:22], simp12891_0[23:23]);
  BUFF I1739 (simp12892_0[8:8], simp12891_0[24:24]);
  C3 I1740 (simp12893_0[0:0], simp12892_0[0:0], simp12892_0[1:1], simp12892_0[2:2]);
  C3 I1741 (simp12893_0[1:1], simp12892_0[3:3], simp12892_0[4:4], simp12892_0[5:5]);
  C3 I1742 (simp12893_0[2:2], simp12892_0[6:6], simp12892_0[7:7], simp12892_0[8:8]);
  C3 I1743 (icomp_4, simp12893_0[0:0], simp12893_0[1:1], simp12893_0[2:2]);
  C2R I1744 (choice_0, icomp_0, nchosen_0, reset);
  C2R I1745 (choice_1, icomp_1, nchosen_0, reset);
  C2R I1746 (choice_2, icomp_2, nchosen_0, reset);
  C2R I1747 (choice_3, icomp_3, nchosen_0, reset);
  C2R I1748 (choice_4, icomp_4, nchosen_0, reset);
  NOR3 I1749 (simp12951_0[0:0], choice_0, choice_1, choice_2);
  NOR2 I1750 (simp12951_0[1:1], choice_3, choice_4);
  NAND2 I1751 (anychoice_0, simp12951_0[0:0], simp12951_0[1:1]);
  NOR2 I1752 (nchosen_0, anychoice_0, o_0a);
  C2R I1753 (i_0a, choice_0, o_0a, reset);
  C2R I1754 (i_1a, choice_1, o_0a, reset);
  C2R I1755 (i_2a, choice_2, o_0a, reset);
  C2R I1756 (i_3a, choice_3, o_0a, reset);
  C2R I1757 (i_4a, choice_4, o_0a, reset);
endmodule

// tko0m5_1nm5b1 TeakO [
//     (1,TeakOConstant 5 1)] [One 0,One 5]
module tko0m5_1nm5b1 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [4:0] o_0r0;
  output [4:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  GND I1 (o_0r0[0:0]);
  BUFF I2 (o_0r0[1:1], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  GND I6 (o_0r1[1:1]);
  GND I7 (o_0r1[2:2]);
  GND I8 (o_0r1[3:3]);
  GND I9 (o_0r1[4:4]);
  BUFF I10 (i_0a, o_0a);
endmodule

// tko0m5_1nm5b2 TeakO [
//     (1,TeakOConstant 5 2)] [One 0,One 5]
module tko0m5_1nm5b2 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [4:0] o_0r0;
  output [4:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[1:1], i_0r);
  GND I1 (o_0r0[1:1]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  GND I6 (o_0r1[0:0]);
  GND I7 (o_0r1[2:2]);
  GND I8 (o_0r1[3:3]);
  GND I9 (o_0r1[4:4]);
  BUFF I10 (i_0a, o_0a);
endmodule

// tko0m5_1nm5b4 TeakO [
//     (1,TeakOConstant 5 4)] [One 0,One 5]
module tko0m5_1nm5b4 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [4:0] o_0r0;
  output [4:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[2:2], i_0r);
  GND I1 (o_0r0[2:2]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  GND I6 (o_0r1[0:0]);
  GND I7 (o_0r1[1:1]);
  GND I8 (o_0r1[3:3]);
  GND I9 (o_0r1[4:4]);
  BUFF I10 (i_0a, o_0a);
endmodule

// tko0m5_1nm5b8 TeakO [
//     (1,TeakOConstant 5 8)] [One 0,One 5]
module tko0m5_1nm5b8 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [4:0] o_0r0;
  output [4:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[3:3], i_0r);
  GND I1 (o_0r0[3:3]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  GND I6 (o_0r1[0:0]);
  GND I7 (o_0r1[1:1]);
  GND I8 (o_0r1[2:2]);
  GND I9 (o_0r1[4:4]);
  BUFF I10 (i_0a, o_0a);
endmodule

// tko0m5_1nm5b10 TeakO [
//     (1,TeakOConstant 5 16)] [One 0,One 5]
module tko0m5_1nm5b10 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [4:0] o_0r0;
  output [4:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[4:4], i_0r);
  GND I1 (o_0r0[4:4]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  GND I6 (o_0r1[0:0]);
  GND I7 (o_0r1[1:1]);
  GND I8 (o_0r1[2:2]);
  GND I9 (o_0r1[3:3]);
  BUFF I10 (i_0a, o_0a);
endmodule

// tkm5x5b TeakM [Many [5,5,5,5,5],One 5]
module tkm5x5b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, i_4r0, i_4r1, i_4a, o_0r0, o_0r1, o_0a, reset);
  input [4:0] i_0r0;
  input [4:0] i_0r1;
  output i_0a;
  input [4:0] i_1r0;
  input [4:0] i_1r1;
  output i_1a;
  input [4:0] i_2r0;
  input [4:0] i_2r1;
  output i_2a;
  input [4:0] i_3r0;
  input [4:0] i_3r1;
  output i_3a;
  input [4:0] i_4r0;
  input [4:0] i_4r1;
  output i_4a;
  output [4:0] o_0r0;
  output [4:0] o_0r1;
  input o_0a;
  input reset;
  wire [4:0] gfint_0;
  wire [4:0] gfint_1;
  wire [4:0] gfint_2;
  wire [4:0] gfint_3;
  wire [4:0] gfint_4;
  wire [4:0] gtint_0;
  wire [4:0] gtint_1;
  wire [4:0] gtint_2;
  wire [4:0] gtint_3;
  wire [4:0] gtint_4;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire choice_4;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire icomp_3;
  wire icomp_4;
  wire nchosen_0;
  wire [1:0] simp221_0;
  wire [1:0] simp231_0;
  wire [1:0] simp241_0;
  wire [1:0] simp251_0;
  wire [1:0] simp261_0;
  wire [1:0] simp271_0;
  wire [1:0] simp281_0;
  wire [1:0] simp291_0;
  wire [1:0] simp301_0;
  wire [1:0] simp311_0;
  wire [4:0] comp0_0;
  wire [1:0] simp881_0;
  wire [4:0] comp1_0;
  wire [1:0] simp951_0;
  wire [4:0] comp2_0;
  wire [1:0] simp1021_0;
  wire [4:0] comp3_0;
  wire [1:0] simp1091_0;
  wire [4:0] comp4_0;
  wire [1:0] simp1161_0;
  wire [1:0] simp1221_0;
  NOR3 I0 (simp221_0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  NOR2 I1 (simp221_0[1:1], gfint_3[0:0], gfint_4[0:0]);
  NAND2 I2 (o_0r0[0:0], simp221_0[0:0], simp221_0[1:1]);
  NOR3 I3 (simp231_0[0:0], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  NOR2 I4 (simp231_0[1:1], gfint_3[1:1], gfint_4[1:1]);
  NAND2 I5 (o_0r0[1:1], simp231_0[0:0], simp231_0[1:1]);
  NOR3 I6 (simp241_0[0:0], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  NOR2 I7 (simp241_0[1:1], gfint_3[2:2], gfint_4[2:2]);
  NAND2 I8 (o_0r0[2:2], simp241_0[0:0], simp241_0[1:1]);
  NOR3 I9 (simp251_0[0:0], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  NOR2 I10 (simp251_0[1:1], gfint_3[3:3], gfint_4[3:3]);
  NAND2 I11 (o_0r0[3:3], simp251_0[0:0], simp251_0[1:1]);
  NOR3 I12 (simp261_0[0:0], gfint_0[4:4], gfint_1[4:4], gfint_2[4:4]);
  NOR2 I13 (simp261_0[1:1], gfint_3[4:4], gfint_4[4:4]);
  NAND2 I14 (o_0r0[4:4], simp261_0[0:0], simp261_0[1:1]);
  NOR3 I15 (simp271_0[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  NOR2 I16 (simp271_0[1:1], gtint_3[0:0], gtint_4[0:0]);
  NAND2 I17 (o_0r1[0:0], simp271_0[0:0], simp271_0[1:1]);
  NOR3 I18 (simp281_0[0:0], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  NOR2 I19 (simp281_0[1:1], gtint_3[1:1], gtint_4[1:1]);
  NAND2 I20 (o_0r1[1:1], simp281_0[0:0], simp281_0[1:1]);
  NOR3 I21 (simp291_0[0:0], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  NOR2 I22 (simp291_0[1:1], gtint_3[2:2], gtint_4[2:2]);
  NAND2 I23 (o_0r1[2:2], simp291_0[0:0], simp291_0[1:1]);
  NOR3 I24 (simp301_0[0:0], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  NOR2 I25 (simp301_0[1:1], gtint_3[3:3], gtint_4[3:3]);
  NAND2 I26 (o_0r1[3:3], simp301_0[0:0], simp301_0[1:1]);
  NOR3 I27 (simp311_0[0:0], gtint_0[4:4], gtint_1[4:4], gtint_2[4:4]);
  NOR2 I28 (simp311_0[1:1], gtint_3[4:4], gtint_4[4:4]);
  NAND2 I29 (o_0r1[4:4], simp311_0[0:0], simp311_0[1:1]);
  AND2 I30 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I31 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I32 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I33 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I34 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I35 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I36 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I37 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I38 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I39 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I40 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I41 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I42 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I43 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AND2 I44 (gtint_2[4:4], choice_2, i_2r1[4:4]);
  AND2 I45 (gtint_3[0:0], choice_3, i_3r1[0:0]);
  AND2 I46 (gtint_3[1:1], choice_3, i_3r1[1:1]);
  AND2 I47 (gtint_3[2:2], choice_3, i_3r1[2:2]);
  AND2 I48 (gtint_3[3:3], choice_3, i_3r1[3:3]);
  AND2 I49 (gtint_3[4:4], choice_3, i_3r1[4:4]);
  AND2 I50 (gtint_4[0:0], choice_4, i_4r1[0:0]);
  AND2 I51 (gtint_4[1:1], choice_4, i_4r1[1:1]);
  AND2 I52 (gtint_4[2:2], choice_4, i_4r1[2:2]);
  AND2 I53 (gtint_4[3:3], choice_4, i_4r1[3:3]);
  AND2 I54 (gtint_4[4:4], choice_4, i_4r1[4:4]);
  AND2 I55 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I56 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I57 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I58 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I59 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I60 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I61 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I62 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I63 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I64 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I65 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I66 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I67 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I68 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AND2 I69 (gfint_2[4:4], choice_2, i_2r0[4:4]);
  AND2 I70 (gfint_3[0:0], choice_3, i_3r0[0:0]);
  AND2 I71 (gfint_3[1:1], choice_3, i_3r0[1:1]);
  AND2 I72 (gfint_3[2:2], choice_3, i_3r0[2:2]);
  AND2 I73 (gfint_3[3:3], choice_3, i_3r0[3:3]);
  AND2 I74 (gfint_3[4:4], choice_3, i_3r0[4:4]);
  AND2 I75 (gfint_4[0:0], choice_4, i_4r0[0:0]);
  AND2 I76 (gfint_4[1:1], choice_4, i_4r0[1:1]);
  AND2 I77 (gfint_4[2:2], choice_4, i_4r0[2:2]);
  AND2 I78 (gfint_4[3:3], choice_4, i_4r0[3:3]);
  AND2 I79 (gfint_4[4:4], choice_4, i_4r0[4:4]);
  OR2 I80 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I81 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I82 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I83 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I84 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  C3 I85 (simp881_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C2 I86 (simp881_0[1:1], comp0_0[3:3], comp0_0[4:4]);
  C2 I87 (icomp_0, simp881_0[0:0], simp881_0[1:1]);
  OR2 I88 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I89 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I90 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I91 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I92 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  C3 I93 (simp951_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C2 I94 (simp951_0[1:1], comp1_0[3:3], comp1_0[4:4]);
  C2 I95 (icomp_1, simp951_0[0:0], simp951_0[1:1]);
  OR2 I96 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I97 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I98 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2 I99 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  OR2 I100 (comp2_0[4:4], i_2r0[4:4], i_2r1[4:4]);
  C3 I101 (simp1021_0[0:0], comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C2 I102 (simp1021_0[1:1], comp2_0[3:3], comp2_0[4:4]);
  C2 I103 (icomp_2, simp1021_0[0:0], simp1021_0[1:1]);
  OR2 I104 (comp3_0[0:0], i_3r0[0:0], i_3r1[0:0]);
  OR2 I105 (comp3_0[1:1], i_3r0[1:1], i_3r1[1:1]);
  OR2 I106 (comp3_0[2:2], i_3r0[2:2], i_3r1[2:2]);
  OR2 I107 (comp3_0[3:3], i_3r0[3:3], i_3r1[3:3]);
  OR2 I108 (comp3_0[4:4], i_3r0[4:4], i_3r1[4:4]);
  C3 I109 (simp1091_0[0:0], comp3_0[0:0], comp3_0[1:1], comp3_0[2:2]);
  C2 I110 (simp1091_0[1:1], comp3_0[3:3], comp3_0[4:4]);
  C2 I111 (icomp_3, simp1091_0[0:0], simp1091_0[1:1]);
  OR2 I112 (comp4_0[0:0], i_4r0[0:0], i_4r1[0:0]);
  OR2 I113 (comp4_0[1:1], i_4r0[1:1], i_4r1[1:1]);
  OR2 I114 (comp4_0[2:2], i_4r0[2:2], i_4r1[2:2]);
  OR2 I115 (comp4_0[3:3], i_4r0[3:3], i_4r1[3:3]);
  OR2 I116 (comp4_0[4:4], i_4r0[4:4], i_4r1[4:4]);
  C3 I117 (simp1161_0[0:0], comp4_0[0:0], comp4_0[1:1], comp4_0[2:2]);
  C2 I118 (simp1161_0[1:1], comp4_0[3:3], comp4_0[4:4]);
  C2 I119 (icomp_4, simp1161_0[0:0], simp1161_0[1:1]);
  C2R I120 (choice_0, icomp_0, nchosen_0, reset);
  C2R I121 (choice_1, icomp_1, nchosen_0, reset);
  C2R I122 (choice_2, icomp_2, nchosen_0, reset);
  C2R I123 (choice_3, icomp_3, nchosen_0, reset);
  C2R I124 (choice_4, icomp_4, nchosen_0, reset);
  NOR3 I125 (simp1221_0[0:0], choice_0, choice_1, choice_2);
  NOR2 I126 (simp1221_0[1:1], choice_3, choice_4);
  NAND2 I127 (anychoice_0, simp1221_0[0:0], simp1221_0[1:1]);
  NOR2 I128 (nchosen_0, anychoice_0, o_0a);
  C2R I129 (i_0a, choice_0, o_0a, reset);
  C2R I130 (i_1a, choice_1, o_0a, reset);
  C2R I131 (i_2a, choice_2, o_0a, reset);
  C2R I132 (i_3a, choice_3, o_0a, reset);
  C2R I133 (i_4a, choice_4, o_0a, reset);
endmodule

// tkj5m0_5 TeakJ [Many [0,5],One 5]
module tkj5m0_5 (i_0r, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  input [4:0] i_1r0;
  input [4:0] i_1r1;
  output i_1a;
  output [4:0] o_0r0;
  output [4:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [4:0] joinf_0;
  wire [4:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_1r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_1r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_1r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_1r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_1r0[4:4]);
  BUFF I5 (joint_0[0:0], i_1r1[0:0]);
  BUFF I6 (joint_0[1:1], i_1r1[1:1]);
  BUFF I7 (joint_0[2:2], i_1r1[2:2]);
  BUFF I8 (joint_0[3:3], i_1r1[3:3]);
  BUFF I9 (joint_0[4:4], i_1r1[4:4]);
  BUFF I10 (icomplete_0, i_0r);
  C2 I11 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I12 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I13 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I14 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I15 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I16 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I17 (o_0r1[1:1], joint_0[1:1]);
  BUFF I18 (o_0r1[2:2], joint_0[2:2]);
  BUFF I19 (o_0r1[3:3], joint_0[3:3]);
  BUFF I20 (o_0r1[4:4], joint_0[4:4]);
  BUFF I21 (i_0a, o_0a);
  BUFF I22 (i_1a, o_0a);
endmodule

// tks5_o0w5_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0 TeakS (0+:5) [([Imp 1 0],0),([Imp 2 0],0),([Imp 4 0],0),([I
//   mp 8 0],0),([Imp 16 0],0)] [One 5,Many [0,0,0,0,0]]
module tks5_o0w5_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, reset);
  input [4:0] i_0r0;
  input [4:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire sel_4;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire gsel_4;
  wire oack_0;
  wire match0_0;
  wire [1:0] simp141_0;
  wire match1_0;
  wire [1:0] simp171_0;
  wire match2_0;
  wire [1:0] simp201_0;
  wire match3_0;
  wire [1:0] simp231_0;
  wire match4_0;
  wire [1:0] simp261_0;
  wire [4:0] comp_0;
  wire [1:0] simp381_0;
  wire [1:0] simp441_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (simp141_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C2 I2 (simp141_0[1:1], i_0r0[3:3], i_0r0[4:4]);
  C2 I3 (match0_0, simp141_0[0:0], simp141_0[1:1]);
  BUFF I4 (sel_1, match1_0);
  C3 I5 (simp171_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C2 I6 (simp171_0[1:1], i_0r0[3:3], i_0r0[4:4]);
  C2 I7 (match1_0, simp171_0[0:0], simp171_0[1:1]);
  BUFF I8 (sel_2, match2_0);
  C3 I9 (simp201_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C2 I10 (simp201_0[1:1], i_0r0[3:3], i_0r0[4:4]);
  C2 I11 (match2_0, simp201_0[0:0], simp201_0[1:1]);
  BUFF I12 (sel_3, match3_0);
  C3 I13 (simp231_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C2 I14 (simp231_0[1:1], i_0r1[3:3], i_0r0[4:4]);
  C2 I15 (match3_0, simp231_0[0:0], simp231_0[1:1]);
  BUFF I16 (sel_4, match4_0);
  C3 I17 (simp261_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C2 I18 (simp261_0[1:1], i_0r0[3:3], i_0r1[4:4]);
  C2 I19 (match4_0, simp261_0[0:0], simp261_0[1:1]);
  C2 I20 (gsel_0, sel_0, icomplete_0);
  C2 I21 (gsel_1, sel_1, icomplete_0);
  C2 I22 (gsel_2, sel_2, icomplete_0);
  C2 I23 (gsel_3, sel_3, icomplete_0);
  C2 I24 (gsel_4, sel_4, icomplete_0);
  OR2 I25 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I26 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I27 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I28 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I29 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  C3 I30 (simp381_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C2 I31 (simp381_0[1:1], comp_0[3:3], comp_0[4:4]);
  C2 I32 (icomplete_0, simp381_0[0:0], simp381_0[1:1]);
  BUFF I33 (o_0r, gsel_0);
  BUFF I34 (o_1r, gsel_1);
  BUFF I35 (o_2r, gsel_2);
  BUFF I36 (o_3r, gsel_3);
  BUFF I37 (o_4r, gsel_4);
  NOR3 I38 (simp441_0[0:0], o_0a, o_1a, o_2a);
  NOR2 I39 (simp441_0[1:1], o_3a, o_4a);
  NAND2 I40 (oack_0, simp441_0[0:0], simp441_0[1:1]);
  C2 I41 (i_0a, oack_0, icomplete_0);
endmodule

// tkf33mo0w0_o0w33 TeakF [0,0] [One 33,Many [0,33]]
module tkf33mo0w0_o0w33 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [32:0] i_0r0;
  input [32:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [32:0] o_1r0;
  output [32:0] o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_1r0[0:0], i_0r0[0:0]);
  BUFF I3 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I4 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I5 (o_1r0[3:3], i_0r0[3:3]);
  BUFF I6 (o_1r0[4:4], i_0r0[4:4]);
  BUFF I7 (o_1r0[5:5], i_0r0[5:5]);
  BUFF I8 (o_1r0[6:6], i_0r0[6:6]);
  BUFF I9 (o_1r0[7:7], i_0r0[7:7]);
  BUFF I10 (o_1r0[8:8], i_0r0[8:8]);
  BUFF I11 (o_1r0[9:9], i_0r0[9:9]);
  BUFF I12 (o_1r0[10:10], i_0r0[10:10]);
  BUFF I13 (o_1r0[11:11], i_0r0[11:11]);
  BUFF I14 (o_1r0[12:12], i_0r0[12:12]);
  BUFF I15 (o_1r0[13:13], i_0r0[13:13]);
  BUFF I16 (o_1r0[14:14], i_0r0[14:14]);
  BUFF I17 (o_1r0[15:15], i_0r0[15:15]);
  BUFF I18 (o_1r0[16:16], i_0r0[16:16]);
  BUFF I19 (o_1r0[17:17], i_0r0[17:17]);
  BUFF I20 (o_1r0[18:18], i_0r0[18:18]);
  BUFF I21 (o_1r0[19:19], i_0r0[19:19]);
  BUFF I22 (o_1r0[20:20], i_0r0[20:20]);
  BUFF I23 (o_1r0[21:21], i_0r0[21:21]);
  BUFF I24 (o_1r0[22:22], i_0r0[22:22]);
  BUFF I25 (o_1r0[23:23], i_0r0[23:23]);
  BUFF I26 (o_1r0[24:24], i_0r0[24:24]);
  BUFF I27 (o_1r0[25:25], i_0r0[25:25]);
  BUFF I28 (o_1r0[26:26], i_0r0[26:26]);
  BUFF I29 (o_1r0[27:27], i_0r0[27:27]);
  BUFF I30 (o_1r0[28:28], i_0r0[28:28]);
  BUFF I31 (o_1r0[29:29], i_0r0[29:29]);
  BUFF I32 (o_1r0[30:30], i_0r0[30:30]);
  BUFF I33 (o_1r0[31:31], i_0r0[31:31]);
  BUFF I34 (o_1r0[32:32], i_0r0[32:32]);
  BUFF I35 (o_1r1[0:0], i_0r1[0:0]);
  BUFF I36 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I37 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I38 (o_1r1[3:3], i_0r1[3:3]);
  BUFF I39 (o_1r1[4:4], i_0r1[4:4]);
  BUFF I40 (o_1r1[5:5], i_0r1[5:5]);
  BUFF I41 (o_1r1[6:6], i_0r1[6:6]);
  BUFF I42 (o_1r1[7:7], i_0r1[7:7]);
  BUFF I43 (o_1r1[8:8], i_0r1[8:8]);
  BUFF I44 (o_1r1[9:9], i_0r1[9:9]);
  BUFF I45 (o_1r1[10:10], i_0r1[10:10]);
  BUFF I46 (o_1r1[11:11], i_0r1[11:11]);
  BUFF I47 (o_1r1[12:12], i_0r1[12:12]);
  BUFF I48 (o_1r1[13:13], i_0r1[13:13]);
  BUFF I49 (o_1r1[14:14], i_0r1[14:14]);
  BUFF I50 (o_1r1[15:15], i_0r1[15:15]);
  BUFF I51 (o_1r1[16:16], i_0r1[16:16]);
  BUFF I52 (o_1r1[17:17], i_0r1[17:17]);
  BUFF I53 (o_1r1[18:18], i_0r1[18:18]);
  BUFF I54 (o_1r1[19:19], i_0r1[19:19]);
  BUFF I55 (o_1r1[20:20], i_0r1[20:20]);
  BUFF I56 (o_1r1[21:21], i_0r1[21:21]);
  BUFF I57 (o_1r1[22:22], i_0r1[22:22]);
  BUFF I58 (o_1r1[23:23], i_0r1[23:23]);
  BUFF I59 (o_1r1[24:24], i_0r1[24:24]);
  BUFF I60 (o_1r1[25:25], i_0r1[25:25]);
  BUFF I61 (o_1r1[26:26], i_0r1[26:26]);
  BUFF I62 (o_1r1[27:27], i_0r1[27:27]);
  BUFF I63 (o_1r1[28:28], i_0r1[28:28]);
  BUFF I64 (o_1r1[29:29], i_0r1[29:29]);
  BUFF I65 (o_1r1[30:30], i_0r1[30:30]);
  BUFF I66 (o_1r1[31:31], i_0r1[31:31]);
  BUFF I67 (o_1r1[32:32], i_0r1[32:32]);
  BUFF I68 (o_0r, icomplete_0);
  C3 I69 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tki TeakI [One 0,One 0]
module tki (i_0r, i_0a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  input reset;
  wire nreset_0;
  wire firsthsa_0;
  wire nfirsthsa_0;
  wire firsthsd_0;
  wire noa_0;
  INV I0 (nreset_0, reset);
  INV I1 (nfirsthsa_0, firsthsa_0);
  INV I2 (noa_0, o_0a);
  AO22 I3 (o_0r, nreset_0, nfirsthsa_0, i_0r, firsthsd_0);
  AO22 I4 (firsthsa_0, nreset_0, o_0a, nreset_0, firsthsa_0);
  AO22 I5 (firsthsd_0, firsthsa_0, noa_0, firsthsa_0, firsthsd_0);
  AND2 I6 (i_0a, o_0a, firsthsd_0);
endmodule

// tkj32m1_31 TeakJ [Many [1,31],One 32]
module tkj32m1_31 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input [30:0] i_1r0;
  input [30:0] i_1r1;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [31:0] joinf_0;
  wire [31:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0);
  BUFF I1 (joinf_0[1:1], i_1r0[0:0]);
  BUFF I2 (joinf_0[2:2], i_1r0[1:1]);
  BUFF I3 (joinf_0[3:3], i_1r0[2:2]);
  BUFF I4 (joinf_0[4:4], i_1r0[3:3]);
  BUFF I5 (joinf_0[5:5], i_1r0[4:4]);
  BUFF I6 (joinf_0[6:6], i_1r0[5:5]);
  BUFF I7 (joinf_0[7:7], i_1r0[6:6]);
  BUFF I8 (joinf_0[8:8], i_1r0[7:7]);
  BUFF I9 (joinf_0[9:9], i_1r0[8:8]);
  BUFF I10 (joinf_0[10:10], i_1r0[9:9]);
  BUFF I11 (joinf_0[11:11], i_1r0[10:10]);
  BUFF I12 (joinf_0[12:12], i_1r0[11:11]);
  BUFF I13 (joinf_0[13:13], i_1r0[12:12]);
  BUFF I14 (joinf_0[14:14], i_1r0[13:13]);
  BUFF I15 (joinf_0[15:15], i_1r0[14:14]);
  BUFF I16 (joinf_0[16:16], i_1r0[15:15]);
  BUFF I17 (joinf_0[17:17], i_1r0[16:16]);
  BUFF I18 (joinf_0[18:18], i_1r0[17:17]);
  BUFF I19 (joinf_0[19:19], i_1r0[18:18]);
  BUFF I20 (joinf_0[20:20], i_1r0[19:19]);
  BUFF I21 (joinf_0[21:21], i_1r0[20:20]);
  BUFF I22 (joinf_0[22:22], i_1r0[21:21]);
  BUFF I23 (joinf_0[23:23], i_1r0[22:22]);
  BUFF I24 (joinf_0[24:24], i_1r0[23:23]);
  BUFF I25 (joinf_0[25:25], i_1r0[24:24]);
  BUFF I26 (joinf_0[26:26], i_1r0[25:25]);
  BUFF I27 (joinf_0[27:27], i_1r0[26:26]);
  BUFF I28 (joinf_0[28:28], i_1r0[27:27]);
  BUFF I29 (joinf_0[29:29], i_1r0[28:28]);
  BUFF I30 (joinf_0[30:30], i_1r0[29:29]);
  BUFF I31 (joinf_0[31:31], i_1r0[30:30]);
  BUFF I32 (joint_0[0:0], i_0r1);
  BUFF I33 (joint_0[1:1], i_1r1[0:0]);
  BUFF I34 (joint_0[2:2], i_1r1[1:1]);
  BUFF I35 (joint_0[3:3], i_1r1[2:2]);
  BUFF I36 (joint_0[4:4], i_1r1[3:3]);
  BUFF I37 (joint_0[5:5], i_1r1[4:4]);
  BUFF I38 (joint_0[6:6], i_1r1[5:5]);
  BUFF I39 (joint_0[7:7], i_1r1[6:6]);
  BUFF I40 (joint_0[8:8], i_1r1[7:7]);
  BUFF I41 (joint_0[9:9], i_1r1[8:8]);
  BUFF I42 (joint_0[10:10], i_1r1[9:9]);
  BUFF I43 (joint_0[11:11], i_1r1[10:10]);
  BUFF I44 (joint_0[12:12], i_1r1[11:11]);
  BUFF I45 (joint_0[13:13], i_1r1[12:12]);
  BUFF I46 (joint_0[14:14], i_1r1[13:13]);
  BUFF I47 (joint_0[15:15], i_1r1[14:14]);
  BUFF I48 (joint_0[16:16], i_1r1[15:15]);
  BUFF I49 (joint_0[17:17], i_1r1[16:16]);
  BUFF I50 (joint_0[18:18], i_1r1[17:17]);
  BUFF I51 (joint_0[19:19], i_1r1[18:18]);
  BUFF I52 (joint_0[20:20], i_1r1[19:19]);
  BUFF I53 (joint_0[21:21], i_1r1[20:20]);
  BUFF I54 (joint_0[22:22], i_1r1[21:21]);
  BUFF I55 (joint_0[23:23], i_1r1[22:22]);
  BUFF I56 (joint_0[24:24], i_1r1[23:23]);
  BUFF I57 (joint_0[25:25], i_1r1[24:24]);
  BUFF I58 (joint_0[26:26], i_1r1[25:25]);
  BUFF I59 (joint_0[27:27], i_1r1[26:26]);
  BUFF I60 (joint_0[28:28], i_1r1[27:27]);
  BUFF I61 (joint_0[29:29], i_1r1[28:28]);
  BUFF I62 (joint_0[30:30], i_1r1[29:29]);
  BUFF I63 (joint_0[31:31], i_1r1[30:30]);
  OR2 I64 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I65 (icomplete_0, dcomplete_0);
  C2 I66 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I67 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I68 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I69 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I70 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I71 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I72 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I73 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I74 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I75 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I76 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I77 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I78 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I79 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I80 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I81 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I82 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I83 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I84 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I85 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I86 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I87 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I88 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I89 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I90 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I91 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I92 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I93 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I94 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I95 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I96 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I97 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I98 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I99 (o_0r1[1:1], joint_0[1:1]);
  BUFF I100 (o_0r1[2:2], joint_0[2:2]);
  BUFF I101 (o_0r1[3:3], joint_0[3:3]);
  BUFF I102 (o_0r1[4:4], joint_0[4:4]);
  BUFF I103 (o_0r1[5:5], joint_0[5:5]);
  BUFF I104 (o_0r1[6:6], joint_0[6:6]);
  BUFF I105 (o_0r1[7:7], joint_0[7:7]);
  BUFF I106 (o_0r1[8:8], joint_0[8:8]);
  BUFF I107 (o_0r1[9:9], joint_0[9:9]);
  BUFF I108 (o_0r1[10:10], joint_0[10:10]);
  BUFF I109 (o_0r1[11:11], joint_0[11:11]);
  BUFF I110 (o_0r1[12:12], joint_0[12:12]);
  BUFF I111 (o_0r1[13:13], joint_0[13:13]);
  BUFF I112 (o_0r1[14:14], joint_0[14:14]);
  BUFF I113 (o_0r1[15:15], joint_0[15:15]);
  BUFF I114 (o_0r1[16:16], joint_0[16:16]);
  BUFF I115 (o_0r1[17:17], joint_0[17:17]);
  BUFF I116 (o_0r1[18:18], joint_0[18:18]);
  BUFF I117 (o_0r1[19:19], joint_0[19:19]);
  BUFF I118 (o_0r1[20:20], joint_0[20:20]);
  BUFF I119 (o_0r1[21:21], joint_0[21:21]);
  BUFF I120 (o_0r1[22:22], joint_0[22:22]);
  BUFF I121 (o_0r1[23:23], joint_0[23:23]);
  BUFF I122 (o_0r1[24:24], joint_0[24:24]);
  BUFF I123 (o_0r1[25:25], joint_0[25:25]);
  BUFF I124 (o_0r1[26:26], joint_0[26:26]);
  BUFF I125 (o_0r1[27:27], joint_0[27:27]);
  BUFF I126 (o_0r1[28:28], joint_0[28:28]);
  BUFF I127 (o_0r1[29:29], joint_0[29:29]);
  BUFF I128 (o_0r1[30:30], joint_0[30:30]);
  BUFF I129 (o_0r1[31:31], joint_0[31:31]);
  BUFF I130 (i_0a, o_0a);
  BUFF I131 (i_1a, o_0a);
endmodule

// tkj32m31_1 TeakJ [Many [31,1],One 32]
module tkj32m31_1 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [30:0] i_0r0;
  input [30:0] i_0r1;
  output i_0a;
  input i_1r0;
  input i_1r1;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [31:0] joinf_0;
  wire [31:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_1r0);
  BUFF I32 (joint_0[0:0], i_0r1[0:0]);
  BUFF I33 (joint_0[1:1], i_0r1[1:1]);
  BUFF I34 (joint_0[2:2], i_0r1[2:2]);
  BUFF I35 (joint_0[3:3], i_0r1[3:3]);
  BUFF I36 (joint_0[4:4], i_0r1[4:4]);
  BUFF I37 (joint_0[5:5], i_0r1[5:5]);
  BUFF I38 (joint_0[6:6], i_0r1[6:6]);
  BUFF I39 (joint_0[7:7], i_0r1[7:7]);
  BUFF I40 (joint_0[8:8], i_0r1[8:8]);
  BUFF I41 (joint_0[9:9], i_0r1[9:9]);
  BUFF I42 (joint_0[10:10], i_0r1[10:10]);
  BUFF I43 (joint_0[11:11], i_0r1[11:11]);
  BUFF I44 (joint_0[12:12], i_0r1[12:12]);
  BUFF I45 (joint_0[13:13], i_0r1[13:13]);
  BUFF I46 (joint_0[14:14], i_0r1[14:14]);
  BUFF I47 (joint_0[15:15], i_0r1[15:15]);
  BUFF I48 (joint_0[16:16], i_0r1[16:16]);
  BUFF I49 (joint_0[17:17], i_0r1[17:17]);
  BUFF I50 (joint_0[18:18], i_0r1[18:18]);
  BUFF I51 (joint_0[19:19], i_0r1[19:19]);
  BUFF I52 (joint_0[20:20], i_0r1[20:20]);
  BUFF I53 (joint_0[21:21], i_0r1[21:21]);
  BUFF I54 (joint_0[22:22], i_0r1[22:22]);
  BUFF I55 (joint_0[23:23], i_0r1[23:23]);
  BUFF I56 (joint_0[24:24], i_0r1[24:24]);
  BUFF I57 (joint_0[25:25], i_0r1[25:25]);
  BUFF I58 (joint_0[26:26], i_0r1[26:26]);
  BUFF I59 (joint_0[27:27], i_0r1[27:27]);
  BUFF I60 (joint_0[28:28], i_0r1[28:28]);
  BUFF I61 (joint_0[29:29], i_0r1[29:29]);
  BUFF I62 (joint_0[30:30], i_0r1[30:30]);
  BUFF I63 (joint_0[31:31], i_1r1);
  OR2 I64 (dcomplete_0, i_1r0, i_1r1);
  BUFF I65 (icomplete_0, dcomplete_0);
  C2 I66 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I67 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I68 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I69 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I70 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I71 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I72 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I73 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I74 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I75 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I76 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I77 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I78 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I79 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I80 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I81 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I82 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I83 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I84 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I85 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I86 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I87 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I88 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I89 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I90 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I91 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I92 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I93 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I94 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I95 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I96 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I97 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I98 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I99 (o_0r1[1:1], joint_0[1:1]);
  BUFF I100 (o_0r1[2:2], joint_0[2:2]);
  BUFF I101 (o_0r1[3:3], joint_0[3:3]);
  BUFF I102 (o_0r1[4:4], joint_0[4:4]);
  BUFF I103 (o_0r1[5:5], joint_0[5:5]);
  BUFF I104 (o_0r1[6:6], joint_0[6:6]);
  BUFF I105 (o_0r1[7:7], joint_0[7:7]);
  BUFF I106 (o_0r1[8:8], joint_0[8:8]);
  BUFF I107 (o_0r1[9:9], joint_0[9:9]);
  BUFF I108 (o_0r1[10:10], joint_0[10:10]);
  BUFF I109 (o_0r1[11:11], joint_0[11:11]);
  BUFF I110 (o_0r1[12:12], joint_0[12:12]);
  BUFF I111 (o_0r1[13:13], joint_0[13:13]);
  BUFF I112 (o_0r1[14:14], joint_0[14:14]);
  BUFF I113 (o_0r1[15:15], joint_0[15:15]);
  BUFF I114 (o_0r1[16:16], joint_0[16:16]);
  BUFF I115 (o_0r1[17:17], joint_0[17:17]);
  BUFF I116 (o_0r1[18:18], joint_0[18:18]);
  BUFF I117 (o_0r1[19:19], joint_0[19:19]);
  BUFF I118 (o_0r1[20:20], joint_0[20:20]);
  BUFF I119 (o_0r1[21:21], joint_0[21:21]);
  BUFF I120 (o_0r1[22:22], joint_0[22:22]);
  BUFF I121 (o_0r1[23:23], joint_0[23:23]);
  BUFF I122 (o_0r1[24:24], joint_0[24:24]);
  BUFF I123 (o_0r1[25:25], joint_0[25:25]);
  BUFF I124 (o_0r1[26:26], joint_0[26:26]);
  BUFF I125 (o_0r1[27:27], joint_0[27:27]);
  BUFF I126 (o_0r1[28:28], joint_0[28:28]);
  BUFF I127 (o_0r1[29:29], joint_0[29:29]);
  BUFF I128 (o_0r1[30:30], joint_0[30:30]);
  BUFF I129 (o_0r1[31:31], joint_0[31:31]);
  BUFF I130 (i_0a, o_0a);
  BUFF I131 (i_1a, o_0a);
endmodule

// tks2_o0w2_0c2o0w0_1o0w0_3o0w0 TeakS (0+:2) [([Imp 0 2],0),([Imp 1 0],0),([Imp 3 0],0)] [One 2,Many [
//   0,0,0]]
module tks2_o0w2_0c2o0w0_1o0w0_3o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire match2_0;
  wire [1:0] comp_0;
  BUFF I0 (sel_0, match0_0);
  BUFF I1 (match0_0, i_0r0[0:0]);
  BUFF I2 (sel_1, match1_0);
  C2 I3 (match1_0, i_0r1[0:0], i_0r0[1:1]);
  BUFF I4 (sel_2, match2_0);
  C2 I5 (match2_0, i_0r1[0:0], i_0r1[1:1]);
  C2 I6 (gsel_0, sel_0, icomplete_0);
  C2 I7 (gsel_1, sel_1, icomplete_0);
  C2 I8 (gsel_2, sel_2, icomplete_0);
  OR2 I9 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I10 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  C2 I11 (icomplete_0, comp_0[0:0], comp_0[1:1]);
  BUFF I12 (o_0r, gsel_0);
  BUFF I13 (o_1r, gsel_1);
  BUFF I14 (o_2r, gsel_2);
  OR3 I15 (oack_0, o_0a, o_1a, o_2a);
  C2 I16 (i_0a, oack_0, icomplete_0);
endmodule

// tkvi32_wo0w32_ro0w32o0w31o1w31o1w31 TeakV "i" 32 [] [0] [0,0,1,1] [Many [32],Many [0],Many [0,0,0,0]
//   ,Many [32,31,31,31]]
module tkvi32_wo0w32_ro0w32o0w31o1w31o1w31 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [30:0] rd_1r0;
  output [30:0] rd_1r1;
  input rd_1a;
  output [30:0] rd_2r0;
  output [30:0] rd_2r1;
  input rd_2a;
  output [30:0] rd_3r0;
  output [30:0] rd_3r1;
  input rd_3a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [2:0] simp6581_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_2r0[0:0], df_0[1:1], rg_2r);
  AND2 I488 (rd_2r0[1:1], df_0[2:2], rg_2r);
  AND2 I489 (rd_2r0[2:2], df_0[3:3], rg_2r);
  AND2 I490 (rd_2r0[3:3], df_0[4:4], rg_2r);
  AND2 I491 (rd_2r0[4:4], df_0[5:5], rg_2r);
  AND2 I492 (rd_2r0[5:5], df_0[6:6], rg_2r);
  AND2 I493 (rd_2r0[6:6], df_0[7:7], rg_2r);
  AND2 I494 (rd_2r0[7:7], df_0[8:8], rg_2r);
  AND2 I495 (rd_2r0[8:8], df_0[9:9], rg_2r);
  AND2 I496 (rd_2r0[9:9], df_0[10:10], rg_2r);
  AND2 I497 (rd_2r0[10:10], df_0[11:11], rg_2r);
  AND2 I498 (rd_2r0[11:11], df_0[12:12], rg_2r);
  AND2 I499 (rd_2r0[12:12], df_0[13:13], rg_2r);
  AND2 I500 (rd_2r0[13:13], df_0[14:14], rg_2r);
  AND2 I501 (rd_2r0[14:14], df_0[15:15], rg_2r);
  AND2 I502 (rd_2r0[15:15], df_0[16:16], rg_2r);
  AND2 I503 (rd_2r0[16:16], df_0[17:17], rg_2r);
  AND2 I504 (rd_2r0[17:17], df_0[18:18], rg_2r);
  AND2 I505 (rd_2r0[18:18], df_0[19:19], rg_2r);
  AND2 I506 (rd_2r0[19:19], df_0[20:20], rg_2r);
  AND2 I507 (rd_2r0[20:20], df_0[21:21], rg_2r);
  AND2 I508 (rd_2r0[21:21], df_0[22:22], rg_2r);
  AND2 I509 (rd_2r0[22:22], df_0[23:23], rg_2r);
  AND2 I510 (rd_2r0[23:23], df_0[24:24], rg_2r);
  AND2 I511 (rd_2r0[24:24], df_0[25:25], rg_2r);
  AND2 I512 (rd_2r0[25:25], df_0[26:26], rg_2r);
  AND2 I513 (rd_2r0[26:26], df_0[27:27], rg_2r);
  AND2 I514 (rd_2r0[27:27], df_0[28:28], rg_2r);
  AND2 I515 (rd_2r0[28:28], df_0[29:29], rg_2r);
  AND2 I516 (rd_2r0[29:29], df_0[30:30], rg_2r);
  AND2 I517 (rd_2r0[30:30], df_0[31:31], rg_2r);
  AND2 I518 (rd_3r0[0:0], df_0[1:1], rg_3r);
  AND2 I519 (rd_3r0[1:1], df_0[2:2], rg_3r);
  AND2 I520 (rd_3r0[2:2], df_0[3:3], rg_3r);
  AND2 I521 (rd_3r0[3:3], df_0[4:4], rg_3r);
  AND2 I522 (rd_3r0[4:4], df_0[5:5], rg_3r);
  AND2 I523 (rd_3r0[5:5], df_0[6:6], rg_3r);
  AND2 I524 (rd_3r0[6:6], df_0[7:7], rg_3r);
  AND2 I525 (rd_3r0[7:7], df_0[8:8], rg_3r);
  AND2 I526 (rd_3r0[8:8], df_0[9:9], rg_3r);
  AND2 I527 (rd_3r0[9:9], df_0[10:10], rg_3r);
  AND2 I528 (rd_3r0[10:10], df_0[11:11], rg_3r);
  AND2 I529 (rd_3r0[11:11], df_0[12:12], rg_3r);
  AND2 I530 (rd_3r0[12:12], df_0[13:13], rg_3r);
  AND2 I531 (rd_3r0[13:13], df_0[14:14], rg_3r);
  AND2 I532 (rd_3r0[14:14], df_0[15:15], rg_3r);
  AND2 I533 (rd_3r0[15:15], df_0[16:16], rg_3r);
  AND2 I534 (rd_3r0[16:16], df_0[17:17], rg_3r);
  AND2 I535 (rd_3r0[17:17], df_0[18:18], rg_3r);
  AND2 I536 (rd_3r0[18:18], df_0[19:19], rg_3r);
  AND2 I537 (rd_3r0[19:19], df_0[20:20], rg_3r);
  AND2 I538 (rd_3r0[20:20], df_0[21:21], rg_3r);
  AND2 I539 (rd_3r0[21:21], df_0[22:22], rg_3r);
  AND2 I540 (rd_3r0[22:22], df_0[23:23], rg_3r);
  AND2 I541 (rd_3r0[23:23], df_0[24:24], rg_3r);
  AND2 I542 (rd_3r0[24:24], df_0[25:25], rg_3r);
  AND2 I543 (rd_3r0[25:25], df_0[26:26], rg_3r);
  AND2 I544 (rd_3r0[26:26], df_0[27:27], rg_3r);
  AND2 I545 (rd_3r0[27:27], df_0[28:28], rg_3r);
  AND2 I546 (rd_3r0[28:28], df_0[29:29], rg_3r);
  AND2 I547 (rd_3r0[29:29], df_0[30:30], rg_3r);
  AND2 I548 (rd_3r0[30:30], df_0[31:31], rg_3r);
  AND2 I549 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I550 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I551 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I552 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I553 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I554 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I555 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I556 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I557 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I558 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I559 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I560 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I561 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I562 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I563 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I564 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I565 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I566 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I567 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I568 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I569 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I570 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I571 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I572 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I573 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I574 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I575 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I576 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I577 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I578 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I579 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I580 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I581 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I582 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I583 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I584 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I585 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I586 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I587 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I588 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I589 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I590 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I591 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I592 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I593 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I594 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I595 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I596 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I597 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I598 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I599 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I600 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I601 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I602 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I603 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I604 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I605 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I606 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I607 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I608 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I609 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I610 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I611 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I612 (rd_2r1[0:0], dt_0[1:1], rg_2r);
  AND2 I613 (rd_2r1[1:1], dt_0[2:2], rg_2r);
  AND2 I614 (rd_2r1[2:2], dt_0[3:3], rg_2r);
  AND2 I615 (rd_2r1[3:3], dt_0[4:4], rg_2r);
  AND2 I616 (rd_2r1[4:4], dt_0[5:5], rg_2r);
  AND2 I617 (rd_2r1[5:5], dt_0[6:6], rg_2r);
  AND2 I618 (rd_2r1[6:6], dt_0[7:7], rg_2r);
  AND2 I619 (rd_2r1[7:7], dt_0[8:8], rg_2r);
  AND2 I620 (rd_2r1[8:8], dt_0[9:9], rg_2r);
  AND2 I621 (rd_2r1[9:9], dt_0[10:10], rg_2r);
  AND2 I622 (rd_2r1[10:10], dt_0[11:11], rg_2r);
  AND2 I623 (rd_2r1[11:11], dt_0[12:12], rg_2r);
  AND2 I624 (rd_2r1[12:12], dt_0[13:13], rg_2r);
  AND2 I625 (rd_2r1[13:13], dt_0[14:14], rg_2r);
  AND2 I626 (rd_2r1[14:14], dt_0[15:15], rg_2r);
  AND2 I627 (rd_2r1[15:15], dt_0[16:16], rg_2r);
  AND2 I628 (rd_2r1[16:16], dt_0[17:17], rg_2r);
  AND2 I629 (rd_2r1[17:17], dt_0[18:18], rg_2r);
  AND2 I630 (rd_2r1[18:18], dt_0[19:19], rg_2r);
  AND2 I631 (rd_2r1[19:19], dt_0[20:20], rg_2r);
  AND2 I632 (rd_2r1[20:20], dt_0[21:21], rg_2r);
  AND2 I633 (rd_2r1[21:21], dt_0[22:22], rg_2r);
  AND2 I634 (rd_2r1[22:22], dt_0[23:23], rg_2r);
  AND2 I635 (rd_2r1[23:23], dt_0[24:24], rg_2r);
  AND2 I636 (rd_2r1[24:24], dt_0[25:25], rg_2r);
  AND2 I637 (rd_2r1[25:25], dt_0[26:26], rg_2r);
  AND2 I638 (rd_2r1[26:26], dt_0[27:27], rg_2r);
  AND2 I639 (rd_2r1[27:27], dt_0[28:28], rg_2r);
  AND2 I640 (rd_2r1[28:28], dt_0[29:29], rg_2r);
  AND2 I641 (rd_2r1[29:29], dt_0[30:30], rg_2r);
  AND2 I642 (rd_2r1[30:30], dt_0[31:31], rg_2r);
  AND2 I643 (rd_3r1[0:0], dt_0[1:1], rg_3r);
  AND2 I644 (rd_3r1[1:1], dt_0[2:2], rg_3r);
  AND2 I645 (rd_3r1[2:2], dt_0[3:3], rg_3r);
  AND2 I646 (rd_3r1[3:3], dt_0[4:4], rg_3r);
  AND2 I647 (rd_3r1[4:4], dt_0[5:5], rg_3r);
  AND2 I648 (rd_3r1[5:5], dt_0[6:6], rg_3r);
  AND2 I649 (rd_3r1[6:6], dt_0[7:7], rg_3r);
  AND2 I650 (rd_3r1[7:7], dt_0[8:8], rg_3r);
  AND2 I651 (rd_3r1[8:8], dt_0[9:9], rg_3r);
  AND2 I652 (rd_3r1[9:9], dt_0[10:10], rg_3r);
  AND2 I653 (rd_3r1[10:10], dt_0[11:11], rg_3r);
  AND2 I654 (rd_3r1[11:11], dt_0[12:12], rg_3r);
  AND2 I655 (rd_3r1[12:12], dt_0[13:13], rg_3r);
  AND2 I656 (rd_3r1[13:13], dt_0[14:14], rg_3r);
  AND2 I657 (rd_3r1[14:14], dt_0[15:15], rg_3r);
  AND2 I658 (rd_3r1[15:15], dt_0[16:16], rg_3r);
  AND2 I659 (rd_3r1[16:16], dt_0[17:17], rg_3r);
  AND2 I660 (rd_3r1[17:17], dt_0[18:18], rg_3r);
  AND2 I661 (rd_3r1[18:18], dt_0[19:19], rg_3r);
  AND2 I662 (rd_3r1[19:19], dt_0[20:20], rg_3r);
  AND2 I663 (rd_3r1[20:20], dt_0[21:21], rg_3r);
  AND2 I664 (rd_3r1[21:21], dt_0[22:22], rg_3r);
  AND2 I665 (rd_3r1[22:22], dt_0[23:23], rg_3r);
  AND2 I666 (rd_3r1[23:23], dt_0[24:24], rg_3r);
  AND2 I667 (rd_3r1[24:24], dt_0[25:25], rg_3r);
  AND2 I668 (rd_3r1[25:25], dt_0[26:26], rg_3r);
  AND2 I669 (rd_3r1[26:26], dt_0[27:27], rg_3r);
  AND2 I670 (rd_3r1[27:27], dt_0[28:28], rg_3r);
  AND2 I671 (rd_3r1[28:28], dt_0[29:29], rg_3r);
  AND2 I672 (rd_3r1[29:29], dt_0[30:30], rg_3r);
  AND2 I673 (rd_3r1[30:30], dt_0[31:31], rg_3r);
  NOR3 I674 (simp6581_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I675 (simp6581_0[1:1], rg_3r, rg_0a, rg_1a);
  NOR2 I676 (simp6581_0[2:2], rg_2a, rg_3a);
  NAND3 I677 (anyread_0, simp6581_0[0:0], simp6581_0[1:1], simp6581_0[2:2]);
  BUFF I678 (wg_0a, wd_0a);
  BUFF I679 (rg_0a, rd_0a);
  BUFF I680 (rg_1a, rd_1a);
  BUFF I681 (rg_2a, rd_2a);
  BUFF I682 (rg_3a, rd_3a);
endmodule

// tkj32m2_30 TeakJ [Many [2,30],One 32]
module tkj32m2_30 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  input [29:0] i_1r0;
  input [29:0] i_1r1;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [31:0] joinf_0;
  wire [31:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_1r0[0:0]);
  BUFF I3 (joinf_0[3:3], i_1r0[1:1]);
  BUFF I4 (joinf_0[4:4], i_1r0[2:2]);
  BUFF I5 (joinf_0[5:5], i_1r0[3:3]);
  BUFF I6 (joinf_0[6:6], i_1r0[4:4]);
  BUFF I7 (joinf_0[7:7], i_1r0[5:5]);
  BUFF I8 (joinf_0[8:8], i_1r0[6:6]);
  BUFF I9 (joinf_0[9:9], i_1r0[7:7]);
  BUFF I10 (joinf_0[10:10], i_1r0[8:8]);
  BUFF I11 (joinf_0[11:11], i_1r0[9:9]);
  BUFF I12 (joinf_0[12:12], i_1r0[10:10]);
  BUFF I13 (joinf_0[13:13], i_1r0[11:11]);
  BUFF I14 (joinf_0[14:14], i_1r0[12:12]);
  BUFF I15 (joinf_0[15:15], i_1r0[13:13]);
  BUFF I16 (joinf_0[16:16], i_1r0[14:14]);
  BUFF I17 (joinf_0[17:17], i_1r0[15:15]);
  BUFF I18 (joinf_0[18:18], i_1r0[16:16]);
  BUFF I19 (joinf_0[19:19], i_1r0[17:17]);
  BUFF I20 (joinf_0[20:20], i_1r0[18:18]);
  BUFF I21 (joinf_0[21:21], i_1r0[19:19]);
  BUFF I22 (joinf_0[22:22], i_1r0[20:20]);
  BUFF I23 (joinf_0[23:23], i_1r0[21:21]);
  BUFF I24 (joinf_0[24:24], i_1r0[22:22]);
  BUFF I25 (joinf_0[25:25], i_1r0[23:23]);
  BUFF I26 (joinf_0[26:26], i_1r0[24:24]);
  BUFF I27 (joinf_0[27:27], i_1r0[25:25]);
  BUFF I28 (joinf_0[28:28], i_1r0[26:26]);
  BUFF I29 (joinf_0[29:29], i_1r0[27:27]);
  BUFF I30 (joinf_0[30:30], i_1r0[28:28]);
  BUFF I31 (joinf_0[31:31], i_1r0[29:29]);
  BUFF I32 (joint_0[0:0], i_0r1[0:0]);
  BUFF I33 (joint_0[1:1], i_0r1[1:1]);
  BUFF I34 (joint_0[2:2], i_1r1[0:0]);
  BUFF I35 (joint_0[3:3], i_1r1[1:1]);
  BUFF I36 (joint_0[4:4], i_1r1[2:2]);
  BUFF I37 (joint_0[5:5], i_1r1[3:3]);
  BUFF I38 (joint_0[6:6], i_1r1[4:4]);
  BUFF I39 (joint_0[7:7], i_1r1[5:5]);
  BUFF I40 (joint_0[8:8], i_1r1[6:6]);
  BUFF I41 (joint_0[9:9], i_1r1[7:7]);
  BUFF I42 (joint_0[10:10], i_1r1[8:8]);
  BUFF I43 (joint_0[11:11], i_1r1[9:9]);
  BUFF I44 (joint_0[12:12], i_1r1[10:10]);
  BUFF I45 (joint_0[13:13], i_1r1[11:11]);
  BUFF I46 (joint_0[14:14], i_1r1[12:12]);
  BUFF I47 (joint_0[15:15], i_1r1[13:13]);
  BUFF I48 (joint_0[16:16], i_1r1[14:14]);
  BUFF I49 (joint_0[17:17], i_1r1[15:15]);
  BUFF I50 (joint_0[18:18], i_1r1[16:16]);
  BUFF I51 (joint_0[19:19], i_1r1[17:17]);
  BUFF I52 (joint_0[20:20], i_1r1[18:18]);
  BUFF I53 (joint_0[21:21], i_1r1[19:19]);
  BUFF I54 (joint_0[22:22], i_1r1[20:20]);
  BUFF I55 (joint_0[23:23], i_1r1[21:21]);
  BUFF I56 (joint_0[24:24], i_1r1[22:22]);
  BUFF I57 (joint_0[25:25], i_1r1[23:23]);
  BUFF I58 (joint_0[26:26], i_1r1[24:24]);
  BUFF I59 (joint_0[27:27], i_1r1[25:25]);
  BUFF I60 (joint_0[28:28], i_1r1[26:26]);
  BUFF I61 (joint_0[29:29], i_1r1[27:27]);
  BUFF I62 (joint_0[30:30], i_1r1[28:28]);
  BUFF I63 (joint_0[31:31], i_1r1[29:29]);
  OR2 I64 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I65 (icomplete_0, dcomplete_0);
  C2 I66 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I67 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I68 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I69 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I70 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I71 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I72 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I73 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I74 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I75 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I76 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I77 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I78 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I79 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I80 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I81 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I82 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I83 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I84 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I85 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I86 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I87 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I88 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I89 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I90 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I91 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I92 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I93 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I94 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I95 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I96 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I97 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I98 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I99 (o_0r1[1:1], joint_0[1:1]);
  BUFF I100 (o_0r1[2:2], joint_0[2:2]);
  BUFF I101 (o_0r1[3:3], joint_0[3:3]);
  BUFF I102 (o_0r1[4:4], joint_0[4:4]);
  BUFF I103 (o_0r1[5:5], joint_0[5:5]);
  BUFF I104 (o_0r1[6:6], joint_0[6:6]);
  BUFF I105 (o_0r1[7:7], joint_0[7:7]);
  BUFF I106 (o_0r1[8:8], joint_0[8:8]);
  BUFF I107 (o_0r1[9:9], joint_0[9:9]);
  BUFF I108 (o_0r1[10:10], joint_0[10:10]);
  BUFF I109 (o_0r1[11:11], joint_0[11:11]);
  BUFF I110 (o_0r1[12:12], joint_0[12:12]);
  BUFF I111 (o_0r1[13:13], joint_0[13:13]);
  BUFF I112 (o_0r1[14:14], joint_0[14:14]);
  BUFF I113 (o_0r1[15:15], joint_0[15:15]);
  BUFF I114 (o_0r1[16:16], joint_0[16:16]);
  BUFF I115 (o_0r1[17:17], joint_0[17:17]);
  BUFF I116 (o_0r1[18:18], joint_0[18:18]);
  BUFF I117 (o_0r1[19:19], joint_0[19:19]);
  BUFF I118 (o_0r1[20:20], joint_0[20:20]);
  BUFF I119 (o_0r1[21:21], joint_0[21:21]);
  BUFF I120 (o_0r1[22:22], joint_0[22:22]);
  BUFF I121 (o_0r1[23:23], joint_0[23:23]);
  BUFF I122 (o_0r1[24:24], joint_0[24:24]);
  BUFF I123 (o_0r1[25:25], joint_0[25:25]);
  BUFF I124 (o_0r1[26:26], joint_0[26:26]);
  BUFF I125 (o_0r1[27:27], joint_0[27:27]);
  BUFF I126 (o_0r1[28:28], joint_0[28:28]);
  BUFF I127 (o_0r1[29:29], joint_0[29:29]);
  BUFF I128 (o_0r1[30:30], joint_0[30:30]);
  BUFF I129 (o_0r1[31:31], joint_0[31:31]);
  BUFF I130 (i_0a, o_0a);
  BUFF I131 (i_1a, o_0a);
endmodule

// tkj32m30_2 TeakJ [Many [30,2],One 32]
module tkj32m30_2 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [29:0] i_0r0;
  input [29:0] i_0r1;
  output i_0a;
  input [1:0] i_1r0;
  input [1:0] i_1r1;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [31:0] joinf_0;
  wire [31:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_1r0[0:0]);
  BUFF I31 (joinf_0[31:31], i_1r0[1:1]);
  BUFF I32 (joint_0[0:0], i_0r1[0:0]);
  BUFF I33 (joint_0[1:1], i_0r1[1:1]);
  BUFF I34 (joint_0[2:2], i_0r1[2:2]);
  BUFF I35 (joint_0[3:3], i_0r1[3:3]);
  BUFF I36 (joint_0[4:4], i_0r1[4:4]);
  BUFF I37 (joint_0[5:5], i_0r1[5:5]);
  BUFF I38 (joint_0[6:6], i_0r1[6:6]);
  BUFF I39 (joint_0[7:7], i_0r1[7:7]);
  BUFF I40 (joint_0[8:8], i_0r1[8:8]);
  BUFF I41 (joint_0[9:9], i_0r1[9:9]);
  BUFF I42 (joint_0[10:10], i_0r1[10:10]);
  BUFF I43 (joint_0[11:11], i_0r1[11:11]);
  BUFF I44 (joint_0[12:12], i_0r1[12:12]);
  BUFF I45 (joint_0[13:13], i_0r1[13:13]);
  BUFF I46 (joint_0[14:14], i_0r1[14:14]);
  BUFF I47 (joint_0[15:15], i_0r1[15:15]);
  BUFF I48 (joint_0[16:16], i_0r1[16:16]);
  BUFF I49 (joint_0[17:17], i_0r1[17:17]);
  BUFF I50 (joint_0[18:18], i_0r1[18:18]);
  BUFF I51 (joint_0[19:19], i_0r1[19:19]);
  BUFF I52 (joint_0[20:20], i_0r1[20:20]);
  BUFF I53 (joint_0[21:21], i_0r1[21:21]);
  BUFF I54 (joint_0[22:22], i_0r1[22:22]);
  BUFF I55 (joint_0[23:23], i_0r1[23:23]);
  BUFF I56 (joint_0[24:24], i_0r1[24:24]);
  BUFF I57 (joint_0[25:25], i_0r1[25:25]);
  BUFF I58 (joint_0[26:26], i_0r1[26:26]);
  BUFF I59 (joint_0[27:27], i_0r1[27:27]);
  BUFF I60 (joint_0[28:28], i_0r1[28:28]);
  BUFF I61 (joint_0[29:29], i_0r1[29:29]);
  BUFF I62 (joint_0[30:30], i_1r1[0:0]);
  BUFF I63 (joint_0[31:31], i_1r1[1:1]);
  OR2 I64 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I65 (icomplete_0, dcomplete_0);
  C2 I66 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I67 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I68 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I69 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I70 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I71 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I72 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I73 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I74 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I75 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I76 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I77 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I78 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I79 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I80 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I81 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I82 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I83 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I84 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I85 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I86 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I87 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I88 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I89 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I90 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I91 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I92 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I93 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I94 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I95 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I96 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I97 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I98 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I99 (o_0r1[1:1], joint_0[1:1]);
  BUFF I100 (o_0r1[2:2], joint_0[2:2]);
  BUFF I101 (o_0r1[3:3], joint_0[3:3]);
  BUFF I102 (o_0r1[4:4], joint_0[4:4]);
  BUFF I103 (o_0r1[5:5], joint_0[5:5]);
  BUFF I104 (o_0r1[6:6], joint_0[6:6]);
  BUFF I105 (o_0r1[7:7], joint_0[7:7]);
  BUFF I106 (o_0r1[8:8], joint_0[8:8]);
  BUFF I107 (o_0r1[9:9], joint_0[9:9]);
  BUFF I108 (o_0r1[10:10], joint_0[10:10]);
  BUFF I109 (o_0r1[11:11], joint_0[11:11]);
  BUFF I110 (o_0r1[12:12], joint_0[12:12]);
  BUFF I111 (o_0r1[13:13], joint_0[13:13]);
  BUFF I112 (o_0r1[14:14], joint_0[14:14]);
  BUFF I113 (o_0r1[15:15], joint_0[15:15]);
  BUFF I114 (o_0r1[16:16], joint_0[16:16]);
  BUFF I115 (o_0r1[17:17], joint_0[17:17]);
  BUFF I116 (o_0r1[18:18], joint_0[18:18]);
  BUFF I117 (o_0r1[19:19], joint_0[19:19]);
  BUFF I118 (o_0r1[20:20], joint_0[20:20]);
  BUFF I119 (o_0r1[21:21], joint_0[21:21]);
  BUFF I120 (o_0r1[22:22], joint_0[22:22]);
  BUFF I121 (o_0r1[23:23], joint_0[23:23]);
  BUFF I122 (o_0r1[24:24], joint_0[24:24]);
  BUFF I123 (o_0r1[25:25], joint_0[25:25]);
  BUFF I124 (o_0r1[26:26], joint_0[26:26]);
  BUFF I125 (o_0r1[27:27], joint_0[27:27]);
  BUFF I126 (o_0r1[28:28], joint_0[28:28]);
  BUFF I127 (o_0r1[29:29], joint_0[29:29]);
  BUFF I128 (o_0r1[30:30], joint_0[30:30]);
  BUFF I129 (o_0r1[31:31], joint_0[31:31]);
  BUFF I130 (i_0a, o_0a);
  BUFF I131 (i_1a, o_0a);
endmodule

// tko0m2_1nm2b3 TeakO [
//     (1,TeakOConstant 2 3)] [One 0,One 2]
module tko0m2_1nm2b3 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  BUFF I1 (o_0r1[1:1], i_0r);
  GND I2 (o_0r0[0:0]);
  GND I3 (o_0r0[1:1]);
  BUFF I4 (i_0a, o_0a);
endmodule

// tkvi32_wo0w32_ro0w32o0w30o2w30o2w30 TeakV "i" 32 [] [0] [0,0,2,2] [Many [32],Many [0],Many [0,0,0,0]
//   ,Many [32,30,30,30]]
module tkvi32_wo0w32_ro0w32o0w30o2w30o2w30 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [29:0] rd_1r0;
  output [29:0] rd_1r1;
  input rd_1a;
  output [29:0] rd_2r0;
  output [29:0] rd_2r1;
  input rd_2a;
  output [29:0] rd_3r0;
  output [29:0] rd_3r1;
  input rd_3a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [2:0] simp6521_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_2r0[0:0], df_0[2:2], rg_2r);
  AND2 I487 (rd_2r0[1:1], df_0[3:3], rg_2r);
  AND2 I488 (rd_2r0[2:2], df_0[4:4], rg_2r);
  AND2 I489 (rd_2r0[3:3], df_0[5:5], rg_2r);
  AND2 I490 (rd_2r0[4:4], df_0[6:6], rg_2r);
  AND2 I491 (rd_2r0[5:5], df_0[7:7], rg_2r);
  AND2 I492 (rd_2r0[6:6], df_0[8:8], rg_2r);
  AND2 I493 (rd_2r0[7:7], df_0[9:9], rg_2r);
  AND2 I494 (rd_2r0[8:8], df_0[10:10], rg_2r);
  AND2 I495 (rd_2r0[9:9], df_0[11:11], rg_2r);
  AND2 I496 (rd_2r0[10:10], df_0[12:12], rg_2r);
  AND2 I497 (rd_2r0[11:11], df_0[13:13], rg_2r);
  AND2 I498 (rd_2r0[12:12], df_0[14:14], rg_2r);
  AND2 I499 (rd_2r0[13:13], df_0[15:15], rg_2r);
  AND2 I500 (rd_2r0[14:14], df_0[16:16], rg_2r);
  AND2 I501 (rd_2r0[15:15], df_0[17:17], rg_2r);
  AND2 I502 (rd_2r0[16:16], df_0[18:18], rg_2r);
  AND2 I503 (rd_2r0[17:17], df_0[19:19], rg_2r);
  AND2 I504 (rd_2r0[18:18], df_0[20:20], rg_2r);
  AND2 I505 (rd_2r0[19:19], df_0[21:21], rg_2r);
  AND2 I506 (rd_2r0[20:20], df_0[22:22], rg_2r);
  AND2 I507 (rd_2r0[21:21], df_0[23:23], rg_2r);
  AND2 I508 (rd_2r0[22:22], df_0[24:24], rg_2r);
  AND2 I509 (rd_2r0[23:23], df_0[25:25], rg_2r);
  AND2 I510 (rd_2r0[24:24], df_0[26:26], rg_2r);
  AND2 I511 (rd_2r0[25:25], df_0[27:27], rg_2r);
  AND2 I512 (rd_2r0[26:26], df_0[28:28], rg_2r);
  AND2 I513 (rd_2r0[27:27], df_0[29:29], rg_2r);
  AND2 I514 (rd_2r0[28:28], df_0[30:30], rg_2r);
  AND2 I515 (rd_2r0[29:29], df_0[31:31], rg_2r);
  AND2 I516 (rd_3r0[0:0], df_0[2:2], rg_3r);
  AND2 I517 (rd_3r0[1:1], df_0[3:3], rg_3r);
  AND2 I518 (rd_3r0[2:2], df_0[4:4], rg_3r);
  AND2 I519 (rd_3r0[3:3], df_0[5:5], rg_3r);
  AND2 I520 (rd_3r0[4:4], df_0[6:6], rg_3r);
  AND2 I521 (rd_3r0[5:5], df_0[7:7], rg_3r);
  AND2 I522 (rd_3r0[6:6], df_0[8:8], rg_3r);
  AND2 I523 (rd_3r0[7:7], df_0[9:9], rg_3r);
  AND2 I524 (rd_3r0[8:8], df_0[10:10], rg_3r);
  AND2 I525 (rd_3r0[9:9], df_0[11:11], rg_3r);
  AND2 I526 (rd_3r0[10:10], df_0[12:12], rg_3r);
  AND2 I527 (rd_3r0[11:11], df_0[13:13], rg_3r);
  AND2 I528 (rd_3r0[12:12], df_0[14:14], rg_3r);
  AND2 I529 (rd_3r0[13:13], df_0[15:15], rg_3r);
  AND2 I530 (rd_3r0[14:14], df_0[16:16], rg_3r);
  AND2 I531 (rd_3r0[15:15], df_0[17:17], rg_3r);
  AND2 I532 (rd_3r0[16:16], df_0[18:18], rg_3r);
  AND2 I533 (rd_3r0[17:17], df_0[19:19], rg_3r);
  AND2 I534 (rd_3r0[18:18], df_0[20:20], rg_3r);
  AND2 I535 (rd_3r0[19:19], df_0[21:21], rg_3r);
  AND2 I536 (rd_3r0[20:20], df_0[22:22], rg_3r);
  AND2 I537 (rd_3r0[21:21], df_0[23:23], rg_3r);
  AND2 I538 (rd_3r0[22:22], df_0[24:24], rg_3r);
  AND2 I539 (rd_3r0[23:23], df_0[25:25], rg_3r);
  AND2 I540 (rd_3r0[24:24], df_0[26:26], rg_3r);
  AND2 I541 (rd_3r0[25:25], df_0[27:27], rg_3r);
  AND2 I542 (rd_3r0[26:26], df_0[28:28], rg_3r);
  AND2 I543 (rd_3r0[27:27], df_0[29:29], rg_3r);
  AND2 I544 (rd_3r0[28:28], df_0[30:30], rg_3r);
  AND2 I545 (rd_3r0[29:29], df_0[31:31], rg_3r);
  AND2 I546 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I547 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I548 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I549 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I550 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I551 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I552 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I553 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I554 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I555 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I556 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I557 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I558 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I559 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I560 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I561 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I562 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I563 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I564 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I565 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I566 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I567 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I568 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I569 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I570 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I571 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I572 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I573 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I574 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I575 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I576 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I577 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I578 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I579 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I580 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I581 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I582 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I583 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I584 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I585 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I586 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I587 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I588 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I589 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I590 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I591 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I592 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I593 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I594 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I595 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I596 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I597 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I598 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I599 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I600 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I601 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I602 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I603 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I604 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I605 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I606 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I607 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I608 (rd_2r1[0:0], dt_0[2:2], rg_2r);
  AND2 I609 (rd_2r1[1:1], dt_0[3:3], rg_2r);
  AND2 I610 (rd_2r1[2:2], dt_0[4:4], rg_2r);
  AND2 I611 (rd_2r1[3:3], dt_0[5:5], rg_2r);
  AND2 I612 (rd_2r1[4:4], dt_0[6:6], rg_2r);
  AND2 I613 (rd_2r1[5:5], dt_0[7:7], rg_2r);
  AND2 I614 (rd_2r1[6:6], dt_0[8:8], rg_2r);
  AND2 I615 (rd_2r1[7:7], dt_0[9:9], rg_2r);
  AND2 I616 (rd_2r1[8:8], dt_0[10:10], rg_2r);
  AND2 I617 (rd_2r1[9:9], dt_0[11:11], rg_2r);
  AND2 I618 (rd_2r1[10:10], dt_0[12:12], rg_2r);
  AND2 I619 (rd_2r1[11:11], dt_0[13:13], rg_2r);
  AND2 I620 (rd_2r1[12:12], dt_0[14:14], rg_2r);
  AND2 I621 (rd_2r1[13:13], dt_0[15:15], rg_2r);
  AND2 I622 (rd_2r1[14:14], dt_0[16:16], rg_2r);
  AND2 I623 (rd_2r1[15:15], dt_0[17:17], rg_2r);
  AND2 I624 (rd_2r1[16:16], dt_0[18:18], rg_2r);
  AND2 I625 (rd_2r1[17:17], dt_0[19:19], rg_2r);
  AND2 I626 (rd_2r1[18:18], dt_0[20:20], rg_2r);
  AND2 I627 (rd_2r1[19:19], dt_0[21:21], rg_2r);
  AND2 I628 (rd_2r1[20:20], dt_0[22:22], rg_2r);
  AND2 I629 (rd_2r1[21:21], dt_0[23:23], rg_2r);
  AND2 I630 (rd_2r1[22:22], dt_0[24:24], rg_2r);
  AND2 I631 (rd_2r1[23:23], dt_0[25:25], rg_2r);
  AND2 I632 (rd_2r1[24:24], dt_0[26:26], rg_2r);
  AND2 I633 (rd_2r1[25:25], dt_0[27:27], rg_2r);
  AND2 I634 (rd_2r1[26:26], dt_0[28:28], rg_2r);
  AND2 I635 (rd_2r1[27:27], dt_0[29:29], rg_2r);
  AND2 I636 (rd_2r1[28:28], dt_0[30:30], rg_2r);
  AND2 I637 (rd_2r1[29:29], dt_0[31:31], rg_2r);
  AND2 I638 (rd_3r1[0:0], dt_0[2:2], rg_3r);
  AND2 I639 (rd_3r1[1:1], dt_0[3:3], rg_3r);
  AND2 I640 (rd_3r1[2:2], dt_0[4:4], rg_3r);
  AND2 I641 (rd_3r1[3:3], dt_0[5:5], rg_3r);
  AND2 I642 (rd_3r1[4:4], dt_0[6:6], rg_3r);
  AND2 I643 (rd_3r1[5:5], dt_0[7:7], rg_3r);
  AND2 I644 (rd_3r1[6:6], dt_0[8:8], rg_3r);
  AND2 I645 (rd_3r1[7:7], dt_0[9:9], rg_3r);
  AND2 I646 (rd_3r1[8:8], dt_0[10:10], rg_3r);
  AND2 I647 (rd_3r1[9:9], dt_0[11:11], rg_3r);
  AND2 I648 (rd_3r1[10:10], dt_0[12:12], rg_3r);
  AND2 I649 (rd_3r1[11:11], dt_0[13:13], rg_3r);
  AND2 I650 (rd_3r1[12:12], dt_0[14:14], rg_3r);
  AND2 I651 (rd_3r1[13:13], dt_0[15:15], rg_3r);
  AND2 I652 (rd_3r1[14:14], dt_0[16:16], rg_3r);
  AND2 I653 (rd_3r1[15:15], dt_0[17:17], rg_3r);
  AND2 I654 (rd_3r1[16:16], dt_0[18:18], rg_3r);
  AND2 I655 (rd_3r1[17:17], dt_0[19:19], rg_3r);
  AND2 I656 (rd_3r1[18:18], dt_0[20:20], rg_3r);
  AND2 I657 (rd_3r1[19:19], dt_0[21:21], rg_3r);
  AND2 I658 (rd_3r1[20:20], dt_0[22:22], rg_3r);
  AND2 I659 (rd_3r1[21:21], dt_0[23:23], rg_3r);
  AND2 I660 (rd_3r1[22:22], dt_0[24:24], rg_3r);
  AND2 I661 (rd_3r1[23:23], dt_0[25:25], rg_3r);
  AND2 I662 (rd_3r1[24:24], dt_0[26:26], rg_3r);
  AND2 I663 (rd_3r1[25:25], dt_0[27:27], rg_3r);
  AND2 I664 (rd_3r1[26:26], dt_0[28:28], rg_3r);
  AND2 I665 (rd_3r1[27:27], dt_0[29:29], rg_3r);
  AND2 I666 (rd_3r1[28:28], dt_0[30:30], rg_3r);
  AND2 I667 (rd_3r1[29:29], dt_0[31:31], rg_3r);
  NOR3 I668 (simp6521_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I669 (simp6521_0[1:1], rg_3r, rg_0a, rg_1a);
  NOR2 I670 (simp6521_0[2:2], rg_2a, rg_3a);
  NAND3 I671 (anyread_0, simp6521_0[0:0], simp6521_0[1:1], simp6521_0[2:2]);
  BUFF I672 (wg_0a, wd_0a);
  BUFF I673 (rg_0a, rd_0a);
  BUFF I674 (rg_1a, rd_1a);
  BUFF I675 (rg_2a, rd_2a);
  BUFF I676 (rg_3a, rd_3a);
endmodule

// tkm4x32b TeakM [Many [32,32,32,32],One 32]
module tkm4x32b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  input [31:0] i_2r0;
  input [31:0] i_2r1;
  output i_2a;
  input [31:0] i_3r0;
  input [31:0] i_3r1;
  output i_3a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire [31:0] gfint_0;
  wire [31:0] gfint_1;
  wire [31:0] gfint_2;
  wire [31:0] gfint_3;
  wire [31:0] gtint_0;
  wire [31:0] gtint_1;
  wire [31:0] gtint_2;
  wire [31:0] gtint_3;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire icomp_3;
  wire nchosen_0;
  wire [1:0] simp181_0;
  wire [1:0] simp191_0;
  wire [1:0] simp201_0;
  wire [1:0] simp211_0;
  wire [1:0] simp221_0;
  wire [1:0] simp231_0;
  wire [1:0] simp241_0;
  wire [1:0] simp251_0;
  wire [1:0] simp261_0;
  wire [1:0] simp271_0;
  wire [1:0] simp281_0;
  wire [1:0] simp291_0;
  wire [1:0] simp301_0;
  wire [1:0] simp311_0;
  wire [1:0] simp321_0;
  wire [1:0] simp331_0;
  wire [1:0] simp341_0;
  wire [1:0] simp351_0;
  wire [1:0] simp361_0;
  wire [1:0] simp371_0;
  wire [1:0] simp381_0;
  wire [1:0] simp391_0;
  wire [1:0] simp401_0;
  wire [1:0] simp411_0;
  wire [1:0] simp421_0;
  wire [1:0] simp431_0;
  wire [1:0] simp441_0;
  wire [1:0] simp451_0;
  wire [1:0] simp461_0;
  wire [1:0] simp471_0;
  wire [1:0] simp481_0;
  wire [1:0] simp491_0;
  wire [1:0] simp501_0;
  wire [1:0] simp511_0;
  wire [1:0] simp521_0;
  wire [1:0] simp531_0;
  wire [1:0] simp541_0;
  wire [1:0] simp551_0;
  wire [1:0] simp561_0;
  wire [1:0] simp571_0;
  wire [1:0] simp581_0;
  wire [1:0] simp591_0;
  wire [1:0] simp601_0;
  wire [1:0] simp611_0;
  wire [1:0] simp621_0;
  wire [1:0] simp631_0;
  wire [1:0] simp641_0;
  wire [1:0] simp651_0;
  wire [1:0] simp661_0;
  wire [1:0] simp671_0;
  wire [1:0] simp681_0;
  wire [1:0] simp691_0;
  wire [1:0] simp701_0;
  wire [1:0] simp711_0;
  wire [1:0] simp721_0;
  wire [1:0] simp731_0;
  wire [1:0] simp741_0;
  wire [1:0] simp751_0;
  wire [1:0] simp761_0;
  wire [1:0] simp771_0;
  wire [1:0] simp781_0;
  wire [1:0] simp791_0;
  wire [1:0] simp801_0;
  wire [1:0] simp811_0;
  wire [31:0] comp0_0;
  wire [10:0] simp3711_0;
  wire [3:0] simp3712_0;
  wire [1:0] simp3713_0;
  wire [31:0] comp1_0;
  wire [10:0] simp4051_0;
  wire [3:0] simp4052_0;
  wire [1:0] simp4053_0;
  wire [31:0] comp2_0;
  wire [10:0] simp4391_0;
  wire [3:0] simp4392_0;
  wire [1:0] simp4393_0;
  wire [31:0] comp3_0;
  wire [10:0] simp4731_0;
  wire [3:0] simp4732_0;
  wire [1:0] simp4733_0;
  wire [1:0] simp4781_0;
  NOR3 I0 (simp181_0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  INV I1 (simp181_0[1:1], gfint_3[0:0]);
  NAND2 I2 (o_0r0[0:0], simp181_0[0:0], simp181_0[1:1]);
  NOR3 I3 (simp191_0[0:0], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  INV I4 (simp191_0[1:1], gfint_3[1:1]);
  NAND2 I5 (o_0r0[1:1], simp191_0[0:0], simp191_0[1:1]);
  NOR3 I6 (simp201_0[0:0], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  INV I7 (simp201_0[1:1], gfint_3[2:2]);
  NAND2 I8 (o_0r0[2:2], simp201_0[0:0], simp201_0[1:1]);
  NOR3 I9 (simp211_0[0:0], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  INV I10 (simp211_0[1:1], gfint_3[3:3]);
  NAND2 I11 (o_0r0[3:3], simp211_0[0:0], simp211_0[1:1]);
  NOR3 I12 (simp221_0[0:0], gfint_0[4:4], gfint_1[4:4], gfint_2[4:4]);
  INV I13 (simp221_0[1:1], gfint_3[4:4]);
  NAND2 I14 (o_0r0[4:4], simp221_0[0:0], simp221_0[1:1]);
  NOR3 I15 (simp231_0[0:0], gfint_0[5:5], gfint_1[5:5], gfint_2[5:5]);
  INV I16 (simp231_0[1:1], gfint_3[5:5]);
  NAND2 I17 (o_0r0[5:5], simp231_0[0:0], simp231_0[1:1]);
  NOR3 I18 (simp241_0[0:0], gfint_0[6:6], gfint_1[6:6], gfint_2[6:6]);
  INV I19 (simp241_0[1:1], gfint_3[6:6]);
  NAND2 I20 (o_0r0[6:6], simp241_0[0:0], simp241_0[1:1]);
  NOR3 I21 (simp251_0[0:0], gfint_0[7:7], gfint_1[7:7], gfint_2[7:7]);
  INV I22 (simp251_0[1:1], gfint_3[7:7]);
  NAND2 I23 (o_0r0[7:7], simp251_0[0:0], simp251_0[1:1]);
  NOR3 I24 (simp261_0[0:0], gfint_0[8:8], gfint_1[8:8], gfint_2[8:8]);
  INV I25 (simp261_0[1:1], gfint_3[8:8]);
  NAND2 I26 (o_0r0[8:8], simp261_0[0:0], simp261_0[1:1]);
  NOR3 I27 (simp271_0[0:0], gfint_0[9:9], gfint_1[9:9], gfint_2[9:9]);
  INV I28 (simp271_0[1:1], gfint_3[9:9]);
  NAND2 I29 (o_0r0[9:9], simp271_0[0:0], simp271_0[1:1]);
  NOR3 I30 (simp281_0[0:0], gfint_0[10:10], gfint_1[10:10], gfint_2[10:10]);
  INV I31 (simp281_0[1:1], gfint_3[10:10]);
  NAND2 I32 (o_0r0[10:10], simp281_0[0:0], simp281_0[1:1]);
  NOR3 I33 (simp291_0[0:0], gfint_0[11:11], gfint_1[11:11], gfint_2[11:11]);
  INV I34 (simp291_0[1:1], gfint_3[11:11]);
  NAND2 I35 (o_0r0[11:11], simp291_0[0:0], simp291_0[1:1]);
  NOR3 I36 (simp301_0[0:0], gfint_0[12:12], gfint_1[12:12], gfint_2[12:12]);
  INV I37 (simp301_0[1:1], gfint_3[12:12]);
  NAND2 I38 (o_0r0[12:12], simp301_0[0:0], simp301_0[1:1]);
  NOR3 I39 (simp311_0[0:0], gfint_0[13:13], gfint_1[13:13], gfint_2[13:13]);
  INV I40 (simp311_0[1:1], gfint_3[13:13]);
  NAND2 I41 (o_0r0[13:13], simp311_0[0:0], simp311_0[1:1]);
  NOR3 I42 (simp321_0[0:0], gfint_0[14:14], gfint_1[14:14], gfint_2[14:14]);
  INV I43 (simp321_0[1:1], gfint_3[14:14]);
  NAND2 I44 (o_0r0[14:14], simp321_0[0:0], simp321_0[1:1]);
  NOR3 I45 (simp331_0[0:0], gfint_0[15:15], gfint_1[15:15], gfint_2[15:15]);
  INV I46 (simp331_0[1:1], gfint_3[15:15]);
  NAND2 I47 (o_0r0[15:15], simp331_0[0:0], simp331_0[1:1]);
  NOR3 I48 (simp341_0[0:0], gfint_0[16:16], gfint_1[16:16], gfint_2[16:16]);
  INV I49 (simp341_0[1:1], gfint_3[16:16]);
  NAND2 I50 (o_0r0[16:16], simp341_0[0:0], simp341_0[1:1]);
  NOR3 I51 (simp351_0[0:0], gfint_0[17:17], gfint_1[17:17], gfint_2[17:17]);
  INV I52 (simp351_0[1:1], gfint_3[17:17]);
  NAND2 I53 (o_0r0[17:17], simp351_0[0:0], simp351_0[1:1]);
  NOR3 I54 (simp361_0[0:0], gfint_0[18:18], gfint_1[18:18], gfint_2[18:18]);
  INV I55 (simp361_0[1:1], gfint_3[18:18]);
  NAND2 I56 (o_0r0[18:18], simp361_0[0:0], simp361_0[1:1]);
  NOR3 I57 (simp371_0[0:0], gfint_0[19:19], gfint_1[19:19], gfint_2[19:19]);
  INV I58 (simp371_0[1:1], gfint_3[19:19]);
  NAND2 I59 (o_0r0[19:19], simp371_0[0:0], simp371_0[1:1]);
  NOR3 I60 (simp381_0[0:0], gfint_0[20:20], gfint_1[20:20], gfint_2[20:20]);
  INV I61 (simp381_0[1:1], gfint_3[20:20]);
  NAND2 I62 (o_0r0[20:20], simp381_0[0:0], simp381_0[1:1]);
  NOR3 I63 (simp391_0[0:0], gfint_0[21:21], gfint_1[21:21], gfint_2[21:21]);
  INV I64 (simp391_0[1:1], gfint_3[21:21]);
  NAND2 I65 (o_0r0[21:21], simp391_0[0:0], simp391_0[1:1]);
  NOR3 I66 (simp401_0[0:0], gfint_0[22:22], gfint_1[22:22], gfint_2[22:22]);
  INV I67 (simp401_0[1:1], gfint_3[22:22]);
  NAND2 I68 (o_0r0[22:22], simp401_0[0:0], simp401_0[1:1]);
  NOR3 I69 (simp411_0[0:0], gfint_0[23:23], gfint_1[23:23], gfint_2[23:23]);
  INV I70 (simp411_0[1:1], gfint_3[23:23]);
  NAND2 I71 (o_0r0[23:23], simp411_0[0:0], simp411_0[1:1]);
  NOR3 I72 (simp421_0[0:0], gfint_0[24:24], gfint_1[24:24], gfint_2[24:24]);
  INV I73 (simp421_0[1:1], gfint_3[24:24]);
  NAND2 I74 (o_0r0[24:24], simp421_0[0:0], simp421_0[1:1]);
  NOR3 I75 (simp431_0[0:0], gfint_0[25:25], gfint_1[25:25], gfint_2[25:25]);
  INV I76 (simp431_0[1:1], gfint_3[25:25]);
  NAND2 I77 (o_0r0[25:25], simp431_0[0:0], simp431_0[1:1]);
  NOR3 I78 (simp441_0[0:0], gfint_0[26:26], gfint_1[26:26], gfint_2[26:26]);
  INV I79 (simp441_0[1:1], gfint_3[26:26]);
  NAND2 I80 (o_0r0[26:26], simp441_0[0:0], simp441_0[1:1]);
  NOR3 I81 (simp451_0[0:0], gfint_0[27:27], gfint_1[27:27], gfint_2[27:27]);
  INV I82 (simp451_0[1:1], gfint_3[27:27]);
  NAND2 I83 (o_0r0[27:27], simp451_0[0:0], simp451_0[1:1]);
  NOR3 I84 (simp461_0[0:0], gfint_0[28:28], gfint_1[28:28], gfint_2[28:28]);
  INV I85 (simp461_0[1:1], gfint_3[28:28]);
  NAND2 I86 (o_0r0[28:28], simp461_0[0:0], simp461_0[1:1]);
  NOR3 I87 (simp471_0[0:0], gfint_0[29:29], gfint_1[29:29], gfint_2[29:29]);
  INV I88 (simp471_0[1:1], gfint_3[29:29]);
  NAND2 I89 (o_0r0[29:29], simp471_0[0:0], simp471_0[1:1]);
  NOR3 I90 (simp481_0[0:0], gfint_0[30:30], gfint_1[30:30], gfint_2[30:30]);
  INV I91 (simp481_0[1:1], gfint_3[30:30]);
  NAND2 I92 (o_0r0[30:30], simp481_0[0:0], simp481_0[1:1]);
  NOR3 I93 (simp491_0[0:0], gfint_0[31:31], gfint_1[31:31], gfint_2[31:31]);
  INV I94 (simp491_0[1:1], gfint_3[31:31]);
  NAND2 I95 (o_0r0[31:31], simp491_0[0:0], simp491_0[1:1]);
  NOR3 I96 (simp501_0[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  INV I97 (simp501_0[1:1], gtint_3[0:0]);
  NAND2 I98 (o_0r1[0:0], simp501_0[0:0], simp501_0[1:1]);
  NOR3 I99 (simp511_0[0:0], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  INV I100 (simp511_0[1:1], gtint_3[1:1]);
  NAND2 I101 (o_0r1[1:1], simp511_0[0:0], simp511_0[1:1]);
  NOR3 I102 (simp521_0[0:0], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  INV I103 (simp521_0[1:1], gtint_3[2:2]);
  NAND2 I104 (o_0r1[2:2], simp521_0[0:0], simp521_0[1:1]);
  NOR3 I105 (simp531_0[0:0], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  INV I106 (simp531_0[1:1], gtint_3[3:3]);
  NAND2 I107 (o_0r1[3:3], simp531_0[0:0], simp531_0[1:1]);
  NOR3 I108 (simp541_0[0:0], gtint_0[4:4], gtint_1[4:4], gtint_2[4:4]);
  INV I109 (simp541_0[1:1], gtint_3[4:4]);
  NAND2 I110 (o_0r1[4:4], simp541_0[0:0], simp541_0[1:1]);
  NOR3 I111 (simp551_0[0:0], gtint_0[5:5], gtint_1[5:5], gtint_2[5:5]);
  INV I112 (simp551_0[1:1], gtint_3[5:5]);
  NAND2 I113 (o_0r1[5:5], simp551_0[0:0], simp551_0[1:1]);
  NOR3 I114 (simp561_0[0:0], gtint_0[6:6], gtint_1[6:6], gtint_2[6:6]);
  INV I115 (simp561_0[1:1], gtint_3[6:6]);
  NAND2 I116 (o_0r1[6:6], simp561_0[0:0], simp561_0[1:1]);
  NOR3 I117 (simp571_0[0:0], gtint_0[7:7], gtint_1[7:7], gtint_2[7:7]);
  INV I118 (simp571_0[1:1], gtint_3[7:7]);
  NAND2 I119 (o_0r1[7:7], simp571_0[0:0], simp571_0[1:1]);
  NOR3 I120 (simp581_0[0:0], gtint_0[8:8], gtint_1[8:8], gtint_2[8:8]);
  INV I121 (simp581_0[1:1], gtint_3[8:8]);
  NAND2 I122 (o_0r1[8:8], simp581_0[0:0], simp581_0[1:1]);
  NOR3 I123 (simp591_0[0:0], gtint_0[9:9], gtint_1[9:9], gtint_2[9:9]);
  INV I124 (simp591_0[1:1], gtint_3[9:9]);
  NAND2 I125 (o_0r1[9:9], simp591_0[0:0], simp591_0[1:1]);
  NOR3 I126 (simp601_0[0:0], gtint_0[10:10], gtint_1[10:10], gtint_2[10:10]);
  INV I127 (simp601_0[1:1], gtint_3[10:10]);
  NAND2 I128 (o_0r1[10:10], simp601_0[0:0], simp601_0[1:1]);
  NOR3 I129 (simp611_0[0:0], gtint_0[11:11], gtint_1[11:11], gtint_2[11:11]);
  INV I130 (simp611_0[1:1], gtint_3[11:11]);
  NAND2 I131 (o_0r1[11:11], simp611_0[0:0], simp611_0[1:1]);
  NOR3 I132 (simp621_0[0:0], gtint_0[12:12], gtint_1[12:12], gtint_2[12:12]);
  INV I133 (simp621_0[1:1], gtint_3[12:12]);
  NAND2 I134 (o_0r1[12:12], simp621_0[0:0], simp621_0[1:1]);
  NOR3 I135 (simp631_0[0:0], gtint_0[13:13], gtint_1[13:13], gtint_2[13:13]);
  INV I136 (simp631_0[1:1], gtint_3[13:13]);
  NAND2 I137 (o_0r1[13:13], simp631_0[0:0], simp631_0[1:1]);
  NOR3 I138 (simp641_0[0:0], gtint_0[14:14], gtint_1[14:14], gtint_2[14:14]);
  INV I139 (simp641_0[1:1], gtint_3[14:14]);
  NAND2 I140 (o_0r1[14:14], simp641_0[0:0], simp641_0[1:1]);
  NOR3 I141 (simp651_0[0:0], gtint_0[15:15], gtint_1[15:15], gtint_2[15:15]);
  INV I142 (simp651_0[1:1], gtint_3[15:15]);
  NAND2 I143 (o_0r1[15:15], simp651_0[0:0], simp651_0[1:1]);
  NOR3 I144 (simp661_0[0:0], gtint_0[16:16], gtint_1[16:16], gtint_2[16:16]);
  INV I145 (simp661_0[1:1], gtint_3[16:16]);
  NAND2 I146 (o_0r1[16:16], simp661_0[0:0], simp661_0[1:1]);
  NOR3 I147 (simp671_0[0:0], gtint_0[17:17], gtint_1[17:17], gtint_2[17:17]);
  INV I148 (simp671_0[1:1], gtint_3[17:17]);
  NAND2 I149 (o_0r1[17:17], simp671_0[0:0], simp671_0[1:1]);
  NOR3 I150 (simp681_0[0:0], gtint_0[18:18], gtint_1[18:18], gtint_2[18:18]);
  INV I151 (simp681_0[1:1], gtint_3[18:18]);
  NAND2 I152 (o_0r1[18:18], simp681_0[0:0], simp681_0[1:1]);
  NOR3 I153 (simp691_0[0:0], gtint_0[19:19], gtint_1[19:19], gtint_2[19:19]);
  INV I154 (simp691_0[1:1], gtint_3[19:19]);
  NAND2 I155 (o_0r1[19:19], simp691_0[0:0], simp691_0[1:1]);
  NOR3 I156 (simp701_0[0:0], gtint_0[20:20], gtint_1[20:20], gtint_2[20:20]);
  INV I157 (simp701_0[1:1], gtint_3[20:20]);
  NAND2 I158 (o_0r1[20:20], simp701_0[0:0], simp701_0[1:1]);
  NOR3 I159 (simp711_0[0:0], gtint_0[21:21], gtint_1[21:21], gtint_2[21:21]);
  INV I160 (simp711_0[1:1], gtint_3[21:21]);
  NAND2 I161 (o_0r1[21:21], simp711_0[0:0], simp711_0[1:1]);
  NOR3 I162 (simp721_0[0:0], gtint_0[22:22], gtint_1[22:22], gtint_2[22:22]);
  INV I163 (simp721_0[1:1], gtint_3[22:22]);
  NAND2 I164 (o_0r1[22:22], simp721_0[0:0], simp721_0[1:1]);
  NOR3 I165 (simp731_0[0:0], gtint_0[23:23], gtint_1[23:23], gtint_2[23:23]);
  INV I166 (simp731_0[1:1], gtint_3[23:23]);
  NAND2 I167 (o_0r1[23:23], simp731_0[0:0], simp731_0[1:1]);
  NOR3 I168 (simp741_0[0:0], gtint_0[24:24], gtint_1[24:24], gtint_2[24:24]);
  INV I169 (simp741_0[1:1], gtint_3[24:24]);
  NAND2 I170 (o_0r1[24:24], simp741_0[0:0], simp741_0[1:1]);
  NOR3 I171 (simp751_0[0:0], gtint_0[25:25], gtint_1[25:25], gtint_2[25:25]);
  INV I172 (simp751_0[1:1], gtint_3[25:25]);
  NAND2 I173 (o_0r1[25:25], simp751_0[0:0], simp751_0[1:1]);
  NOR3 I174 (simp761_0[0:0], gtint_0[26:26], gtint_1[26:26], gtint_2[26:26]);
  INV I175 (simp761_0[1:1], gtint_3[26:26]);
  NAND2 I176 (o_0r1[26:26], simp761_0[0:0], simp761_0[1:1]);
  NOR3 I177 (simp771_0[0:0], gtint_0[27:27], gtint_1[27:27], gtint_2[27:27]);
  INV I178 (simp771_0[1:1], gtint_3[27:27]);
  NAND2 I179 (o_0r1[27:27], simp771_0[0:0], simp771_0[1:1]);
  NOR3 I180 (simp781_0[0:0], gtint_0[28:28], gtint_1[28:28], gtint_2[28:28]);
  INV I181 (simp781_0[1:1], gtint_3[28:28]);
  NAND2 I182 (o_0r1[28:28], simp781_0[0:0], simp781_0[1:1]);
  NOR3 I183 (simp791_0[0:0], gtint_0[29:29], gtint_1[29:29], gtint_2[29:29]);
  INV I184 (simp791_0[1:1], gtint_3[29:29]);
  NAND2 I185 (o_0r1[29:29], simp791_0[0:0], simp791_0[1:1]);
  NOR3 I186 (simp801_0[0:0], gtint_0[30:30], gtint_1[30:30], gtint_2[30:30]);
  INV I187 (simp801_0[1:1], gtint_3[30:30]);
  NAND2 I188 (o_0r1[30:30], simp801_0[0:0], simp801_0[1:1]);
  NOR3 I189 (simp811_0[0:0], gtint_0[31:31], gtint_1[31:31], gtint_2[31:31]);
  INV I190 (simp811_0[1:1], gtint_3[31:31]);
  NAND2 I191 (o_0r1[31:31], simp811_0[0:0], simp811_0[1:1]);
  AND2 I192 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I193 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I194 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I195 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I196 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I197 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I198 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I199 (gtint_0[7:7], choice_0, i_0r1[7:7]);
  AND2 I200 (gtint_0[8:8], choice_0, i_0r1[8:8]);
  AND2 I201 (gtint_0[9:9], choice_0, i_0r1[9:9]);
  AND2 I202 (gtint_0[10:10], choice_0, i_0r1[10:10]);
  AND2 I203 (gtint_0[11:11], choice_0, i_0r1[11:11]);
  AND2 I204 (gtint_0[12:12], choice_0, i_0r1[12:12]);
  AND2 I205 (gtint_0[13:13], choice_0, i_0r1[13:13]);
  AND2 I206 (gtint_0[14:14], choice_0, i_0r1[14:14]);
  AND2 I207 (gtint_0[15:15], choice_0, i_0r1[15:15]);
  AND2 I208 (gtint_0[16:16], choice_0, i_0r1[16:16]);
  AND2 I209 (gtint_0[17:17], choice_0, i_0r1[17:17]);
  AND2 I210 (gtint_0[18:18], choice_0, i_0r1[18:18]);
  AND2 I211 (gtint_0[19:19], choice_0, i_0r1[19:19]);
  AND2 I212 (gtint_0[20:20], choice_0, i_0r1[20:20]);
  AND2 I213 (gtint_0[21:21], choice_0, i_0r1[21:21]);
  AND2 I214 (gtint_0[22:22], choice_0, i_0r1[22:22]);
  AND2 I215 (gtint_0[23:23], choice_0, i_0r1[23:23]);
  AND2 I216 (gtint_0[24:24], choice_0, i_0r1[24:24]);
  AND2 I217 (gtint_0[25:25], choice_0, i_0r1[25:25]);
  AND2 I218 (gtint_0[26:26], choice_0, i_0r1[26:26]);
  AND2 I219 (gtint_0[27:27], choice_0, i_0r1[27:27]);
  AND2 I220 (gtint_0[28:28], choice_0, i_0r1[28:28]);
  AND2 I221 (gtint_0[29:29], choice_0, i_0r1[29:29]);
  AND2 I222 (gtint_0[30:30], choice_0, i_0r1[30:30]);
  AND2 I223 (gtint_0[31:31], choice_0, i_0r1[31:31]);
  AND2 I224 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I225 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I226 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I227 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I228 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I229 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I230 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I231 (gtint_1[7:7], choice_1, i_1r1[7:7]);
  AND2 I232 (gtint_1[8:8], choice_1, i_1r1[8:8]);
  AND2 I233 (gtint_1[9:9], choice_1, i_1r1[9:9]);
  AND2 I234 (gtint_1[10:10], choice_1, i_1r1[10:10]);
  AND2 I235 (gtint_1[11:11], choice_1, i_1r1[11:11]);
  AND2 I236 (gtint_1[12:12], choice_1, i_1r1[12:12]);
  AND2 I237 (gtint_1[13:13], choice_1, i_1r1[13:13]);
  AND2 I238 (gtint_1[14:14], choice_1, i_1r1[14:14]);
  AND2 I239 (gtint_1[15:15], choice_1, i_1r1[15:15]);
  AND2 I240 (gtint_1[16:16], choice_1, i_1r1[16:16]);
  AND2 I241 (gtint_1[17:17], choice_1, i_1r1[17:17]);
  AND2 I242 (gtint_1[18:18], choice_1, i_1r1[18:18]);
  AND2 I243 (gtint_1[19:19], choice_1, i_1r1[19:19]);
  AND2 I244 (gtint_1[20:20], choice_1, i_1r1[20:20]);
  AND2 I245 (gtint_1[21:21], choice_1, i_1r1[21:21]);
  AND2 I246 (gtint_1[22:22], choice_1, i_1r1[22:22]);
  AND2 I247 (gtint_1[23:23], choice_1, i_1r1[23:23]);
  AND2 I248 (gtint_1[24:24], choice_1, i_1r1[24:24]);
  AND2 I249 (gtint_1[25:25], choice_1, i_1r1[25:25]);
  AND2 I250 (gtint_1[26:26], choice_1, i_1r1[26:26]);
  AND2 I251 (gtint_1[27:27], choice_1, i_1r1[27:27]);
  AND2 I252 (gtint_1[28:28], choice_1, i_1r1[28:28]);
  AND2 I253 (gtint_1[29:29], choice_1, i_1r1[29:29]);
  AND2 I254 (gtint_1[30:30], choice_1, i_1r1[30:30]);
  AND2 I255 (gtint_1[31:31], choice_1, i_1r1[31:31]);
  AND2 I256 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I257 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I258 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I259 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AND2 I260 (gtint_2[4:4], choice_2, i_2r1[4:4]);
  AND2 I261 (gtint_2[5:5], choice_2, i_2r1[5:5]);
  AND2 I262 (gtint_2[6:6], choice_2, i_2r1[6:6]);
  AND2 I263 (gtint_2[7:7], choice_2, i_2r1[7:7]);
  AND2 I264 (gtint_2[8:8], choice_2, i_2r1[8:8]);
  AND2 I265 (gtint_2[9:9], choice_2, i_2r1[9:9]);
  AND2 I266 (gtint_2[10:10], choice_2, i_2r1[10:10]);
  AND2 I267 (gtint_2[11:11], choice_2, i_2r1[11:11]);
  AND2 I268 (gtint_2[12:12], choice_2, i_2r1[12:12]);
  AND2 I269 (gtint_2[13:13], choice_2, i_2r1[13:13]);
  AND2 I270 (gtint_2[14:14], choice_2, i_2r1[14:14]);
  AND2 I271 (gtint_2[15:15], choice_2, i_2r1[15:15]);
  AND2 I272 (gtint_2[16:16], choice_2, i_2r1[16:16]);
  AND2 I273 (gtint_2[17:17], choice_2, i_2r1[17:17]);
  AND2 I274 (gtint_2[18:18], choice_2, i_2r1[18:18]);
  AND2 I275 (gtint_2[19:19], choice_2, i_2r1[19:19]);
  AND2 I276 (gtint_2[20:20], choice_2, i_2r1[20:20]);
  AND2 I277 (gtint_2[21:21], choice_2, i_2r1[21:21]);
  AND2 I278 (gtint_2[22:22], choice_2, i_2r1[22:22]);
  AND2 I279 (gtint_2[23:23], choice_2, i_2r1[23:23]);
  AND2 I280 (gtint_2[24:24], choice_2, i_2r1[24:24]);
  AND2 I281 (gtint_2[25:25], choice_2, i_2r1[25:25]);
  AND2 I282 (gtint_2[26:26], choice_2, i_2r1[26:26]);
  AND2 I283 (gtint_2[27:27], choice_2, i_2r1[27:27]);
  AND2 I284 (gtint_2[28:28], choice_2, i_2r1[28:28]);
  AND2 I285 (gtint_2[29:29], choice_2, i_2r1[29:29]);
  AND2 I286 (gtint_2[30:30], choice_2, i_2r1[30:30]);
  AND2 I287 (gtint_2[31:31], choice_2, i_2r1[31:31]);
  AND2 I288 (gtint_3[0:0], choice_3, i_3r1[0:0]);
  AND2 I289 (gtint_3[1:1], choice_3, i_3r1[1:1]);
  AND2 I290 (gtint_3[2:2], choice_3, i_3r1[2:2]);
  AND2 I291 (gtint_3[3:3], choice_3, i_3r1[3:3]);
  AND2 I292 (gtint_3[4:4], choice_3, i_3r1[4:4]);
  AND2 I293 (gtint_3[5:5], choice_3, i_3r1[5:5]);
  AND2 I294 (gtint_3[6:6], choice_3, i_3r1[6:6]);
  AND2 I295 (gtint_3[7:7], choice_3, i_3r1[7:7]);
  AND2 I296 (gtint_3[8:8], choice_3, i_3r1[8:8]);
  AND2 I297 (gtint_3[9:9], choice_3, i_3r1[9:9]);
  AND2 I298 (gtint_3[10:10], choice_3, i_3r1[10:10]);
  AND2 I299 (gtint_3[11:11], choice_3, i_3r1[11:11]);
  AND2 I300 (gtint_3[12:12], choice_3, i_3r1[12:12]);
  AND2 I301 (gtint_3[13:13], choice_3, i_3r1[13:13]);
  AND2 I302 (gtint_3[14:14], choice_3, i_3r1[14:14]);
  AND2 I303 (gtint_3[15:15], choice_3, i_3r1[15:15]);
  AND2 I304 (gtint_3[16:16], choice_3, i_3r1[16:16]);
  AND2 I305 (gtint_3[17:17], choice_3, i_3r1[17:17]);
  AND2 I306 (gtint_3[18:18], choice_3, i_3r1[18:18]);
  AND2 I307 (gtint_3[19:19], choice_3, i_3r1[19:19]);
  AND2 I308 (gtint_3[20:20], choice_3, i_3r1[20:20]);
  AND2 I309 (gtint_3[21:21], choice_3, i_3r1[21:21]);
  AND2 I310 (gtint_3[22:22], choice_3, i_3r1[22:22]);
  AND2 I311 (gtint_3[23:23], choice_3, i_3r1[23:23]);
  AND2 I312 (gtint_3[24:24], choice_3, i_3r1[24:24]);
  AND2 I313 (gtint_3[25:25], choice_3, i_3r1[25:25]);
  AND2 I314 (gtint_3[26:26], choice_3, i_3r1[26:26]);
  AND2 I315 (gtint_3[27:27], choice_3, i_3r1[27:27]);
  AND2 I316 (gtint_3[28:28], choice_3, i_3r1[28:28]);
  AND2 I317 (gtint_3[29:29], choice_3, i_3r1[29:29]);
  AND2 I318 (gtint_3[30:30], choice_3, i_3r1[30:30]);
  AND2 I319 (gtint_3[31:31], choice_3, i_3r1[31:31]);
  AND2 I320 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I321 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I322 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I323 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I324 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I325 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I326 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I327 (gfint_0[7:7], choice_0, i_0r0[7:7]);
  AND2 I328 (gfint_0[8:8], choice_0, i_0r0[8:8]);
  AND2 I329 (gfint_0[9:9], choice_0, i_0r0[9:9]);
  AND2 I330 (gfint_0[10:10], choice_0, i_0r0[10:10]);
  AND2 I331 (gfint_0[11:11], choice_0, i_0r0[11:11]);
  AND2 I332 (gfint_0[12:12], choice_0, i_0r0[12:12]);
  AND2 I333 (gfint_0[13:13], choice_0, i_0r0[13:13]);
  AND2 I334 (gfint_0[14:14], choice_0, i_0r0[14:14]);
  AND2 I335 (gfint_0[15:15], choice_0, i_0r0[15:15]);
  AND2 I336 (gfint_0[16:16], choice_0, i_0r0[16:16]);
  AND2 I337 (gfint_0[17:17], choice_0, i_0r0[17:17]);
  AND2 I338 (gfint_0[18:18], choice_0, i_0r0[18:18]);
  AND2 I339 (gfint_0[19:19], choice_0, i_0r0[19:19]);
  AND2 I340 (gfint_0[20:20], choice_0, i_0r0[20:20]);
  AND2 I341 (gfint_0[21:21], choice_0, i_0r0[21:21]);
  AND2 I342 (gfint_0[22:22], choice_0, i_0r0[22:22]);
  AND2 I343 (gfint_0[23:23], choice_0, i_0r0[23:23]);
  AND2 I344 (gfint_0[24:24], choice_0, i_0r0[24:24]);
  AND2 I345 (gfint_0[25:25], choice_0, i_0r0[25:25]);
  AND2 I346 (gfint_0[26:26], choice_0, i_0r0[26:26]);
  AND2 I347 (gfint_0[27:27], choice_0, i_0r0[27:27]);
  AND2 I348 (gfint_0[28:28], choice_0, i_0r0[28:28]);
  AND2 I349 (gfint_0[29:29], choice_0, i_0r0[29:29]);
  AND2 I350 (gfint_0[30:30], choice_0, i_0r0[30:30]);
  AND2 I351 (gfint_0[31:31], choice_0, i_0r0[31:31]);
  AND2 I352 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I353 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I354 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I355 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I356 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I357 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I358 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I359 (gfint_1[7:7], choice_1, i_1r0[7:7]);
  AND2 I360 (gfint_1[8:8], choice_1, i_1r0[8:8]);
  AND2 I361 (gfint_1[9:9], choice_1, i_1r0[9:9]);
  AND2 I362 (gfint_1[10:10], choice_1, i_1r0[10:10]);
  AND2 I363 (gfint_1[11:11], choice_1, i_1r0[11:11]);
  AND2 I364 (gfint_1[12:12], choice_1, i_1r0[12:12]);
  AND2 I365 (gfint_1[13:13], choice_1, i_1r0[13:13]);
  AND2 I366 (gfint_1[14:14], choice_1, i_1r0[14:14]);
  AND2 I367 (gfint_1[15:15], choice_1, i_1r0[15:15]);
  AND2 I368 (gfint_1[16:16], choice_1, i_1r0[16:16]);
  AND2 I369 (gfint_1[17:17], choice_1, i_1r0[17:17]);
  AND2 I370 (gfint_1[18:18], choice_1, i_1r0[18:18]);
  AND2 I371 (gfint_1[19:19], choice_1, i_1r0[19:19]);
  AND2 I372 (gfint_1[20:20], choice_1, i_1r0[20:20]);
  AND2 I373 (gfint_1[21:21], choice_1, i_1r0[21:21]);
  AND2 I374 (gfint_1[22:22], choice_1, i_1r0[22:22]);
  AND2 I375 (gfint_1[23:23], choice_1, i_1r0[23:23]);
  AND2 I376 (gfint_1[24:24], choice_1, i_1r0[24:24]);
  AND2 I377 (gfint_1[25:25], choice_1, i_1r0[25:25]);
  AND2 I378 (gfint_1[26:26], choice_1, i_1r0[26:26]);
  AND2 I379 (gfint_1[27:27], choice_1, i_1r0[27:27]);
  AND2 I380 (gfint_1[28:28], choice_1, i_1r0[28:28]);
  AND2 I381 (gfint_1[29:29], choice_1, i_1r0[29:29]);
  AND2 I382 (gfint_1[30:30], choice_1, i_1r0[30:30]);
  AND2 I383 (gfint_1[31:31], choice_1, i_1r0[31:31]);
  AND2 I384 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I385 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I386 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I387 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AND2 I388 (gfint_2[4:4], choice_2, i_2r0[4:4]);
  AND2 I389 (gfint_2[5:5], choice_2, i_2r0[5:5]);
  AND2 I390 (gfint_2[6:6], choice_2, i_2r0[6:6]);
  AND2 I391 (gfint_2[7:7], choice_2, i_2r0[7:7]);
  AND2 I392 (gfint_2[8:8], choice_2, i_2r0[8:8]);
  AND2 I393 (gfint_2[9:9], choice_2, i_2r0[9:9]);
  AND2 I394 (gfint_2[10:10], choice_2, i_2r0[10:10]);
  AND2 I395 (gfint_2[11:11], choice_2, i_2r0[11:11]);
  AND2 I396 (gfint_2[12:12], choice_2, i_2r0[12:12]);
  AND2 I397 (gfint_2[13:13], choice_2, i_2r0[13:13]);
  AND2 I398 (gfint_2[14:14], choice_2, i_2r0[14:14]);
  AND2 I399 (gfint_2[15:15], choice_2, i_2r0[15:15]);
  AND2 I400 (gfint_2[16:16], choice_2, i_2r0[16:16]);
  AND2 I401 (gfint_2[17:17], choice_2, i_2r0[17:17]);
  AND2 I402 (gfint_2[18:18], choice_2, i_2r0[18:18]);
  AND2 I403 (gfint_2[19:19], choice_2, i_2r0[19:19]);
  AND2 I404 (gfint_2[20:20], choice_2, i_2r0[20:20]);
  AND2 I405 (gfint_2[21:21], choice_2, i_2r0[21:21]);
  AND2 I406 (gfint_2[22:22], choice_2, i_2r0[22:22]);
  AND2 I407 (gfint_2[23:23], choice_2, i_2r0[23:23]);
  AND2 I408 (gfint_2[24:24], choice_2, i_2r0[24:24]);
  AND2 I409 (gfint_2[25:25], choice_2, i_2r0[25:25]);
  AND2 I410 (gfint_2[26:26], choice_2, i_2r0[26:26]);
  AND2 I411 (gfint_2[27:27], choice_2, i_2r0[27:27]);
  AND2 I412 (gfint_2[28:28], choice_2, i_2r0[28:28]);
  AND2 I413 (gfint_2[29:29], choice_2, i_2r0[29:29]);
  AND2 I414 (gfint_2[30:30], choice_2, i_2r0[30:30]);
  AND2 I415 (gfint_2[31:31], choice_2, i_2r0[31:31]);
  AND2 I416 (gfint_3[0:0], choice_3, i_3r0[0:0]);
  AND2 I417 (gfint_3[1:1], choice_3, i_3r0[1:1]);
  AND2 I418 (gfint_3[2:2], choice_3, i_3r0[2:2]);
  AND2 I419 (gfint_3[3:3], choice_3, i_3r0[3:3]);
  AND2 I420 (gfint_3[4:4], choice_3, i_3r0[4:4]);
  AND2 I421 (gfint_3[5:5], choice_3, i_3r0[5:5]);
  AND2 I422 (gfint_3[6:6], choice_3, i_3r0[6:6]);
  AND2 I423 (gfint_3[7:7], choice_3, i_3r0[7:7]);
  AND2 I424 (gfint_3[8:8], choice_3, i_3r0[8:8]);
  AND2 I425 (gfint_3[9:9], choice_3, i_3r0[9:9]);
  AND2 I426 (gfint_3[10:10], choice_3, i_3r0[10:10]);
  AND2 I427 (gfint_3[11:11], choice_3, i_3r0[11:11]);
  AND2 I428 (gfint_3[12:12], choice_3, i_3r0[12:12]);
  AND2 I429 (gfint_3[13:13], choice_3, i_3r0[13:13]);
  AND2 I430 (gfint_3[14:14], choice_3, i_3r0[14:14]);
  AND2 I431 (gfint_3[15:15], choice_3, i_3r0[15:15]);
  AND2 I432 (gfint_3[16:16], choice_3, i_3r0[16:16]);
  AND2 I433 (gfint_3[17:17], choice_3, i_3r0[17:17]);
  AND2 I434 (gfint_3[18:18], choice_3, i_3r0[18:18]);
  AND2 I435 (gfint_3[19:19], choice_3, i_3r0[19:19]);
  AND2 I436 (gfint_3[20:20], choice_3, i_3r0[20:20]);
  AND2 I437 (gfint_3[21:21], choice_3, i_3r0[21:21]);
  AND2 I438 (gfint_3[22:22], choice_3, i_3r0[22:22]);
  AND2 I439 (gfint_3[23:23], choice_3, i_3r0[23:23]);
  AND2 I440 (gfint_3[24:24], choice_3, i_3r0[24:24]);
  AND2 I441 (gfint_3[25:25], choice_3, i_3r0[25:25]);
  AND2 I442 (gfint_3[26:26], choice_3, i_3r0[26:26]);
  AND2 I443 (gfint_3[27:27], choice_3, i_3r0[27:27]);
  AND2 I444 (gfint_3[28:28], choice_3, i_3r0[28:28]);
  AND2 I445 (gfint_3[29:29], choice_3, i_3r0[29:29]);
  AND2 I446 (gfint_3[30:30], choice_3, i_3r0[30:30]);
  AND2 I447 (gfint_3[31:31], choice_3, i_3r0[31:31]);
  OR2 I448 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I449 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I450 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I451 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I452 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I453 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I454 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I455 (comp0_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I456 (comp0_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I457 (comp0_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I458 (comp0_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I459 (comp0_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I460 (comp0_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I461 (comp0_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I462 (comp0_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I463 (comp0_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I464 (comp0_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I465 (comp0_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I466 (comp0_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I467 (comp0_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I468 (comp0_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I469 (comp0_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I470 (comp0_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I471 (comp0_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I472 (comp0_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I473 (comp0_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I474 (comp0_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I475 (comp0_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I476 (comp0_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I477 (comp0_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I478 (comp0_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I479 (comp0_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  C3 I480 (simp3711_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I481 (simp3711_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I482 (simp3711_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I483 (simp3711_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I484 (simp3711_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I485 (simp3711_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I486 (simp3711_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I487 (simp3711_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I488 (simp3711_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I489 (simp3711_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I490 (simp3711_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I491 (simp3712_0[0:0], simp3711_0[0:0], simp3711_0[1:1], simp3711_0[2:2]);
  C3 I492 (simp3712_0[1:1], simp3711_0[3:3], simp3711_0[4:4], simp3711_0[5:5]);
  C3 I493 (simp3712_0[2:2], simp3711_0[6:6], simp3711_0[7:7], simp3711_0[8:8]);
  C2 I494 (simp3712_0[3:3], simp3711_0[9:9], simp3711_0[10:10]);
  C3 I495 (simp3713_0[0:0], simp3712_0[0:0], simp3712_0[1:1], simp3712_0[2:2]);
  BUFF I496 (simp3713_0[1:1], simp3712_0[3:3]);
  C2 I497 (icomp_0, simp3713_0[0:0], simp3713_0[1:1]);
  OR2 I498 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I499 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I500 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I501 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I502 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I503 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I504 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  OR2 I505 (comp1_0[7:7], i_1r0[7:7], i_1r1[7:7]);
  OR2 I506 (comp1_0[8:8], i_1r0[8:8], i_1r1[8:8]);
  OR2 I507 (comp1_0[9:9], i_1r0[9:9], i_1r1[9:9]);
  OR2 I508 (comp1_0[10:10], i_1r0[10:10], i_1r1[10:10]);
  OR2 I509 (comp1_0[11:11], i_1r0[11:11], i_1r1[11:11]);
  OR2 I510 (comp1_0[12:12], i_1r0[12:12], i_1r1[12:12]);
  OR2 I511 (comp1_0[13:13], i_1r0[13:13], i_1r1[13:13]);
  OR2 I512 (comp1_0[14:14], i_1r0[14:14], i_1r1[14:14]);
  OR2 I513 (comp1_0[15:15], i_1r0[15:15], i_1r1[15:15]);
  OR2 I514 (comp1_0[16:16], i_1r0[16:16], i_1r1[16:16]);
  OR2 I515 (comp1_0[17:17], i_1r0[17:17], i_1r1[17:17]);
  OR2 I516 (comp1_0[18:18], i_1r0[18:18], i_1r1[18:18]);
  OR2 I517 (comp1_0[19:19], i_1r0[19:19], i_1r1[19:19]);
  OR2 I518 (comp1_0[20:20], i_1r0[20:20], i_1r1[20:20]);
  OR2 I519 (comp1_0[21:21], i_1r0[21:21], i_1r1[21:21]);
  OR2 I520 (comp1_0[22:22], i_1r0[22:22], i_1r1[22:22]);
  OR2 I521 (comp1_0[23:23], i_1r0[23:23], i_1r1[23:23]);
  OR2 I522 (comp1_0[24:24], i_1r0[24:24], i_1r1[24:24]);
  OR2 I523 (comp1_0[25:25], i_1r0[25:25], i_1r1[25:25]);
  OR2 I524 (comp1_0[26:26], i_1r0[26:26], i_1r1[26:26]);
  OR2 I525 (comp1_0[27:27], i_1r0[27:27], i_1r1[27:27]);
  OR2 I526 (comp1_0[28:28], i_1r0[28:28], i_1r1[28:28]);
  OR2 I527 (comp1_0[29:29], i_1r0[29:29], i_1r1[29:29]);
  OR2 I528 (comp1_0[30:30], i_1r0[30:30], i_1r1[30:30]);
  OR2 I529 (comp1_0[31:31], i_1r0[31:31], i_1r1[31:31]);
  C3 I530 (simp4051_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I531 (simp4051_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  C3 I532 (simp4051_0[2:2], comp1_0[6:6], comp1_0[7:7], comp1_0[8:8]);
  C3 I533 (simp4051_0[3:3], comp1_0[9:9], comp1_0[10:10], comp1_0[11:11]);
  C3 I534 (simp4051_0[4:4], comp1_0[12:12], comp1_0[13:13], comp1_0[14:14]);
  C3 I535 (simp4051_0[5:5], comp1_0[15:15], comp1_0[16:16], comp1_0[17:17]);
  C3 I536 (simp4051_0[6:6], comp1_0[18:18], comp1_0[19:19], comp1_0[20:20]);
  C3 I537 (simp4051_0[7:7], comp1_0[21:21], comp1_0[22:22], comp1_0[23:23]);
  C3 I538 (simp4051_0[8:8], comp1_0[24:24], comp1_0[25:25], comp1_0[26:26]);
  C3 I539 (simp4051_0[9:9], comp1_0[27:27], comp1_0[28:28], comp1_0[29:29]);
  C2 I540 (simp4051_0[10:10], comp1_0[30:30], comp1_0[31:31]);
  C3 I541 (simp4052_0[0:0], simp4051_0[0:0], simp4051_0[1:1], simp4051_0[2:2]);
  C3 I542 (simp4052_0[1:1], simp4051_0[3:3], simp4051_0[4:4], simp4051_0[5:5]);
  C3 I543 (simp4052_0[2:2], simp4051_0[6:6], simp4051_0[7:7], simp4051_0[8:8]);
  C2 I544 (simp4052_0[3:3], simp4051_0[9:9], simp4051_0[10:10]);
  C3 I545 (simp4053_0[0:0], simp4052_0[0:0], simp4052_0[1:1], simp4052_0[2:2]);
  BUFF I546 (simp4053_0[1:1], simp4052_0[3:3]);
  C2 I547 (icomp_1, simp4053_0[0:0], simp4053_0[1:1]);
  OR2 I548 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I549 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I550 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2 I551 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  OR2 I552 (comp2_0[4:4], i_2r0[4:4], i_2r1[4:4]);
  OR2 I553 (comp2_0[5:5], i_2r0[5:5], i_2r1[5:5]);
  OR2 I554 (comp2_0[6:6], i_2r0[6:6], i_2r1[6:6]);
  OR2 I555 (comp2_0[7:7], i_2r0[7:7], i_2r1[7:7]);
  OR2 I556 (comp2_0[8:8], i_2r0[8:8], i_2r1[8:8]);
  OR2 I557 (comp2_0[9:9], i_2r0[9:9], i_2r1[9:9]);
  OR2 I558 (comp2_0[10:10], i_2r0[10:10], i_2r1[10:10]);
  OR2 I559 (comp2_0[11:11], i_2r0[11:11], i_2r1[11:11]);
  OR2 I560 (comp2_0[12:12], i_2r0[12:12], i_2r1[12:12]);
  OR2 I561 (comp2_0[13:13], i_2r0[13:13], i_2r1[13:13]);
  OR2 I562 (comp2_0[14:14], i_2r0[14:14], i_2r1[14:14]);
  OR2 I563 (comp2_0[15:15], i_2r0[15:15], i_2r1[15:15]);
  OR2 I564 (comp2_0[16:16], i_2r0[16:16], i_2r1[16:16]);
  OR2 I565 (comp2_0[17:17], i_2r0[17:17], i_2r1[17:17]);
  OR2 I566 (comp2_0[18:18], i_2r0[18:18], i_2r1[18:18]);
  OR2 I567 (comp2_0[19:19], i_2r0[19:19], i_2r1[19:19]);
  OR2 I568 (comp2_0[20:20], i_2r0[20:20], i_2r1[20:20]);
  OR2 I569 (comp2_0[21:21], i_2r0[21:21], i_2r1[21:21]);
  OR2 I570 (comp2_0[22:22], i_2r0[22:22], i_2r1[22:22]);
  OR2 I571 (comp2_0[23:23], i_2r0[23:23], i_2r1[23:23]);
  OR2 I572 (comp2_0[24:24], i_2r0[24:24], i_2r1[24:24]);
  OR2 I573 (comp2_0[25:25], i_2r0[25:25], i_2r1[25:25]);
  OR2 I574 (comp2_0[26:26], i_2r0[26:26], i_2r1[26:26]);
  OR2 I575 (comp2_0[27:27], i_2r0[27:27], i_2r1[27:27]);
  OR2 I576 (comp2_0[28:28], i_2r0[28:28], i_2r1[28:28]);
  OR2 I577 (comp2_0[29:29], i_2r0[29:29], i_2r1[29:29]);
  OR2 I578 (comp2_0[30:30], i_2r0[30:30], i_2r1[30:30]);
  OR2 I579 (comp2_0[31:31], i_2r0[31:31], i_2r1[31:31]);
  C3 I580 (simp4391_0[0:0], comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C3 I581 (simp4391_0[1:1], comp2_0[3:3], comp2_0[4:4], comp2_0[5:5]);
  C3 I582 (simp4391_0[2:2], comp2_0[6:6], comp2_0[7:7], comp2_0[8:8]);
  C3 I583 (simp4391_0[3:3], comp2_0[9:9], comp2_0[10:10], comp2_0[11:11]);
  C3 I584 (simp4391_0[4:4], comp2_0[12:12], comp2_0[13:13], comp2_0[14:14]);
  C3 I585 (simp4391_0[5:5], comp2_0[15:15], comp2_0[16:16], comp2_0[17:17]);
  C3 I586 (simp4391_0[6:6], comp2_0[18:18], comp2_0[19:19], comp2_0[20:20]);
  C3 I587 (simp4391_0[7:7], comp2_0[21:21], comp2_0[22:22], comp2_0[23:23]);
  C3 I588 (simp4391_0[8:8], comp2_0[24:24], comp2_0[25:25], comp2_0[26:26]);
  C3 I589 (simp4391_0[9:9], comp2_0[27:27], comp2_0[28:28], comp2_0[29:29]);
  C2 I590 (simp4391_0[10:10], comp2_0[30:30], comp2_0[31:31]);
  C3 I591 (simp4392_0[0:0], simp4391_0[0:0], simp4391_0[1:1], simp4391_0[2:2]);
  C3 I592 (simp4392_0[1:1], simp4391_0[3:3], simp4391_0[4:4], simp4391_0[5:5]);
  C3 I593 (simp4392_0[2:2], simp4391_0[6:6], simp4391_0[7:7], simp4391_0[8:8]);
  C2 I594 (simp4392_0[3:3], simp4391_0[9:9], simp4391_0[10:10]);
  C3 I595 (simp4393_0[0:0], simp4392_0[0:0], simp4392_0[1:1], simp4392_0[2:2]);
  BUFF I596 (simp4393_0[1:1], simp4392_0[3:3]);
  C2 I597 (icomp_2, simp4393_0[0:0], simp4393_0[1:1]);
  OR2 I598 (comp3_0[0:0], i_3r0[0:0], i_3r1[0:0]);
  OR2 I599 (comp3_0[1:1], i_3r0[1:1], i_3r1[1:1]);
  OR2 I600 (comp3_0[2:2], i_3r0[2:2], i_3r1[2:2]);
  OR2 I601 (comp3_0[3:3], i_3r0[3:3], i_3r1[3:3]);
  OR2 I602 (comp3_0[4:4], i_3r0[4:4], i_3r1[4:4]);
  OR2 I603 (comp3_0[5:5], i_3r0[5:5], i_3r1[5:5]);
  OR2 I604 (comp3_0[6:6], i_3r0[6:6], i_3r1[6:6]);
  OR2 I605 (comp3_0[7:7], i_3r0[7:7], i_3r1[7:7]);
  OR2 I606 (comp3_0[8:8], i_3r0[8:8], i_3r1[8:8]);
  OR2 I607 (comp3_0[9:9], i_3r0[9:9], i_3r1[9:9]);
  OR2 I608 (comp3_0[10:10], i_3r0[10:10], i_3r1[10:10]);
  OR2 I609 (comp3_0[11:11], i_3r0[11:11], i_3r1[11:11]);
  OR2 I610 (comp3_0[12:12], i_3r0[12:12], i_3r1[12:12]);
  OR2 I611 (comp3_0[13:13], i_3r0[13:13], i_3r1[13:13]);
  OR2 I612 (comp3_0[14:14], i_3r0[14:14], i_3r1[14:14]);
  OR2 I613 (comp3_0[15:15], i_3r0[15:15], i_3r1[15:15]);
  OR2 I614 (comp3_0[16:16], i_3r0[16:16], i_3r1[16:16]);
  OR2 I615 (comp3_0[17:17], i_3r0[17:17], i_3r1[17:17]);
  OR2 I616 (comp3_0[18:18], i_3r0[18:18], i_3r1[18:18]);
  OR2 I617 (comp3_0[19:19], i_3r0[19:19], i_3r1[19:19]);
  OR2 I618 (comp3_0[20:20], i_3r0[20:20], i_3r1[20:20]);
  OR2 I619 (comp3_0[21:21], i_3r0[21:21], i_3r1[21:21]);
  OR2 I620 (comp3_0[22:22], i_3r0[22:22], i_3r1[22:22]);
  OR2 I621 (comp3_0[23:23], i_3r0[23:23], i_3r1[23:23]);
  OR2 I622 (comp3_0[24:24], i_3r0[24:24], i_3r1[24:24]);
  OR2 I623 (comp3_0[25:25], i_3r0[25:25], i_3r1[25:25]);
  OR2 I624 (comp3_0[26:26], i_3r0[26:26], i_3r1[26:26]);
  OR2 I625 (comp3_0[27:27], i_3r0[27:27], i_3r1[27:27]);
  OR2 I626 (comp3_0[28:28], i_3r0[28:28], i_3r1[28:28]);
  OR2 I627 (comp3_0[29:29], i_3r0[29:29], i_3r1[29:29]);
  OR2 I628 (comp3_0[30:30], i_3r0[30:30], i_3r1[30:30]);
  OR2 I629 (comp3_0[31:31], i_3r0[31:31], i_3r1[31:31]);
  C3 I630 (simp4731_0[0:0], comp3_0[0:0], comp3_0[1:1], comp3_0[2:2]);
  C3 I631 (simp4731_0[1:1], comp3_0[3:3], comp3_0[4:4], comp3_0[5:5]);
  C3 I632 (simp4731_0[2:2], comp3_0[6:6], comp3_0[7:7], comp3_0[8:8]);
  C3 I633 (simp4731_0[3:3], comp3_0[9:9], comp3_0[10:10], comp3_0[11:11]);
  C3 I634 (simp4731_0[4:4], comp3_0[12:12], comp3_0[13:13], comp3_0[14:14]);
  C3 I635 (simp4731_0[5:5], comp3_0[15:15], comp3_0[16:16], comp3_0[17:17]);
  C3 I636 (simp4731_0[6:6], comp3_0[18:18], comp3_0[19:19], comp3_0[20:20]);
  C3 I637 (simp4731_0[7:7], comp3_0[21:21], comp3_0[22:22], comp3_0[23:23]);
  C3 I638 (simp4731_0[8:8], comp3_0[24:24], comp3_0[25:25], comp3_0[26:26]);
  C3 I639 (simp4731_0[9:9], comp3_0[27:27], comp3_0[28:28], comp3_0[29:29]);
  C2 I640 (simp4731_0[10:10], comp3_0[30:30], comp3_0[31:31]);
  C3 I641 (simp4732_0[0:0], simp4731_0[0:0], simp4731_0[1:1], simp4731_0[2:2]);
  C3 I642 (simp4732_0[1:1], simp4731_0[3:3], simp4731_0[4:4], simp4731_0[5:5]);
  C3 I643 (simp4732_0[2:2], simp4731_0[6:6], simp4731_0[7:7], simp4731_0[8:8]);
  C2 I644 (simp4732_0[3:3], simp4731_0[9:9], simp4731_0[10:10]);
  C3 I645 (simp4733_0[0:0], simp4732_0[0:0], simp4732_0[1:1], simp4732_0[2:2]);
  BUFF I646 (simp4733_0[1:1], simp4732_0[3:3]);
  C2 I647 (icomp_3, simp4733_0[0:0], simp4733_0[1:1]);
  C2R I648 (choice_0, icomp_0, nchosen_0, reset);
  C2R I649 (choice_1, icomp_1, nchosen_0, reset);
  C2R I650 (choice_2, icomp_2, nchosen_0, reset);
  C2R I651 (choice_3, icomp_3, nchosen_0, reset);
  NOR3 I652 (simp4781_0[0:0], choice_0, choice_1, choice_2);
  INV I653 (simp4781_0[1:1], choice_3);
  NAND2 I654 (anychoice_0, simp4781_0[0:0], simp4781_0[1:1]);
  NOR2 I655 (nchosen_0, anychoice_0, o_0a);
  C2R I656 (i_0a, choice_0, o_0a, reset);
  C2R I657 (i_1a, choice_1, o_0a, reset);
  C2R I658 (i_2a, choice_2, o_0a, reset);
  C2R I659 (i_3a, choice_3, o_0a, reset);
endmodule

// tko0m4_1nm4b0 TeakO [
//     (1,TeakOConstant 4 0)] [One 0,One 4]
module tko0m4_1nm4b0 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r);
  BUFF I1 (o_0r0[1:1], i_0r);
  BUFF I2 (o_0r0[2:2], i_0r);
  BUFF I3 (o_0r0[3:3], i_0r);
  GND I4 (o_0r1[0:0]);
  GND I5 (o_0r1[1:1]);
  GND I6 (o_0r1[2:2]);
  GND I7 (o_0r1[3:3]);
  BUFF I8 (i_0a, o_0a);
endmodule

// tkj32m4_28 TeakJ [Many [4,28],One 32]
module tkj32m4_28 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  input [27:0] i_1r0;
  input [27:0] i_1r1;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [31:0] joinf_0;
  wire [31:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_1r0[0:0]);
  BUFF I5 (joinf_0[5:5], i_1r0[1:1]);
  BUFF I6 (joinf_0[6:6], i_1r0[2:2]);
  BUFF I7 (joinf_0[7:7], i_1r0[3:3]);
  BUFF I8 (joinf_0[8:8], i_1r0[4:4]);
  BUFF I9 (joinf_0[9:9], i_1r0[5:5]);
  BUFF I10 (joinf_0[10:10], i_1r0[6:6]);
  BUFF I11 (joinf_0[11:11], i_1r0[7:7]);
  BUFF I12 (joinf_0[12:12], i_1r0[8:8]);
  BUFF I13 (joinf_0[13:13], i_1r0[9:9]);
  BUFF I14 (joinf_0[14:14], i_1r0[10:10]);
  BUFF I15 (joinf_0[15:15], i_1r0[11:11]);
  BUFF I16 (joinf_0[16:16], i_1r0[12:12]);
  BUFF I17 (joinf_0[17:17], i_1r0[13:13]);
  BUFF I18 (joinf_0[18:18], i_1r0[14:14]);
  BUFF I19 (joinf_0[19:19], i_1r0[15:15]);
  BUFF I20 (joinf_0[20:20], i_1r0[16:16]);
  BUFF I21 (joinf_0[21:21], i_1r0[17:17]);
  BUFF I22 (joinf_0[22:22], i_1r0[18:18]);
  BUFF I23 (joinf_0[23:23], i_1r0[19:19]);
  BUFF I24 (joinf_0[24:24], i_1r0[20:20]);
  BUFF I25 (joinf_0[25:25], i_1r0[21:21]);
  BUFF I26 (joinf_0[26:26], i_1r0[22:22]);
  BUFF I27 (joinf_0[27:27], i_1r0[23:23]);
  BUFF I28 (joinf_0[28:28], i_1r0[24:24]);
  BUFF I29 (joinf_0[29:29], i_1r0[25:25]);
  BUFF I30 (joinf_0[30:30], i_1r0[26:26]);
  BUFF I31 (joinf_0[31:31], i_1r0[27:27]);
  BUFF I32 (joint_0[0:0], i_0r1[0:0]);
  BUFF I33 (joint_0[1:1], i_0r1[1:1]);
  BUFF I34 (joint_0[2:2], i_0r1[2:2]);
  BUFF I35 (joint_0[3:3], i_0r1[3:3]);
  BUFF I36 (joint_0[4:4], i_1r1[0:0]);
  BUFF I37 (joint_0[5:5], i_1r1[1:1]);
  BUFF I38 (joint_0[6:6], i_1r1[2:2]);
  BUFF I39 (joint_0[7:7], i_1r1[3:3]);
  BUFF I40 (joint_0[8:8], i_1r1[4:4]);
  BUFF I41 (joint_0[9:9], i_1r1[5:5]);
  BUFF I42 (joint_0[10:10], i_1r1[6:6]);
  BUFF I43 (joint_0[11:11], i_1r1[7:7]);
  BUFF I44 (joint_0[12:12], i_1r1[8:8]);
  BUFF I45 (joint_0[13:13], i_1r1[9:9]);
  BUFF I46 (joint_0[14:14], i_1r1[10:10]);
  BUFF I47 (joint_0[15:15], i_1r1[11:11]);
  BUFF I48 (joint_0[16:16], i_1r1[12:12]);
  BUFF I49 (joint_0[17:17], i_1r1[13:13]);
  BUFF I50 (joint_0[18:18], i_1r1[14:14]);
  BUFF I51 (joint_0[19:19], i_1r1[15:15]);
  BUFF I52 (joint_0[20:20], i_1r1[16:16]);
  BUFF I53 (joint_0[21:21], i_1r1[17:17]);
  BUFF I54 (joint_0[22:22], i_1r1[18:18]);
  BUFF I55 (joint_0[23:23], i_1r1[19:19]);
  BUFF I56 (joint_0[24:24], i_1r1[20:20]);
  BUFF I57 (joint_0[25:25], i_1r1[21:21]);
  BUFF I58 (joint_0[26:26], i_1r1[22:22]);
  BUFF I59 (joint_0[27:27], i_1r1[23:23]);
  BUFF I60 (joint_0[28:28], i_1r1[24:24]);
  BUFF I61 (joint_0[29:29], i_1r1[25:25]);
  BUFF I62 (joint_0[30:30], i_1r1[26:26]);
  BUFF I63 (joint_0[31:31], i_1r1[27:27]);
  OR2 I64 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I65 (icomplete_0, dcomplete_0);
  C2 I66 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I67 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I68 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I69 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I70 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I71 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I72 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I73 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I74 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I75 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I76 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I77 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I78 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I79 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I80 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I81 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I82 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I83 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I84 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I85 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I86 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I87 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I88 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I89 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I90 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I91 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I92 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I93 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I94 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I95 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I96 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I97 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I98 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I99 (o_0r1[1:1], joint_0[1:1]);
  BUFF I100 (o_0r1[2:2], joint_0[2:2]);
  BUFF I101 (o_0r1[3:3], joint_0[3:3]);
  BUFF I102 (o_0r1[4:4], joint_0[4:4]);
  BUFF I103 (o_0r1[5:5], joint_0[5:5]);
  BUFF I104 (o_0r1[6:6], joint_0[6:6]);
  BUFF I105 (o_0r1[7:7], joint_0[7:7]);
  BUFF I106 (o_0r1[8:8], joint_0[8:8]);
  BUFF I107 (o_0r1[9:9], joint_0[9:9]);
  BUFF I108 (o_0r1[10:10], joint_0[10:10]);
  BUFF I109 (o_0r1[11:11], joint_0[11:11]);
  BUFF I110 (o_0r1[12:12], joint_0[12:12]);
  BUFF I111 (o_0r1[13:13], joint_0[13:13]);
  BUFF I112 (o_0r1[14:14], joint_0[14:14]);
  BUFF I113 (o_0r1[15:15], joint_0[15:15]);
  BUFF I114 (o_0r1[16:16], joint_0[16:16]);
  BUFF I115 (o_0r1[17:17], joint_0[17:17]);
  BUFF I116 (o_0r1[18:18], joint_0[18:18]);
  BUFF I117 (o_0r1[19:19], joint_0[19:19]);
  BUFF I118 (o_0r1[20:20], joint_0[20:20]);
  BUFF I119 (o_0r1[21:21], joint_0[21:21]);
  BUFF I120 (o_0r1[22:22], joint_0[22:22]);
  BUFF I121 (o_0r1[23:23], joint_0[23:23]);
  BUFF I122 (o_0r1[24:24], joint_0[24:24]);
  BUFF I123 (o_0r1[25:25], joint_0[25:25]);
  BUFF I124 (o_0r1[26:26], joint_0[26:26]);
  BUFF I125 (o_0r1[27:27], joint_0[27:27]);
  BUFF I126 (o_0r1[28:28], joint_0[28:28]);
  BUFF I127 (o_0r1[29:29], joint_0[29:29]);
  BUFF I128 (o_0r1[30:30], joint_0[30:30]);
  BUFF I129 (o_0r1[31:31], joint_0[31:31]);
  BUFF I130 (i_0a, o_0a);
  BUFF I131 (i_1a, o_0a);
endmodule

// tkj32m28_4 TeakJ [Many [28,4],One 32]
module tkj32m28_4 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [27:0] i_0r0;
  input [27:0] i_0r1;
  output i_0a;
  input [3:0] i_1r0;
  input [3:0] i_1r1;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [31:0] joinf_0;
  wire [31:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_1r0[0:0]);
  BUFF I29 (joinf_0[29:29], i_1r0[1:1]);
  BUFF I30 (joinf_0[30:30], i_1r0[2:2]);
  BUFF I31 (joinf_0[31:31], i_1r0[3:3]);
  BUFF I32 (joint_0[0:0], i_0r1[0:0]);
  BUFF I33 (joint_0[1:1], i_0r1[1:1]);
  BUFF I34 (joint_0[2:2], i_0r1[2:2]);
  BUFF I35 (joint_0[3:3], i_0r1[3:3]);
  BUFF I36 (joint_0[4:4], i_0r1[4:4]);
  BUFF I37 (joint_0[5:5], i_0r1[5:5]);
  BUFF I38 (joint_0[6:6], i_0r1[6:6]);
  BUFF I39 (joint_0[7:7], i_0r1[7:7]);
  BUFF I40 (joint_0[8:8], i_0r1[8:8]);
  BUFF I41 (joint_0[9:9], i_0r1[9:9]);
  BUFF I42 (joint_0[10:10], i_0r1[10:10]);
  BUFF I43 (joint_0[11:11], i_0r1[11:11]);
  BUFF I44 (joint_0[12:12], i_0r1[12:12]);
  BUFF I45 (joint_0[13:13], i_0r1[13:13]);
  BUFF I46 (joint_0[14:14], i_0r1[14:14]);
  BUFF I47 (joint_0[15:15], i_0r1[15:15]);
  BUFF I48 (joint_0[16:16], i_0r1[16:16]);
  BUFF I49 (joint_0[17:17], i_0r1[17:17]);
  BUFF I50 (joint_0[18:18], i_0r1[18:18]);
  BUFF I51 (joint_0[19:19], i_0r1[19:19]);
  BUFF I52 (joint_0[20:20], i_0r1[20:20]);
  BUFF I53 (joint_0[21:21], i_0r1[21:21]);
  BUFF I54 (joint_0[22:22], i_0r1[22:22]);
  BUFF I55 (joint_0[23:23], i_0r1[23:23]);
  BUFF I56 (joint_0[24:24], i_0r1[24:24]);
  BUFF I57 (joint_0[25:25], i_0r1[25:25]);
  BUFF I58 (joint_0[26:26], i_0r1[26:26]);
  BUFF I59 (joint_0[27:27], i_0r1[27:27]);
  BUFF I60 (joint_0[28:28], i_1r1[0:0]);
  BUFF I61 (joint_0[29:29], i_1r1[1:1]);
  BUFF I62 (joint_0[30:30], i_1r1[2:2]);
  BUFF I63 (joint_0[31:31], i_1r1[3:3]);
  OR2 I64 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I65 (icomplete_0, dcomplete_0);
  C2 I66 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I67 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I68 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I69 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I70 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I71 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I72 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I73 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I74 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I75 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I76 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I77 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I78 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I79 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I80 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I81 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I82 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I83 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I84 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I85 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I86 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I87 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I88 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I89 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I90 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I91 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I92 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I93 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I94 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I95 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I96 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I97 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I98 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I99 (o_0r1[1:1], joint_0[1:1]);
  BUFF I100 (o_0r1[2:2], joint_0[2:2]);
  BUFF I101 (o_0r1[3:3], joint_0[3:3]);
  BUFF I102 (o_0r1[4:4], joint_0[4:4]);
  BUFF I103 (o_0r1[5:5], joint_0[5:5]);
  BUFF I104 (o_0r1[6:6], joint_0[6:6]);
  BUFF I105 (o_0r1[7:7], joint_0[7:7]);
  BUFF I106 (o_0r1[8:8], joint_0[8:8]);
  BUFF I107 (o_0r1[9:9], joint_0[9:9]);
  BUFF I108 (o_0r1[10:10], joint_0[10:10]);
  BUFF I109 (o_0r1[11:11], joint_0[11:11]);
  BUFF I110 (o_0r1[12:12], joint_0[12:12]);
  BUFF I111 (o_0r1[13:13], joint_0[13:13]);
  BUFF I112 (o_0r1[14:14], joint_0[14:14]);
  BUFF I113 (o_0r1[15:15], joint_0[15:15]);
  BUFF I114 (o_0r1[16:16], joint_0[16:16]);
  BUFF I115 (o_0r1[17:17], joint_0[17:17]);
  BUFF I116 (o_0r1[18:18], joint_0[18:18]);
  BUFF I117 (o_0r1[19:19], joint_0[19:19]);
  BUFF I118 (o_0r1[20:20], joint_0[20:20]);
  BUFF I119 (o_0r1[21:21], joint_0[21:21]);
  BUFF I120 (o_0r1[22:22], joint_0[22:22]);
  BUFF I121 (o_0r1[23:23], joint_0[23:23]);
  BUFF I122 (o_0r1[24:24], joint_0[24:24]);
  BUFF I123 (o_0r1[25:25], joint_0[25:25]);
  BUFF I124 (o_0r1[26:26], joint_0[26:26]);
  BUFF I125 (o_0r1[27:27], joint_0[27:27]);
  BUFF I126 (o_0r1[28:28], joint_0[28:28]);
  BUFF I127 (o_0r1[29:29], joint_0[29:29]);
  BUFF I128 (o_0r1[30:30], joint_0[30:30]);
  BUFF I129 (o_0r1[31:31], joint_0[31:31]);
  BUFF I130 (i_0a, o_0a);
  BUFF I131 (i_1a, o_0a);
endmodule

// tko0m4_1nm4bf TeakO [
//     (1,TeakOConstant 4 15)] [One 0,One 4]
module tko0m4_1nm4bf (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  BUFF I1 (o_0r1[1:1], i_0r);
  BUFF I2 (o_0r1[2:2], i_0r);
  BUFF I3 (o_0r1[3:3], i_0r);
  GND I4 (o_0r0[0:0]);
  GND I5 (o_0r0[1:1]);
  GND I6 (o_0r0[2:2]);
  GND I7 (o_0r0[3:3]);
  BUFF I8 (i_0a, o_0a);
endmodule

// tkvi32_wo0w32_ro0w32o0w28o4w28o4w28 TeakV "i" 32 [] [0] [0,0,4,4] [Many [32],Many [0],Many [0,0,0,0]
//   ,Many [32,28,28,28]]
module tkvi32_wo0w32_ro0w32o0w28o4w28o4w28 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [27:0] rd_1r0;
  output [27:0] rd_1r1;
  input rd_1a;
  output [27:0] rd_2r0;
  output [27:0] rd_2r1;
  input rd_2a;
  output [27:0] rd_3r0;
  output [27:0] rd_3r1;
  input rd_3a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [2:0] simp6401_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_2r0[0:0], df_0[4:4], rg_2r);
  AND2 I485 (rd_2r0[1:1], df_0[5:5], rg_2r);
  AND2 I486 (rd_2r0[2:2], df_0[6:6], rg_2r);
  AND2 I487 (rd_2r0[3:3], df_0[7:7], rg_2r);
  AND2 I488 (rd_2r0[4:4], df_0[8:8], rg_2r);
  AND2 I489 (rd_2r0[5:5], df_0[9:9], rg_2r);
  AND2 I490 (rd_2r0[6:6], df_0[10:10], rg_2r);
  AND2 I491 (rd_2r0[7:7], df_0[11:11], rg_2r);
  AND2 I492 (rd_2r0[8:8], df_0[12:12], rg_2r);
  AND2 I493 (rd_2r0[9:9], df_0[13:13], rg_2r);
  AND2 I494 (rd_2r0[10:10], df_0[14:14], rg_2r);
  AND2 I495 (rd_2r0[11:11], df_0[15:15], rg_2r);
  AND2 I496 (rd_2r0[12:12], df_0[16:16], rg_2r);
  AND2 I497 (rd_2r0[13:13], df_0[17:17], rg_2r);
  AND2 I498 (rd_2r0[14:14], df_0[18:18], rg_2r);
  AND2 I499 (rd_2r0[15:15], df_0[19:19], rg_2r);
  AND2 I500 (rd_2r0[16:16], df_0[20:20], rg_2r);
  AND2 I501 (rd_2r0[17:17], df_0[21:21], rg_2r);
  AND2 I502 (rd_2r0[18:18], df_0[22:22], rg_2r);
  AND2 I503 (rd_2r0[19:19], df_0[23:23], rg_2r);
  AND2 I504 (rd_2r0[20:20], df_0[24:24], rg_2r);
  AND2 I505 (rd_2r0[21:21], df_0[25:25], rg_2r);
  AND2 I506 (rd_2r0[22:22], df_0[26:26], rg_2r);
  AND2 I507 (rd_2r0[23:23], df_0[27:27], rg_2r);
  AND2 I508 (rd_2r0[24:24], df_0[28:28], rg_2r);
  AND2 I509 (rd_2r0[25:25], df_0[29:29], rg_2r);
  AND2 I510 (rd_2r0[26:26], df_0[30:30], rg_2r);
  AND2 I511 (rd_2r0[27:27], df_0[31:31], rg_2r);
  AND2 I512 (rd_3r0[0:0], df_0[4:4], rg_3r);
  AND2 I513 (rd_3r0[1:1], df_0[5:5], rg_3r);
  AND2 I514 (rd_3r0[2:2], df_0[6:6], rg_3r);
  AND2 I515 (rd_3r0[3:3], df_0[7:7], rg_3r);
  AND2 I516 (rd_3r0[4:4], df_0[8:8], rg_3r);
  AND2 I517 (rd_3r0[5:5], df_0[9:9], rg_3r);
  AND2 I518 (rd_3r0[6:6], df_0[10:10], rg_3r);
  AND2 I519 (rd_3r0[7:7], df_0[11:11], rg_3r);
  AND2 I520 (rd_3r0[8:8], df_0[12:12], rg_3r);
  AND2 I521 (rd_3r0[9:9], df_0[13:13], rg_3r);
  AND2 I522 (rd_3r0[10:10], df_0[14:14], rg_3r);
  AND2 I523 (rd_3r0[11:11], df_0[15:15], rg_3r);
  AND2 I524 (rd_3r0[12:12], df_0[16:16], rg_3r);
  AND2 I525 (rd_3r0[13:13], df_0[17:17], rg_3r);
  AND2 I526 (rd_3r0[14:14], df_0[18:18], rg_3r);
  AND2 I527 (rd_3r0[15:15], df_0[19:19], rg_3r);
  AND2 I528 (rd_3r0[16:16], df_0[20:20], rg_3r);
  AND2 I529 (rd_3r0[17:17], df_0[21:21], rg_3r);
  AND2 I530 (rd_3r0[18:18], df_0[22:22], rg_3r);
  AND2 I531 (rd_3r0[19:19], df_0[23:23], rg_3r);
  AND2 I532 (rd_3r0[20:20], df_0[24:24], rg_3r);
  AND2 I533 (rd_3r0[21:21], df_0[25:25], rg_3r);
  AND2 I534 (rd_3r0[22:22], df_0[26:26], rg_3r);
  AND2 I535 (rd_3r0[23:23], df_0[27:27], rg_3r);
  AND2 I536 (rd_3r0[24:24], df_0[28:28], rg_3r);
  AND2 I537 (rd_3r0[25:25], df_0[29:29], rg_3r);
  AND2 I538 (rd_3r0[26:26], df_0[30:30], rg_3r);
  AND2 I539 (rd_3r0[27:27], df_0[31:31], rg_3r);
  AND2 I540 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I541 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I542 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I543 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I544 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I545 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I546 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I547 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I548 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I549 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I550 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I551 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I552 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I553 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I554 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I555 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I556 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I557 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I558 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I559 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I560 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I561 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I562 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I563 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I564 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I565 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I566 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I567 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I568 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I569 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I570 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I571 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I572 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I573 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I574 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I575 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I576 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I577 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I578 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I579 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I580 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I581 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I582 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I583 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I584 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I585 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I586 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I587 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I588 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I589 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I590 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I591 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I592 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I593 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I594 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I595 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I596 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I597 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I598 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I599 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I600 (rd_2r1[0:0], dt_0[4:4], rg_2r);
  AND2 I601 (rd_2r1[1:1], dt_0[5:5], rg_2r);
  AND2 I602 (rd_2r1[2:2], dt_0[6:6], rg_2r);
  AND2 I603 (rd_2r1[3:3], dt_0[7:7], rg_2r);
  AND2 I604 (rd_2r1[4:4], dt_0[8:8], rg_2r);
  AND2 I605 (rd_2r1[5:5], dt_0[9:9], rg_2r);
  AND2 I606 (rd_2r1[6:6], dt_0[10:10], rg_2r);
  AND2 I607 (rd_2r1[7:7], dt_0[11:11], rg_2r);
  AND2 I608 (rd_2r1[8:8], dt_0[12:12], rg_2r);
  AND2 I609 (rd_2r1[9:9], dt_0[13:13], rg_2r);
  AND2 I610 (rd_2r1[10:10], dt_0[14:14], rg_2r);
  AND2 I611 (rd_2r1[11:11], dt_0[15:15], rg_2r);
  AND2 I612 (rd_2r1[12:12], dt_0[16:16], rg_2r);
  AND2 I613 (rd_2r1[13:13], dt_0[17:17], rg_2r);
  AND2 I614 (rd_2r1[14:14], dt_0[18:18], rg_2r);
  AND2 I615 (rd_2r1[15:15], dt_0[19:19], rg_2r);
  AND2 I616 (rd_2r1[16:16], dt_0[20:20], rg_2r);
  AND2 I617 (rd_2r1[17:17], dt_0[21:21], rg_2r);
  AND2 I618 (rd_2r1[18:18], dt_0[22:22], rg_2r);
  AND2 I619 (rd_2r1[19:19], dt_0[23:23], rg_2r);
  AND2 I620 (rd_2r1[20:20], dt_0[24:24], rg_2r);
  AND2 I621 (rd_2r1[21:21], dt_0[25:25], rg_2r);
  AND2 I622 (rd_2r1[22:22], dt_0[26:26], rg_2r);
  AND2 I623 (rd_2r1[23:23], dt_0[27:27], rg_2r);
  AND2 I624 (rd_2r1[24:24], dt_0[28:28], rg_2r);
  AND2 I625 (rd_2r1[25:25], dt_0[29:29], rg_2r);
  AND2 I626 (rd_2r1[26:26], dt_0[30:30], rg_2r);
  AND2 I627 (rd_2r1[27:27], dt_0[31:31], rg_2r);
  AND2 I628 (rd_3r1[0:0], dt_0[4:4], rg_3r);
  AND2 I629 (rd_3r1[1:1], dt_0[5:5], rg_3r);
  AND2 I630 (rd_3r1[2:2], dt_0[6:6], rg_3r);
  AND2 I631 (rd_3r1[3:3], dt_0[7:7], rg_3r);
  AND2 I632 (rd_3r1[4:4], dt_0[8:8], rg_3r);
  AND2 I633 (rd_3r1[5:5], dt_0[9:9], rg_3r);
  AND2 I634 (rd_3r1[6:6], dt_0[10:10], rg_3r);
  AND2 I635 (rd_3r1[7:7], dt_0[11:11], rg_3r);
  AND2 I636 (rd_3r1[8:8], dt_0[12:12], rg_3r);
  AND2 I637 (rd_3r1[9:9], dt_0[13:13], rg_3r);
  AND2 I638 (rd_3r1[10:10], dt_0[14:14], rg_3r);
  AND2 I639 (rd_3r1[11:11], dt_0[15:15], rg_3r);
  AND2 I640 (rd_3r1[12:12], dt_0[16:16], rg_3r);
  AND2 I641 (rd_3r1[13:13], dt_0[17:17], rg_3r);
  AND2 I642 (rd_3r1[14:14], dt_0[18:18], rg_3r);
  AND2 I643 (rd_3r1[15:15], dt_0[19:19], rg_3r);
  AND2 I644 (rd_3r1[16:16], dt_0[20:20], rg_3r);
  AND2 I645 (rd_3r1[17:17], dt_0[21:21], rg_3r);
  AND2 I646 (rd_3r1[18:18], dt_0[22:22], rg_3r);
  AND2 I647 (rd_3r1[19:19], dt_0[23:23], rg_3r);
  AND2 I648 (rd_3r1[20:20], dt_0[24:24], rg_3r);
  AND2 I649 (rd_3r1[21:21], dt_0[25:25], rg_3r);
  AND2 I650 (rd_3r1[22:22], dt_0[26:26], rg_3r);
  AND2 I651 (rd_3r1[23:23], dt_0[27:27], rg_3r);
  AND2 I652 (rd_3r1[24:24], dt_0[28:28], rg_3r);
  AND2 I653 (rd_3r1[25:25], dt_0[29:29], rg_3r);
  AND2 I654 (rd_3r1[26:26], dt_0[30:30], rg_3r);
  AND2 I655 (rd_3r1[27:27], dt_0[31:31], rg_3r);
  NOR3 I656 (simp6401_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I657 (simp6401_0[1:1], rg_3r, rg_0a, rg_1a);
  NOR2 I658 (simp6401_0[2:2], rg_2a, rg_3a);
  NAND3 I659 (anyread_0, simp6401_0[0:0], simp6401_0[1:1], simp6401_0[2:2]);
  BUFF I660 (wg_0a, wd_0a);
  BUFF I661 (rg_0a, rd_0a);
  BUFF I662 (rg_1a, rd_1a);
  BUFF I663 (rg_2a, rd_2a);
  BUFF I664 (rg_3a, rd_3a);
endmodule

// tko0m8_1nm8b0 TeakO [
//     (1,TeakOConstant 8 0)] [One 0,One 8]
module tko0m8_1nm8b0 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [7:0] o_0r0;
  output [7:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r);
  BUFF I1 (o_0r0[1:1], i_0r);
  BUFF I2 (o_0r0[2:2], i_0r);
  BUFF I3 (o_0r0[3:3], i_0r);
  BUFF I4 (o_0r0[4:4], i_0r);
  BUFF I5 (o_0r0[5:5], i_0r);
  BUFF I6 (o_0r0[6:6], i_0r);
  BUFF I7 (o_0r0[7:7], i_0r);
  GND I8 (o_0r1[0:0]);
  GND I9 (o_0r1[1:1]);
  GND I10 (o_0r1[2:2]);
  GND I11 (o_0r1[3:3]);
  GND I12 (o_0r1[4:4]);
  GND I13 (o_0r1[5:5]);
  GND I14 (o_0r1[6:6]);
  GND I15 (o_0r1[7:7]);
  BUFF I16 (i_0a, o_0a);
endmodule

// tkj32m8_24 TeakJ [Many [8,24],One 32]
module tkj32m8_24 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [7:0] i_0r0;
  input [7:0] i_0r1;
  output i_0a;
  input [23:0] i_1r0;
  input [23:0] i_1r1;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [31:0] joinf_0;
  wire [31:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_1r0[0:0]);
  BUFF I9 (joinf_0[9:9], i_1r0[1:1]);
  BUFF I10 (joinf_0[10:10], i_1r0[2:2]);
  BUFF I11 (joinf_0[11:11], i_1r0[3:3]);
  BUFF I12 (joinf_0[12:12], i_1r0[4:4]);
  BUFF I13 (joinf_0[13:13], i_1r0[5:5]);
  BUFF I14 (joinf_0[14:14], i_1r0[6:6]);
  BUFF I15 (joinf_0[15:15], i_1r0[7:7]);
  BUFF I16 (joinf_0[16:16], i_1r0[8:8]);
  BUFF I17 (joinf_0[17:17], i_1r0[9:9]);
  BUFF I18 (joinf_0[18:18], i_1r0[10:10]);
  BUFF I19 (joinf_0[19:19], i_1r0[11:11]);
  BUFF I20 (joinf_0[20:20], i_1r0[12:12]);
  BUFF I21 (joinf_0[21:21], i_1r0[13:13]);
  BUFF I22 (joinf_0[22:22], i_1r0[14:14]);
  BUFF I23 (joinf_0[23:23], i_1r0[15:15]);
  BUFF I24 (joinf_0[24:24], i_1r0[16:16]);
  BUFF I25 (joinf_0[25:25], i_1r0[17:17]);
  BUFF I26 (joinf_0[26:26], i_1r0[18:18]);
  BUFF I27 (joinf_0[27:27], i_1r0[19:19]);
  BUFF I28 (joinf_0[28:28], i_1r0[20:20]);
  BUFF I29 (joinf_0[29:29], i_1r0[21:21]);
  BUFF I30 (joinf_0[30:30], i_1r0[22:22]);
  BUFF I31 (joinf_0[31:31], i_1r0[23:23]);
  BUFF I32 (joint_0[0:0], i_0r1[0:0]);
  BUFF I33 (joint_0[1:1], i_0r1[1:1]);
  BUFF I34 (joint_0[2:2], i_0r1[2:2]);
  BUFF I35 (joint_0[3:3], i_0r1[3:3]);
  BUFF I36 (joint_0[4:4], i_0r1[4:4]);
  BUFF I37 (joint_0[5:5], i_0r1[5:5]);
  BUFF I38 (joint_0[6:6], i_0r1[6:6]);
  BUFF I39 (joint_0[7:7], i_0r1[7:7]);
  BUFF I40 (joint_0[8:8], i_1r1[0:0]);
  BUFF I41 (joint_0[9:9], i_1r1[1:1]);
  BUFF I42 (joint_0[10:10], i_1r1[2:2]);
  BUFF I43 (joint_0[11:11], i_1r1[3:3]);
  BUFF I44 (joint_0[12:12], i_1r1[4:4]);
  BUFF I45 (joint_0[13:13], i_1r1[5:5]);
  BUFF I46 (joint_0[14:14], i_1r1[6:6]);
  BUFF I47 (joint_0[15:15], i_1r1[7:7]);
  BUFF I48 (joint_0[16:16], i_1r1[8:8]);
  BUFF I49 (joint_0[17:17], i_1r1[9:9]);
  BUFF I50 (joint_0[18:18], i_1r1[10:10]);
  BUFF I51 (joint_0[19:19], i_1r1[11:11]);
  BUFF I52 (joint_0[20:20], i_1r1[12:12]);
  BUFF I53 (joint_0[21:21], i_1r1[13:13]);
  BUFF I54 (joint_0[22:22], i_1r1[14:14]);
  BUFF I55 (joint_0[23:23], i_1r1[15:15]);
  BUFF I56 (joint_0[24:24], i_1r1[16:16]);
  BUFF I57 (joint_0[25:25], i_1r1[17:17]);
  BUFF I58 (joint_0[26:26], i_1r1[18:18]);
  BUFF I59 (joint_0[27:27], i_1r1[19:19]);
  BUFF I60 (joint_0[28:28], i_1r1[20:20]);
  BUFF I61 (joint_0[29:29], i_1r1[21:21]);
  BUFF I62 (joint_0[30:30], i_1r1[22:22]);
  BUFF I63 (joint_0[31:31], i_1r1[23:23]);
  OR2 I64 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I65 (icomplete_0, dcomplete_0);
  C2 I66 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I67 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I68 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I69 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I70 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I71 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I72 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I73 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I74 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I75 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I76 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I77 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I78 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I79 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I80 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I81 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I82 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I83 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I84 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I85 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I86 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I87 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I88 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I89 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I90 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I91 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I92 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I93 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I94 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I95 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I96 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I97 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I98 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I99 (o_0r1[1:1], joint_0[1:1]);
  BUFF I100 (o_0r1[2:2], joint_0[2:2]);
  BUFF I101 (o_0r1[3:3], joint_0[3:3]);
  BUFF I102 (o_0r1[4:4], joint_0[4:4]);
  BUFF I103 (o_0r1[5:5], joint_0[5:5]);
  BUFF I104 (o_0r1[6:6], joint_0[6:6]);
  BUFF I105 (o_0r1[7:7], joint_0[7:7]);
  BUFF I106 (o_0r1[8:8], joint_0[8:8]);
  BUFF I107 (o_0r1[9:9], joint_0[9:9]);
  BUFF I108 (o_0r1[10:10], joint_0[10:10]);
  BUFF I109 (o_0r1[11:11], joint_0[11:11]);
  BUFF I110 (o_0r1[12:12], joint_0[12:12]);
  BUFF I111 (o_0r1[13:13], joint_0[13:13]);
  BUFF I112 (o_0r1[14:14], joint_0[14:14]);
  BUFF I113 (o_0r1[15:15], joint_0[15:15]);
  BUFF I114 (o_0r1[16:16], joint_0[16:16]);
  BUFF I115 (o_0r1[17:17], joint_0[17:17]);
  BUFF I116 (o_0r1[18:18], joint_0[18:18]);
  BUFF I117 (o_0r1[19:19], joint_0[19:19]);
  BUFF I118 (o_0r1[20:20], joint_0[20:20]);
  BUFF I119 (o_0r1[21:21], joint_0[21:21]);
  BUFF I120 (o_0r1[22:22], joint_0[22:22]);
  BUFF I121 (o_0r1[23:23], joint_0[23:23]);
  BUFF I122 (o_0r1[24:24], joint_0[24:24]);
  BUFF I123 (o_0r1[25:25], joint_0[25:25]);
  BUFF I124 (o_0r1[26:26], joint_0[26:26]);
  BUFF I125 (o_0r1[27:27], joint_0[27:27]);
  BUFF I126 (o_0r1[28:28], joint_0[28:28]);
  BUFF I127 (o_0r1[29:29], joint_0[29:29]);
  BUFF I128 (o_0r1[30:30], joint_0[30:30]);
  BUFF I129 (o_0r1[31:31], joint_0[31:31]);
  BUFF I130 (i_0a, o_0a);
  BUFF I131 (i_1a, o_0a);
endmodule

// tkj32m24_8 TeakJ [Many [24,8],One 32]
module tkj32m24_8 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [23:0] i_0r0;
  input [23:0] i_0r1;
  output i_0a;
  input [7:0] i_1r0;
  input [7:0] i_1r1;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [31:0] joinf_0;
  wire [31:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_1r0[0:0]);
  BUFF I25 (joinf_0[25:25], i_1r0[1:1]);
  BUFF I26 (joinf_0[26:26], i_1r0[2:2]);
  BUFF I27 (joinf_0[27:27], i_1r0[3:3]);
  BUFF I28 (joinf_0[28:28], i_1r0[4:4]);
  BUFF I29 (joinf_0[29:29], i_1r0[5:5]);
  BUFF I30 (joinf_0[30:30], i_1r0[6:6]);
  BUFF I31 (joinf_0[31:31], i_1r0[7:7]);
  BUFF I32 (joint_0[0:0], i_0r1[0:0]);
  BUFF I33 (joint_0[1:1], i_0r1[1:1]);
  BUFF I34 (joint_0[2:2], i_0r1[2:2]);
  BUFF I35 (joint_0[3:3], i_0r1[3:3]);
  BUFF I36 (joint_0[4:4], i_0r1[4:4]);
  BUFF I37 (joint_0[5:5], i_0r1[5:5]);
  BUFF I38 (joint_0[6:6], i_0r1[6:6]);
  BUFF I39 (joint_0[7:7], i_0r1[7:7]);
  BUFF I40 (joint_0[8:8], i_0r1[8:8]);
  BUFF I41 (joint_0[9:9], i_0r1[9:9]);
  BUFF I42 (joint_0[10:10], i_0r1[10:10]);
  BUFF I43 (joint_0[11:11], i_0r1[11:11]);
  BUFF I44 (joint_0[12:12], i_0r1[12:12]);
  BUFF I45 (joint_0[13:13], i_0r1[13:13]);
  BUFF I46 (joint_0[14:14], i_0r1[14:14]);
  BUFF I47 (joint_0[15:15], i_0r1[15:15]);
  BUFF I48 (joint_0[16:16], i_0r1[16:16]);
  BUFF I49 (joint_0[17:17], i_0r1[17:17]);
  BUFF I50 (joint_0[18:18], i_0r1[18:18]);
  BUFF I51 (joint_0[19:19], i_0r1[19:19]);
  BUFF I52 (joint_0[20:20], i_0r1[20:20]);
  BUFF I53 (joint_0[21:21], i_0r1[21:21]);
  BUFF I54 (joint_0[22:22], i_0r1[22:22]);
  BUFF I55 (joint_0[23:23], i_0r1[23:23]);
  BUFF I56 (joint_0[24:24], i_1r1[0:0]);
  BUFF I57 (joint_0[25:25], i_1r1[1:1]);
  BUFF I58 (joint_0[26:26], i_1r1[2:2]);
  BUFF I59 (joint_0[27:27], i_1r1[3:3]);
  BUFF I60 (joint_0[28:28], i_1r1[4:4]);
  BUFF I61 (joint_0[29:29], i_1r1[5:5]);
  BUFF I62 (joint_0[30:30], i_1r1[6:6]);
  BUFF I63 (joint_0[31:31], i_1r1[7:7]);
  OR2 I64 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I65 (icomplete_0, dcomplete_0);
  C2 I66 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I67 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I68 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I69 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I70 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I71 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I72 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I73 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I74 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I75 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I76 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I77 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I78 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I79 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I80 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I81 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I82 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I83 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I84 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I85 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I86 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I87 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I88 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I89 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I90 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I91 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I92 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I93 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I94 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I95 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I96 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I97 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I98 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I99 (o_0r1[1:1], joint_0[1:1]);
  BUFF I100 (o_0r1[2:2], joint_0[2:2]);
  BUFF I101 (o_0r1[3:3], joint_0[3:3]);
  BUFF I102 (o_0r1[4:4], joint_0[4:4]);
  BUFF I103 (o_0r1[5:5], joint_0[5:5]);
  BUFF I104 (o_0r1[6:6], joint_0[6:6]);
  BUFF I105 (o_0r1[7:7], joint_0[7:7]);
  BUFF I106 (o_0r1[8:8], joint_0[8:8]);
  BUFF I107 (o_0r1[9:9], joint_0[9:9]);
  BUFF I108 (o_0r1[10:10], joint_0[10:10]);
  BUFF I109 (o_0r1[11:11], joint_0[11:11]);
  BUFF I110 (o_0r1[12:12], joint_0[12:12]);
  BUFF I111 (o_0r1[13:13], joint_0[13:13]);
  BUFF I112 (o_0r1[14:14], joint_0[14:14]);
  BUFF I113 (o_0r1[15:15], joint_0[15:15]);
  BUFF I114 (o_0r1[16:16], joint_0[16:16]);
  BUFF I115 (o_0r1[17:17], joint_0[17:17]);
  BUFF I116 (o_0r1[18:18], joint_0[18:18]);
  BUFF I117 (o_0r1[19:19], joint_0[19:19]);
  BUFF I118 (o_0r1[20:20], joint_0[20:20]);
  BUFF I119 (o_0r1[21:21], joint_0[21:21]);
  BUFF I120 (o_0r1[22:22], joint_0[22:22]);
  BUFF I121 (o_0r1[23:23], joint_0[23:23]);
  BUFF I122 (o_0r1[24:24], joint_0[24:24]);
  BUFF I123 (o_0r1[25:25], joint_0[25:25]);
  BUFF I124 (o_0r1[26:26], joint_0[26:26]);
  BUFF I125 (o_0r1[27:27], joint_0[27:27]);
  BUFF I126 (o_0r1[28:28], joint_0[28:28]);
  BUFF I127 (o_0r1[29:29], joint_0[29:29]);
  BUFF I128 (o_0r1[30:30], joint_0[30:30]);
  BUFF I129 (o_0r1[31:31], joint_0[31:31]);
  BUFF I130 (i_0a, o_0a);
  BUFF I131 (i_1a, o_0a);
endmodule

// tko0m8_1nm8bff TeakO [
//     (1,TeakOConstant 8 255)] [One 0,One 8]
module tko0m8_1nm8bff (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [7:0] o_0r0;
  output [7:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  BUFF I1 (o_0r1[1:1], i_0r);
  BUFF I2 (o_0r1[2:2], i_0r);
  BUFF I3 (o_0r1[3:3], i_0r);
  BUFF I4 (o_0r1[4:4], i_0r);
  BUFF I5 (o_0r1[5:5], i_0r);
  BUFF I6 (o_0r1[6:6], i_0r);
  BUFF I7 (o_0r1[7:7], i_0r);
  GND I8 (o_0r0[0:0]);
  GND I9 (o_0r0[1:1]);
  GND I10 (o_0r0[2:2]);
  GND I11 (o_0r0[3:3]);
  GND I12 (o_0r0[4:4]);
  GND I13 (o_0r0[5:5]);
  GND I14 (o_0r0[6:6]);
  GND I15 (o_0r0[7:7]);
  BUFF I16 (i_0a, o_0a);
endmodule

// tkvi32_wo0w32_ro0w32o0w24o8w24o8w24 TeakV "i" 32 [] [0] [0,0,8,8] [Many [32],Many [0],Many [0,0,0,0]
//   ,Many [32,24,24,24]]
module tkvi32_wo0w32_ro0w32o0w24o8w24o8w24 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [23:0] rd_1r0;
  output [23:0] rd_1r1;
  input rd_1a;
  output [23:0] rd_2r0;
  output [23:0] rd_2r1;
  input rd_2a;
  output [23:0] rd_3r0;
  output [23:0] rd_3r1;
  input rd_3a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [2:0] simp6161_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_2r0[0:0], df_0[8:8], rg_2r);
  AND2 I481 (rd_2r0[1:1], df_0[9:9], rg_2r);
  AND2 I482 (rd_2r0[2:2], df_0[10:10], rg_2r);
  AND2 I483 (rd_2r0[3:3], df_0[11:11], rg_2r);
  AND2 I484 (rd_2r0[4:4], df_0[12:12], rg_2r);
  AND2 I485 (rd_2r0[5:5], df_0[13:13], rg_2r);
  AND2 I486 (rd_2r0[6:6], df_0[14:14], rg_2r);
  AND2 I487 (rd_2r0[7:7], df_0[15:15], rg_2r);
  AND2 I488 (rd_2r0[8:8], df_0[16:16], rg_2r);
  AND2 I489 (rd_2r0[9:9], df_0[17:17], rg_2r);
  AND2 I490 (rd_2r0[10:10], df_0[18:18], rg_2r);
  AND2 I491 (rd_2r0[11:11], df_0[19:19], rg_2r);
  AND2 I492 (rd_2r0[12:12], df_0[20:20], rg_2r);
  AND2 I493 (rd_2r0[13:13], df_0[21:21], rg_2r);
  AND2 I494 (rd_2r0[14:14], df_0[22:22], rg_2r);
  AND2 I495 (rd_2r0[15:15], df_0[23:23], rg_2r);
  AND2 I496 (rd_2r0[16:16], df_0[24:24], rg_2r);
  AND2 I497 (rd_2r0[17:17], df_0[25:25], rg_2r);
  AND2 I498 (rd_2r0[18:18], df_0[26:26], rg_2r);
  AND2 I499 (rd_2r0[19:19], df_0[27:27], rg_2r);
  AND2 I500 (rd_2r0[20:20], df_0[28:28], rg_2r);
  AND2 I501 (rd_2r0[21:21], df_0[29:29], rg_2r);
  AND2 I502 (rd_2r0[22:22], df_0[30:30], rg_2r);
  AND2 I503 (rd_2r0[23:23], df_0[31:31], rg_2r);
  AND2 I504 (rd_3r0[0:0], df_0[8:8], rg_3r);
  AND2 I505 (rd_3r0[1:1], df_0[9:9], rg_3r);
  AND2 I506 (rd_3r0[2:2], df_0[10:10], rg_3r);
  AND2 I507 (rd_3r0[3:3], df_0[11:11], rg_3r);
  AND2 I508 (rd_3r0[4:4], df_0[12:12], rg_3r);
  AND2 I509 (rd_3r0[5:5], df_0[13:13], rg_3r);
  AND2 I510 (rd_3r0[6:6], df_0[14:14], rg_3r);
  AND2 I511 (rd_3r0[7:7], df_0[15:15], rg_3r);
  AND2 I512 (rd_3r0[8:8], df_0[16:16], rg_3r);
  AND2 I513 (rd_3r0[9:9], df_0[17:17], rg_3r);
  AND2 I514 (rd_3r0[10:10], df_0[18:18], rg_3r);
  AND2 I515 (rd_3r0[11:11], df_0[19:19], rg_3r);
  AND2 I516 (rd_3r0[12:12], df_0[20:20], rg_3r);
  AND2 I517 (rd_3r0[13:13], df_0[21:21], rg_3r);
  AND2 I518 (rd_3r0[14:14], df_0[22:22], rg_3r);
  AND2 I519 (rd_3r0[15:15], df_0[23:23], rg_3r);
  AND2 I520 (rd_3r0[16:16], df_0[24:24], rg_3r);
  AND2 I521 (rd_3r0[17:17], df_0[25:25], rg_3r);
  AND2 I522 (rd_3r0[18:18], df_0[26:26], rg_3r);
  AND2 I523 (rd_3r0[19:19], df_0[27:27], rg_3r);
  AND2 I524 (rd_3r0[20:20], df_0[28:28], rg_3r);
  AND2 I525 (rd_3r0[21:21], df_0[29:29], rg_3r);
  AND2 I526 (rd_3r0[22:22], df_0[30:30], rg_3r);
  AND2 I527 (rd_3r0[23:23], df_0[31:31], rg_3r);
  AND2 I528 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I529 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I530 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I531 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I532 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I533 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I534 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I535 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I536 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I537 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I538 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I539 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I540 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I541 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I542 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I543 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I544 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I545 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I546 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I547 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I548 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I549 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I550 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I551 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I552 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I553 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I554 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I555 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I556 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I557 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I558 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I559 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I560 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I561 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I562 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I563 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I564 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I565 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I566 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I567 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I568 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I569 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I570 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I571 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I572 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I573 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I574 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I575 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I576 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I577 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I578 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I579 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I580 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I581 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I582 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I583 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[8:8], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[9:9], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[10:10], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[11:11], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[12:12], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[13:13], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[14:14], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[15:15], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[16:16], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[17:17], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[18:18], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[19:19], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[20:20], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[21:21], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[22:22], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[23:23], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[24:24], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[25:25], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[26:26], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[27:27], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[28:28], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[29:29], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[30:30], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[31:31], rg_2r);
  AND2 I608 (rd_3r1[0:0], dt_0[8:8], rg_3r);
  AND2 I609 (rd_3r1[1:1], dt_0[9:9], rg_3r);
  AND2 I610 (rd_3r1[2:2], dt_0[10:10], rg_3r);
  AND2 I611 (rd_3r1[3:3], dt_0[11:11], rg_3r);
  AND2 I612 (rd_3r1[4:4], dt_0[12:12], rg_3r);
  AND2 I613 (rd_3r1[5:5], dt_0[13:13], rg_3r);
  AND2 I614 (rd_3r1[6:6], dt_0[14:14], rg_3r);
  AND2 I615 (rd_3r1[7:7], dt_0[15:15], rg_3r);
  AND2 I616 (rd_3r1[8:8], dt_0[16:16], rg_3r);
  AND2 I617 (rd_3r1[9:9], dt_0[17:17], rg_3r);
  AND2 I618 (rd_3r1[10:10], dt_0[18:18], rg_3r);
  AND2 I619 (rd_3r1[11:11], dt_0[19:19], rg_3r);
  AND2 I620 (rd_3r1[12:12], dt_0[20:20], rg_3r);
  AND2 I621 (rd_3r1[13:13], dt_0[21:21], rg_3r);
  AND2 I622 (rd_3r1[14:14], dt_0[22:22], rg_3r);
  AND2 I623 (rd_3r1[15:15], dt_0[23:23], rg_3r);
  AND2 I624 (rd_3r1[16:16], dt_0[24:24], rg_3r);
  AND2 I625 (rd_3r1[17:17], dt_0[25:25], rg_3r);
  AND2 I626 (rd_3r1[18:18], dt_0[26:26], rg_3r);
  AND2 I627 (rd_3r1[19:19], dt_0[27:27], rg_3r);
  AND2 I628 (rd_3r1[20:20], dt_0[28:28], rg_3r);
  AND2 I629 (rd_3r1[21:21], dt_0[29:29], rg_3r);
  AND2 I630 (rd_3r1[22:22], dt_0[30:30], rg_3r);
  AND2 I631 (rd_3r1[23:23], dt_0[31:31], rg_3r);
  NOR3 I632 (simp6161_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I633 (simp6161_0[1:1], rg_3r, rg_0a, rg_1a);
  NOR2 I634 (simp6161_0[2:2], rg_2a, rg_3a);
  NAND3 I635 (anyread_0, simp6161_0[0:0], simp6161_0[1:1], simp6161_0[2:2]);
  BUFF I636 (wg_0a, wd_0a);
  BUFF I637 (rg_0a, rd_0a);
  BUFF I638 (rg_1a, rd_1a);
  BUFF I639 (rg_2a, rd_2a);
  BUFF I640 (rg_3a, rd_3a);
endmodule

// tko0m16_1nm16b0 TeakO [
//     (1,TeakOConstant 16 0)] [One 0,One 16]
module tko0m16_1nm16b0 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [15:0] o_0r0;
  output [15:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r0[0:0], i_0r);
  BUFF I1 (o_0r0[1:1], i_0r);
  BUFF I2 (o_0r0[2:2], i_0r);
  BUFF I3 (o_0r0[3:3], i_0r);
  BUFF I4 (o_0r0[4:4], i_0r);
  BUFF I5 (o_0r0[5:5], i_0r);
  BUFF I6 (o_0r0[6:6], i_0r);
  BUFF I7 (o_0r0[7:7], i_0r);
  BUFF I8 (o_0r0[8:8], i_0r);
  BUFF I9 (o_0r0[9:9], i_0r);
  BUFF I10 (o_0r0[10:10], i_0r);
  BUFF I11 (o_0r0[11:11], i_0r);
  BUFF I12 (o_0r0[12:12], i_0r);
  BUFF I13 (o_0r0[13:13], i_0r);
  BUFF I14 (o_0r0[14:14], i_0r);
  BUFF I15 (o_0r0[15:15], i_0r);
  GND I16 (o_0r1[0:0]);
  GND I17 (o_0r1[1:1]);
  GND I18 (o_0r1[2:2]);
  GND I19 (o_0r1[3:3]);
  GND I20 (o_0r1[4:4]);
  GND I21 (o_0r1[5:5]);
  GND I22 (o_0r1[6:6]);
  GND I23 (o_0r1[7:7]);
  GND I24 (o_0r1[8:8]);
  GND I25 (o_0r1[9:9]);
  GND I26 (o_0r1[10:10]);
  GND I27 (o_0r1[11:11]);
  GND I28 (o_0r1[12:12]);
  GND I29 (o_0r1[13:13]);
  GND I30 (o_0r1[14:14]);
  GND I31 (o_0r1[15:15]);
  BUFF I32 (i_0a, o_0a);
endmodule

// tkj32m16_16 TeakJ [Many [16,16],One 32]
module tkj32m16_16 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [15:0] i_0r0;
  input [15:0] i_0r1;
  output i_0a;
  input [15:0] i_1r0;
  input [15:0] i_1r1;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [31:0] joinf_0;
  wire [31:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_1r0[0:0]);
  BUFF I17 (joinf_0[17:17], i_1r0[1:1]);
  BUFF I18 (joinf_0[18:18], i_1r0[2:2]);
  BUFF I19 (joinf_0[19:19], i_1r0[3:3]);
  BUFF I20 (joinf_0[20:20], i_1r0[4:4]);
  BUFF I21 (joinf_0[21:21], i_1r0[5:5]);
  BUFF I22 (joinf_0[22:22], i_1r0[6:6]);
  BUFF I23 (joinf_0[23:23], i_1r0[7:7]);
  BUFF I24 (joinf_0[24:24], i_1r0[8:8]);
  BUFF I25 (joinf_0[25:25], i_1r0[9:9]);
  BUFF I26 (joinf_0[26:26], i_1r0[10:10]);
  BUFF I27 (joinf_0[27:27], i_1r0[11:11]);
  BUFF I28 (joinf_0[28:28], i_1r0[12:12]);
  BUFF I29 (joinf_0[29:29], i_1r0[13:13]);
  BUFF I30 (joinf_0[30:30], i_1r0[14:14]);
  BUFF I31 (joinf_0[31:31], i_1r0[15:15]);
  BUFF I32 (joint_0[0:0], i_0r1[0:0]);
  BUFF I33 (joint_0[1:1], i_0r1[1:1]);
  BUFF I34 (joint_0[2:2], i_0r1[2:2]);
  BUFF I35 (joint_0[3:3], i_0r1[3:3]);
  BUFF I36 (joint_0[4:4], i_0r1[4:4]);
  BUFF I37 (joint_0[5:5], i_0r1[5:5]);
  BUFF I38 (joint_0[6:6], i_0r1[6:6]);
  BUFF I39 (joint_0[7:7], i_0r1[7:7]);
  BUFF I40 (joint_0[8:8], i_0r1[8:8]);
  BUFF I41 (joint_0[9:9], i_0r1[9:9]);
  BUFF I42 (joint_0[10:10], i_0r1[10:10]);
  BUFF I43 (joint_0[11:11], i_0r1[11:11]);
  BUFF I44 (joint_0[12:12], i_0r1[12:12]);
  BUFF I45 (joint_0[13:13], i_0r1[13:13]);
  BUFF I46 (joint_0[14:14], i_0r1[14:14]);
  BUFF I47 (joint_0[15:15], i_0r1[15:15]);
  BUFF I48 (joint_0[16:16], i_1r1[0:0]);
  BUFF I49 (joint_0[17:17], i_1r1[1:1]);
  BUFF I50 (joint_0[18:18], i_1r1[2:2]);
  BUFF I51 (joint_0[19:19], i_1r1[3:3]);
  BUFF I52 (joint_0[20:20], i_1r1[4:4]);
  BUFF I53 (joint_0[21:21], i_1r1[5:5]);
  BUFF I54 (joint_0[22:22], i_1r1[6:6]);
  BUFF I55 (joint_0[23:23], i_1r1[7:7]);
  BUFF I56 (joint_0[24:24], i_1r1[8:8]);
  BUFF I57 (joint_0[25:25], i_1r1[9:9]);
  BUFF I58 (joint_0[26:26], i_1r1[10:10]);
  BUFF I59 (joint_0[27:27], i_1r1[11:11]);
  BUFF I60 (joint_0[28:28], i_1r1[12:12]);
  BUFF I61 (joint_0[29:29], i_1r1[13:13]);
  BUFF I62 (joint_0[30:30], i_1r1[14:14]);
  BUFF I63 (joint_0[31:31], i_1r1[15:15]);
  OR2 I64 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I65 (icomplete_0, dcomplete_0);
  C2 I66 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I67 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I68 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I69 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I70 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I71 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I72 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I73 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I74 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I75 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I76 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I77 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I78 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I79 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I80 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I81 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I82 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I83 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I84 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I85 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I86 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I87 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I88 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I89 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I90 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I91 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I92 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I93 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I94 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I95 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I96 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I97 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I98 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I99 (o_0r1[1:1], joint_0[1:1]);
  BUFF I100 (o_0r1[2:2], joint_0[2:2]);
  BUFF I101 (o_0r1[3:3], joint_0[3:3]);
  BUFF I102 (o_0r1[4:4], joint_0[4:4]);
  BUFF I103 (o_0r1[5:5], joint_0[5:5]);
  BUFF I104 (o_0r1[6:6], joint_0[6:6]);
  BUFF I105 (o_0r1[7:7], joint_0[7:7]);
  BUFF I106 (o_0r1[8:8], joint_0[8:8]);
  BUFF I107 (o_0r1[9:9], joint_0[9:9]);
  BUFF I108 (o_0r1[10:10], joint_0[10:10]);
  BUFF I109 (o_0r1[11:11], joint_0[11:11]);
  BUFF I110 (o_0r1[12:12], joint_0[12:12]);
  BUFF I111 (o_0r1[13:13], joint_0[13:13]);
  BUFF I112 (o_0r1[14:14], joint_0[14:14]);
  BUFF I113 (o_0r1[15:15], joint_0[15:15]);
  BUFF I114 (o_0r1[16:16], joint_0[16:16]);
  BUFF I115 (o_0r1[17:17], joint_0[17:17]);
  BUFF I116 (o_0r1[18:18], joint_0[18:18]);
  BUFF I117 (o_0r1[19:19], joint_0[19:19]);
  BUFF I118 (o_0r1[20:20], joint_0[20:20]);
  BUFF I119 (o_0r1[21:21], joint_0[21:21]);
  BUFF I120 (o_0r1[22:22], joint_0[22:22]);
  BUFF I121 (o_0r1[23:23], joint_0[23:23]);
  BUFF I122 (o_0r1[24:24], joint_0[24:24]);
  BUFF I123 (o_0r1[25:25], joint_0[25:25]);
  BUFF I124 (o_0r1[26:26], joint_0[26:26]);
  BUFF I125 (o_0r1[27:27], joint_0[27:27]);
  BUFF I126 (o_0r1[28:28], joint_0[28:28]);
  BUFF I127 (o_0r1[29:29], joint_0[29:29]);
  BUFF I128 (o_0r1[30:30], joint_0[30:30]);
  BUFF I129 (o_0r1[31:31], joint_0[31:31]);
  BUFF I130 (i_0a, o_0a);
  BUFF I131 (i_1a, o_0a);
endmodule

// tko0m16_1nm16bffff TeakO [
//     (1,TeakOConstant 16 65535)] [One 0,One 16]
module tko0m16_1nm16bffff (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [15:0] o_0r0;
  output [15:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  BUFF I1 (o_0r1[1:1], i_0r);
  BUFF I2 (o_0r1[2:2], i_0r);
  BUFF I3 (o_0r1[3:3], i_0r);
  BUFF I4 (o_0r1[4:4], i_0r);
  BUFF I5 (o_0r1[5:5], i_0r);
  BUFF I6 (o_0r1[6:6], i_0r);
  BUFF I7 (o_0r1[7:7], i_0r);
  BUFF I8 (o_0r1[8:8], i_0r);
  BUFF I9 (o_0r1[9:9], i_0r);
  BUFF I10 (o_0r1[10:10], i_0r);
  BUFF I11 (o_0r1[11:11], i_0r);
  BUFF I12 (o_0r1[12:12], i_0r);
  BUFF I13 (o_0r1[13:13], i_0r);
  BUFF I14 (o_0r1[14:14], i_0r);
  BUFF I15 (o_0r1[15:15], i_0r);
  GND I16 (o_0r0[0:0]);
  GND I17 (o_0r0[1:1]);
  GND I18 (o_0r0[2:2]);
  GND I19 (o_0r0[3:3]);
  GND I20 (o_0r0[4:4]);
  GND I21 (o_0r0[5:5]);
  GND I22 (o_0r0[6:6]);
  GND I23 (o_0r0[7:7]);
  GND I24 (o_0r0[8:8]);
  GND I25 (o_0r0[9:9]);
  GND I26 (o_0r0[10:10]);
  GND I27 (o_0r0[11:11]);
  GND I28 (o_0r0[12:12]);
  GND I29 (o_0r0[13:13]);
  GND I30 (o_0r0[14:14]);
  GND I31 (o_0r0[15:15]);
  BUFF I32 (i_0a, o_0a);
endmodule

// tkvi32_wo0w32_ro0w32o0w16o16w16o16w16 TeakV "i" 32 [] [0] [0,0,16,16] [Many [32],Many [0],Many [0,0,
//   0,0],Many [32,16,16,16]]
module tkvi32_wo0w32_ro0w32o0w16o16w16o16w16 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [15:0] rd_1r0;
  output [15:0] rd_1r1;
  input rd_1a;
  output [15:0] rd_2r0;
  output [15:0] rd_2r1;
  input rd_2a;
  output [15:0] rd_3r0;
  output [15:0] rd_3r1;
  input rd_3a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [2:0] simp5681_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_2r0[0:0], df_0[16:16], rg_2r);
  AND2 I473 (rd_2r0[1:1], df_0[17:17], rg_2r);
  AND2 I474 (rd_2r0[2:2], df_0[18:18], rg_2r);
  AND2 I475 (rd_2r0[3:3], df_0[19:19], rg_2r);
  AND2 I476 (rd_2r0[4:4], df_0[20:20], rg_2r);
  AND2 I477 (rd_2r0[5:5], df_0[21:21], rg_2r);
  AND2 I478 (rd_2r0[6:6], df_0[22:22], rg_2r);
  AND2 I479 (rd_2r0[7:7], df_0[23:23], rg_2r);
  AND2 I480 (rd_2r0[8:8], df_0[24:24], rg_2r);
  AND2 I481 (rd_2r0[9:9], df_0[25:25], rg_2r);
  AND2 I482 (rd_2r0[10:10], df_0[26:26], rg_2r);
  AND2 I483 (rd_2r0[11:11], df_0[27:27], rg_2r);
  AND2 I484 (rd_2r0[12:12], df_0[28:28], rg_2r);
  AND2 I485 (rd_2r0[13:13], df_0[29:29], rg_2r);
  AND2 I486 (rd_2r0[14:14], df_0[30:30], rg_2r);
  AND2 I487 (rd_2r0[15:15], df_0[31:31], rg_2r);
  AND2 I488 (rd_3r0[0:0], df_0[16:16], rg_3r);
  AND2 I489 (rd_3r0[1:1], df_0[17:17], rg_3r);
  AND2 I490 (rd_3r0[2:2], df_0[18:18], rg_3r);
  AND2 I491 (rd_3r0[3:3], df_0[19:19], rg_3r);
  AND2 I492 (rd_3r0[4:4], df_0[20:20], rg_3r);
  AND2 I493 (rd_3r0[5:5], df_0[21:21], rg_3r);
  AND2 I494 (rd_3r0[6:6], df_0[22:22], rg_3r);
  AND2 I495 (rd_3r0[7:7], df_0[23:23], rg_3r);
  AND2 I496 (rd_3r0[8:8], df_0[24:24], rg_3r);
  AND2 I497 (rd_3r0[9:9], df_0[25:25], rg_3r);
  AND2 I498 (rd_3r0[10:10], df_0[26:26], rg_3r);
  AND2 I499 (rd_3r0[11:11], df_0[27:27], rg_3r);
  AND2 I500 (rd_3r0[12:12], df_0[28:28], rg_3r);
  AND2 I501 (rd_3r0[13:13], df_0[29:29], rg_3r);
  AND2 I502 (rd_3r0[14:14], df_0[30:30], rg_3r);
  AND2 I503 (rd_3r0[15:15], df_0[31:31], rg_3r);
  AND2 I504 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I505 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I506 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I507 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I508 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I509 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I510 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I511 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I512 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I513 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I514 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I515 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I516 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I517 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I518 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I519 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I520 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I521 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I522 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I523 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I524 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I525 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I526 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I527 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I528 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I529 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I530 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I531 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I532 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I533 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I534 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I535 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I536 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I537 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I538 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I539 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I540 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I541 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I542 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I543 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I544 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I545 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I546 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I547 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I548 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I549 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I550 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I551 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I552 (rd_2r1[0:0], dt_0[16:16], rg_2r);
  AND2 I553 (rd_2r1[1:1], dt_0[17:17], rg_2r);
  AND2 I554 (rd_2r1[2:2], dt_0[18:18], rg_2r);
  AND2 I555 (rd_2r1[3:3], dt_0[19:19], rg_2r);
  AND2 I556 (rd_2r1[4:4], dt_0[20:20], rg_2r);
  AND2 I557 (rd_2r1[5:5], dt_0[21:21], rg_2r);
  AND2 I558 (rd_2r1[6:6], dt_0[22:22], rg_2r);
  AND2 I559 (rd_2r1[7:7], dt_0[23:23], rg_2r);
  AND2 I560 (rd_2r1[8:8], dt_0[24:24], rg_2r);
  AND2 I561 (rd_2r1[9:9], dt_0[25:25], rg_2r);
  AND2 I562 (rd_2r1[10:10], dt_0[26:26], rg_2r);
  AND2 I563 (rd_2r1[11:11], dt_0[27:27], rg_2r);
  AND2 I564 (rd_2r1[12:12], dt_0[28:28], rg_2r);
  AND2 I565 (rd_2r1[13:13], dt_0[29:29], rg_2r);
  AND2 I566 (rd_2r1[14:14], dt_0[30:30], rg_2r);
  AND2 I567 (rd_2r1[15:15], dt_0[31:31], rg_2r);
  AND2 I568 (rd_3r1[0:0], dt_0[16:16], rg_3r);
  AND2 I569 (rd_3r1[1:1], dt_0[17:17], rg_3r);
  AND2 I570 (rd_3r1[2:2], dt_0[18:18], rg_3r);
  AND2 I571 (rd_3r1[3:3], dt_0[19:19], rg_3r);
  AND2 I572 (rd_3r1[4:4], dt_0[20:20], rg_3r);
  AND2 I573 (rd_3r1[5:5], dt_0[21:21], rg_3r);
  AND2 I574 (rd_3r1[6:6], dt_0[22:22], rg_3r);
  AND2 I575 (rd_3r1[7:7], dt_0[23:23], rg_3r);
  AND2 I576 (rd_3r1[8:8], dt_0[24:24], rg_3r);
  AND2 I577 (rd_3r1[9:9], dt_0[25:25], rg_3r);
  AND2 I578 (rd_3r1[10:10], dt_0[26:26], rg_3r);
  AND2 I579 (rd_3r1[11:11], dt_0[27:27], rg_3r);
  AND2 I580 (rd_3r1[12:12], dt_0[28:28], rg_3r);
  AND2 I581 (rd_3r1[13:13], dt_0[29:29], rg_3r);
  AND2 I582 (rd_3r1[14:14], dt_0[30:30], rg_3r);
  AND2 I583 (rd_3r1[15:15], dt_0[31:31], rg_3r);
  NOR3 I584 (simp5681_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I585 (simp5681_0[1:1], rg_3r, rg_0a, rg_1a);
  NOR2 I586 (simp5681_0[2:2], rg_2a, rg_3a);
  NAND3 I587 (anyread_0, simp5681_0[0:0], simp5681_0[1:1], simp5681_0[2:2]);
  BUFF I588 (wg_0a, wd_0a);
  BUFF I589 (rg_0a, rd_0a);
  BUFF I590 (rg_1a, rd_1a);
  BUFF I591 (rg_2a, rd_2a);
  BUFF I592 (rg_3a, rd_3a);
endmodule

// tkvdistanceI5_wo0w5_ro0w1o1w1o2w1o3w1o4w1 TeakV "distanceI" 5 [] [0] [0,1,2,3,4] [Many [5],Many [0],
//   Many [0,0,0,0,0],Many [1,1,1,1,1]]
module tkvdistanceI5_wo0w5_ro0w1o1w1o2w1o3w1o4w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, reset);
  input [4:0] wg_0r0;
  input [4:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  output rd_1r0;
  output rd_1r1;
  input rd_1a;
  output rd_2r0;
  output rd_2r1;
  input rd_2a;
  output rd_3r0;
  output rd_3r1;
  input rd_3a;
  output rd_4r0;
  output rd_4r1;
  input rd_4a;
  input reset;
  wire [4:0] wf_0;
  wire [4:0] wt_0;
  wire [4:0] df_0;
  wire [4:0] dt_0;
  wire wc_0;
  wire [4:0] wacks_0;
  wire [4:0] wenr_0;
  wire [4:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [4:0] drlgf_0;
  wire [4:0] drlgt_0;
  wire [4:0] comp0_0;
  wire [1:0] simp491_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [4:0] conwgit_0;
  wire [4:0] conwgif_0;
  wire conwig_0;
  wire [1:0] simp831_0;
  wire [3:0] simp941_0;
  wire [1:0] simp942_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I7 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I8 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I9 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I10 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I11 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I12 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I13 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I14 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I15 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  NOR2 I16 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I17 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I18 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I19 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I20 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR3 I21 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I22 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I23 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I24 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I25 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  AO22 I26 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I27 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I28 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I29 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I30 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  OR2 I31 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I32 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I33 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I34 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I35 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  C3 I36 (simp491_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C2 I37 (simp491_0[1:1], comp0_0[3:3], comp0_0[4:4]);
  C2 I38 (wc_0, simp491_0[0:0], simp491_0[1:1]);
  AND2 I39 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I40 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I41 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I42 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I43 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I44 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I45 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I46 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I47 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I48 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  BUFF I49 (conwigc_0, wc_0);
  AO22 I50 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I51 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I52 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I53 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I54 (wenr_0[0:0], wc_0);
  BUFF I55 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I56 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I57 (wenr_0[1:1], wc_0);
  BUFF I58 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I59 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I60 (wenr_0[2:2], wc_0);
  BUFF I61 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I62 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I63 (wenr_0[3:3], wc_0);
  BUFF I64 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I65 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I66 (wenr_0[4:4], wc_0);
  C3 I67 (simp831_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I68 (simp831_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C2 I69 (wd_0r, simp831_0[0:0], simp831_0[1:1]);
  AND2 I70 (rd_0r0, df_0[0:0], rg_0r);
  AND2 I71 (rd_1r0, df_0[1:1], rg_1r);
  AND2 I72 (rd_2r0, df_0[2:2], rg_2r);
  AND2 I73 (rd_3r0, df_0[3:3], rg_3r);
  AND2 I74 (rd_4r0, df_0[4:4], rg_4r);
  AND2 I75 (rd_0r1, dt_0[0:0], rg_0r);
  AND2 I76 (rd_1r1, dt_0[1:1], rg_1r);
  AND2 I77 (rd_2r1, dt_0[2:2], rg_2r);
  AND2 I78 (rd_3r1, dt_0[3:3], rg_3r);
  AND2 I79 (rd_4r1, dt_0[4:4], rg_4r);
  NOR3 I80 (simp941_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I81 (simp941_0[1:1], rg_3r, rg_4r, rg_0a);
  NOR3 I82 (simp941_0[2:2], rg_1a, rg_2a, rg_3a);
  INV I83 (simp941_0[3:3], rg_4a);
  NAND3 I84 (simp942_0[0:0], simp941_0[0:0], simp941_0[1:1], simp941_0[2:2]);
  INV I85 (simp942_0[1:1], simp941_0[3:3]);
  OR2 I86 (anyread_0, simp942_0[0:0], simp942_0[1:1]);
  BUFF I87 (wg_0a, wd_0a);
  BUFF I88 (rg_0a, rd_0a);
  BUFF I89 (rg_1a, rd_1a);
  BUFF I90 (rg_2a, rd_2a);
  BUFF I91 (rg_3a, rd_3a);
  BUFF I92 (rg_4a, rd_4a);
endmodule

// tkvshift2_wo0w2_ro0w2o0w2o0w2o0w2o0w2 TeakV "shift" 2 [] [0] [0,0,0,0,0] [Many [2],Many [0],Many [0,
//   0,0,0,0],Many [2,2,2,2,2]]
module tkvshift2_wo0w2_ro0w2o0w2o0w2o0w2o0w2 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, reset);
  input [1:0] wg_0r0;
  input [1:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  output [1:0] rd_0r0;
  output [1:0] rd_0r1;
  input rd_0a;
  output [1:0] rd_1r0;
  output [1:0] rd_1r1;
  input rd_1a;
  output [1:0] rd_2r0;
  output [1:0] rd_2r1;
  input rd_2a;
  output [1:0] rd_3r0;
  output [1:0] rd_3r1;
  input rd_3a;
  output [1:0] rd_4r0;
  output [1:0] rd_4r1;
  input rd_4a;
  input reset;
  wire [1:0] wf_0;
  wire [1:0] wt_0;
  wire [1:0] df_0;
  wire [1:0] dt_0;
  wire wc_0;
  wire [1:0] wacks_0;
  wire [1:0] wenr_0;
  wire [1:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [1:0] drlgf_0;
  wire [1:0] drlgt_0;
  wire [1:0] comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [1:0] conwgit_0;
  wire [1:0] conwgif_0;
  wire conwig_0;
  wire [3:0] simp681_0;
  wire [1:0] simp682_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I4 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I5 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I6 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  NOR2 I7 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I8 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR3 I9 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I10 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  AO22 I11 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I12 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  OR2 I13 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I14 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  C2 I15 (wc_0, comp0_0[0:0], comp0_0[1:1]);
  AND2 I16 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I17 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I18 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I19 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  BUFF I20 (conwigc_0, wc_0);
  AO22 I21 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I22 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I23 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I24 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I25 (wenr_0[0:0], wc_0);
  BUFF I26 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I27 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I28 (wenr_0[1:1], wc_0);
  C3 I29 (wd_0r, conwig_0, wacks_0[0:0], wacks_0[1:1]);
  AND2 I30 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I31 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I32 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I33 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I34 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I35 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I36 (rd_3r0[0:0], df_0[0:0], rg_3r);
  AND2 I37 (rd_3r0[1:1], df_0[1:1], rg_3r);
  AND2 I38 (rd_4r0[0:0], df_0[0:0], rg_4r);
  AND2 I39 (rd_4r0[1:1], df_0[1:1], rg_4r);
  AND2 I40 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I41 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I42 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I43 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I44 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I45 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I46 (rd_3r1[0:0], dt_0[0:0], rg_3r);
  AND2 I47 (rd_3r1[1:1], dt_0[1:1], rg_3r);
  AND2 I48 (rd_4r1[0:0], dt_0[0:0], rg_4r);
  AND2 I49 (rd_4r1[1:1], dt_0[1:1], rg_4r);
  NOR3 I50 (simp681_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I51 (simp681_0[1:1], rg_3r, rg_4r, rg_0a);
  NOR3 I52 (simp681_0[2:2], rg_1a, rg_2a, rg_3a);
  INV I53 (simp681_0[3:3], rg_4a);
  NAND3 I54 (simp682_0[0:0], simp681_0[0:0], simp681_0[1:1], simp681_0[2:2]);
  INV I55 (simp682_0[1:1], simp681_0[3:3]);
  OR2 I56 (anyread_0, simp682_0[0:0], simp682_0[1:1]);
  BUFF I57 (wg_0a, wd_0a);
  BUFF I58 (rg_0a, rd_0a);
  BUFF I59 (rg_1a, rd_1a);
  BUFF I60 (rg_2a, rd_2a);
  BUFF I61 (rg_3a, rd_3a);
  BUFF I62 (rg_4a, rd_4a);
endmodule

// tkj2m2_0 TeakJ [Many [2,0],One 2]
module tkj2m2_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [1:0] joinf_0;
  wire [1:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joint_0[0:0], i_0r1[0:0]);
  BUFF I3 (joint_0[1:1], i_0r1[1:1]);
  BUFF I4 (icomplete_0, i_1r);
  C2 I5 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I6 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I7 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I8 (o_0r1[1:1], joint_0[1:1]);
  BUFF I9 (i_0a, o_0a);
  BUFF I10 (i_1a, o_0a);
endmodule

// tkj5m5_0 TeakJ [Many [5,0],One 5]
module tkj5m5_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [4:0] i_0r0;
  input [4:0] i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  output [4:0] o_0r0;
  output [4:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [4:0] joinf_0;
  wire [4:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joint_0[0:0], i_0r1[0:0]);
  BUFF I6 (joint_0[1:1], i_0r1[1:1]);
  BUFF I7 (joint_0[2:2], i_0r1[2:2]);
  BUFF I8 (joint_0[3:3], i_0r1[3:3]);
  BUFF I9 (joint_0[4:4], i_0r1[4:4]);
  BUFF I10 (icomplete_0, i_1r);
  C2 I11 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I12 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I13 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I14 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I15 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I16 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I17 (o_0r1[1:1], joint_0[1:1]);
  BUFF I18 (o_0r1[2:2], joint_0[2:2]);
  BUFF I19 (o_0r1[3:3], joint_0[3:3]);
  BUFF I20 (o_0r1[4:4], joint_0[4:4]);
  BUFF I21 (i_0a, o_0a);
  BUFF I22 (i_1a, o_0a);
endmodule

// tko32m32_1noti0w32b TeakO [
//     (1,TeakOp TeakOpNot [(0,0+:32)])] [One 32,One 32]
module tko32m32_1noti0w32b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r0[0:0]);
  BUFF I1 (o_0r0[0:0], i_0r1[0:0]);
  BUFF I2 (o_0r1[1:1], i_0r0[1:1]);
  BUFF I3 (o_0r0[1:1], i_0r1[1:1]);
  BUFF I4 (o_0r1[2:2], i_0r0[2:2]);
  BUFF I5 (o_0r0[2:2], i_0r1[2:2]);
  BUFF I6 (o_0r1[3:3], i_0r0[3:3]);
  BUFF I7 (o_0r0[3:3], i_0r1[3:3]);
  BUFF I8 (o_0r1[4:4], i_0r0[4:4]);
  BUFF I9 (o_0r0[4:4], i_0r1[4:4]);
  BUFF I10 (o_0r1[5:5], i_0r0[5:5]);
  BUFF I11 (o_0r0[5:5], i_0r1[5:5]);
  BUFF I12 (o_0r1[6:6], i_0r0[6:6]);
  BUFF I13 (o_0r0[6:6], i_0r1[6:6]);
  BUFF I14 (o_0r1[7:7], i_0r0[7:7]);
  BUFF I15 (o_0r0[7:7], i_0r1[7:7]);
  BUFF I16 (o_0r1[8:8], i_0r0[8:8]);
  BUFF I17 (o_0r0[8:8], i_0r1[8:8]);
  BUFF I18 (o_0r1[9:9], i_0r0[9:9]);
  BUFF I19 (o_0r0[9:9], i_0r1[9:9]);
  BUFF I20 (o_0r1[10:10], i_0r0[10:10]);
  BUFF I21 (o_0r0[10:10], i_0r1[10:10]);
  BUFF I22 (o_0r1[11:11], i_0r0[11:11]);
  BUFF I23 (o_0r0[11:11], i_0r1[11:11]);
  BUFF I24 (o_0r1[12:12], i_0r0[12:12]);
  BUFF I25 (o_0r0[12:12], i_0r1[12:12]);
  BUFF I26 (o_0r1[13:13], i_0r0[13:13]);
  BUFF I27 (o_0r0[13:13], i_0r1[13:13]);
  BUFF I28 (o_0r1[14:14], i_0r0[14:14]);
  BUFF I29 (o_0r0[14:14], i_0r1[14:14]);
  BUFF I30 (o_0r1[15:15], i_0r0[15:15]);
  BUFF I31 (o_0r0[15:15], i_0r1[15:15]);
  BUFF I32 (o_0r1[16:16], i_0r0[16:16]);
  BUFF I33 (o_0r0[16:16], i_0r1[16:16]);
  BUFF I34 (o_0r1[17:17], i_0r0[17:17]);
  BUFF I35 (o_0r0[17:17], i_0r1[17:17]);
  BUFF I36 (o_0r1[18:18], i_0r0[18:18]);
  BUFF I37 (o_0r0[18:18], i_0r1[18:18]);
  BUFF I38 (o_0r1[19:19], i_0r0[19:19]);
  BUFF I39 (o_0r0[19:19], i_0r1[19:19]);
  BUFF I40 (o_0r1[20:20], i_0r0[20:20]);
  BUFF I41 (o_0r0[20:20], i_0r1[20:20]);
  BUFF I42 (o_0r1[21:21], i_0r0[21:21]);
  BUFF I43 (o_0r0[21:21], i_0r1[21:21]);
  BUFF I44 (o_0r1[22:22], i_0r0[22:22]);
  BUFF I45 (o_0r0[22:22], i_0r1[22:22]);
  BUFF I46 (o_0r1[23:23], i_0r0[23:23]);
  BUFF I47 (o_0r0[23:23], i_0r1[23:23]);
  BUFF I48 (o_0r1[24:24], i_0r0[24:24]);
  BUFF I49 (o_0r0[24:24], i_0r1[24:24]);
  BUFF I50 (o_0r1[25:25], i_0r0[25:25]);
  BUFF I51 (o_0r0[25:25], i_0r1[25:25]);
  BUFF I52 (o_0r1[26:26], i_0r0[26:26]);
  BUFF I53 (o_0r0[26:26], i_0r1[26:26]);
  BUFF I54 (o_0r1[27:27], i_0r0[27:27]);
  BUFF I55 (o_0r0[27:27], i_0r1[27:27]);
  BUFF I56 (o_0r1[28:28], i_0r0[28:28]);
  BUFF I57 (o_0r0[28:28], i_0r1[28:28]);
  BUFF I58 (o_0r1[29:29], i_0r0[29:29]);
  BUFF I59 (o_0r0[29:29], i_0r1[29:29]);
  BUFF I60 (o_0r1[30:30], i_0r0[30:30]);
  BUFF I61 (o_0r0[30:30], i_0r1[30:30]);
  BUFF I62 (o_0r1[31:31], i_0r0[31:31]);
  BUFF I63 (o_0r0[31:31], i_0r1[31:31]);
  BUFF I64 (i_0a, o_0a);
endmodule

// tks6_o0w6_0c38m1c3em2c3cm24m2cm34m3co0w0_4mcm14m1co0w0 TeakS (0+:6) [([Imp 0 56,Imp 1 62,Imp 2 60,Im
//   p 36 0,Imp 44 0,Imp 52 0,Imp 60 0],0),([Imp 4 0,Imp 12 0,Imp 20 0,Imp 28 0],0)] [One 6,Many [0,0]]
module tks6_o0w6_0c38m1c3em2c3cm24m2cm34m3co0w0_4mcm14m1co0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input [5:0] i_0r0;
  input [5:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire [6:0] match0_0;
  wire [2:0] simp71_0;
  wire [1:0] simp111_0;
  wire [1:0] simp121_0;
  wire [1:0] simp131_0;
  wire [1:0] simp141_0;
  wire [3:0] match1_0;
  wire [1:0] simp161_0;
  wire [1:0] simp171_0;
  wire [1:0] simp181_0;
  wire [1:0] simp191_0;
  wire [1:0] simp201_0;
  wire [5:0] comp_0;
  wire [1:0] simp301_0;
  NOR3 I0 (simp71_0[0:0], match0_0[0:0], match0_0[1:1], match0_0[2:2]);
  NOR3 I1 (simp71_0[1:1], match0_0[3:3], match0_0[4:4], match0_0[5:5]);
  INV I2 (simp71_0[2:2], match0_0[6:6]);
  NAND3 I3 (sel_0, simp71_0[0:0], simp71_0[1:1], simp71_0[2:2]);
  C3 I4 (match0_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I5 (match0_0[1:1], i_0r1[0:0]);
  C2 I6 (match0_0[2:2], i_0r0[0:0], i_0r1[1:1]);
  C3 I7 (simp111_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I8 (simp111_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I9 (match0_0[3:3], simp111_0[0:0], simp111_0[1:1]);
  C3 I10 (simp121_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I11 (simp121_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I12 (match0_0[4:4], simp121_0[0:0], simp121_0[1:1]);
  C3 I13 (simp131_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I14 (simp131_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I15 (match0_0[5:5], simp131_0[0:0], simp131_0[1:1]);
  C3 I16 (simp141_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I17 (simp141_0[1:1], i_0r1[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I18 (match0_0[6:6], simp141_0[0:0], simp141_0[1:1]);
  NOR3 I19 (simp161_0[0:0], match1_0[0:0], match1_0[1:1], match1_0[2:2]);
  INV I20 (simp161_0[1:1], match1_0[3:3]);
  NAND2 I21 (sel_1, simp161_0[0:0], simp161_0[1:1]);
  C3 I22 (simp171_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I23 (simp171_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I24 (match1_0[0:0], simp171_0[0:0], simp171_0[1:1]);
  C3 I25 (simp181_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I26 (simp181_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I27 (match1_0[1:1], simp181_0[0:0], simp181_0[1:1]);
  C3 I28 (simp191_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I29 (simp191_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I30 (match1_0[2:2], simp191_0[0:0], simp191_0[1:1]);
  C3 I31 (simp201_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I32 (simp201_0[1:1], i_0r1[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I33 (match1_0[3:3], simp201_0[0:0], simp201_0[1:1]);
  C2 I34 (gsel_0, sel_0, icomplete_0);
  C2 I35 (gsel_1, sel_1, icomplete_0);
  OR2 I36 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I37 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I38 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I39 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I40 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I41 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  C3 I42 (simp301_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I43 (simp301_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C2 I44 (icomplete_0, simp301_0[0:0], simp301_0[1:1]);
  BUFF I45 (o_0r, gsel_0);
  BUFF I46 (o_1r, gsel_1);
  OR2 I47 (oack_0, o_0a, o_1a);
  C2 I48 (i_0a, oack_0, icomplete_0);
endmodule

// tks6_o0w6_0c30m1c3em2c3cm24m28m2cm34m38m3co0w0_4m14o0w0_8m18o0w0_cm1co0w0 TeakS (0+:6) [([Imp 0 48,I
//   mp 1 62,Imp 2 60,Imp 36 0,Imp 40 0,Imp 44 0,Imp 52 0,Imp 56 0,Imp 60 0],0),([Imp 4 0,Imp 20 0],0),([
//   Imp 8 0,Imp 24 0],0),([Imp 12 0,Imp 28 0],0)] [One 6,Many [0,0,0,0]]
module tks6_o0w6_0c30m1c3em2c3cm24m28m2cm34m38m3co0w0_4m14o0w0_8m18o0w0_cm1co0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, reset);
  input [5:0] i_0r0;
  input [5:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire oack_0;
  wire [8:0] match0_0;
  wire [2:0] simp111_0;
  wire [1:0] simp121_0;
  wire [1:0] simp151_0;
  wire [1:0] simp161_0;
  wire [1:0] simp171_0;
  wire [1:0] simp181_0;
  wire [1:0] simp191_0;
  wire [1:0] simp201_0;
  wire [1:0] match1_0;
  wire [1:0] simp231_0;
  wire [1:0] simp241_0;
  wire [1:0] match2_0;
  wire [1:0] simp271_0;
  wire [1:0] simp281_0;
  wire [1:0] match3_0;
  wire [1:0] simp311_0;
  wire [1:0] simp321_0;
  wire [5:0] comp_0;
  wire [1:0] simp441_0;
  wire [1:0] simp491_0;
  NOR3 I0 (simp111_0[0:0], match0_0[0:0], match0_0[1:1], match0_0[2:2]);
  NOR3 I1 (simp111_0[1:1], match0_0[3:3], match0_0[4:4], match0_0[5:5]);
  NOR3 I2 (simp111_0[2:2], match0_0[6:6], match0_0[7:7], match0_0[8:8]);
  NAND3 I3 (sel_0, simp111_0[0:0], simp111_0[1:1], simp111_0[2:2]);
  C3 I4 (simp121_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I5 (simp121_0[1:1], i_0r0[3:3]);
  C2 I6 (match0_0[0:0], simp121_0[0:0], simp121_0[1:1]);
  BUFF I7 (match0_0[1:1], i_0r1[0:0]);
  C2 I8 (match0_0[2:2], i_0r0[0:0], i_0r1[1:1]);
  C3 I9 (simp151_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I10 (simp151_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I11 (match0_0[3:3], simp151_0[0:0], simp151_0[1:1]);
  C3 I12 (simp161_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I13 (simp161_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I14 (match0_0[4:4], simp161_0[0:0], simp161_0[1:1]);
  C3 I15 (simp171_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I16 (simp171_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I17 (match0_0[5:5], simp171_0[0:0], simp171_0[1:1]);
  C3 I18 (simp181_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I19 (simp181_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I20 (match0_0[6:6], simp181_0[0:0], simp181_0[1:1]);
  C3 I21 (simp191_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I22 (simp191_0[1:1], i_0r1[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I23 (match0_0[7:7], simp191_0[0:0], simp191_0[1:1]);
  C3 I24 (simp201_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I25 (simp201_0[1:1], i_0r1[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I26 (match0_0[8:8], simp201_0[0:0], simp201_0[1:1]);
  OR2 I27 (sel_1, match1_0[0:0], match1_0[1:1]);
  C3 I28 (simp231_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I29 (simp231_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I30 (match1_0[0:0], simp231_0[0:0], simp231_0[1:1]);
  C3 I31 (simp241_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I32 (simp241_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I33 (match1_0[1:1], simp241_0[0:0], simp241_0[1:1]);
  OR2 I34 (sel_2, match2_0[0:0], match2_0[1:1]);
  C3 I35 (simp271_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I36 (simp271_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I37 (match2_0[0:0], simp271_0[0:0], simp271_0[1:1]);
  C3 I38 (simp281_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I39 (simp281_0[1:1], i_0r1[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I40 (match2_0[1:1], simp281_0[0:0], simp281_0[1:1]);
  OR2 I41 (sel_3, match3_0[0:0], match3_0[1:1]);
  C3 I42 (simp311_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I43 (simp311_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I44 (match3_0[0:0], simp311_0[0:0], simp311_0[1:1]);
  C3 I45 (simp321_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I46 (simp321_0[1:1], i_0r1[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I47 (match3_0[1:1], simp321_0[0:0], simp321_0[1:1]);
  C2 I48 (gsel_0, sel_0, icomplete_0);
  C2 I49 (gsel_1, sel_1, icomplete_0);
  C2 I50 (gsel_2, sel_2, icomplete_0);
  C2 I51 (gsel_3, sel_3, icomplete_0);
  OR2 I52 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I53 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I54 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I55 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I56 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I57 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  C3 I58 (simp441_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I59 (simp441_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C2 I60 (icomplete_0, simp441_0[0:0], simp441_0[1:1]);
  BUFF I61 (o_0r, gsel_0);
  BUFF I62 (o_1r, gsel_1);
  BUFF I63 (o_2r, gsel_2);
  BUFF I64 (o_3r, gsel_3);
  NOR3 I65 (simp491_0[0:0], o_0a, o_1a, o_2a);
  INV I66 (simp491_0[1:1], o_3a);
  NAND2 I67 (oack_0, simp491_0[0:0], simp491_0[1:1]);
  C2 I68 (i_0a, oack_0, icomplete_0);
endmodule

// tkj33m1_32 TeakJ [Many [1,32],One 33]
module tkj33m1_32 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [32:0] joinf_0;
  wire [32:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0);
  BUFF I1 (joinf_0[1:1], i_1r0[0:0]);
  BUFF I2 (joinf_0[2:2], i_1r0[1:1]);
  BUFF I3 (joinf_0[3:3], i_1r0[2:2]);
  BUFF I4 (joinf_0[4:4], i_1r0[3:3]);
  BUFF I5 (joinf_0[5:5], i_1r0[4:4]);
  BUFF I6 (joinf_0[6:6], i_1r0[5:5]);
  BUFF I7 (joinf_0[7:7], i_1r0[6:6]);
  BUFF I8 (joinf_0[8:8], i_1r0[7:7]);
  BUFF I9 (joinf_0[9:9], i_1r0[8:8]);
  BUFF I10 (joinf_0[10:10], i_1r0[9:9]);
  BUFF I11 (joinf_0[11:11], i_1r0[10:10]);
  BUFF I12 (joinf_0[12:12], i_1r0[11:11]);
  BUFF I13 (joinf_0[13:13], i_1r0[12:12]);
  BUFF I14 (joinf_0[14:14], i_1r0[13:13]);
  BUFF I15 (joinf_0[15:15], i_1r0[14:14]);
  BUFF I16 (joinf_0[16:16], i_1r0[15:15]);
  BUFF I17 (joinf_0[17:17], i_1r0[16:16]);
  BUFF I18 (joinf_0[18:18], i_1r0[17:17]);
  BUFF I19 (joinf_0[19:19], i_1r0[18:18]);
  BUFF I20 (joinf_0[20:20], i_1r0[19:19]);
  BUFF I21 (joinf_0[21:21], i_1r0[20:20]);
  BUFF I22 (joinf_0[22:22], i_1r0[21:21]);
  BUFF I23 (joinf_0[23:23], i_1r0[22:22]);
  BUFF I24 (joinf_0[24:24], i_1r0[23:23]);
  BUFF I25 (joinf_0[25:25], i_1r0[24:24]);
  BUFF I26 (joinf_0[26:26], i_1r0[25:25]);
  BUFF I27 (joinf_0[27:27], i_1r0[26:26]);
  BUFF I28 (joinf_0[28:28], i_1r0[27:27]);
  BUFF I29 (joinf_0[29:29], i_1r0[28:28]);
  BUFF I30 (joinf_0[30:30], i_1r0[29:29]);
  BUFF I31 (joinf_0[31:31], i_1r0[30:30]);
  BUFF I32 (joinf_0[32:32], i_1r0[31:31]);
  BUFF I33 (joint_0[0:0], i_0r1);
  BUFF I34 (joint_0[1:1], i_1r1[0:0]);
  BUFF I35 (joint_0[2:2], i_1r1[1:1]);
  BUFF I36 (joint_0[3:3], i_1r1[2:2]);
  BUFF I37 (joint_0[4:4], i_1r1[3:3]);
  BUFF I38 (joint_0[5:5], i_1r1[4:4]);
  BUFF I39 (joint_0[6:6], i_1r1[5:5]);
  BUFF I40 (joint_0[7:7], i_1r1[6:6]);
  BUFF I41 (joint_0[8:8], i_1r1[7:7]);
  BUFF I42 (joint_0[9:9], i_1r1[8:8]);
  BUFF I43 (joint_0[10:10], i_1r1[9:9]);
  BUFF I44 (joint_0[11:11], i_1r1[10:10]);
  BUFF I45 (joint_0[12:12], i_1r1[11:11]);
  BUFF I46 (joint_0[13:13], i_1r1[12:12]);
  BUFF I47 (joint_0[14:14], i_1r1[13:13]);
  BUFF I48 (joint_0[15:15], i_1r1[14:14]);
  BUFF I49 (joint_0[16:16], i_1r1[15:15]);
  BUFF I50 (joint_0[17:17], i_1r1[16:16]);
  BUFF I51 (joint_0[18:18], i_1r1[17:17]);
  BUFF I52 (joint_0[19:19], i_1r1[18:18]);
  BUFF I53 (joint_0[20:20], i_1r1[19:19]);
  BUFF I54 (joint_0[21:21], i_1r1[20:20]);
  BUFF I55 (joint_0[22:22], i_1r1[21:21]);
  BUFF I56 (joint_0[23:23], i_1r1[22:22]);
  BUFF I57 (joint_0[24:24], i_1r1[23:23]);
  BUFF I58 (joint_0[25:25], i_1r1[24:24]);
  BUFF I59 (joint_0[26:26], i_1r1[25:25]);
  BUFF I60 (joint_0[27:27], i_1r1[26:26]);
  BUFF I61 (joint_0[28:28], i_1r1[27:27]);
  BUFF I62 (joint_0[29:29], i_1r1[28:28]);
  BUFF I63 (joint_0[30:30], i_1r1[29:29]);
  BUFF I64 (joint_0[31:31], i_1r1[30:30]);
  BUFF I65 (joint_0[32:32], i_1r1[31:31]);
  OR2 I66 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I67 (icomplete_0, dcomplete_0);
  C2 I68 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I69 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I70 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I71 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I72 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I73 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I74 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I75 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I76 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I77 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I78 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I79 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I80 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I81 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I82 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I83 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I84 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I85 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I86 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I87 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I88 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I89 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I90 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I91 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I92 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I93 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I94 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I95 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I96 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I97 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I98 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I99 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I100 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I101 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I102 (o_0r1[1:1], joint_0[1:1]);
  BUFF I103 (o_0r1[2:2], joint_0[2:2]);
  BUFF I104 (o_0r1[3:3], joint_0[3:3]);
  BUFF I105 (o_0r1[4:4], joint_0[4:4]);
  BUFF I106 (o_0r1[5:5], joint_0[5:5]);
  BUFF I107 (o_0r1[6:6], joint_0[6:6]);
  BUFF I108 (o_0r1[7:7], joint_0[7:7]);
  BUFF I109 (o_0r1[8:8], joint_0[8:8]);
  BUFF I110 (o_0r1[9:9], joint_0[9:9]);
  BUFF I111 (o_0r1[10:10], joint_0[10:10]);
  BUFF I112 (o_0r1[11:11], joint_0[11:11]);
  BUFF I113 (o_0r1[12:12], joint_0[12:12]);
  BUFF I114 (o_0r1[13:13], joint_0[13:13]);
  BUFF I115 (o_0r1[14:14], joint_0[14:14]);
  BUFF I116 (o_0r1[15:15], joint_0[15:15]);
  BUFF I117 (o_0r1[16:16], joint_0[16:16]);
  BUFF I118 (o_0r1[17:17], joint_0[17:17]);
  BUFF I119 (o_0r1[18:18], joint_0[18:18]);
  BUFF I120 (o_0r1[19:19], joint_0[19:19]);
  BUFF I121 (o_0r1[20:20], joint_0[20:20]);
  BUFF I122 (o_0r1[21:21], joint_0[21:21]);
  BUFF I123 (o_0r1[22:22], joint_0[22:22]);
  BUFF I124 (o_0r1[23:23], joint_0[23:23]);
  BUFF I125 (o_0r1[24:24], joint_0[24:24]);
  BUFF I126 (o_0r1[25:25], joint_0[25:25]);
  BUFF I127 (o_0r1[26:26], joint_0[26:26]);
  BUFF I128 (o_0r1[27:27], joint_0[27:27]);
  BUFF I129 (o_0r1[28:28], joint_0[28:28]);
  BUFF I130 (o_0r1[29:29], joint_0[29:29]);
  BUFF I131 (o_0r1[30:30], joint_0[30:30]);
  BUFF I132 (o_0r1[31:31], joint_0[31:31]);
  BUFF I133 (o_0r1[32:32], joint_0[32:32]);
  BUFF I134 (i_0a, o_0a);
  BUFF I135 (i_1a, o_0a);
endmodule

// tkj66m33_33 TeakJ [Many [33,33],One 66]
module tkj66m33_33 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [32:0] i_0r0;
  input [32:0] i_0r1;
  output i_0a;
  input [32:0] i_1r0;
  input [32:0] i_1r1;
  output i_1a;
  output [65:0] o_0r0;
  output [65:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [65:0] joinf_0;
  wire [65:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joinf_0[32:32], i_0r0[32:32]);
  BUFF I33 (joinf_0[33:33], i_1r0[0:0]);
  BUFF I34 (joinf_0[34:34], i_1r0[1:1]);
  BUFF I35 (joinf_0[35:35], i_1r0[2:2]);
  BUFF I36 (joinf_0[36:36], i_1r0[3:3]);
  BUFF I37 (joinf_0[37:37], i_1r0[4:4]);
  BUFF I38 (joinf_0[38:38], i_1r0[5:5]);
  BUFF I39 (joinf_0[39:39], i_1r0[6:6]);
  BUFF I40 (joinf_0[40:40], i_1r0[7:7]);
  BUFF I41 (joinf_0[41:41], i_1r0[8:8]);
  BUFF I42 (joinf_0[42:42], i_1r0[9:9]);
  BUFF I43 (joinf_0[43:43], i_1r0[10:10]);
  BUFF I44 (joinf_0[44:44], i_1r0[11:11]);
  BUFF I45 (joinf_0[45:45], i_1r0[12:12]);
  BUFF I46 (joinf_0[46:46], i_1r0[13:13]);
  BUFF I47 (joinf_0[47:47], i_1r0[14:14]);
  BUFF I48 (joinf_0[48:48], i_1r0[15:15]);
  BUFF I49 (joinf_0[49:49], i_1r0[16:16]);
  BUFF I50 (joinf_0[50:50], i_1r0[17:17]);
  BUFF I51 (joinf_0[51:51], i_1r0[18:18]);
  BUFF I52 (joinf_0[52:52], i_1r0[19:19]);
  BUFF I53 (joinf_0[53:53], i_1r0[20:20]);
  BUFF I54 (joinf_0[54:54], i_1r0[21:21]);
  BUFF I55 (joinf_0[55:55], i_1r0[22:22]);
  BUFF I56 (joinf_0[56:56], i_1r0[23:23]);
  BUFF I57 (joinf_0[57:57], i_1r0[24:24]);
  BUFF I58 (joinf_0[58:58], i_1r0[25:25]);
  BUFF I59 (joinf_0[59:59], i_1r0[26:26]);
  BUFF I60 (joinf_0[60:60], i_1r0[27:27]);
  BUFF I61 (joinf_0[61:61], i_1r0[28:28]);
  BUFF I62 (joinf_0[62:62], i_1r0[29:29]);
  BUFF I63 (joinf_0[63:63], i_1r0[30:30]);
  BUFF I64 (joinf_0[64:64], i_1r0[31:31]);
  BUFF I65 (joinf_0[65:65], i_1r0[32:32]);
  BUFF I66 (joint_0[0:0], i_0r1[0:0]);
  BUFF I67 (joint_0[1:1], i_0r1[1:1]);
  BUFF I68 (joint_0[2:2], i_0r1[2:2]);
  BUFF I69 (joint_0[3:3], i_0r1[3:3]);
  BUFF I70 (joint_0[4:4], i_0r1[4:4]);
  BUFF I71 (joint_0[5:5], i_0r1[5:5]);
  BUFF I72 (joint_0[6:6], i_0r1[6:6]);
  BUFF I73 (joint_0[7:7], i_0r1[7:7]);
  BUFF I74 (joint_0[8:8], i_0r1[8:8]);
  BUFF I75 (joint_0[9:9], i_0r1[9:9]);
  BUFF I76 (joint_0[10:10], i_0r1[10:10]);
  BUFF I77 (joint_0[11:11], i_0r1[11:11]);
  BUFF I78 (joint_0[12:12], i_0r1[12:12]);
  BUFF I79 (joint_0[13:13], i_0r1[13:13]);
  BUFF I80 (joint_0[14:14], i_0r1[14:14]);
  BUFF I81 (joint_0[15:15], i_0r1[15:15]);
  BUFF I82 (joint_0[16:16], i_0r1[16:16]);
  BUFF I83 (joint_0[17:17], i_0r1[17:17]);
  BUFF I84 (joint_0[18:18], i_0r1[18:18]);
  BUFF I85 (joint_0[19:19], i_0r1[19:19]);
  BUFF I86 (joint_0[20:20], i_0r1[20:20]);
  BUFF I87 (joint_0[21:21], i_0r1[21:21]);
  BUFF I88 (joint_0[22:22], i_0r1[22:22]);
  BUFF I89 (joint_0[23:23], i_0r1[23:23]);
  BUFF I90 (joint_0[24:24], i_0r1[24:24]);
  BUFF I91 (joint_0[25:25], i_0r1[25:25]);
  BUFF I92 (joint_0[26:26], i_0r1[26:26]);
  BUFF I93 (joint_0[27:27], i_0r1[27:27]);
  BUFF I94 (joint_0[28:28], i_0r1[28:28]);
  BUFF I95 (joint_0[29:29], i_0r1[29:29]);
  BUFF I96 (joint_0[30:30], i_0r1[30:30]);
  BUFF I97 (joint_0[31:31], i_0r1[31:31]);
  BUFF I98 (joint_0[32:32], i_0r1[32:32]);
  BUFF I99 (joint_0[33:33], i_1r1[0:0]);
  BUFF I100 (joint_0[34:34], i_1r1[1:1]);
  BUFF I101 (joint_0[35:35], i_1r1[2:2]);
  BUFF I102 (joint_0[36:36], i_1r1[3:3]);
  BUFF I103 (joint_0[37:37], i_1r1[4:4]);
  BUFF I104 (joint_0[38:38], i_1r1[5:5]);
  BUFF I105 (joint_0[39:39], i_1r1[6:6]);
  BUFF I106 (joint_0[40:40], i_1r1[7:7]);
  BUFF I107 (joint_0[41:41], i_1r1[8:8]);
  BUFF I108 (joint_0[42:42], i_1r1[9:9]);
  BUFF I109 (joint_0[43:43], i_1r1[10:10]);
  BUFF I110 (joint_0[44:44], i_1r1[11:11]);
  BUFF I111 (joint_0[45:45], i_1r1[12:12]);
  BUFF I112 (joint_0[46:46], i_1r1[13:13]);
  BUFF I113 (joint_0[47:47], i_1r1[14:14]);
  BUFF I114 (joint_0[48:48], i_1r1[15:15]);
  BUFF I115 (joint_0[49:49], i_1r1[16:16]);
  BUFF I116 (joint_0[50:50], i_1r1[17:17]);
  BUFF I117 (joint_0[51:51], i_1r1[18:18]);
  BUFF I118 (joint_0[52:52], i_1r1[19:19]);
  BUFF I119 (joint_0[53:53], i_1r1[20:20]);
  BUFF I120 (joint_0[54:54], i_1r1[21:21]);
  BUFF I121 (joint_0[55:55], i_1r1[22:22]);
  BUFF I122 (joint_0[56:56], i_1r1[23:23]);
  BUFF I123 (joint_0[57:57], i_1r1[24:24]);
  BUFF I124 (joint_0[58:58], i_1r1[25:25]);
  BUFF I125 (joint_0[59:59], i_1r1[26:26]);
  BUFF I126 (joint_0[60:60], i_1r1[27:27]);
  BUFF I127 (joint_0[61:61], i_1r1[28:28]);
  BUFF I128 (joint_0[62:62], i_1r1[29:29]);
  BUFF I129 (joint_0[63:63], i_1r1[30:30]);
  BUFF I130 (joint_0[64:64], i_1r1[31:31]);
  BUFF I131 (joint_0[65:65], i_1r1[32:32]);
  OR2 I132 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I133 (icomplete_0, dcomplete_0);
  C2 I134 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I135 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I136 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I137 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I138 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I139 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I140 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I141 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I142 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I143 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I144 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I145 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I146 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I147 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I148 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I149 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I150 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I151 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I152 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I153 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I154 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I155 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I156 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I157 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I158 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I159 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I160 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I161 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I162 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I163 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I164 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I165 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I166 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I167 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I168 (o_0r0[33:33], joinf_0[33:33]);
  BUFF I169 (o_0r0[34:34], joinf_0[34:34]);
  BUFF I170 (o_0r0[35:35], joinf_0[35:35]);
  BUFF I171 (o_0r0[36:36], joinf_0[36:36]);
  BUFF I172 (o_0r0[37:37], joinf_0[37:37]);
  BUFF I173 (o_0r0[38:38], joinf_0[38:38]);
  BUFF I174 (o_0r0[39:39], joinf_0[39:39]);
  BUFF I175 (o_0r0[40:40], joinf_0[40:40]);
  BUFF I176 (o_0r0[41:41], joinf_0[41:41]);
  BUFF I177 (o_0r0[42:42], joinf_0[42:42]);
  BUFF I178 (o_0r0[43:43], joinf_0[43:43]);
  BUFF I179 (o_0r0[44:44], joinf_0[44:44]);
  BUFF I180 (o_0r0[45:45], joinf_0[45:45]);
  BUFF I181 (o_0r0[46:46], joinf_0[46:46]);
  BUFF I182 (o_0r0[47:47], joinf_0[47:47]);
  BUFF I183 (o_0r0[48:48], joinf_0[48:48]);
  BUFF I184 (o_0r0[49:49], joinf_0[49:49]);
  BUFF I185 (o_0r0[50:50], joinf_0[50:50]);
  BUFF I186 (o_0r0[51:51], joinf_0[51:51]);
  BUFF I187 (o_0r0[52:52], joinf_0[52:52]);
  BUFF I188 (o_0r0[53:53], joinf_0[53:53]);
  BUFF I189 (o_0r0[54:54], joinf_0[54:54]);
  BUFF I190 (o_0r0[55:55], joinf_0[55:55]);
  BUFF I191 (o_0r0[56:56], joinf_0[56:56]);
  BUFF I192 (o_0r0[57:57], joinf_0[57:57]);
  BUFF I193 (o_0r0[58:58], joinf_0[58:58]);
  BUFF I194 (o_0r0[59:59], joinf_0[59:59]);
  BUFF I195 (o_0r0[60:60], joinf_0[60:60]);
  BUFF I196 (o_0r0[61:61], joinf_0[61:61]);
  BUFF I197 (o_0r0[62:62], joinf_0[62:62]);
  BUFF I198 (o_0r0[63:63], joinf_0[63:63]);
  BUFF I199 (o_0r0[64:64], joinf_0[64:64]);
  BUFF I200 (o_0r0[65:65], joinf_0[65:65]);
  BUFF I201 (o_0r1[1:1], joint_0[1:1]);
  BUFF I202 (o_0r1[2:2], joint_0[2:2]);
  BUFF I203 (o_0r1[3:3], joint_0[3:3]);
  BUFF I204 (o_0r1[4:4], joint_0[4:4]);
  BUFF I205 (o_0r1[5:5], joint_0[5:5]);
  BUFF I206 (o_0r1[6:6], joint_0[6:6]);
  BUFF I207 (o_0r1[7:7], joint_0[7:7]);
  BUFF I208 (o_0r1[8:8], joint_0[8:8]);
  BUFF I209 (o_0r1[9:9], joint_0[9:9]);
  BUFF I210 (o_0r1[10:10], joint_0[10:10]);
  BUFF I211 (o_0r1[11:11], joint_0[11:11]);
  BUFF I212 (o_0r1[12:12], joint_0[12:12]);
  BUFF I213 (o_0r1[13:13], joint_0[13:13]);
  BUFF I214 (o_0r1[14:14], joint_0[14:14]);
  BUFF I215 (o_0r1[15:15], joint_0[15:15]);
  BUFF I216 (o_0r1[16:16], joint_0[16:16]);
  BUFF I217 (o_0r1[17:17], joint_0[17:17]);
  BUFF I218 (o_0r1[18:18], joint_0[18:18]);
  BUFF I219 (o_0r1[19:19], joint_0[19:19]);
  BUFF I220 (o_0r1[20:20], joint_0[20:20]);
  BUFF I221 (o_0r1[21:21], joint_0[21:21]);
  BUFF I222 (o_0r1[22:22], joint_0[22:22]);
  BUFF I223 (o_0r1[23:23], joint_0[23:23]);
  BUFF I224 (o_0r1[24:24], joint_0[24:24]);
  BUFF I225 (o_0r1[25:25], joint_0[25:25]);
  BUFF I226 (o_0r1[26:26], joint_0[26:26]);
  BUFF I227 (o_0r1[27:27], joint_0[27:27]);
  BUFF I228 (o_0r1[28:28], joint_0[28:28]);
  BUFF I229 (o_0r1[29:29], joint_0[29:29]);
  BUFF I230 (o_0r1[30:30], joint_0[30:30]);
  BUFF I231 (o_0r1[31:31], joint_0[31:31]);
  BUFF I232 (o_0r1[32:32], joint_0[32:32]);
  BUFF I233 (o_0r1[33:33], joint_0[33:33]);
  BUFF I234 (o_0r1[34:34], joint_0[34:34]);
  BUFF I235 (o_0r1[35:35], joint_0[35:35]);
  BUFF I236 (o_0r1[36:36], joint_0[36:36]);
  BUFF I237 (o_0r1[37:37], joint_0[37:37]);
  BUFF I238 (o_0r1[38:38], joint_0[38:38]);
  BUFF I239 (o_0r1[39:39], joint_0[39:39]);
  BUFF I240 (o_0r1[40:40], joint_0[40:40]);
  BUFF I241 (o_0r1[41:41], joint_0[41:41]);
  BUFF I242 (o_0r1[42:42], joint_0[42:42]);
  BUFF I243 (o_0r1[43:43], joint_0[43:43]);
  BUFF I244 (o_0r1[44:44], joint_0[44:44]);
  BUFF I245 (o_0r1[45:45], joint_0[45:45]);
  BUFF I246 (o_0r1[46:46], joint_0[46:46]);
  BUFF I247 (o_0r1[47:47], joint_0[47:47]);
  BUFF I248 (o_0r1[48:48], joint_0[48:48]);
  BUFF I249 (o_0r1[49:49], joint_0[49:49]);
  BUFF I250 (o_0r1[50:50], joint_0[50:50]);
  BUFF I251 (o_0r1[51:51], joint_0[51:51]);
  BUFF I252 (o_0r1[52:52], joint_0[52:52]);
  BUFF I253 (o_0r1[53:53], joint_0[53:53]);
  BUFF I254 (o_0r1[54:54], joint_0[54:54]);
  BUFF I255 (o_0r1[55:55], joint_0[55:55]);
  BUFF I256 (o_0r1[56:56], joint_0[56:56]);
  BUFF I257 (o_0r1[57:57], joint_0[57:57]);
  BUFF I258 (o_0r1[58:58], joint_0[58:58]);
  BUFF I259 (o_0r1[59:59], joint_0[59:59]);
  BUFF I260 (o_0r1[60:60], joint_0[60:60]);
  BUFF I261 (o_0r1[61:61], joint_0[61:61]);
  BUFF I262 (o_0r1[62:62], joint_0[62:62]);
  BUFF I263 (o_0r1[63:63], joint_0[63:63]);
  BUFF I264 (o_0r1[64:64], joint_0[64:64]);
  BUFF I265 (o_0r1[65:65], joint_0[65:65]);
  BUFF I266 (i_0a, o_0a);
  BUFF I267 (i_1a, o_0a);
endmodule

// tko66m34_1api0w33b_2api33w33b_3nm1b0_4apt1o0w33bt3o0w1b_5nm1b0_6apt2o0w33bt5o0w1b_7addt4o0w34bt6o0w3
//   4b TeakO [
//     (1,TeakOAppend 1 [(0,0+:33)]),
//     (2,TeakOAppend 1 [(0,33+:33)]),
//     (3,TeakOConstant 1 0),
//     (4,TeakOAppend 1 [(1,0+:33),(3,0+:1)]),
//     (5,TeakOConstant 1 0),
//     (6,TeakOAppend 1 [(2,0+:33),(5,0+:1)]),
//     (7,TeakOp TeakOpAdd [(4,0+:34),(6,0+:34)])] [One 66,One 34]
module tko66m34_1api0w33b_2api33w33b_3nm1b0_4apt1o0w33bt3o0w1b_5nm1b0_6apt2o0w33bt5o0w1b_7addt4o0w34bt6o0w34b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [65:0] i_0r0;
  input [65:0] i_0r1;
  output i_0a;
  output [33:0] o_0r0;
  output [33:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [65:0] gocomp_0;
  wire [21:0] simp681_0;
  wire [7:0] simp682_0;
  wire [2:0] simp683_0;
  wire [32:0] termf_1;
  wire [32:0] termf_2;
  wire termf_3;
  wire [33:0] termf_4;
  wire termf_5;
  wire [33:0] termf_6;
  wire [32:0] termt_1;
  wire [32:0] termt_2;
  wire termt_3;
  wire [33:0] termt_4;
  wire termt_5;
  wire [33:0] termt_6;
  wire [33:0] cf7__0;
  wire [33:0] ct7__0;
  wire [3:0] ha7__0;
  wire [7:0] fa7_1min_0;
  wire [1:0] simp3751_0;
  wire [1:0] simp3761_0;
  wire [7:0] fa7_2min_0;
  wire [1:0] simp3881_0;
  wire [1:0] simp3891_0;
  wire [7:0] fa7_3min_0;
  wire [1:0] simp4011_0;
  wire [1:0] simp4021_0;
  wire [7:0] fa7_4min_0;
  wire [1:0] simp4141_0;
  wire [1:0] simp4151_0;
  wire [7:0] fa7_5min_0;
  wire [1:0] simp4271_0;
  wire [1:0] simp4281_0;
  wire [7:0] fa7_6min_0;
  wire [1:0] simp4401_0;
  wire [1:0] simp4411_0;
  wire [7:0] fa7_7min_0;
  wire [1:0] simp4531_0;
  wire [1:0] simp4541_0;
  wire [7:0] fa7_8min_0;
  wire [1:0] simp4661_0;
  wire [1:0] simp4671_0;
  wire [7:0] fa7_9min_0;
  wire [1:0] simp4791_0;
  wire [1:0] simp4801_0;
  wire [7:0] fa7_10min_0;
  wire [1:0] simp4921_0;
  wire [1:0] simp4931_0;
  wire [7:0] fa7_11min_0;
  wire [1:0] simp5051_0;
  wire [1:0] simp5061_0;
  wire [7:0] fa7_12min_0;
  wire [1:0] simp5181_0;
  wire [1:0] simp5191_0;
  wire [7:0] fa7_13min_0;
  wire [1:0] simp5311_0;
  wire [1:0] simp5321_0;
  wire [7:0] fa7_14min_0;
  wire [1:0] simp5441_0;
  wire [1:0] simp5451_0;
  wire [7:0] fa7_15min_0;
  wire [1:0] simp5571_0;
  wire [1:0] simp5581_0;
  wire [7:0] fa7_16min_0;
  wire [1:0] simp5701_0;
  wire [1:0] simp5711_0;
  wire [7:0] fa7_17min_0;
  wire [1:0] simp5831_0;
  wire [1:0] simp5841_0;
  wire [7:0] fa7_18min_0;
  wire [1:0] simp5961_0;
  wire [1:0] simp5971_0;
  wire [7:0] fa7_19min_0;
  wire [1:0] simp6091_0;
  wire [1:0] simp6101_0;
  wire [7:0] fa7_20min_0;
  wire [1:0] simp6221_0;
  wire [1:0] simp6231_0;
  wire [7:0] fa7_21min_0;
  wire [1:0] simp6351_0;
  wire [1:0] simp6361_0;
  wire [7:0] fa7_22min_0;
  wire [1:0] simp6481_0;
  wire [1:0] simp6491_0;
  wire [7:0] fa7_23min_0;
  wire [1:0] simp6611_0;
  wire [1:0] simp6621_0;
  wire [7:0] fa7_24min_0;
  wire [1:0] simp6741_0;
  wire [1:0] simp6751_0;
  wire [7:0] fa7_25min_0;
  wire [1:0] simp6871_0;
  wire [1:0] simp6881_0;
  wire [7:0] fa7_26min_0;
  wire [1:0] simp7001_0;
  wire [1:0] simp7011_0;
  wire [7:0] fa7_27min_0;
  wire [1:0] simp7131_0;
  wire [1:0] simp7141_0;
  wire [7:0] fa7_28min_0;
  wire [1:0] simp7261_0;
  wire [1:0] simp7271_0;
  wire [7:0] fa7_29min_0;
  wire [1:0] simp7391_0;
  wire [1:0] simp7401_0;
  wire [7:0] fa7_30min_0;
  wire [1:0] simp7521_0;
  wire [1:0] simp7531_0;
  wire [7:0] fa7_31min_0;
  wire [1:0] simp7651_0;
  wire [1:0] simp7661_0;
  wire [7:0] fa7_32min_0;
  wire [1:0] simp7781_0;
  wire [1:0] simp7791_0;
  wire [7:0] fa7_33min_0;
  wire [1:0] simp7911_0;
  wire [1:0] simp7921_0;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I30 (gocomp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I31 (gocomp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I32 (gocomp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  OR2 I33 (gocomp_0[33:33], i_0r0[33:33], i_0r1[33:33]);
  OR2 I34 (gocomp_0[34:34], i_0r0[34:34], i_0r1[34:34]);
  OR2 I35 (gocomp_0[35:35], i_0r0[35:35], i_0r1[35:35]);
  OR2 I36 (gocomp_0[36:36], i_0r0[36:36], i_0r1[36:36]);
  OR2 I37 (gocomp_0[37:37], i_0r0[37:37], i_0r1[37:37]);
  OR2 I38 (gocomp_0[38:38], i_0r0[38:38], i_0r1[38:38]);
  OR2 I39 (gocomp_0[39:39], i_0r0[39:39], i_0r1[39:39]);
  OR2 I40 (gocomp_0[40:40], i_0r0[40:40], i_0r1[40:40]);
  OR2 I41 (gocomp_0[41:41], i_0r0[41:41], i_0r1[41:41]);
  OR2 I42 (gocomp_0[42:42], i_0r0[42:42], i_0r1[42:42]);
  OR2 I43 (gocomp_0[43:43], i_0r0[43:43], i_0r1[43:43]);
  OR2 I44 (gocomp_0[44:44], i_0r0[44:44], i_0r1[44:44]);
  OR2 I45 (gocomp_0[45:45], i_0r0[45:45], i_0r1[45:45]);
  OR2 I46 (gocomp_0[46:46], i_0r0[46:46], i_0r1[46:46]);
  OR2 I47 (gocomp_0[47:47], i_0r0[47:47], i_0r1[47:47]);
  OR2 I48 (gocomp_0[48:48], i_0r0[48:48], i_0r1[48:48]);
  OR2 I49 (gocomp_0[49:49], i_0r0[49:49], i_0r1[49:49]);
  OR2 I50 (gocomp_0[50:50], i_0r0[50:50], i_0r1[50:50]);
  OR2 I51 (gocomp_0[51:51], i_0r0[51:51], i_0r1[51:51]);
  OR2 I52 (gocomp_0[52:52], i_0r0[52:52], i_0r1[52:52]);
  OR2 I53 (gocomp_0[53:53], i_0r0[53:53], i_0r1[53:53]);
  OR2 I54 (gocomp_0[54:54], i_0r0[54:54], i_0r1[54:54]);
  OR2 I55 (gocomp_0[55:55], i_0r0[55:55], i_0r1[55:55]);
  OR2 I56 (gocomp_0[56:56], i_0r0[56:56], i_0r1[56:56]);
  OR2 I57 (gocomp_0[57:57], i_0r0[57:57], i_0r1[57:57]);
  OR2 I58 (gocomp_0[58:58], i_0r0[58:58], i_0r1[58:58]);
  OR2 I59 (gocomp_0[59:59], i_0r0[59:59], i_0r1[59:59]);
  OR2 I60 (gocomp_0[60:60], i_0r0[60:60], i_0r1[60:60]);
  OR2 I61 (gocomp_0[61:61], i_0r0[61:61], i_0r1[61:61]);
  OR2 I62 (gocomp_0[62:62], i_0r0[62:62], i_0r1[62:62]);
  OR2 I63 (gocomp_0[63:63], i_0r0[63:63], i_0r1[63:63]);
  OR2 I64 (gocomp_0[64:64], i_0r0[64:64], i_0r1[64:64]);
  OR2 I65 (gocomp_0[65:65], i_0r0[65:65], i_0r1[65:65]);
  C3 I66 (simp681_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  C3 I67 (simp681_0[1:1], gocomp_0[3:3], gocomp_0[4:4], gocomp_0[5:5]);
  C3 I68 (simp681_0[2:2], gocomp_0[6:6], gocomp_0[7:7], gocomp_0[8:8]);
  C3 I69 (simp681_0[3:3], gocomp_0[9:9], gocomp_0[10:10], gocomp_0[11:11]);
  C3 I70 (simp681_0[4:4], gocomp_0[12:12], gocomp_0[13:13], gocomp_0[14:14]);
  C3 I71 (simp681_0[5:5], gocomp_0[15:15], gocomp_0[16:16], gocomp_0[17:17]);
  C3 I72 (simp681_0[6:6], gocomp_0[18:18], gocomp_0[19:19], gocomp_0[20:20]);
  C3 I73 (simp681_0[7:7], gocomp_0[21:21], gocomp_0[22:22], gocomp_0[23:23]);
  C3 I74 (simp681_0[8:8], gocomp_0[24:24], gocomp_0[25:25], gocomp_0[26:26]);
  C3 I75 (simp681_0[9:9], gocomp_0[27:27], gocomp_0[28:28], gocomp_0[29:29]);
  C3 I76 (simp681_0[10:10], gocomp_0[30:30], gocomp_0[31:31], gocomp_0[32:32]);
  C3 I77 (simp681_0[11:11], gocomp_0[33:33], gocomp_0[34:34], gocomp_0[35:35]);
  C3 I78 (simp681_0[12:12], gocomp_0[36:36], gocomp_0[37:37], gocomp_0[38:38]);
  C3 I79 (simp681_0[13:13], gocomp_0[39:39], gocomp_0[40:40], gocomp_0[41:41]);
  C3 I80 (simp681_0[14:14], gocomp_0[42:42], gocomp_0[43:43], gocomp_0[44:44]);
  C3 I81 (simp681_0[15:15], gocomp_0[45:45], gocomp_0[46:46], gocomp_0[47:47]);
  C3 I82 (simp681_0[16:16], gocomp_0[48:48], gocomp_0[49:49], gocomp_0[50:50]);
  C3 I83 (simp681_0[17:17], gocomp_0[51:51], gocomp_0[52:52], gocomp_0[53:53]);
  C3 I84 (simp681_0[18:18], gocomp_0[54:54], gocomp_0[55:55], gocomp_0[56:56]);
  C3 I85 (simp681_0[19:19], gocomp_0[57:57], gocomp_0[58:58], gocomp_0[59:59]);
  C3 I86 (simp681_0[20:20], gocomp_0[60:60], gocomp_0[61:61], gocomp_0[62:62]);
  C3 I87 (simp681_0[21:21], gocomp_0[63:63], gocomp_0[64:64], gocomp_0[65:65]);
  C3 I88 (simp682_0[0:0], simp681_0[0:0], simp681_0[1:1], simp681_0[2:2]);
  C3 I89 (simp682_0[1:1], simp681_0[3:3], simp681_0[4:4], simp681_0[5:5]);
  C3 I90 (simp682_0[2:2], simp681_0[6:6], simp681_0[7:7], simp681_0[8:8]);
  C3 I91 (simp682_0[3:3], simp681_0[9:9], simp681_0[10:10], simp681_0[11:11]);
  C3 I92 (simp682_0[4:4], simp681_0[12:12], simp681_0[13:13], simp681_0[14:14]);
  C3 I93 (simp682_0[5:5], simp681_0[15:15], simp681_0[16:16], simp681_0[17:17]);
  C3 I94 (simp682_0[6:6], simp681_0[18:18], simp681_0[19:19], simp681_0[20:20]);
  BUFF I95 (simp682_0[7:7], simp681_0[21:21]);
  C3 I96 (simp683_0[0:0], simp682_0[0:0], simp682_0[1:1], simp682_0[2:2]);
  C3 I97 (simp683_0[1:1], simp682_0[3:3], simp682_0[4:4], simp682_0[5:5]);
  C2 I98 (simp683_0[2:2], simp682_0[6:6], simp682_0[7:7]);
  C3 I99 (go_0, simp683_0[0:0], simp683_0[1:1], simp683_0[2:2]);
  BUFF I100 (termf_1[0:0], i_0r0[0:0]);
  BUFF I101 (termf_1[1:1], i_0r0[1:1]);
  BUFF I102 (termf_1[2:2], i_0r0[2:2]);
  BUFF I103 (termf_1[3:3], i_0r0[3:3]);
  BUFF I104 (termf_1[4:4], i_0r0[4:4]);
  BUFF I105 (termf_1[5:5], i_0r0[5:5]);
  BUFF I106 (termf_1[6:6], i_0r0[6:6]);
  BUFF I107 (termf_1[7:7], i_0r0[7:7]);
  BUFF I108 (termf_1[8:8], i_0r0[8:8]);
  BUFF I109 (termf_1[9:9], i_0r0[9:9]);
  BUFF I110 (termf_1[10:10], i_0r0[10:10]);
  BUFF I111 (termf_1[11:11], i_0r0[11:11]);
  BUFF I112 (termf_1[12:12], i_0r0[12:12]);
  BUFF I113 (termf_1[13:13], i_0r0[13:13]);
  BUFF I114 (termf_1[14:14], i_0r0[14:14]);
  BUFF I115 (termf_1[15:15], i_0r0[15:15]);
  BUFF I116 (termf_1[16:16], i_0r0[16:16]);
  BUFF I117 (termf_1[17:17], i_0r0[17:17]);
  BUFF I118 (termf_1[18:18], i_0r0[18:18]);
  BUFF I119 (termf_1[19:19], i_0r0[19:19]);
  BUFF I120 (termf_1[20:20], i_0r0[20:20]);
  BUFF I121 (termf_1[21:21], i_0r0[21:21]);
  BUFF I122 (termf_1[22:22], i_0r0[22:22]);
  BUFF I123 (termf_1[23:23], i_0r0[23:23]);
  BUFF I124 (termf_1[24:24], i_0r0[24:24]);
  BUFF I125 (termf_1[25:25], i_0r0[25:25]);
  BUFF I126 (termf_1[26:26], i_0r0[26:26]);
  BUFF I127 (termf_1[27:27], i_0r0[27:27]);
  BUFF I128 (termf_1[28:28], i_0r0[28:28]);
  BUFF I129 (termf_1[29:29], i_0r0[29:29]);
  BUFF I130 (termf_1[30:30], i_0r0[30:30]);
  BUFF I131 (termf_1[31:31], i_0r0[31:31]);
  BUFF I132 (termf_1[32:32], i_0r0[32:32]);
  BUFF I133 (termt_1[0:0], i_0r1[0:0]);
  BUFF I134 (termt_1[1:1], i_0r1[1:1]);
  BUFF I135 (termt_1[2:2], i_0r1[2:2]);
  BUFF I136 (termt_1[3:3], i_0r1[3:3]);
  BUFF I137 (termt_1[4:4], i_0r1[4:4]);
  BUFF I138 (termt_1[5:5], i_0r1[5:5]);
  BUFF I139 (termt_1[6:6], i_0r1[6:6]);
  BUFF I140 (termt_1[7:7], i_0r1[7:7]);
  BUFF I141 (termt_1[8:8], i_0r1[8:8]);
  BUFF I142 (termt_1[9:9], i_0r1[9:9]);
  BUFF I143 (termt_1[10:10], i_0r1[10:10]);
  BUFF I144 (termt_1[11:11], i_0r1[11:11]);
  BUFF I145 (termt_1[12:12], i_0r1[12:12]);
  BUFF I146 (termt_1[13:13], i_0r1[13:13]);
  BUFF I147 (termt_1[14:14], i_0r1[14:14]);
  BUFF I148 (termt_1[15:15], i_0r1[15:15]);
  BUFF I149 (termt_1[16:16], i_0r1[16:16]);
  BUFF I150 (termt_1[17:17], i_0r1[17:17]);
  BUFF I151 (termt_1[18:18], i_0r1[18:18]);
  BUFF I152 (termt_1[19:19], i_0r1[19:19]);
  BUFF I153 (termt_1[20:20], i_0r1[20:20]);
  BUFF I154 (termt_1[21:21], i_0r1[21:21]);
  BUFF I155 (termt_1[22:22], i_0r1[22:22]);
  BUFF I156 (termt_1[23:23], i_0r1[23:23]);
  BUFF I157 (termt_1[24:24], i_0r1[24:24]);
  BUFF I158 (termt_1[25:25], i_0r1[25:25]);
  BUFF I159 (termt_1[26:26], i_0r1[26:26]);
  BUFF I160 (termt_1[27:27], i_0r1[27:27]);
  BUFF I161 (termt_1[28:28], i_0r1[28:28]);
  BUFF I162 (termt_1[29:29], i_0r1[29:29]);
  BUFF I163 (termt_1[30:30], i_0r1[30:30]);
  BUFF I164 (termt_1[31:31], i_0r1[31:31]);
  BUFF I165 (termt_1[32:32], i_0r1[32:32]);
  BUFF I166 (termf_2[0:0], i_0r0[33:33]);
  BUFF I167 (termf_2[1:1], i_0r0[34:34]);
  BUFF I168 (termf_2[2:2], i_0r0[35:35]);
  BUFF I169 (termf_2[3:3], i_0r0[36:36]);
  BUFF I170 (termf_2[4:4], i_0r0[37:37]);
  BUFF I171 (termf_2[5:5], i_0r0[38:38]);
  BUFF I172 (termf_2[6:6], i_0r0[39:39]);
  BUFF I173 (termf_2[7:7], i_0r0[40:40]);
  BUFF I174 (termf_2[8:8], i_0r0[41:41]);
  BUFF I175 (termf_2[9:9], i_0r0[42:42]);
  BUFF I176 (termf_2[10:10], i_0r0[43:43]);
  BUFF I177 (termf_2[11:11], i_0r0[44:44]);
  BUFF I178 (termf_2[12:12], i_0r0[45:45]);
  BUFF I179 (termf_2[13:13], i_0r0[46:46]);
  BUFF I180 (termf_2[14:14], i_0r0[47:47]);
  BUFF I181 (termf_2[15:15], i_0r0[48:48]);
  BUFF I182 (termf_2[16:16], i_0r0[49:49]);
  BUFF I183 (termf_2[17:17], i_0r0[50:50]);
  BUFF I184 (termf_2[18:18], i_0r0[51:51]);
  BUFF I185 (termf_2[19:19], i_0r0[52:52]);
  BUFF I186 (termf_2[20:20], i_0r0[53:53]);
  BUFF I187 (termf_2[21:21], i_0r0[54:54]);
  BUFF I188 (termf_2[22:22], i_0r0[55:55]);
  BUFF I189 (termf_2[23:23], i_0r0[56:56]);
  BUFF I190 (termf_2[24:24], i_0r0[57:57]);
  BUFF I191 (termf_2[25:25], i_0r0[58:58]);
  BUFF I192 (termf_2[26:26], i_0r0[59:59]);
  BUFF I193 (termf_2[27:27], i_0r0[60:60]);
  BUFF I194 (termf_2[28:28], i_0r0[61:61]);
  BUFF I195 (termf_2[29:29], i_0r0[62:62]);
  BUFF I196 (termf_2[30:30], i_0r0[63:63]);
  BUFF I197 (termf_2[31:31], i_0r0[64:64]);
  BUFF I198 (termf_2[32:32], i_0r0[65:65]);
  BUFF I199 (termt_2[0:0], i_0r1[33:33]);
  BUFF I200 (termt_2[1:1], i_0r1[34:34]);
  BUFF I201 (termt_2[2:2], i_0r1[35:35]);
  BUFF I202 (termt_2[3:3], i_0r1[36:36]);
  BUFF I203 (termt_2[4:4], i_0r1[37:37]);
  BUFF I204 (termt_2[5:5], i_0r1[38:38]);
  BUFF I205 (termt_2[6:6], i_0r1[39:39]);
  BUFF I206 (termt_2[7:7], i_0r1[40:40]);
  BUFF I207 (termt_2[8:8], i_0r1[41:41]);
  BUFF I208 (termt_2[9:9], i_0r1[42:42]);
  BUFF I209 (termt_2[10:10], i_0r1[43:43]);
  BUFF I210 (termt_2[11:11], i_0r1[44:44]);
  BUFF I211 (termt_2[12:12], i_0r1[45:45]);
  BUFF I212 (termt_2[13:13], i_0r1[46:46]);
  BUFF I213 (termt_2[14:14], i_0r1[47:47]);
  BUFF I214 (termt_2[15:15], i_0r1[48:48]);
  BUFF I215 (termt_2[16:16], i_0r1[49:49]);
  BUFF I216 (termt_2[17:17], i_0r1[50:50]);
  BUFF I217 (termt_2[18:18], i_0r1[51:51]);
  BUFF I218 (termt_2[19:19], i_0r1[52:52]);
  BUFF I219 (termt_2[20:20], i_0r1[53:53]);
  BUFF I220 (termt_2[21:21], i_0r1[54:54]);
  BUFF I221 (termt_2[22:22], i_0r1[55:55]);
  BUFF I222 (termt_2[23:23], i_0r1[56:56]);
  BUFF I223 (termt_2[24:24], i_0r1[57:57]);
  BUFF I224 (termt_2[25:25], i_0r1[58:58]);
  BUFF I225 (termt_2[26:26], i_0r1[59:59]);
  BUFF I226 (termt_2[27:27], i_0r1[60:60]);
  BUFF I227 (termt_2[28:28], i_0r1[61:61]);
  BUFF I228 (termt_2[29:29], i_0r1[62:62]);
  BUFF I229 (termt_2[30:30], i_0r1[63:63]);
  BUFF I230 (termt_2[31:31], i_0r1[64:64]);
  BUFF I231 (termt_2[32:32], i_0r1[65:65]);
  BUFF I232 (termf_3, go_0);
  GND I233 (termt_3);
  BUFF I234 (termf_4[0:0], termf_1[0:0]);
  BUFF I235 (termf_4[1:1], termf_1[1:1]);
  BUFF I236 (termf_4[2:2], termf_1[2:2]);
  BUFF I237 (termf_4[3:3], termf_1[3:3]);
  BUFF I238 (termf_4[4:4], termf_1[4:4]);
  BUFF I239 (termf_4[5:5], termf_1[5:5]);
  BUFF I240 (termf_4[6:6], termf_1[6:6]);
  BUFF I241 (termf_4[7:7], termf_1[7:7]);
  BUFF I242 (termf_4[8:8], termf_1[8:8]);
  BUFF I243 (termf_4[9:9], termf_1[9:9]);
  BUFF I244 (termf_4[10:10], termf_1[10:10]);
  BUFF I245 (termf_4[11:11], termf_1[11:11]);
  BUFF I246 (termf_4[12:12], termf_1[12:12]);
  BUFF I247 (termf_4[13:13], termf_1[13:13]);
  BUFF I248 (termf_4[14:14], termf_1[14:14]);
  BUFF I249 (termf_4[15:15], termf_1[15:15]);
  BUFF I250 (termf_4[16:16], termf_1[16:16]);
  BUFF I251 (termf_4[17:17], termf_1[17:17]);
  BUFF I252 (termf_4[18:18], termf_1[18:18]);
  BUFF I253 (termf_4[19:19], termf_1[19:19]);
  BUFF I254 (termf_4[20:20], termf_1[20:20]);
  BUFF I255 (termf_4[21:21], termf_1[21:21]);
  BUFF I256 (termf_4[22:22], termf_1[22:22]);
  BUFF I257 (termf_4[23:23], termf_1[23:23]);
  BUFF I258 (termf_4[24:24], termf_1[24:24]);
  BUFF I259 (termf_4[25:25], termf_1[25:25]);
  BUFF I260 (termf_4[26:26], termf_1[26:26]);
  BUFF I261 (termf_4[27:27], termf_1[27:27]);
  BUFF I262 (termf_4[28:28], termf_1[28:28]);
  BUFF I263 (termf_4[29:29], termf_1[29:29]);
  BUFF I264 (termf_4[30:30], termf_1[30:30]);
  BUFF I265 (termf_4[31:31], termf_1[31:31]);
  BUFF I266 (termf_4[32:32], termf_1[32:32]);
  BUFF I267 (termf_4[33:33], termf_3);
  BUFF I268 (termt_4[0:0], termt_1[0:0]);
  BUFF I269 (termt_4[1:1], termt_1[1:1]);
  BUFF I270 (termt_4[2:2], termt_1[2:2]);
  BUFF I271 (termt_4[3:3], termt_1[3:3]);
  BUFF I272 (termt_4[4:4], termt_1[4:4]);
  BUFF I273 (termt_4[5:5], termt_1[5:5]);
  BUFF I274 (termt_4[6:6], termt_1[6:6]);
  BUFF I275 (termt_4[7:7], termt_1[7:7]);
  BUFF I276 (termt_4[8:8], termt_1[8:8]);
  BUFF I277 (termt_4[9:9], termt_1[9:9]);
  BUFF I278 (termt_4[10:10], termt_1[10:10]);
  BUFF I279 (termt_4[11:11], termt_1[11:11]);
  BUFF I280 (termt_4[12:12], termt_1[12:12]);
  BUFF I281 (termt_4[13:13], termt_1[13:13]);
  BUFF I282 (termt_4[14:14], termt_1[14:14]);
  BUFF I283 (termt_4[15:15], termt_1[15:15]);
  BUFF I284 (termt_4[16:16], termt_1[16:16]);
  BUFF I285 (termt_4[17:17], termt_1[17:17]);
  BUFF I286 (termt_4[18:18], termt_1[18:18]);
  BUFF I287 (termt_4[19:19], termt_1[19:19]);
  BUFF I288 (termt_4[20:20], termt_1[20:20]);
  BUFF I289 (termt_4[21:21], termt_1[21:21]);
  BUFF I290 (termt_4[22:22], termt_1[22:22]);
  BUFF I291 (termt_4[23:23], termt_1[23:23]);
  BUFF I292 (termt_4[24:24], termt_1[24:24]);
  BUFF I293 (termt_4[25:25], termt_1[25:25]);
  BUFF I294 (termt_4[26:26], termt_1[26:26]);
  BUFF I295 (termt_4[27:27], termt_1[27:27]);
  BUFF I296 (termt_4[28:28], termt_1[28:28]);
  BUFF I297 (termt_4[29:29], termt_1[29:29]);
  BUFF I298 (termt_4[30:30], termt_1[30:30]);
  BUFF I299 (termt_4[31:31], termt_1[31:31]);
  BUFF I300 (termt_4[32:32], termt_1[32:32]);
  BUFF I301 (termt_4[33:33], termt_3);
  BUFF I302 (termf_5, go_0);
  GND I303 (termt_5);
  BUFF I304 (termf_6[0:0], termf_2[0:0]);
  BUFF I305 (termf_6[1:1], termf_2[1:1]);
  BUFF I306 (termf_6[2:2], termf_2[2:2]);
  BUFF I307 (termf_6[3:3], termf_2[3:3]);
  BUFF I308 (termf_6[4:4], termf_2[4:4]);
  BUFF I309 (termf_6[5:5], termf_2[5:5]);
  BUFF I310 (termf_6[6:6], termf_2[6:6]);
  BUFF I311 (termf_6[7:7], termf_2[7:7]);
  BUFF I312 (termf_6[8:8], termf_2[8:8]);
  BUFF I313 (termf_6[9:9], termf_2[9:9]);
  BUFF I314 (termf_6[10:10], termf_2[10:10]);
  BUFF I315 (termf_6[11:11], termf_2[11:11]);
  BUFF I316 (termf_6[12:12], termf_2[12:12]);
  BUFF I317 (termf_6[13:13], termf_2[13:13]);
  BUFF I318 (termf_6[14:14], termf_2[14:14]);
  BUFF I319 (termf_6[15:15], termf_2[15:15]);
  BUFF I320 (termf_6[16:16], termf_2[16:16]);
  BUFF I321 (termf_6[17:17], termf_2[17:17]);
  BUFF I322 (termf_6[18:18], termf_2[18:18]);
  BUFF I323 (termf_6[19:19], termf_2[19:19]);
  BUFF I324 (termf_6[20:20], termf_2[20:20]);
  BUFF I325 (termf_6[21:21], termf_2[21:21]);
  BUFF I326 (termf_6[22:22], termf_2[22:22]);
  BUFF I327 (termf_6[23:23], termf_2[23:23]);
  BUFF I328 (termf_6[24:24], termf_2[24:24]);
  BUFF I329 (termf_6[25:25], termf_2[25:25]);
  BUFF I330 (termf_6[26:26], termf_2[26:26]);
  BUFF I331 (termf_6[27:27], termf_2[27:27]);
  BUFF I332 (termf_6[28:28], termf_2[28:28]);
  BUFF I333 (termf_6[29:29], termf_2[29:29]);
  BUFF I334 (termf_6[30:30], termf_2[30:30]);
  BUFF I335 (termf_6[31:31], termf_2[31:31]);
  BUFF I336 (termf_6[32:32], termf_2[32:32]);
  BUFF I337 (termf_6[33:33], termf_5);
  BUFF I338 (termt_6[0:0], termt_2[0:0]);
  BUFF I339 (termt_6[1:1], termt_2[1:1]);
  BUFF I340 (termt_6[2:2], termt_2[2:2]);
  BUFF I341 (termt_6[3:3], termt_2[3:3]);
  BUFF I342 (termt_6[4:4], termt_2[4:4]);
  BUFF I343 (termt_6[5:5], termt_2[5:5]);
  BUFF I344 (termt_6[6:6], termt_2[6:6]);
  BUFF I345 (termt_6[7:7], termt_2[7:7]);
  BUFF I346 (termt_6[8:8], termt_2[8:8]);
  BUFF I347 (termt_6[9:9], termt_2[9:9]);
  BUFF I348 (termt_6[10:10], termt_2[10:10]);
  BUFF I349 (termt_6[11:11], termt_2[11:11]);
  BUFF I350 (termt_6[12:12], termt_2[12:12]);
  BUFF I351 (termt_6[13:13], termt_2[13:13]);
  BUFF I352 (termt_6[14:14], termt_2[14:14]);
  BUFF I353 (termt_6[15:15], termt_2[15:15]);
  BUFF I354 (termt_6[16:16], termt_2[16:16]);
  BUFF I355 (termt_6[17:17], termt_2[17:17]);
  BUFF I356 (termt_6[18:18], termt_2[18:18]);
  BUFF I357 (termt_6[19:19], termt_2[19:19]);
  BUFF I358 (termt_6[20:20], termt_2[20:20]);
  BUFF I359 (termt_6[21:21], termt_2[21:21]);
  BUFF I360 (termt_6[22:22], termt_2[22:22]);
  BUFF I361 (termt_6[23:23], termt_2[23:23]);
  BUFF I362 (termt_6[24:24], termt_2[24:24]);
  BUFF I363 (termt_6[25:25], termt_2[25:25]);
  BUFF I364 (termt_6[26:26], termt_2[26:26]);
  BUFF I365 (termt_6[27:27], termt_2[27:27]);
  BUFF I366 (termt_6[28:28], termt_2[28:28]);
  BUFF I367 (termt_6[29:29], termt_2[29:29]);
  BUFF I368 (termt_6[30:30], termt_2[30:30]);
  BUFF I369 (termt_6[31:31], termt_2[31:31]);
  BUFF I370 (termt_6[32:32], termt_2[32:32]);
  BUFF I371 (termt_6[33:33], termt_5);
  C2 I372 (ha7__0[0:0], termf_6[0:0], termf_4[0:0]);
  C2 I373 (ha7__0[1:1], termf_6[0:0], termt_4[0:0]);
  C2 I374 (ha7__0[2:2], termt_6[0:0], termf_4[0:0]);
  C2 I375 (ha7__0[3:3], termt_6[0:0], termt_4[0:0]);
  OR3 I376 (cf7__0[0:0], ha7__0[0:0], ha7__0[1:1], ha7__0[2:2]);
  BUFF I377 (ct7__0[0:0], ha7__0[3:3]);
  OR2 I378 (o_0r0[0:0], ha7__0[0:0], ha7__0[3:3]);
  OR2 I379 (o_0r1[0:0], ha7__0[1:1], ha7__0[2:2]);
  C3 I380 (fa7_1min_0[0:0], cf7__0[0:0], termf_6[1:1], termf_4[1:1]);
  C3 I381 (fa7_1min_0[1:1], cf7__0[0:0], termf_6[1:1], termt_4[1:1]);
  C3 I382 (fa7_1min_0[2:2], cf7__0[0:0], termt_6[1:1], termf_4[1:1]);
  C3 I383 (fa7_1min_0[3:3], cf7__0[0:0], termt_6[1:1], termt_4[1:1]);
  C3 I384 (fa7_1min_0[4:4], ct7__0[0:0], termf_6[1:1], termf_4[1:1]);
  C3 I385 (fa7_1min_0[5:5], ct7__0[0:0], termf_6[1:1], termt_4[1:1]);
  C3 I386 (fa7_1min_0[6:6], ct7__0[0:0], termt_6[1:1], termf_4[1:1]);
  C3 I387 (fa7_1min_0[7:7], ct7__0[0:0], termt_6[1:1], termt_4[1:1]);
  NOR3 I388 (simp3751_0[0:0], fa7_1min_0[0:0], fa7_1min_0[3:3], fa7_1min_0[5:5]);
  INV I389 (simp3751_0[1:1], fa7_1min_0[6:6]);
  NAND2 I390 (o_0r0[1:1], simp3751_0[0:0], simp3751_0[1:1]);
  NOR3 I391 (simp3761_0[0:0], fa7_1min_0[1:1], fa7_1min_0[2:2], fa7_1min_0[4:4]);
  INV I392 (simp3761_0[1:1], fa7_1min_0[7:7]);
  NAND2 I393 (o_0r1[1:1], simp3761_0[0:0], simp3761_0[1:1]);
  AO222 I394 (ct7__0[1:1], termt_4[1:1], termt_6[1:1], termt_4[1:1], ct7__0[0:0], termt_6[1:1], ct7__0[0:0]);
  AO222 I395 (cf7__0[1:1], termf_4[1:1], termf_6[1:1], termf_4[1:1], cf7__0[0:0], termf_6[1:1], cf7__0[0:0]);
  C3 I396 (fa7_2min_0[0:0], cf7__0[1:1], termf_6[2:2], termf_4[2:2]);
  C3 I397 (fa7_2min_0[1:1], cf7__0[1:1], termf_6[2:2], termt_4[2:2]);
  C3 I398 (fa7_2min_0[2:2], cf7__0[1:1], termt_6[2:2], termf_4[2:2]);
  C3 I399 (fa7_2min_0[3:3], cf7__0[1:1], termt_6[2:2], termt_4[2:2]);
  C3 I400 (fa7_2min_0[4:4], ct7__0[1:1], termf_6[2:2], termf_4[2:2]);
  C3 I401 (fa7_2min_0[5:5], ct7__0[1:1], termf_6[2:2], termt_4[2:2]);
  C3 I402 (fa7_2min_0[6:6], ct7__0[1:1], termt_6[2:2], termf_4[2:2]);
  C3 I403 (fa7_2min_0[7:7], ct7__0[1:1], termt_6[2:2], termt_4[2:2]);
  NOR3 I404 (simp3881_0[0:0], fa7_2min_0[0:0], fa7_2min_0[3:3], fa7_2min_0[5:5]);
  INV I405 (simp3881_0[1:1], fa7_2min_0[6:6]);
  NAND2 I406 (o_0r0[2:2], simp3881_0[0:0], simp3881_0[1:1]);
  NOR3 I407 (simp3891_0[0:0], fa7_2min_0[1:1], fa7_2min_0[2:2], fa7_2min_0[4:4]);
  INV I408 (simp3891_0[1:1], fa7_2min_0[7:7]);
  NAND2 I409 (o_0r1[2:2], simp3891_0[0:0], simp3891_0[1:1]);
  AO222 I410 (ct7__0[2:2], termt_4[2:2], termt_6[2:2], termt_4[2:2], ct7__0[1:1], termt_6[2:2], ct7__0[1:1]);
  AO222 I411 (cf7__0[2:2], termf_4[2:2], termf_6[2:2], termf_4[2:2], cf7__0[1:1], termf_6[2:2], cf7__0[1:1]);
  C3 I412 (fa7_3min_0[0:0], cf7__0[2:2], termf_6[3:3], termf_4[3:3]);
  C3 I413 (fa7_3min_0[1:1], cf7__0[2:2], termf_6[3:3], termt_4[3:3]);
  C3 I414 (fa7_3min_0[2:2], cf7__0[2:2], termt_6[3:3], termf_4[3:3]);
  C3 I415 (fa7_3min_0[3:3], cf7__0[2:2], termt_6[3:3], termt_4[3:3]);
  C3 I416 (fa7_3min_0[4:4], ct7__0[2:2], termf_6[3:3], termf_4[3:3]);
  C3 I417 (fa7_3min_0[5:5], ct7__0[2:2], termf_6[3:3], termt_4[3:3]);
  C3 I418 (fa7_3min_0[6:6], ct7__0[2:2], termt_6[3:3], termf_4[3:3]);
  C3 I419 (fa7_3min_0[7:7], ct7__0[2:2], termt_6[3:3], termt_4[3:3]);
  NOR3 I420 (simp4011_0[0:0], fa7_3min_0[0:0], fa7_3min_0[3:3], fa7_3min_0[5:5]);
  INV I421 (simp4011_0[1:1], fa7_3min_0[6:6]);
  NAND2 I422 (o_0r0[3:3], simp4011_0[0:0], simp4011_0[1:1]);
  NOR3 I423 (simp4021_0[0:0], fa7_3min_0[1:1], fa7_3min_0[2:2], fa7_3min_0[4:4]);
  INV I424 (simp4021_0[1:1], fa7_3min_0[7:7]);
  NAND2 I425 (o_0r1[3:3], simp4021_0[0:0], simp4021_0[1:1]);
  AO222 I426 (ct7__0[3:3], termt_4[3:3], termt_6[3:3], termt_4[3:3], ct7__0[2:2], termt_6[3:3], ct7__0[2:2]);
  AO222 I427 (cf7__0[3:3], termf_4[3:3], termf_6[3:3], termf_4[3:3], cf7__0[2:2], termf_6[3:3], cf7__0[2:2]);
  C3 I428 (fa7_4min_0[0:0], cf7__0[3:3], termf_6[4:4], termf_4[4:4]);
  C3 I429 (fa7_4min_0[1:1], cf7__0[3:3], termf_6[4:4], termt_4[4:4]);
  C3 I430 (fa7_4min_0[2:2], cf7__0[3:3], termt_6[4:4], termf_4[4:4]);
  C3 I431 (fa7_4min_0[3:3], cf7__0[3:3], termt_6[4:4], termt_4[4:4]);
  C3 I432 (fa7_4min_0[4:4], ct7__0[3:3], termf_6[4:4], termf_4[4:4]);
  C3 I433 (fa7_4min_0[5:5], ct7__0[3:3], termf_6[4:4], termt_4[4:4]);
  C3 I434 (fa7_4min_0[6:6], ct7__0[3:3], termt_6[4:4], termf_4[4:4]);
  C3 I435 (fa7_4min_0[7:7], ct7__0[3:3], termt_6[4:4], termt_4[4:4]);
  NOR3 I436 (simp4141_0[0:0], fa7_4min_0[0:0], fa7_4min_0[3:3], fa7_4min_0[5:5]);
  INV I437 (simp4141_0[1:1], fa7_4min_0[6:6]);
  NAND2 I438 (o_0r0[4:4], simp4141_0[0:0], simp4141_0[1:1]);
  NOR3 I439 (simp4151_0[0:0], fa7_4min_0[1:1], fa7_4min_0[2:2], fa7_4min_0[4:4]);
  INV I440 (simp4151_0[1:1], fa7_4min_0[7:7]);
  NAND2 I441 (o_0r1[4:4], simp4151_0[0:0], simp4151_0[1:1]);
  AO222 I442 (ct7__0[4:4], termt_4[4:4], termt_6[4:4], termt_4[4:4], ct7__0[3:3], termt_6[4:4], ct7__0[3:3]);
  AO222 I443 (cf7__0[4:4], termf_4[4:4], termf_6[4:4], termf_4[4:4], cf7__0[3:3], termf_6[4:4], cf7__0[3:3]);
  C3 I444 (fa7_5min_0[0:0], cf7__0[4:4], termf_6[5:5], termf_4[5:5]);
  C3 I445 (fa7_5min_0[1:1], cf7__0[4:4], termf_6[5:5], termt_4[5:5]);
  C3 I446 (fa7_5min_0[2:2], cf7__0[4:4], termt_6[5:5], termf_4[5:5]);
  C3 I447 (fa7_5min_0[3:3], cf7__0[4:4], termt_6[5:5], termt_4[5:5]);
  C3 I448 (fa7_5min_0[4:4], ct7__0[4:4], termf_6[5:5], termf_4[5:5]);
  C3 I449 (fa7_5min_0[5:5], ct7__0[4:4], termf_6[5:5], termt_4[5:5]);
  C3 I450 (fa7_5min_0[6:6], ct7__0[4:4], termt_6[5:5], termf_4[5:5]);
  C3 I451 (fa7_5min_0[7:7], ct7__0[4:4], termt_6[5:5], termt_4[5:5]);
  NOR3 I452 (simp4271_0[0:0], fa7_5min_0[0:0], fa7_5min_0[3:3], fa7_5min_0[5:5]);
  INV I453 (simp4271_0[1:1], fa7_5min_0[6:6]);
  NAND2 I454 (o_0r0[5:5], simp4271_0[0:0], simp4271_0[1:1]);
  NOR3 I455 (simp4281_0[0:0], fa7_5min_0[1:1], fa7_5min_0[2:2], fa7_5min_0[4:4]);
  INV I456 (simp4281_0[1:1], fa7_5min_0[7:7]);
  NAND2 I457 (o_0r1[5:5], simp4281_0[0:0], simp4281_0[1:1]);
  AO222 I458 (ct7__0[5:5], termt_4[5:5], termt_6[5:5], termt_4[5:5], ct7__0[4:4], termt_6[5:5], ct7__0[4:4]);
  AO222 I459 (cf7__0[5:5], termf_4[5:5], termf_6[5:5], termf_4[5:5], cf7__0[4:4], termf_6[5:5], cf7__0[4:4]);
  C3 I460 (fa7_6min_0[0:0], cf7__0[5:5], termf_6[6:6], termf_4[6:6]);
  C3 I461 (fa7_6min_0[1:1], cf7__0[5:5], termf_6[6:6], termt_4[6:6]);
  C3 I462 (fa7_6min_0[2:2], cf7__0[5:5], termt_6[6:6], termf_4[6:6]);
  C3 I463 (fa7_6min_0[3:3], cf7__0[5:5], termt_6[6:6], termt_4[6:6]);
  C3 I464 (fa7_6min_0[4:4], ct7__0[5:5], termf_6[6:6], termf_4[6:6]);
  C3 I465 (fa7_6min_0[5:5], ct7__0[5:5], termf_6[6:6], termt_4[6:6]);
  C3 I466 (fa7_6min_0[6:6], ct7__0[5:5], termt_6[6:6], termf_4[6:6]);
  C3 I467 (fa7_6min_0[7:7], ct7__0[5:5], termt_6[6:6], termt_4[6:6]);
  NOR3 I468 (simp4401_0[0:0], fa7_6min_0[0:0], fa7_6min_0[3:3], fa7_6min_0[5:5]);
  INV I469 (simp4401_0[1:1], fa7_6min_0[6:6]);
  NAND2 I470 (o_0r0[6:6], simp4401_0[0:0], simp4401_0[1:1]);
  NOR3 I471 (simp4411_0[0:0], fa7_6min_0[1:1], fa7_6min_0[2:2], fa7_6min_0[4:4]);
  INV I472 (simp4411_0[1:1], fa7_6min_0[7:7]);
  NAND2 I473 (o_0r1[6:6], simp4411_0[0:0], simp4411_0[1:1]);
  AO222 I474 (ct7__0[6:6], termt_4[6:6], termt_6[6:6], termt_4[6:6], ct7__0[5:5], termt_6[6:6], ct7__0[5:5]);
  AO222 I475 (cf7__0[6:6], termf_4[6:6], termf_6[6:6], termf_4[6:6], cf7__0[5:5], termf_6[6:6], cf7__0[5:5]);
  C3 I476 (fa7_7min_0[0:0], cf7__0[6:6], termf_6[7:7], termf_4[7:7]);
  C3 I477 (fa7_7min_0[1:1], cf7__0[6:6], termf_6[7:7], termt_4[7:7]);
  C3 I478 (fa7_7min_0[2:2], cf7__0[6:6], termt_6[7:7], termf_4[7:7]);
  C3 I479 (fa7_7min_0[3:3], cf7__0[6:6], termt_6[7:7], termt_4[7:7]);
  C3 I480 (fa7_7min_0[4:4], ct7__0[6:6], termf_6[7:7], termf_4[7:7]);
  C3 I481 (fa7_7min_0[5:5], ct7__0[6:6], termf_6[7:7], termt_4[7:7]);
  C3 I482 (fa7_7min_0[6:6], ct7__0[6:6], termt_6[7:7], termf_4[7:7]);
  C3 I483 (fa7_7min_0[7:7], ct7__0[6:6], termt_6[7:7], termt_4[7:7]);
  NOR3 I484 (simp4531_0[0:0], fa7_7min_0[0:0], fa7_7min_0[3:3], fa7_7min_0[5:5]);
  INV I485 (simp4531_0[1:1], fa7_7min_0[6:6]);
  NAND2 I486 (o_0r0[7:7], simp4531_0[0:0], simp4531_0[1:1]);
  NOR3 I487 (simp4541_0[0:0], fa7_7min_0[1:1], fa7_7min_0[2:2], fa7_7min_0[4:4]);
  INV I488 (simp4541_0[1:1], fa7_7min_0[7:7]);
  NAND2 I489 (o_0r1[7:7], simp4541_0[0:0], simp4541_0[1:1]);
  AO222 I490 (ct7__0[7:7], termt_4[7:7], termt_6[7:7], termt_4[7:7], ct7__0[6:6], termt_6[7:7], ct7__0[6:6]);
  AO222 I491 (cf7__0[7:7], termf_4[7:7], termf_6[7:7], termf_4[7:7], cf7__0[6:6], termf_6[7:7], cf7__0[6:6]);
  C3 I492 (fa7_8min_0[0:0], cf7__0[7:7], termf_6[8:8], termf_4[8:8]);
  C3 I493 (fa7_8min_0[1:1], cf7__0[7:7], termf_6[8:8], termt_4[8:8]);
  C3 I494 (fa7_8min_0[2:2], cf7__0[7:7], termt_6[8:8], termf_4[8:8]);
  C3 I495 (fa7_8min_0[3:3], cf7__0[7:7], termt_6[8:8], termt_4[8:8]);
  C3 I496 (fa7_8min_0[4:4], ct7__0[7:7], termf_6[8:8], termf_4[8:8]);
  C3 I497 (fa7_8min_0[5:5], ct7__0[7:7], termf_6[8:8], termt_4[8:8]);
  C3 I498 (fa7_8min_0[6:6], ct7__0[7:7], termt_6[8:8], termf_4[8:8]);
  C3 I499 (fa7_8min_0[7:7], ct7__0[7:7], termt_6[8:8], termt_4[8:8]);
  NOR3 I500 (simp4661_0[0:0], fa7_8min_0[0:0], fa7_8min_0[3:3], fa7_8min_0[5:5]);
  INV I501 (simp4661_0[1:1], fa7_8min_0[6:6]);
  NAND2 I502 (o_0r0[8:8], simp4661_0[0:0], simp4661_0[1:1]);
  NOR3 I503 (simp4671_0[0:0], fa7_8min_0[1:1], fa7_8min_0[2:2], fa7_8min_0[4:4]);
  INV I504 (simp4671_0[1:1], fa7_8min_0[7:7]);
  NAND2 I505 (o_0r1[8:8], simp4671_0[0:0], simp4671_0[1:1]);
  AO222 I506 (ct7__0[8:8], termt_4[8:8], termt_6[8:8], termt_4[8:8], ct7__0[7:7], termt_6[8:8], ct7__0[7:7]);
  AO222 I507 (cf7__0[8:8], termf_4[8:8], termf_6[8:8], termf_4[8:8], cf7__0[7:7], termf_6[8:8], cf7__0[7:7]);
  C3 I508 (fa7_9min_0[0:0], cf7__0[8:8], termf_6[9:9], termf_4[9:9]);
  C3 I509 (fa7_9min_0[1:1], cf7__0[8:8], termf_6[9:9], termt_4[9:9]);
  C3 I510 (fa7_9min_0[2:2], cf7__0[8:8], termt_6[9:9], termf_4[9:9]);
  C3 I511 (fa7_9min_0[3:3], cf7__0[8:8], termt_6[9:9], termt_4[9:9]);
  C3 I512 (fa7_9min_0[4:4], ct7__0[8:8], termf_6[9:9], termf_4[9:9]);
  C3 I513 (fa7_9min_0[5:5], ct7__0[8:8], termf_6[9:9], termt_4[9:9]);
  C3 I514 (fa7_9min_0[6:6], ct7__0[8:8], termt_6[9:9], termf_4[9:9]);
  C3 I515 (fa7_9min_0[7:7], ct7__0[8:8], termt_6[9:9], termt_4[9:9]);
  NOR3 I516 (simp4791_0[0:0], fa7_9min_0[0:0], fa7_9min_0[3:3], fa7_9min_0[5:5]);
  INV I517 (simp4791_0[1:1], fa7_9min_0[6:6]);
  NAND2 I518 (o_0r0[9:9], simp4791_0[0:0], simp4791_0[1:1]);
  NOR3 I519 (simp4801_0[0:0], fa7_9min_0[1:1], fa7_9min_0[2:2], fa7_9min_0[4:4]);
  INV I520 (simp4801_0[1:1], fa7_9min_0[7:7]);
  NAND2 I521 (o_0r1[9:9], simp4801_0[0:0], simp4801_0[1:1]);
  AO222 I522 (ct7__0[9:9], termt_4[9:9], termt_6[9:9], termt_4[9:9], ct7__0[8:8], termt_6[9:9], ct7__0[8:8]);
  AO222 I523 (cf7__0[9:9], termf_4[9:9], termf_6[9:9], termf_4[9:9], cf7__0[8:8], termf_6[9:9], cf7__0[8:8]);
  C3 I524 (fa7_10min_0[0:0], cf7__0[9:9], termf_6[10:10], termf_4[10:10]);
  C3 I525 (fa7_10min_0[1:1], cf7__0[9:9], termf_6[10:10], termt_4[10:10]);
  C3 I526 (fa7_10min_0[2:2], cf7__0[9:9], termt_6[10:10], termf_4[10:10]);
  C3 I527 (fa7_10min_0[3:3], cf7__0[9:9], termt_6[10:10], termt_4[10:10]);
  C3 I528 (fa7_10min_0[4:4], ct7__0[9:9], termf_6[10:10], termf_4[10:10]);
  C3 I529 (fa7_10min_0[5:5], ct7__0[9:9], termf_6[10:10], termt_4[10:10]);
  C3 I530 (fa7_10min_0[6:6], ct7__0[9:9], termt_6[10:10], termf_4[10:10]);
  C3 I531 (fa7_10min_0[7:7], ct7__0[9:9], termt_6[10:10], termt_4[10:10]);
  NOR3 I532 (simp4921_0[0:0], fa7_10min_0[0:0], fa7_10min_0[3:3], fa7_10min_0[5:5]);
  INV I533 (simp4921_0[1:1], fa7_10min_0[6:6]);
  NAND2 I534 (o_0r0[10:10], simp4921_0[0:0], simp4921_0[1:1]);
  NOR3 I535 (simp4931_0[0:0], fa7_10min_0[1:1], fa7_10min_0[2:2], fa7_10min_0[4:4]);
  INV I536 (simp4931_0[1:1], fa7_10min_0[7:7]);
  NAND2 I537 (o_0r1[10:10], simp4931_0[0:0], simp4931_0[1:1]);
  AO222 I538 (ct7__0[10:10], termt_4[10:10], termt_6[10:10], termt_4[10:10], ct7__0[9:9], termt_6[10:10], ct7__0[9:9]);
  AO222 I539 (cf7__0[10:10], termf_4[10:10], termf_6[10:10], termf_4[10:10], cf7__0[9:9], termf_6[10:10], cf7__0[9:9]);
  C3 I540 (fa7_11min_0[0:0], cf7__0[10:10], termf_6[11:11], termf_4[11:11]);
  C3 I541 (fa7_11min_0[1:1], cf7__0[10:10], termf_6[11:11], termt_4[11:11]);
  C3 I542 (fa7_11min_0[2:2], cf7__0[10:10], termt_6[11:11], termf_4[11:11]);
  C3 I543 (fa7_11min_0[3:3], cf7__0[10:10], termt_6[11:11], termt_4[11:11]);
  C3 I544 (fa7_11min_0[4:4], ct7__0[10:10], termf_6[11:11], termf_4[11:11]);
  C3 I545 (fa7_11min_0[5:5], ct7__0[10:10], termf_6[11:11], termt_4[11:11]);
  C3 I546 (fa7_11min_0[6:6], ct7__0[10:10], termt_6[11:11], termf_4[11:11]);
  C3 I547 (fa7_11min_0[7:7], ct7__0[10:10], termt_6[11:11], termt_4[11:11]);
  NOR3 I548 (simp5051_0[0:0], fa7_11min_0[0:0], fa7_11min_0[3:3], fa7_11min_0[5:5]);
  INV I549 (simp5051_0[1:1], fa7_11min_0[6:6]);
  NAND2 I550 (o_0r0[11:11], simp5051_0[0:0], simp5051_0[1:1]);
  NOR3 I551 (simp5061_0[0:0], fa7_11min_0[1:1], fa7_11min_0[2:2], fa7_11min_0[4:4]);
  INV I552 (simp5061_0[1:1], fa7_11min_0[7:7]);
  NAND2 I553 (o_0r1[11:11], simp5061_0[0:0], simp5061_0[1:1]);
  AO222 I554 (ct7__0[11:11], termt_4[11:11], termt_6[11:11], termt_4[11:11], ct7__0[10:10], termt_6[11:11], ct7__0[10:10]);
  AO222 I555 (cf7__0[11:11], termf_4[11:11], termf_6[11:11], termf_4[11:11], cf7__0[10:10], termf_6[11:11], cf7__0[10:10]);
  C3 I556 (fa7_12min_0[0:0], cf7__0[11:11], termf_6[12:12], termf_4[12:12]);
  C3 I557 (fa7_12min_0[1:1], cf7__0[11:11], termf_6[12:12], termt_4[12:12]);
  C3 I558 (fa7_12min_0[2:2], cf7__0[11:11], termt_6[12:12], termf_4[12:12]);
  C3 I559 (fa7_12min_0[3:3], cf7__0[11:11], termt_6[12:12], termt_4[12:12]);
  C3 I560 (fa7_12min_0[4:4], ct7__0[11:11], termf_6[12:12], termf_4[12:12]);
  C3 I561 (fa7_12min_0[5:5], ct7__0[11:11], termf_6[12:12], termt_4[12:12]);
  C3 I562 (fa7_12min_0[6:6], ct7__0[11:11], termt_6[12:12], termf_4[12:12]);
  C3 I563 (fa7_12min_0[7:7], ct7__0[11:11], termt_6[12:12], termt_4[12:12]);
  NOR3 I564 (simp5181_0[0:0], fa7_12min_0[0:0], fa7_12min_0[3:3], fa7_12min_0[5:5]);
  INV I565 (simp5181_0[1:1], fa7_12min_0[6:6]);
  NAND2 I566 (o_0r0[12:12], simp5181_0[0:0], simp5181_0[1:1]);
  NOR3 I567 (simp5191_0[0:0], fa7_12min_0[1:1], fa7_12min_0[2:2], fa7_12min_0[4:4]);
  INV I568 (simp5191_0[1:1], fa7_12min_0[7:7]);
  NAND2 I569 (o_0r1[12:12], simp5191_0[0:0], simp5191_0[1:1]);
  AO222 I570 (ct7__0[12:12], termt_4[12:12], termt_6[12:12], termt_4[12:12], ct7__0[11:11], termt_6[12:12], ct7__0[11:11]);
  AO222 I571 (cf7__0[12:12], termf_4[12:12], termf_6[12:12], termf_4[12:12], cf7__0[11:11], termf_6[12:12], cf7__0[11:11]);
  C3 I572 (fa7_13min_0[0:0], cf7__0[12:12], termf_6[13:13], termf_4[13:13]);
  C3 I573 (fa7_13min_0[1:1], cf7__0[12:12], termf_6[13:13], termt_4[13:13]);
  C3 I574 (fa7_13min_0[2:2], cf7__0[12:12], termt_6[13:13], termf_4[13:13]);
  C3 I575 (fa7_13min_0[3:3], cf7__0[12:12], termt_6[13:13], termt_4[13:13]);
  C3 I576 (fa7_13min_0[4:4], ct7__0[12:12], termf_6[13:13], termf_4[13:13]);
  C3 I577 (fa7_13min_0[5:5], ct7__0[12:12], termf_6[13:13], termt_4[13:13]);
  C3 I578 (fa7_13min_0[6:6], ct7__0[12:12], termt_6[13:13], termf_4[13:13]);
  C3 I579 (fa7_13min_0[7:7], ct7__0[12:12], termt_6[13:13], termt_4[13:13]);
  NOR3 I580 (simp5311_0[0:0], fa7_13min_0[0:0], fa7_13min_0[3:3], fa7_13min_0[5:5]);
  INV I581 (simp5311_0[1:1], fa7_13min_0[6:6]);
  NAND2 I582 (o_0r0[13:13], simp5311_0[0:0], simp5311_0[1:1]);
  NOR3 I583 (simp5321_0[0:0], fa7_13min_0[1:1], fa7_13min_0[2:2], fa7_13min_0[4:4]);
  INV I584 (simp5321_0[1:1], fa7_13min_0[7:7]);
  NAND2 I585 (o_0r1[13:13], simp5321_0[0:0], simp5321_0[1:1]);
  AO222 I586 (ct7__0[13:13], termt_4[13:13], termt_6[13:13], termt_4[13:13], ct7__0[12:12], termt_6[13:13], ct7__0[12:12]);
  AO222 I587 (cf7__0[13:13], termf_4[13:13], termf_6[13:13], termf_4[13:13], cf7__0[12:12], termf_6[13:13], cf7__0[12:12]);
  C3 I588 (fa7_14min_0[0:0], cf7__0[13:13], termf_6[14:14], termf_4[14:14]);
  C3 I589 (fa7_14min_0[1:1], cf7__0[13:13], termf_6[14:14], termt_4[14:14]);
  C3 I590 (fa7_14min_0[2:2], cf7__0[13:13], termt_6[14:14], termf_4[14:14]);
  C3 I591 (fa7_14min_0[3:3], cf7__0[13:13], termt_6[14:14], termt_4[14:14]);
  C3 I592 (fa7_14min_0[4:4], ct7__0[13:13], termf_6[14:14], termf_4[14:14]);
  C3 I593 (fa7_14min_0[5:5], ct7__0[13:13], termf_6[14:14], termt_4[14:14]);
  C3 I594 (fa7_14min_0[6:6], ct7__0[13:13], termt_6[14:14], termf_4[14:14]);
  C3 I595 (fa7_14min_0[7:7], ct7__0[13:13], termt_6[14:14], termt_4[14:14]);
  NOR3 I596 (simp5441_0[0:0], fa7_14min_0[0:0], fa7_14min_0[3:3], fa7_14min_0[5:5]);
  INV I597 (simp5441_0[1:1], fa7_14min_0[6:6]);
  NAND2 I598 (o_0r0[14:14], simp5441_0[0:0], simp5441_0[1:1]);
  NOR3 I599 (simp5451_0[0:0], fa7_14min_0[1:1], fa7_14min_0[2:2], fa7_14min_0[4:4]);
  INV I600 (simp5451_0[1:1], fa7_14min_0[7:7]);
  NAND2 I601 (o_0r1[14:14], simp5451_0[0:0], simp5451_0[1:1]);
  AO222 I602 (ct7__0[14:14], termt_4[14:14], termt_6[14:14], termt_4[14:14], ct7__0[13:13], termt_6[14:14], ct7__0[13:13]);
  AO222 I603 (cf7__0[14:14], termf_4[14:14], termf_6[14:14], termf_4[14:14], cf7__0[13:13], termf_6[14:14], cf7__0[13:13]);
  C3 I604 (fa7_15min_0[0:0], cf7__0[14:14], termf_6[15:15], termf_4[15:15]);
  C3 I605 (fa7_15min_0[1:1], cf7__0[14:14], termf_6[15:15], termt_4[15:15]);
  C3 I606 (fa7_15min_0[2:2], cf7__0[14:14], termt_6[15:15], termf_4[15:15]);
  C3 I607 (fa7_15min_0[3:3], cf7__0[14:14], termt_6[15:15], termt_4[15:15]);
  C3 I608 (fa7_15min_0[4:4], ct7__0[14:14], termf_6[15:15], termf_4[15:15]);
  C3 I609 (fa7_15min_0[5:5], ct7__0[14:14], termf_6[15:15], termt_4[15:15]);
  C3 I610 (fa7_15min_0[6:6], ct7__0[14:14], termt_6[15:15], termf_4[15:15]);
  C3 I611 (fa7_15min_0[7:7], ct7__0[14:14], termt_6[15:15], termt_4[15:15]);
  NOR3 I612 (simp5571_0[0:0], fa7_15min_0[0:0], fa7_15min_0[3:3], fa7_15min_0[5:5]);
  INV I613 (simp5571_0[1:1], fa7_15min_0[6:6]);
  NAND2 I614 (o_0r0[15:15], simp5571_0[0:0], simp5571_0[1:1]);
  NOR3 I615 (simp5581_0[0:0], fa7_15min_0[1:1], fa7_15min_0[2:2], fa7_15min_0[4:4]);
  INV I616 (simp5581_0[1:1], fa7_15min_0[7:7]);
  NAND2 I617 (o_0r1[15:15], simp5581_0[0:0], simp5581_0[1:1]);
  AO222 I618 (ct7__0[15:15], termt_4[15:15], termt_6[15:15], termt_4[15:15], ct7__0[14:14], termt_6[15:15], ct7__0[14:14]);
  AO222 I619 (cf7__0[15:15], termf_4[15:15], termf_6[15:15], termf_4[15:15], cf7__0[14:14], termf_6[15:15], cf7__0[14:14]);
  C3 I620 (fa7_16min_0[0:0], cf7__0[15:15], termf_6[16:16], termf_4[16:16]);
  C3 I621 (fa7_16min_0[1:1], cf7__0[15:15], termf_6[16:16], termt_4[16:16]);
  C3 I622 (fa7_16min_0[2:2], cf7__0[15:15], termt_6[16:16], termf_4[16:16]);
  C3 I623 (fa7_16min_0[3:3], cf7__0[15:15], termt_6[16:16], termt_4[16:16]);
  C3 I624 (fa7_16min_0[4:4], ct7__0[15:15], termf_6[16:16], termf_4[16:16]);
  C3 I625 (fa7_16min_0[5:5], ct7__0[15:15], termf_6[16:16], termt_4[16:16]);
  C3 I626 (fa7_16min_0[6:6], ct7__0[15:15], termt_6[16:16], termf_4[16:16]);
  C3 I627 (fa7_16min_0[7:7], ct7__0[15:15], termt_6[16:16], termt_4[16:16]);
  NOR3 I628 (simp5701_0[0:0], fa7_16min_0[0:0], fa7_16min_0[3:3], fa7_16min_0[5:5]);
  INV I629 (simp5701_0[1:1], fa7_16min_0[6:6]);
  NAND2 I630 (o_0r0[16:16], simp5701_0[0:0], simp5701_0[1:1]);
  NOR3 I631 (simp5711_0[0:0], fa7_16min_0[1:1], fa7_16min_0[2:2], fa7_16min_0[4:4]);
  INV I632 (simp5711_0[1:1], fa7_16min_0[7:7]);
  NAND2 I633 (o_0r1[16:16], simp5711_0[0:0], simp5711_0[1:1]);
  AO222 I634 (ct7__0[16:16], termt_4[16:16], termt_6[16:16], termt_4[16:16], ct7__0[15:15], termt_6[16:16], ct7__0[15:15]);
  AO222 I635 (cf7__0[16:16], termf_4[16:16], termf_6[16:16], termf_4[16:16], cf7__0[15:15], termf_6[16:16], cf7__0[15:15]);
  C3 I636 (fa7_17min_0[0:0], cf7__0[16:16], termf_6[17:17], termf_4[17:17]);
  C3 I637 (fa7_17min_0[1:1], cf7__0[16:16], termf_6[17:17], termt_4[17:17]);
  C3 I638 (fa7_17min_0[2:2], cf7__0[16:16], termt_6[17:17], termf_4[17:17]);
  C3 I639 (fa7_17min_0[3:3], cf7__0[16:16], termt_6[17:17], termt_4[17:17]);
  C3 I640 (fa7_17min_0[4:4], ct7__0[16:16], termf_6[17:17], termf_4[17:17]);
  C3 I641 (fa7_17min_0[5:5], ct7__0[16:16], termf_6[17:17], termt_4[17:17]);
  C3 I642 (fa7_17min_0[6:6], ct7__0[16:16], termt_6[17:17], termf_4[17:17]);
  C3 I643 (fa7_17min_0[7:7], ct7__0[16:16], termt_6[17:17], termt_4[17:17]);
  NOR3 I644 (simp5831_0[0:0], fa7_17min_0[0:0], fa7_17min_0[3:3], fa7_17min_0[5:5]);
  INV I645 (simp5831_0[1:1], fa7_17min_0[6:6]);
  NAND2 I646 (o_0r0[17:17], simp5831_0[0:0], simp5831_0[1:1]);
  NOR3 I647 (simp5841_0[0:0], fa7_17min_0[1:1], fa7_17min_0[2:2], fa7_17min_0[4:4]);
  INV I648 (simp5841_0[1:1], fa7_17min_0[7:7]);
  NAND2 I649 (o_0r1[17:17], simp5841_0[0:0], simp5841_0[1:1]);
  AO222 I650 (ct7__0[17:17], termt_4[17:17], termt_6[17:17], termt_4[17:17], ct7__0[16:16], termt_6[17:17], ct7__0[16:16]);
  AO222 I651 (cf7__0[17:17], termf_4[17:17], termf_6[17:17], termf_4[17:17], cf7__0[16:16], termf_6[17:17], cf7__0[16:16]);
  C3 I652 (fa7_18min_0[0:0], cf7__0[17:17], termf_6[18:18], termf_4[18:18]);
  C3 I653 (fa7_18min_0[1:1], cf7__0[17:17], termf_6[18:18], termt_4[18:18]);
  C3 I654 (fa7_18min_0[2:2], cf7__0[17:17], termt_6[18:18], termf_4[18:18]);
  C3 I655 (fa7_18min_0[3:3], cf7__0[17:17], termt_6[18:18], termt_4[18:18]);
  C3 I656 (fa7_18min_0[4:4], ct7__0[17:17], termf_6[18:18], termf_4[18:18]);
  C3 I657 (fa7_18min_0[5:5], ct7__0[17:17], termf_6[18:18], termt_4[18:18]);
  C3 I658 (fa7_18min_0[6:6], ct7__0[17:17], termt_6[18:18], termf_4[18:18]);
  C3 I659 (fa7_18min_0[7:7], ct7__0[17:17], termt_6[18:18], termt_4[18:18]);
  NOR3 I660 (simp5961_0[0:0], fa7_18min_0[0:0], fa7_18min_0[3:3], fa7_18min_0[5:5]);
  INV I661 (simp5961_0[1:1], fa7_18min_0[6:6]);
  NAND2 I662 (o_0r0[18:18], simp5961_0[0:0], simp5961_0[1:1]);
  NOR3 I663 (simp5971_0[0:0], fa7_18min_0[1:1], fa7_18min_0[2:2], fa7_18min_0[4:4]);
  INV I664 (simp5971_0[1:1], fa7_18min_0[7:7]);
  NAND2 I665 (o_0r1[18:18], simp5971_0[0:0], simp5971_0[1:1]);
  AO222 I666 (ct7__0[18:18], termt_4[18:18], termt_6[18:18], termt_4[18:18], ct7__0[17:17], termt_6[18:18], ct7__0[17:17]);
  AO222 I667 (cf7__0[18:18], termf_4[18:18], termf_6[18:18], termf_4[18:18], cf7__0[17:17], termf_6[18:18], cf7__0[17:17]);
  C3 I668 (fa7_19min_0[0:0], cf7__0[18:18], termf_6[19:19], termf_4[19:19]);
  C3 I669 (fa7_19min_0[1:1], cf7__0[18:18], termf_6[19:19], termt_4[19:19]);
  C3 I670 (fa7_19min_0[2:2], cf7__0[18:18], termt_6[19:19], termf_4[19:19]);
  C3 I671 (fa7_19min_0[3:3], cf7__0[18:18], termt_6[19:19], termt_4[19:19]);
  C3 I672 (fa7_19min_0[4:4], ct7__0[18:18], termf_6[19:19], termf_4[19:19]);
  C3 I673 (fa7_19min_0[5:5], ct7__0[18:18], termf_6[19:19], termt_4[19:19]);
  C3 I674 (fa7_19min_0[6:6], ct7__0[18:18], termt_6[19:19], termf_4[19:19]);
  C3 I675 (fa7_19min_0[7:7], ct7__0[18:18], termt_6[19:19], termt_4[19:19]);
  NOR3 I676 (simp6091_0[0:0], fa7_19min_0[0:0], fa7_19min_0[3:3], fa7_19min_0[5:5]);
  INV I677 (simp6091_0[1:1], fa7_19min_0[6:6]);
  NAND2 I678 (o_0r0[19:19], simp6091_0[0:0], simp6091_0[1:1]);
  NOR3 I679 (simp6101_0[0:0], fa7_19min_0[1:1], fa7_19min_0[2:2], fa7_19min_0[4:4]);
  INV I680 (simp6101_0[1:1], fa7_19min_0[7:7]);
  NAND2 I681 (o_0r1[19:19], simp6101_0[0:0], simp6101_0[1:1]);
  AO222 I682 (ct7__0[19:19], termt_4[19:19], termt_6[19:19], termt_4[19:19], ct7__0[18:18], termt_6[19:19], ct7__0[18:18]);
  AO222 I683 (cf7__0[19:19], termf_4[19:19], termf_6[19:19], termf_4[19:19], cf7__0[18:18], termf_6[19:19], cf7__0[18:18]);
  C3 I684 (fa7_20min_0[0:0], cf7__0[19:19], termf_6[20:20], termf_4[20:20]);
  C3 I685 (fa7_20min_0[1:1], cf7__0[19:19], termf_6[20:20], termt_4[20:20]);
  C3 I686 (fa7_20min_0[2:2], cf7__0[19:19], termt_6[20:20], termf_4[20:20]);
  C3 I687 (fa7_20min_0[3:3], cf7__0[19:19], termt_6[20:20], termt_4[20:20]);
  C3 I688 (fa7_20min_0[4:4], ct7__0[19:19], termf_6[20:20], termf_4[20:20]);
  C3 I689 (fa7_20min_0[5:5], ct7__0[19:19], termf_6[20:20], termt_4[20:20]);
  C3 I690 (fa7_20min_0[6:6], ct7__0[19:19], termt_6[20:20], termf_4[20:20]);
  C3 I691 (fa7_20min_0[7:7], ct7__0[19:19], termt_6[20:20], termt_4[20:20]);
  NOR3 I692 (simp6221_0[0:0], fa7_20min_0[0:0], fa7_20min_0[3:3], fa7_20min_0[5:5]);
  INV I693 (simp6221_0[1:1], fa7_20min_0[6:6]);
  NAND2 I694 (o_0r0[20:20], simp6221_0[0:0], simp6221_0[1:1]);
  NOR3 I695 (simp6231_0[0:0], fa7_20min_0[1:1], fa7_20min_0[2:2], fa7_20min_0[4:4]);
  INV I696 (simp6231_0[1:1], fa7_20min_0[7:7]);
  NAND2 I697 (o_0r1[20:20], simp6231_0[0:0], simp6231_0[1:1]);
  AO222 I698 (ct7__0[20:20], termt_4[20:20], termt_6[20:20], termt_4[20:20], ct7__0[19:19], termt_6[20:20], ct7__0[19:19]);
  AO222 I699 (cf7__0[20:20], termf_4[20:20], termf_6[20:20], termf_4[20:20], cf7__0[19:19], termf_6[20:20], cf7__0[19:19]);
  C3 I700 (fa7_21min_0[0:0], cf7__0[20:20], termf_6[21:21], termf_4[21:21]);
  C3 I701 (fa7_21min_0[1:1], cf7__0[20:20], termf_6[21:21], termt_4[21:21]);
  C3 I702 (fa7_21min_0[2:2], cf7__0[20:20], termt_6[21:21], termf_4[21:21]);
  C3 I703 (fa7_21min_0[3:3], cf7__0[20:20], termt_6[21:21], termt_4[21:21]);
  C3 I704 (fa7_21min_0[4:4], ct7__0[20:20], termf_6[21:21], termf_4[21:21]);
  C3 I705 (fa7_21min_0[5:5], ct7__0[20:20], termf_6[21:21], termt_4[21:21]);
  C3 I706 (fa7_21min_0[6:6], ct7__0[20:20], termt_6[21:21], termf_4[21:21]);
  C3 I707 (fa7_21min_0[7:7], ct7__0[20:20], termt_6[21:21], termt_4[21:21]);
  NOR3 I708 (simp6351_0[0:0], fa7_21min_0[0:0], fa7_21min_0[3:3], fa7_21min_0[5:5]);
  INV I709 (simp6351_0[1:1], fa7_21min_0[6:6]);
  NAND2 I710 (o_0r0[21:21], simp6351_0[0:0], simp6351_0[1:1]);
  NOR3 I711 (simp6361_0[0:0], fa7_21min_0[1:1], fa7_21min_0[2:2], fa7_21min_0[4:4]);
  INV I712 (simp6361_0[1:1], fa7_21min_0[7:7]);
  NAND2 I713 (o_0r1[21:21], simp6361_0[0:0], simp6361_0[1:1]);
  AO222 I714 (ct7__0[21:21], termt_4[21:21], termt_6[21:21], termt_4[21:21], ct7__0[20:20], termt_6[21:21], ct7__0[20:20]);
  AO222 I715 (cf7__0[21:21], termf_4[21:21], termf_6[21:21], termf_4[21:21], cf7__0[20:20], termf_6[21:21], cf7__0[20:20]);
  C3 I716 (fa7_22min_0[0:0], cf7__0[21:21], termf_6[22:22], termf_4[22:22]);
  C3 I717 (fa7_22min_0[1:1], cf7__0[21:21], termf_6[22:22], termt_4[22:22]);
  C3 I718 (fa7_22min_0[2:2], cf7__0[21:21], termt_6[22:22], termf_4[22:22]);
  C3 I719 (fa7_22min_0[3:3], cf7__0[21:21], termt_6[22:22], termt_4[22:22]);
  C3 I720 (fa7_22min_0[4:4], ct7__0[21:21], termf_6[22:22], termf_4[22:22]);
  C3 I721 (fa7_22min_0[5:5], ct7__0[21:21], termf_6[22:22], termt_4[22:22]);
  C3 I722 (fa7_22min_0[6:6], ct7__0[21:21], termt_6[22:22], termf_4[22:22]);
  C3 I723 (fa7_22min_0[7:7], ct7__0[21:21], termt_6[22:22], termt_4[22:22]);
  NOR3 I724 (simp6481_0[0:0], fa7_22min_0[0:0], fa7_22min_0[3:3], fa7_22min_0[5:5]);
  INV I725 (simp6481_0[1:1], fa7_22min_0[6:6]);
  NAND2 I726 (o_0r0[22:22], simp6481_0[0:0], simp6481_0[1:1]);
  NOR3 I727 (simp6491_0[0:0], fa7_22min_0[1:1], fa7_22min_0[2:2], fa7_22min_0[4:4]);
  INV I728 (simp6491_0[1:1], fa7_22min_0[7:7]);
  NAND2 I729 (o_0r1[22:22], simp6491_0[0:0], simp6491_0[1:1]);
  AO222 I730 (ct7__0[22:22], termt_4[22:22], termt_6[22:22], termt_4[22:22], ct7__0[21:21], termt_6[22:22], ct7__0[21:21]);
  AO222 I731 (cf7__0[22:22], termf_4[22:22], termf_6[22:22], termf_4[22:22], cf7__0[21:21], termf_6[22:22], cf7__0[21:21]);
  C3 I732 (fa7_23min_0[0:0], cf7__0[22:22], termf_6[23:23], termf_4[23:23]);
  C3 I733 (fa7_23min_0[1:1], cf7__0[22:22], termf_6[23:23], termt_4[23:23]);
  C3 I734 (fa7_23min_0[2:2], cf7__0[22:22], termt_6[23:23], termf_4[23:23]);
  C3 I735 (fa7_23min_0[3:3], cf7__0[22:22], termt_6[23:23], termt_4[23:23]);
  C3 I736 (fa7_23min_0[4:4], ct7__0[22:22], termf_6[23:23], termf_4[23:23]);
  C3 I737 (fa7_23min_0[5:5], ct7__0[22:22], termf_6[23:23], termt_4[23:23]);
  C3 I738 (fa7_23min_0[6:6], ct7__0[22:22], termt_6[23:23], termf_4[23:23]);
  C3 I739 (fa7_23min_0[7:7], ct7__0[22:22], termt_6[23:23], termt_4[23:23]);
  NOR3 I740 (simp6611_0[0:0], fa7_23min_0[0:0], fa7_23min_0[3:3], fa7_23min_0[5:5]);
  INV I741 (simp6611_0[1:1], fa7_23min_0[6:6]);
  NAND2 I742 (o_0r0[23:23], simp6611_0[0:0], simp6611_0[1:1]);
  NOR3 I743 (simp6621_0[0:0], fa7_23min_0[1:1], fa7_23min_0[2:2], fa7_23min_0[4:4]);
  INV I744 (simp6621_0[1:1], fa7_23min_0[7:7]);
  NAND2 I745 (o_0r1[23:23], simp6621_0[0:0], simp6621_0[1:1]);
  AO222 I746 (ct7__0[23:23], termt_4[23:23], termt_6[23:23], termt_4[23:23], ct7__0[22:22], termt_6[23:23], ct7__0[22:22]);
  AO222 I747 (cf7__0[23:23], termf_4[23:23], termf_6[23:23], termf_4[23:23], cf7__0[22:22], termf_6[23:23], cf7__0[22:22]);
  C3 I748 (fa7_24min_0[0:0], cf7__0[23:23], termf_6[24:24], termf_4[24:24]);
  C3 I749 (fa7_24min_0[1:1], cf7__0[23:23], termf_6[24:24], termt_4[24:24]);
  C3 I750 (fa7_24min_0[2:2], cf7__0[23:23], termt_6[24:24], termf_4[24:24]);
  C3 I751 (fa7_24min_0[3:3], cf7__0[23:23], termt_6[24:24], termt_4[24:24]);
  C3 I752 (fa7_24min_0[4:4], ct7__0[23:23], termf_6[24:24], termf_4[24:24]);
  C3 I753 (fa7_24min_0[5:5], ct7__0[23:23], termf_6[24:24], termt_4[24:24]);
  C3 I754 (fa7_24min_0[6:6], ct7__0[23:23], termt_6[24:24], termf_4[24:24]);
  C3 I755 (fa7_24min_0[7:7], ct7__0[23:23], termt_6[24:24], termt_4[24:24]);
  NOR3 I756 (simp6741_0[0:0], fa7_24min_0[0:0], fa7_24min_0[3:3], fa7_24min_0[5:5]);
  INV I757 (simp6741_0[1:1], fa7_24min_0[6:6]);
  NAND2 I758 (o_0r0[24:24], simp6741_0[0:0], simp6741_0[1:1]);
  NOR3 I759 (simp6751_0[0:0], fa7_24min_0[1:1], fa7_24min_0[2:2], fa7_24min_0[4:4]);
  INV I760 (simp6751_0[1:1], fa7_24min_0[7:7]);
  NAND2 I761 (o_0r1[24:24], simp6751_0[0:0], simp6751_0[1:1]);
  AO222 I762 (ct7__0[24:24], termt_4[24:24], termt_6[24:24], termt_4[24:24], ct7__0[23:23], termt_6[24:24], ct7__0[23:23]);
  AO222 I763 (cf7__0[24:24], termf_4[24:24], termf_6[24:24], termf_4[24:24], cf7__0[23:23], termf_6[24:24], cf7__0[23:23]);
  C3 I764 (fa7_25min_0[0:0], cf7__0[24:24], termf_6[25:25], termf_4[25:25]);
  C3 I765 (fa7_25min_0[1:1], cf7__0[24:24], termf_6[25:25], termt_4[25:25]);
  C3 I766 (fa7_25min_0[2:2], cf7__0[24:24], termt_6[25:25], termf_4[25:25]);
  C3 I767 (fa7_25min_0[3:3], cf7__0[24:24], termt_6[25:25], termt_4[25:25]);
  C3 I768 (fa7_25min_0[4:4], ct7__0[24:24], termf_6[25:25], termf_4[25:25]);
  C3 I769 (fa7_25min_0[5:5], ct7__0[24:24], termf_6[25:25], termt_4[25:25]);
  C3 I770 (fa7_25min_0[6:6], ct7__0[24:24], termt_6[25:25], termf_4[25:25]);
  C3 I771 (fa7_25min_0[7:7], ct7__0[24:24], termt_6[25:25], termt_4[25:25]);
  NOR3 I772 (simp6871_0[0:0], fa7_25min_0[0:0], fa7_25min_0[3:3], fa7_25min_0[5:5]);
  INV I773 (simp6871_0[1:1], fa7_25min_0[6:6]);
  NAND2 I774 (o_0r0[25:25], simp6871_0[0:0], simp6871_0[1:1]);
  NOR3 I775 (simp6881_0[0:0], fa7_25min_0[1:1], fa7_25min_0[2:2], fa7_25min_0[4:4]);
  INV I776 (simp6881_0[1:1], fa7_25min_0[7:7]);
  NAND2 I777 (o_0r1[25:25], simp6881_0[0:0], simp6881_0[1:1]);
  AO222 I778 (ct7__0[25:25], termt_4[25:25], termt_6[25:25], termt_4[25:25], ct7__0[24:24], termt_6[25:25], ct7__0[24:24]);
  AO222 I779 (cf7__0[25:25], termf_4[25:25], termf_6[25:25], termf_4[25:25], cf7__0[24:24], termf_6[25:25], cf7__0[24:24]);
  C3 I780 (fa7_26min_0[0:0], cf7__0[25:25], termf_6[26:26], termf_4[26:26]);
  C3 I781 (fa7_26min_0[1:1], cf7__0[25:25], termf_6[26:26], termt_4[26:26]);
  C3 I782 (fa7_26min_0[2:2], cf7__0[25:25], termt_6[26:26], termf_4[26:26]);
  C3 I783 (fa7_26min_0[3:3], cf7__0[25:25], termt_6[26:26], termt_4[26:26]);
  C3 I784 (fa7_26min_0[4:4], ct7__0[25:25], termf_6[26:26], termf_4[26:26]);
  C3 I785 (fa7_26min_0[5:5], ct7__0[25:25], termf_6[26:26], termt_4[26:26]);
  C3 I786 (fa7_26min_0[6:6], ct7__0[25:25], termt_6[26:26], termf_4[26:26]);
  C3 I787 (fa7_26min_0[7:7], ct7__0[25:25], termt_6[26:26], termt_4[26:26]);
  NOR3 I788 (simp7001_0[0:0], fa7_26min_0[0:0], fa7_26min_0[3:3], fa7_26min_0[5:5]);
  INV I789 (simp7001_0[1:1], fa7_26min_0[6:6]);
  NAND2 I790 (o_0r0[26:26], simp7001_0[0:0], simp7001_0[1:1]);
  NOR3 I791 (simp7011_0[0:0], fa7_26min_0[1:1], fa7_26min_0[2:2], fa7_26min_0[4:4]);
  INV I792 (simp7011_0[1:1], fa7_26min_0[7:7]);
  NAND2 I793 (o_0r1[26:26], simp7011_0[0:0], simp7011_0[1:1]);
  AO222 I794 (ct7__0[26:26], termt_4[26:26], termt_6[26:26], termt_4[26:26], ct7__0[25:25], termt_6[26:26], ct7__0[25:25]);
  AO222 I795 (cf7__0[26:26], termf_4[26:26], termf_6[26:26], termf_4[26:26], cf7__0[25:25], termf_6[26:26], cf7__0[25:25]);
  C3 I796 (fa7_27min_0[0:0], cf7__0[26:26], termf_6[27:27], termf_4[27:27]);
  C3 I797 (fa7_27min_0[1:1], cf7__0[26:26], termf_6[27:27], termt_4[27:27]);
  C3 I798 (fa7_27min_0[2:2], cf7__0[26:26], termt_6[27:27], termf_4[27:27]);
  C3 I799 (fa7_27min_0[3:3], cf7__0[26:26], termt_6[27:27], termt_4[27:27]);
  C3 I800 (fa7_27min_0[4:4], ct7__0[26:26], termf_6[27:27], termf_4[27:27]);
  C3 I801 (fa7_27min_0[5:5], ct7__0[26:26], termf_6[27:27], termt_4[27:27]);
  C3 I802 (fa7_27min_0[6:6], ct7__0[26:26], termt_6[27:27], termf_4[27:27]);
  C3 I803 (fa7_27min_0[7:7], ct7__0[26:26], termt_6[27:27], termt_4[27:27]);
  NOR3 I804 (simp7131_0[0:0], fa7_27min_0[0:0], fa7_27min_0[3:3], fa7_27min_0[5:5]);
  INV I805 (simp7131_0[1:1], fa7_27min_0[6:6]);
  NAND2 I806 (o_0r0[27:27], simp7131_0[0:0], simp7131_0[1:1]);
  NOR3 I807 (simp7141_0[0:0], fa7_27min_0[1:1], fa7_27min_0[2:2], fa7_27min_0[4:4]);
  INV I808 (simp7141_0[1:1], fa7_27min_0[7:7]);
  NAND2 I809 (o_0r1[27:27], simp7141_0[0:0], simp7141_0[1:1]);
  AO222 I810 (ct7__0[27:27], termt_4[27:27], termt_6[27:27], termt_4[27:27], ct7__0[26:26], termt_6[27:27], ct7__0[26:26]);
  AO222 I811 (cf7__0[27:27], termf_4[27:27], termf_6[27:27], termf_4[27:27], cf7__0[26:26], termf_6[27:27], cf7__0[26:26]);
  C3 I812 (fa7_28min_0[0:0], cf7__0[27:27], termf_6[28:28], termf_4[28:28]);
  C3 I813 (fa7_28min_0[1:1], cf7__0[27:27], termf_6[28:28], termt_4[28:28]);
  C3 I814 (fa7_28min_0[2:2], cf7__0[27:27], termt_6[28:28], termf_4[28:28]);
  C3 I815 (fa7_28min_0[3:3], cf7__0[27:27], termt_6[28:28], termt_4[28:28]);
  C3 I816 (fa7_28min_0[4:4], ct7__0[27:27], termf_6[28:28], termf_4[28:28]);
  C3 I817 (fa7_28min_0[5:5], ct7__0[27:27], termf_6[28:28], termt_4[28:28]);
  C3 I818 (fa7_28min_0[6:6], ct7__0[27:27], termt_6[28:28], termf_4[28:28]);
  C3 I819 (fa7_28min_0[7:7], ct7__0[27:27], termt_6[28:28], termt_4[28:28]);
  NOR3 I820 (simp7261_0[0:0], fa7_28min_0[0:0], fa7_28min_0[3:3], fa7_28min_0[5:5]);
  INV I821 (simp7261_0[1:1], fa7_28min_0[6:6]);
  NAND2 I822 (o_0r0[28:28], simp7261_0[0:0], simp7261_0[1:1]);
  NOR3 I823 (simp7271_0[0:0], fa7_28min_0[1:1], fa7_28min_0[2:2], fa7_28min_0[4:4]);
  INV I824 (simp7271_0[1:1], fa7_28min_0[7:7]);
  NAND2 I825 (o_0r1[28:28], simp7271_0[0:0], simp7271_0[1:1]);
  AO222 I826 (ct7__0[28:28], termt_4[28:28], termt_6[28:28], termt_4[28:28], ct7__0[27:27], termt_6[28:28], ct7__0[27:27]);
  AO222 I827 (cf7__0[28:28], termf_4[28:28], termf_6[28:28], termf_4[28:28], cf7__0[27:27], termf_6[28:28], cf7__0[27:27]);
  C3 I828 (fa7_29min_0[0:0], cf7__0[28:28], termf_6[29:29], termf_4[29:29]);
  C3 I829 (fa7_29min_0[1:1], cf7__0[28:28], termf_6[29:29], termt_4[29:29]);
  C3 I830 (fa7_29min_0[2:2], cf7__0[28:28], termt_6[29:29], termf_4[29:29]);
  C3 I831 (fa7_29min_0[3:3], cf7__0[28:28], termt_6[29:29], termt_4[29:29]);
  C3 I832 (fa7_29min_0[4:4], ct7__0[28:28], termf_6[29:29], termf_4[29:29]);
  C3 I833 (fa7_29min_0[5:5], ct7__0[28:28], termf_6[29:29], termt_4[29:29]);
  C3 I834 (fa7_29min_0[6:6], ct7__0[28:28], termt_6[29:29], termf_4[29:29]);
  C3 I835 (fa7_29min_0[7:7], ct7__0[28:28], termt_6[29:29], termt_4[29:29]);
  NOR3 I836 (simp7391_0[0:0], fa7_29min_0[0:0], fa7_29min_0[3:3], fa7_29min_0[5:5]);
  INV I837 (simp7391_0[1:1], fa7_29min_0[6:6]);
  NAND2 I838 (o_0r0[29:29], simp7391_0[0:0], simp7391_0[1:1]);
  NOR3 I839 (simp7401_0[0:0], fa7_29min_0[1:1], fa7_29min_0[2:2], fa7_29min_0[4:4]);
  INV I840 (simp7401_0[1:1], fa7_29min_0[7:7]);
  NAND2 I841 (o_0r1[29:29], simp7401_0[0:0], simp7401_0[1:1]);
  AO222 I842 (ct7__0[29:29], termt_4[29:29], termt_6[29:29], termt_4[29:29], ct7__0[28:28], termt_6[29:29], ct7__0[28:28]);
  AO222 I843 (cf7__0[29:29], termf_4[29:29], termf_6[29:29], termf_4[29:29], cf7__0[28:28], termf_6[29:29], cf7__0[28:28]);
  C3 I844 (fa7_30min_0[0:0], cf7__0[29:29], termf_6[30:30], termf_4[30:30]);
  C3 I845 (fa7_30min_0[1:1], cf7__0[29:29], termf_6[30:30], termt_4[30:30]);
  C3 I846 (fa7_30min_0[2:2], cf7__0[29:29], termt_6[30:30], termf_4[30:30]);
  C3 I847 (fa7_30min_0[3:3], cf7__0[29:29], termt_6[30:30], termt_4[30:30]);
  C3 I848 (fa7_30min_0[4:4], ct7__0[29:29], termf_6[30:30], termf_4[30:30]);
  C3 I849 (fa7_30min_0[5:5], ct7__0[29:29], termf_6[30:30], termt_4[30:30]);
  C3 I850 (fa7_30min_0[6:6], ct7__0[29:29], termt_6[30:30], termf_4[30:30]);
  C3 I851 (fa7_30min_0[7:7], ct7__0[29:29], termt_6[30:30], termt_4[30:30]);
  NOR3 I852 (simp7521_0[0:0], fa7_30min_0[0:0], fa7_30min_0[3:3], fa7_30min_0[5:5]);
  INV I853 (simp7521_0[1:1], fa7_30min_0[6:6]);
  NAND2 I854 (o_0r0[30:30], simp7521_0[0:0], simp7521_0[1:1]);
  NOR3 I855 (simp7531_0[0:0], fa7_30min_0[1:1], fa7_30min_0[2:2], fa7_30min_0[4:4]);
  INV I856 (simp7531_0[1:1], fa7_30min_0[7:7]);
  NAND2 I857 (o_0r1[30:30], simp7531_0[0:0], simp7531_0[1:1]);
  AO222 I858 (ct7__0[30:30], termt_4[30:30], termt_6[30:30], termt_4[30:30], ct7__0[29:29], termt_6[30:30], ct7__0[29:29]);
  AO222 I859 (cf7__0[30:30], termf_4[30:30], termf_6[30:30], termf_4[30:30], cf7__0[29:29], termf_6[30:30], cf7__0[29:29]);
  C3 I860 (fa7_31min_0[0:0], cf7__0[30:30], termf_6[31:31], termf_4[31:31]);
  C3 I861 (fa7_31min_0[1:1], cf7__0[30:30], termf_6[31:31], termt_4[31:31]);
  C3 I862 (fa7_31min_0[2:2], cf7__0[30:30], termt_6[31:31], termf_4[31:31]);
  C3 I863 (fa7_31min_0[3:3], cf7__0[30:30], termt_6[31:31], termt_4[31:31]);
  C3 I864 (fa7_31min_0[4:4], ct7__0[30:30], termf_6[31:31], termf_4[31:31]);
  C3 I865 (fa7_31min_0[5:5], ct7__0[30:30], termf_6[31:31], termt_4[31:31]);
  C3 I866 (fa7_31min_0[6:6], ct7__0[30:30], termt_6[31:31], termf_4[31:31]);
  C3 I867 (fa7_31min_0[7:7], ct7__0[30:30], termt_6[31:31], termt_4[31:31]);
  NOR3 I868 (simp7651_0[0:0], fa7_31min_0[0:0], fa7_31min_0[3:3], fa7_31min_0[5:5]);
  INV I869 (simp7651_0[1:1], fa7_31min_0[6:6]);
  NAND2 I870 (o_0r0[31:31], simp7651_0[0:0], simp7651_0[1:1]);
  NOR3 I871 (simp7661_0[0:0], fa7_31min_0[1:1], fa7_31min_0[2:2], fa7_31min_0[4:4]);
  INV I872 (simp7661_0[1:1], fa7_31min_0[7:7]);
  NAND2 I873 (o_0r1[31:31], simp7661_0[0:0], simp7661_0[1:1]);
  AO222 I874 (ct7__0[31:31], termt_4[31:31], termt_6[31:31], termt_4[31:31], ct7__0[30:30], termt_6[31:31], ct7__0[30:30]);
  AO222 I875 (cf7__0[31:31], termf_4[31:31], termf_6[31:31], termf_4[31:31], cf7__0[30:30], termf_6[31:31], cf7__0[30:30]);
  C3 I876 (fa7_32min_0[0:0], cf7__0[31:31], termf_6[32:32], termf_4[32:32]);
  C3 I877 (fa7_32min_0[1:1], cf7__0[31:31], termf_6[32:32], termt_4[32:32]);
  C3 I878 (fa7_32min_0[2:2], cf7__0[31:31], termt_6[32:32], termf_4[32:32]);
  C3 I879 (fa7_32min_0[3:3], cf7__0[31:31], termt_6[32:32], termt_4[32:32]);
  C3 I880 (fa7_32min_0[4:4], ct7__0[31:31], termf_6[32:32], termf_4[32:32]);
  C3 I881 (fa7_32min_0[5:5], ct7__0[31:31], termf_6[32:32], termt_4[32:32]);
  C3 I882 (fa7_32min_0[6:6], ct7__0[31:31], termt_6[32:32], termf_4[32:32]);
  C3 I883 (fa7_32min_0[7:7], ct7__0[31:31], termt_6[32:32], termt_4[32:32]);
  NOR3 I884 (simp7781_0[0:0], fa7_32min_0[0:0], fa7_32min_0[3:3], fa7_32min_0[5:5]);
  INV I885 (simp7781_0[1:1], fa7_32min_0[6:6]);
  NAND2 I886 (o_0r0[32:32], simp7781_0[0:0], simp7781_0[1:1]);
  NOR3 I887 (simp7791_0[0:0], fa7_32min_0[1:1], fa7_32min_0[2:2], fa7_32min_0[4:4]);
  INV I888 (simp7791_0[1:1], fa7_32min_0[7:7]);
  NAND2 I889 (o_0r1[32:32], simp7791_0[0:0], simp7791_0[1:1]);
  AO222 I890 (ct7__0[32:32], termt_4[32:32], termt_6[32:32], termt_4[32:32], ct7__0[31:31], termt_6[32:32], ct7__0[31:31]);
  AO222 I891 (cf7__0[32:32], termf_4[32:32], termf_6[32:32], termf_4[32:32], cf7__0[31:31], termf_6[32:32], cf7__0[31:31]);
  C3 I892 (fa7_33min_0[0:0], cf7__0[32:32], termf_6[33:33], termf_4[33:33]);
  C3 I893 (fa7_33min_0[1:1], cf7__0[32:32], termf_6[33:33], termt_4[33:33]);
  C3 I894 (fa7_33min_0[2:2], cf7__0[32:32], termt_6[33:33], termf_4[33:33]);
  C3 I895 (fa7_33min_0[3:3], cf7__0[32:32], termt_6[33:33], termt_4[33:33]);
  C3 I896 (fa7_33min_0[4:4], ct7__0[32:32], termf_6[33:33], termf_4[33:33]);
  C3 I897 (fa7_33min_0[5:5], ct7__0[32:32], termf_6[33:33], termt_4[33:33]);
  C3 I898 (fa7_33min_0[6:6], ct7__0[32:32], termt_6[33:33], termf_4[33:33]);
  C3 I899 (fa7_33min_0[7:7], ct7__0[32:32], termt_6[33:33], termt_4[33:33]);
  NOR3 I900 (simp7911_0[0:0], fa7_33min_0[0:0], fa7_33min_0[3:3], fa7_33min_0[5:5]);
  INV I901 (simp7911_0[1:1], fa7_33min_0[6:6]);
  NAND2 I902 (o_0r0[33:33], simp7911_0[0:0], simp7911_0[1:1]);
  NOR3 I903 (simp7921_0[0:0], fa7_33min_0[1:1], fa7_33min_0[2:2], fa7_33min_0[4:4]);
  INV I904 (simp7921_0[1:1], fa7_33min_0[7:7]);
  NAND2 I905 (o_0r1[33:33], simp7921_0[0:0], simp7921_0[1:1]);
  AO222 I906 (ct7__0[33:33], termt_4[33:33], termt_6[33:33], termt_4[33:33], ct7__0[32:32], termt_6[33:33], ct7__0[32:32]);
  AO222 I907 (cf7__0[33:33], termf_4[33:33], termf_6[33:33], termf_4[33:33], cf7__0[32:32], termf_6[33:33], cf7__0[32:32]);
  BUFF I908 (i_0a, o_0a);
endmodule

// tkf34mo1w33 TeakF [1] [One 34,Many [33]]
module tkf34mo1w33 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [33:0] i_0r0;
  input [33:0] i_0r1;
  output i_0a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  wire ucomplete_0;
  wire comp_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (comp_0, i_0r0[0:0], i_0r1[0:0]);
  BUFF I2 (ucomplete_0, comp_0);
  C2 I3 (acomplete_0, ucomplete_0, icomplete_0);
  C2 I4 (o_0r0[0:0], i_0r0[1:1], icomplete_0);
  BUFF I5 (o_0r0[1:1], i_0r0[2:2]);
  BUFF I6 (o_0r0[2:2], i_0r0[3:3]);
  BUFF I7 (o_0r0[3:3], i_0r0[4:4]);
  BUFF I8 (o_0r0[4:4], i_0r0[5:5]);
  BUFF I9 (o_0r0[5:5], i_0r0[6:6]);
  BUFF I10 (o_0r0[6:6], i_0r0[7:7]);
  BUFF I11 (o_0r0[7:7], i_0r0[8:8]);
  BUFF I12 (o_0r0[8:8], i_0r0[9:9]);
  BUFF I13 (o_0r0[9:9], i_0r0[10:10]);
  BUFF I14 (o_0r0[10:10], i_0r0[11:11]);
  BUFF I15 (o_0r0[11:11], i_0r0[12:12]);
  BUFF I16 (o_0r0[12:12], i_0r0[13:13]);
  BUFF I17 (o_0r0[13:13], i_0r0[14:14]);
  BUFF I18 (o_0r0[14:14], i_0r0[15:15]);
  BUFF I19 (o_0r0[15:15], i_0r0[16:16]);
  BUFF I20 (o_0r0[16:16], i_0r0[17:17]);
  BUFF I21 (o_0r0[17:17], i_0r0[18:18]);
  BUFF I22 (o_0r0[18:18], i_0r0[19:19]);
  BUFF I23 (o_0r0[19:19], i_0r0[20:20]);
  BUFF I24 (o_0r0[20:20], i_0r0[21:21]);
  BUFF I25 (o_0r0[21:21], i_0r0[22:22]);
  BUFF I26 (o_0r0[22:22], i_0r0[23:23]);
  BUFF I27 (o_0r0[23:23], i_0r0[24:24]);
  BUFF I28 (o_0r0[24:24], i_0r0[25:25]);
  BUFF I29 (o_0r0[25:25], i_0r0[26:26]);
  BUFF I30 (o_0r0[26:26], i_0r0[27:27]);
  BUFF I31 (o_0r0[27:27], i_0r0[28:28]);
  BUFF I32 (o_0r0[28:28], i_0r0[29:29]);
  BUFF I33 (o_0r0[29:29], i_0r0[30:30]);
  BUFF I34 (o_0r0[30:30], i_0r0[31:31]);
  BUFF I35 (o_0r0[31:31], i_0r0[32:32]);
  BUFF I36 (o_0r0[32:32], i_0r0[33:33]);
  C2 I37 (o_0r1[0:0], i_0r1[1:1], icomplete_0);
  BUFF I38 (o_0r1[1:1], i_0r1[2:2]);
  BUFF I39 (o_0r1[2:2], i_0r1[3:3]);
  BUFF I40 (o_0r1[3:3], i_0r1[4:4]);
  BUFF I41 (o_0r1[4:4], i_0r1[5:5]);
  BUFF I42 (o_0r1[5:5], i_0r1[6:6]);
  BUFF I43 (o_0r1[6:6], i_0r1[7:7]);
  BUFF I44 (o_0r1[7:7], i_0r1[8:8]);
  BUFF I45 (o_0r1[8:8], i_0r1[9:9]);
  BUFF I46 (o_0r1[9:9], i_0r1[10:10]);
  BUFF I47 (o_0r1[10:10], i_0r1[11:11]);
  BUFF I48 (o_0r1[11:11], i_0r1[12:12]);
  BUFF I49 (o_0r1[12:12], i_0r1[13:13]);
  BUFF I50 (o_0r1[13:13], i_0r1[14:14]);
  BUFF I51 (o_0r1[14:14], i_0r1[15:15]);
  BUFF I52 (o_0r1[15:15], i_0r1[16:16]);
  BUFF I53 (o_0r1[16:16], i_0r1[17:17]);
  BUFF I54 (o_0r1[17:17], i_0r1[18:18]);
  BUFF I55 (o_0r1[18:18], i_0r1[19:19]);
  BUFF I56 (o_0r1[19:19], i_0r1[20:20]);
  BUFF I57 (o_0r1[20:20], i_0r1[21:21]);
  BUFF I58 (o_0r1[21:21], i_0r1[22:22]);
  BUFF I59 (o_0r1[22:22], i_0r1[23:23]);
  BUFF I60 (o_0r1[23:23], i_0r1[24:24]);
  BUFF I61 (o_0r1[24:24], i_0r1[25:25]);
  BUFF I62 (o_0r1[25:25], i_0r1[26:26]);
  BUFF I63 (o_0r1[26:26], i_0r1[27:27]);
  BUFF I64 (o_0r1[27:27], i_0r1[28:28]);
  BUFF I65 (o_0r1[28:28], i_0r1[29:29]);
  BUFF I66 (o_0r1[29:29], i_0r1[30:30]);
  BUFF I67 (o_0r1[30:30], i_0r1[31:31]);
  BUFF I68 (o_0r1[31:31], i_0r1[32:32]);
  BUFF I69 (o_0r1[32:32], i_0r1[33:33]);
  C2 I70 (i_0a, acomplete_0, o_0a);
endmodule

// tkf0mo0w0_o0w0_o0w0_o0w0 TeakF [0,0,0,0] [One 0,Many [0,0,0,0]]
module tkf0mo0w0_o0w0_o0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  input reset;
  wire [1:0] simp11_0;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  BUFF I2 (o_2r, i_0r);
  BUFF I3 (o_3r, i_0r);
  C3 I4 (simp11_0[0:0], o_0a, o_1a, o_2a);
  BUFF I5 (simp11_0[1:1], o_3a);
  C2 I6 (i_0a, simp11_0[0:0], simp11_0[1:1]);
endmodule

// tkj64m32_32 TeakJ [Many [32,32],One 64]
module tkj64m32_32 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  output [63:0] o_0r0;
  output [63:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [63:0] joinf_0;
  wire [63:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joinf_0[32:32], i_1r0[0:0]);
  BUFF I33 (joinf_0[33:33], i_1r0[1:1]);
  BUFF I34 (joinf_0[34:34], i_1r0[2:2]);
  BUFF I35 (joinf_0[35:35], i_1r0[3:3]);
  BUFF I36 (joinf_0[36:36], i_1r0[4:4]);
  BUFF I37 (joinf_0[37:37], i_1r0[5:5]);
  BUFF I38 (joinf_0[38:38], i_1r0[6:6]);
  BUFF I39 (joinf_0[39:39], i_1r0[7:7]);
  BUFF I40 (joinf_0[40:40], i_1r0[8:8]);
  BUFF I41 (joinf_0[41:41], i_1r0[9:9]);
  BUFF I42 (joinf_0[42:42], i_1r0[10:10]);
  BUFF I43 (joinf_0[43:43], i_1r0[11:11]);
  BUFF I44 (joinf_0[44:44], i_1r0[12:12]);
  BUFF I45 (joinf_0[45:45], i_1r0[13:13]);
  BUFF I46 (joinf_0[46:46], i_1r0[14:14]);
  BUFF I47 (joinf_0[47:47], i_1r0[15:15]);
  BUFF I48 (joinf_0[48:48], i_1r0[16:16]);
  BUFF I49 (joinf_0[49:49], i_1r0[17:17]);
  BUFF I50 (joinf_0[50:50], i_1r0[18:18]);
  BUFF I51 (joinf_0[51:51], i_1r0[19:19]);
  BUFF I52 (joinf_0[52:52], i_1r0[20:20]);
  BUFF I53 (joinf_0[53:53], i_1r0[21:21]);
  BUFF I54 (joinf_0[54:54], i_1r0[22:22]);
  BUFF I55 (joinf_0[55:55], i_1r0[23:23]);
  BUFF I56 (joinf_0[56:56], i_1r0[24:24]);
  BUFF I57 (joinf_0[57:57], i_1r0[25:25]);
  BUFF I58 (joinf_0[58:58], i_1r0[26:26]);
  BUFF I59 (joinf_0[59:59], i_1r0[27:27]);
  BUFF I60 (joinf_0[60:60], i_1r0[28:28]);
  BUFF I61 (joinf_0[61:61], i_1r0[29:29]);
  BUFF I62 (joinf_0[62:62], i_1r0[30:30]);
  BUFF I63 (joinf_0[63:63], i_1r0[31:31]);
  BUFF I64 (joint_0[0:0], i_0r1[0:0]);
  BUFF I65 (joint_0[1:1], i_0r1[1:1]);
  BUFF I66 (joint_0[2:2], i_0r1[2:2]);
  BUFF I67 (joint_0[3:3], i_0r1[3:3]);
  BUFF I68 (joint_0[4:4], i_0r1[4:4]);
  BUFF I69 (joint_0[5:5], i_0r1[5:5]);
  BUFF I70 (joint_0[6:6], i_0r1[6:6]);
  BUFF I71 (joint_0[7:7], i_0r1[7:7]);
  BUFF I72 (joint_0[8:8], i_0r1[8:8]);
  BUFF I73 (joint_0[9:9], i_0r1[9:9]);
  BUFF I74 (joint_0[10:10], i_0r1[10:10]);
  BUFF I75 (joint_0[11:11], i_0r1[11:11]);
  BUFF I76 (joint_0[12:12], i_0r1[12:12]);
  BUFF I77 (joint_0[13:13], i_0r1[13:13]);
  BUFF I78 (joint_0[14:14], i_0r1[14:14]);
  BUFF I79 (joint_0[15:15], i_0r1[15:15]);
  BUFF I80 (joint_0[16:16], i_0r1[16:16]);
  BUFF I81 (joint_0[17:17], i_0r1[17:17]);
  BUFF I82 (joint_0[18:18], i_0r1[18:18]);
  BUFF I83 (joint_0[19:19], i_0r1[19:19]);
  BUFF I84 (joint_0[20:20], i_0r1[20:20]);
  BUFF I85 (joint_0[21:21], i_0r1[21:21]);
  BUFF I86 (joint_0[22:22], i_0r1[22:22]);
  BUFF I87 (joint_0[23:23], i_0r1[23:23]);
  BUFF I88 (joint_0[24:24], i_0r1[24:24]);
  BUFF I89 (joint_0[25:25], i_0r1[25:25]);
  BUFF I90 (joint_0[26:26], i_0r1[26:26]);
  BUFF I91 (joint_0[27:27], i_0r1[27:27]);
  BUFF I92 (joint_0[28:28], i_0r1[28:28]);
  BUFF I93 (joint_0[29:29], i_0r1[29:29]);
  BUFF I94 (joint_0[30:30], i_0r1[30:30]);
  BUFF I95 (joint_0[31:31], i_0r1[31:31]);
  BUFF I96 (joint_0[32:32], i_1r1[0:0]);
  BUFF I97 (joint_0[33:33], i_1r1[1:1]);
  BUFF I98 (joint_0[34:34], i_1r1[2:2]);
  BUFF I99 (joint_0[35:35], i_1r1[3:3]);
  BUFF I100 (joint_0[36:36], i_1r1[4:4]);
  BUFF I101 (joint_0[37:37], i_1r1[5:5]);
  BUFF I102 (joint_0[38:38], i_1r1[6:6]);
  BUFF I103 (joint_0[39:39], i_1r1[7:7]);
  BUFF I104 (joint_0[40:40], i_1r1[8:8]);
  BUFF I105 (joint_0[41:41], i_1r1[9:9]);
  BUFF I106 (joint_0[42:42], i_1r1[10:10]);
  BUFF I107 (joint_0[43:43], i_1r1[11:11]);
  BUFF I108 (joint_0[44:44], i_1r1[12:12]);
  BUFF I109 (joint_0[45:45], i_1r1[13:13]);
  BUFF I110 (joint_0[46:46], i_1r1[14:14]);
  BUFF I111 (joint_0[47:47], i_1r1[15:15]);
  BUFF I112 (joint_0[48:48], i_1r1[16:16]);
  BUFF I113 (joint_0[49:49], i_1r1[17:17]);
  BUFF I114 (joint_0[50:50], i_1r1[18:18]);
  BUFF I115 (joint_0[51:51], i_1r1[19:19]);
  BUFF I116 (joint_0[52:52], i_1r1[20:20]);
  BUFF I117 (joint_0[53:53], i_1r1[21:21]);
  BUFF I118 (joint_0[54:54], i_1r1[22:22]);
  BUFF I119 (joint_0[55:55], i_1r1[23:23]);
  BUFF I120 (joint_0[56:56], i_1r1[24:24]);
  BUFF I121 (joint_0[57:57], i_1r1[25:25]);
  BUFF I122 (joint_0[58:58], i_1r1[26:26]);
  BUFF I123 (joint_0[59:59], i_1r1[27:27]);
  BUFF I124 (joint_0[60:60], i_1r1[28:28]);
  BUFF I125 (joint_0[61:61], i_1r1[29:29]);
  BUFF I126 (joint_0[62:62], i_1r1[30:30]);
  BUFF I127 (joint_0[63:63], i_1r1[31:31]);
  OR2 I128 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I129 (icomplete_0, dcomplete_0);
  C2 I130 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I131 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I132 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I133 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I134 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I135 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I136 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I137 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I138 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I139 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I140 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I141 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I142 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I143 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I144 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I145 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I146 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I147 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I148 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I149 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I150 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I151 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I152 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I153 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I154 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I155 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I156 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I157 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I158 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I159 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I160 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I161 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I162 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I163 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I164 (o_0r0[33:33], joinf_0[33:33]);
  BUFF I165 (o_0r0[34:34], joinf_0[34:34]);
  BUFF I166 (o_0r0[35:35], joinf_0[35:35]);
  BUFF I167 (o_0r0[36:36], joinf_0[36:36]);
  BUFF I168 (o_0r0[37:37], joinf_0[37:37]);
  BUFF I169 (o_0r0[38:38], joinf_0[38:38]);
  BUFF I170 (o_0r0[39:39], joinf_0[39:39]);
  BUFF I171 (o_0r0[40:40], joinf_0[40:40]);
  BUFF I172 (o_0r0[41:41], joinf_0[41:41]);
  BUFF I173 (o_0r0[42:42], joinf_0[42:42]);
  BUFF I174 (o_0r0[43:43], joinf_0[43:43]);
  BUFF I175 (o_0r0[44:44], joinf_0[44:44]);
  BUFF I176 (o_0r0[45:45], joinf_0[45:45]);
  BUFF I177 (o_0r0[46:46], joinf_0[46:46]);
  BUFF I178 (o_0r0[47:47], joinf_0[47:47]);
  BUFF I179 (o_0r0[48:48], joinf_0[48:48]);
  BUFF I180 (o_0r0[49:49], joinf_0[49:49]);
  BUFF I181 (o_0r0[50:50], joinf_0[50:50]);
  BUFF I182 (o_0r0[51:51], joinf_0[51:51]);
  BUFF I183 (o_0r0[52:52], joinf_0[52:52]);
  BUFF I184 (o_0r0[53:53], joinf_0[53:53]);
  BUFF I185 (o_0r0[54:54], joinf_0[54:54]);
  BUFF I186 (o_0r0[55:55], joinf_0[55:55]);
  BUFF I187 (o_0r0[56:56], joinf_0[56:56]);
  BUFF I188 (o_0r0[57:57], joinf_0[57:57]);
  BUFF I189 (o_0r0[58:58], joinf_0[58:58]);
  BUFF I190 (o_0r0[59:59], joinf_0[59:59]);
  BUFF I191 (o_0r0[60:60], joinf_0[60:60]);
  BUFF I192 (o_0r0[61:61], joinf_0[61:61]);
  BUFF I193 (o_0r0[62:62], joinf_0[62:62]);
  BUFF I194 (o_0r0[63:63], joinf_0[63:63]);
  BUFF I195 (o_0r1[1:1], joint_0[1:1]);
  BUFF I196 (o_0r1[2:2], joint_0[2:2]);
  BUFF I197 (o_0r1[3:3], joint_0[3:3]);
  BUFF I198 (o_0r1[4:4], joint_0[4:4]);
  BUFF I199 (o_0r1[5:5], joint_0[5:5]);
  BUFF I200 (o_0r1[6:6], joint_0[6:6]);
  BUFF I201 (o_0r1[7:7], joint_0[7:7]);
  BUFF I202 (o_0r1[8:8], joint_0[8:8]);
  BUFF I203 (o_0r1[9:9], joint_0[9:9]);
  BUFF I204 (o_0r1[10:10], joint_0[10:10]);
  BUFF I205 (o_0r1[11:11], joint_0[11:11]);
  BUFF I206 (o_0r1[12:12], joint_0[12:12]);
  BUFF I207 (o_0r1[13:13], joint_0[13:13]);
  BUFF I208 (o_0r1[14:14], joint_0[14:14]);
  BUFF I209 (o_0r1[15:15], joint_0[15:15]);
  BUFF I210 (o_0r1[16:16], joint_0[16:16]);
  BUFF I211 (o_0r1[17:17], joint_0[17:17]);
  BUFF I212 (o_0r1[18:18], joint_0[18:18]);
  BUFF I213 (o_0r1[19:19], joint_0[19:19]);
  BUFF I214 (o_0r1[20:20], joint_0[20:20]);
  BUFF I215 (o_0r1[21:21], joint_0[21:21]);
  BUFF I216 (o_0r1[22:22], joint_0[22:22]);
  BUFF I217 (o_0r1[23:23], joint_0[23:23]);
  BUFF I218 (o_0r1[24:24], joint_0[24:24]);
  BUFF I219 (o_0r1[25:25], joint_0[25:25]);
  BUFF I220 (o_0r1[26:26], joint_0[26:26]);
  BUFF I221 (o_0r1[27:27], joint_0[27:27]);
  BUFF I222 (o_0r1[28:28], joint_0[28:28]);
  BUFF I223 (o_0r1[29:29], joint_0[29:29]);
  BUFF I224 (o_0r1[30:30], joint_0[30:30]);
  BUFF I225 (o_0r1[31:31], joint_0[31:31]);
  BUFF I226 (o_0r1[32:32], joint_0[32:32]);
  BUFF I227 (o_0r1[33:33], joint_0[33:33]);
  BUFF I228 (o_0r1[34:34], joint_0[34:34]);
  BUFF I229 (o_0r1[35:35], joint_0[35:35]);
  BUFF I230 (o_0r1[36:36], joint_0[36:36]);
  BUFF I231 (o_0r1[37:37], joint_0[37:37]);
  BUFF I232 (o_0r1[38:38], joint_0[38:38]);
  BUFF I233 (o_0r1[39:39], joint_0[39:39]);
  BUFF I234 (o_0r1[40:40], joint_0[40:40]);
  BUFF I235 (o_0r1[41:41], joint_0[41:41]);
  BUFF I236 (o_0r1[42:42], joint_0[42:42]);
  BUFF I237 (o_0r1[43:43], joint_0[43:43]);
  BUFF I238 (o_0r1[44:44], joint_0[44:44]);
  BUFF I239 (o_0r1[45:45], joint_0[45:45]);
  BUFF I240 (o_0r1[46:46], joint_0[46:46]);
  BUFF I241 (o_0r1[47:47], joint_0[47:47]);
  BUFF I242 (o_0r1[48:48], joint_0[48:48]);
  BUFF I243 (o_0r1[49:49], joint_0[49:49]);
  BUFF I244 (o_0r1[50:50], joint_0[50:50]);
  BUFF I245 (o_0r1[51:51], joint_0[51:51]);
  BUFF I246 (o_0r1[52:52], joint_0[52:52]);
  BUFF I247 (o_0r1[53:53], joint_0[53:53]);
  BUFF I248 (o_0r1[54:54], joint_0[54:54]);
  BUFF I249 (o_0r1[55:55], joint_0[55:55]);
  BUFF I250 (o_0r1[56:56], joint_0[56:56]);
  BUFF I251 (o_0r1[57:57], joint_0[57:57]);
  BUFF I252 (o_0r1[58:58], joint_0[58:58]);
  BUFF I253 (o_0r1[59:59], joint_0[59:59]);
  BUFF I254 (o_0r1[60:60], joint_0[60:60]);
  BUFF I255 (o_0r1[61:61], joint_0[61:61]);
  BUFF I256 (o_0r1[62:62], joint_0[62:62]);
  BUFF I257 (o_0r1[63:63], joint_0[63:63]);
  BUFF I258 (i_0a, o_0a);
  BUFF I259 (i_1a, o_0a);
endmodule

// tko64m32_1api0w32b_2api32w32b_3andt1o0w32bt2o0w32b TeakO [
//     (1,TeakOAppend 1 [(0,0+:32)]),
//     (2,TeakOAppend 1 [(0,32+:32)]),
//     (3,TeakOp TeakOpAnd [(1,0+:32),(2,0+:32)])] [One 64,One 32]
module tko64m32_1api0w32b_2api32w32b_3andt1o0w32bt2o0w32b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [63:0] i_0r0;
  input [63:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire [31:0] termf_1;
  wire [31:0] termf_2;
  wire [31:0] termt_1;
  wire [31:0] termt_2;
  wire [3:0] op3_0_0;
  wire [3:0] op3_1_0;
  wire [3:0] op3_2_0;
  wire [3:0] op3_3_0;
  wire [3:0] op3_4_0;
  wire [3:0] op3_5_0;
  wire [3:0] op3_6_0;
  wire [3:0] op3_7_0;
  wire [3:0] op3_8_0;
  wire [3:0] op3_9_0;
  wire [3:0] op3_10_0;
  wire [3:0] op3_11_0;
  wire [3:0] op3_12_0;
  wire [3:0] op3_13_0;
  wire [3:0] op3_14_0;
  wire [3:0] op3_15_0;
  wire [3:0] op3_16_0;
  wire [3:0] op3_17_0;
  wire [3:0] op3_18_0;
  wire [3:0] op3_19_0;
  wire [3:0] op3_20_0;
  wire [3:0] op3_21_0;
  wire [3:0] op3_22_0;
  wire [3:0] op3_23_0;
  wire [3:0] op3_24_0;
  wire [3:0] op3_25_0;
  wire [3:0] op3_26_0;
  wire [3:0] op3_27_0;
  wire [3:0] op3_28_0;
  wire [3:0] op3_29_0;
  wire [3:0] op3_30_0;
  wire [3:0] op3_31_0;
  BUFF I0 (termf_1[0:0], i_0r0[0:0]);
  BUFF I1 (termf_1[1:1], i_0r0[1:1]);
  BUFF I2 (termf_1[2:2], i_0r0[2:2]);
  BUFF I3 (termf_1[3:3], i_0r0[3:3]);
  BUFF I4 (termf_1[4:4], i_0r0[4:4]);
  BUFF I5 (termf_1[5:5], i_0r0[5:5]);
  BUFF I6 (termf_1[6:6], i_0r0[6:6]);
  BUFF I7 (termf_1[7:7], i_0r0[7:7]);
  BUFF I8 (termf_1[8:8], i_0r0[8:8]);
  BUFF I9 (termf_1[9:9], i_0r0[9:9]);
  BUFF I10 (termf_1[10:10], i_0r0[10:10]);
  BUFF I11 (termf_1[11:11], i_0r0[11:11]);
  BUFF I12 (termf_1[12:12], i_0r0[12:12]);
  BUFF I13 (termf_1[13:13], i_0r0[13:13]);
  BUFF I14 (termf_1[14:14], i_0r0[14:14]);
  BUFF I15 (termf_1[15:15], i_0r0[15:15]);
  BUFF I16 (termf_1[16:16], i_0r0[16:16]);
  BUFF I17 (termf_1[17:17], i_0r0[17:17]);
  BUFF I18 (termf_1[18:18], i_0r0[18:18]);
  BUFF I19 (termf_1[19:19], i_0r0[19:19]);
  BUFF I20 (termf_1[20:20], i_0r0[20:20]);
  BUFF I21 (termf_1[21:21], i_0r0[21:21]);
  BUFF I22 (termf_1[22:22], i_0r0[22:22]);
  BUFF I23 (termf_1[23:23], i_0r0[23:23]);
  BUFF I24 (termf_1[24:24], i_0r0[24:24]);
  BUFF I25 (termf_1[25:25], i_0r0[25:25]);
  BUFF I26 (termf_1[26:26], i_0r0[26:26]);
  BUFF I27 (termf_1[27:27], i_0r0[27:27]);
  BUFF I28 (termf_1[28:28], i_0r0[28:28]);
  BUFF I29 (termf_1[29:29], i_0r0[29:29]);
  BUFF I30 (termf_1[30:30], i_0r0[30:30]);
  BUFF I31 (termf_1[31:31], i_0r0[31:31]);
  BUFF I32 (termt_1[0:0], i_0r1[0:0]);
  BUFF I33 (termt_1[1:1], i_0r1[1:1]);
  BUFF I34 (termt_1[2:2], i_0r1[2:2]);
  BUFF I35 (termt_1[3:3], i_0r1[3:3]);
  BUFF I36 (termt_1[4:4], i_0r1[4:4]);
  BUFF I37 (termt_1[5:5], i_0r1[5:5]);
  BUFF I38 (termt_1[6:6], i_0r1[6:6]);
  BUFF I39 (termt_1[7:7], i_0r1[7:7]);
  BUFF I40 (termt_1[8:8], i_0r1[8:8]);
  BUFF I41 (termt_1[9:9], i_0r1[9:9]);
  BUFF I42 (termt_1[10:10], i_0r1[10:10]);
  BUFF I43 (termt_1[11:11], i_0r1[11:11]);
  BUFF I44 (termt_1[12:12], i_0r1[12:12]);
  BUFF I45 (termt_1[13:13], i_0r1[13:13]);
  BUFF I46 (termt_1[14:14], i_0r1[14:14]);
  BUFF I47 (termt_1[15:15], i_0r1[15:15]);
  BUFF I48 (termt_1[16:16], i_0r1[16:16]);
  BUFF I49 (termt_1[17:17], i_0r1[17:17]);
  BUFF I50 (termt_1[18:18], i_0r1[18:18]);
  BUFF I51 (termt_1[19:19], i_0r1[19:19]);
  BUFF I52 (termt_1[20:20], i_0r1[20:20]);
  BUFF I53 (termt_1[21:21], i_0r1[21:21]);
  BUFF I54 (termt_1[22:22], i_0r1[22:22]);
  BUFF I55 (termt_1[23:23], i_0r1[23:23]);
  BUFF I56 (termt_1[24:24], i_0r1[24:24]);
  BUFF I57 (termt_1[25:25], i_0r1[25:25]);
  BUFF I58 (termt_1[26:26], i_0r1[26:26]);
  BUFF I59 (termt_1[27:27], i_0r1[27:27]);
  BUFF I60 (termt_1[28:28], i_0r1[28:28]);
  BUFF I61 (termt_1[29:29], i_0r1[29:29]);
  BUFF I62 (termt_1[30:30], i_0r1[30:30]);
  BUFF I63 (termt_1[31:31], i_0r1[31:31]);
  BUFF I64 (termf_2[0:0], i_0r0[32:32]);
  BUFF I65 (termf_2[1:1], i_0r0[33:33]);
  BUFF I66 (termf_2[2:2], i_0r0[34:34]);
  BUFF I67 (termf_2[3:3], i_0r0[35:35]);
  BUFF I68 (termf_2[4:4], i_0r0[36:36]);
  BUFF I69 (termf_2[5:5], i_0r0[37:37]);
  BUFF I70 (termf_2[6:6], i_0r0[38:38]);
  BUFF I71 (termf_2[7:7], i_0r0[39:39]);
  BUFF I72 (termf_2[8:8], i_0r0[40:40]);
  BUFF I73 (termf_2[9:9], i_0r0[41:41]);
  BUFF I74 (termf_2[10:10], i_0r0[42:42]);
  BUFF I75 (termf_2[11:11], i_0r0[43:43]);
  BUFF I76 (termf_2[12:12], i_0r0[44:44]);
  BUFF I77 (termf_2[13:13], i_0r0[45:45]);
  BUFF I78 (termf_2[14:14], i_0r0[46:46]);
  BUFF I79 (termf_2[15:15], i_0r0[47:47]);
  BUFF I80 (termf_2[16:16], i_0r0[48:48]);
  BUFF I81 (termf_2[17:17], i_0r0[49:49]);
  BUFF I82 (termf_2[18:18], i_0r0[50:50]);
  BUFF I83 (termf_2[19:19], i_0r0[51:51]);
  BUFF I84 (termf_2[20:20], i_0r0[52:52]);
  BUFF I85 (termf_2[21:21], i_0r0[53:53]);
  BUFF I86 (termf_2[22:22], i_0r0[54:54]);
  BUFF I87 (termf_2[23:23], i_0r0[55:55]);
  BUFF I88 (termf_2[24:24], i_0r0[56:56]);
  BUFF I89 (termf_2[25:25], i_0r0[57:57]);
  BUFF I90 (termf_2[26:26], i_0r0[58:58]);
  BUFF I91 (termf_2[27:27], i_0r0[59:59]);
  BUFF I92 (termf_2[28:28], i_0r0[60:60]);
  BUFF I93 (termf_2[29:29], i_0r0[61:61]);
  BUFF I94 (termf_2[30:30], i_0r0[62:62]);
  BUFF I95 (termf_2[31:31], i_0r0[63:63]);
  BUFF I96 (termt_2[0:0], i_0r1[32:32]);
  BUFF I97 (termt_2[1:1], i_0r1[33:33]);
  BUFF I98 (termt_2[2:2], i_0r1[34:34]);
  BUFF I99 (termt_2[3:3], i_0r1[35:35]);
  BUFF I100 (termt_2[4:4], i_0r1[36:36]);
  BUFF I101 (termt_2[5:5], i_0r1[37:37]);
  BUFF I102 (termt_2[6:6], i_0r1[38:38]);
  BUFF I103 (termt_2[7:7], i_0r1[39:39]);
  BUFF I104 (termt_2[8:8], i_0r1[40:40]);
  BUFF I105 (termt_2[9:9], i_0r1[41:41]);
  BUFF I106 (termt_2[10:10], i_0r1[42:42]);
  BUFF I107 (termt_2[11:11], i_0r1[43:43]);
  BUFF I108 (termt_2[12:12], i_0r1[44:44]);
  BUFF I109 (termt_2[13:13], i_0r1[45:45]);
  BUFF I110 (termt_2[14:14], i_0r1[46:46]);
  BUFF I111 (termt_2[15:15], i_0r1[47:47]);
  BUFF I112 (termt_2[16:16], i_0r1[48:48]);
  BUFF I113 (termt_2[17:17], i_0r1[49:49]);
  BUFF I114 (termt_2[18:18], i_0r1[50:50]);
  BUFF I115 (termt_2[19:19], i_0r1[51:51]);
  BUFF I116 (termt_2[20:20], i_0r1[52:52]);
  BUFF I117 (termt_2[21:21], i_0r1[53:53]);
  BUFF I118 (termt_2[22:22], i_0r1[54:54]);
  BUFF I119 (termt_2[23:23], i_0r1[55:55]);
  BUFF I120 (termt_2[24:24], i_0r1[56:56]);
  BUFF I121 (termt_2[25:25], i_0r1[57:57]);
  BUFF I122 (termt_2[26:26], i_0r1[58:58]);
  BUFF I123 (termt_2[27:27], i_0r1[59:59]);
  BUFF I124 (termt_2[28:28], i_0r1[60:60]);
  BUFF I125 (termt_2[29:29], i_0r1[61:61]);
  BUFF I126 (termt_2[30:30], i_0r1[62:62]);
  BUFF I127 (termt_2[31:31], i_0r1[63:63]);
  C2 I128 (op3_0_0[0:0], termf_2[0:0], termf_1[0:0]);
  C2 I129 (op3_0_0[1:1], termf_2[0:0], termt_1[0:0]);
  C2 I130 (op3_0_0[2:2], termt_2[0:0], termf_1[0:0]);
  C2 I131 (op3_0_0[3:3], termt_2[0:0], termt_1[0:0]);
  OR3 I132 (o_0r0[0:0], op3_0_0[0:0], op3_0_0[1:1], op3_0_0[2:2]);
  BUFF I133 (o_0r1[0:0], op3_0_0[3:3]);
  C2 I134 (op3_1_0[0:0], termf_2[1:1], termf_1[1:1]);
  C2 I135 (op3_1_0[1:1], termf_2[1:1], termt_1[1:1]);
  C2 I136 (op3_1_0[2:2], termt_2[1:1], termf_1[1:1]);
  C2 I137 (op3_1_0[3:3], termt_2[1:1], termt_1[1:1]);
  OR3 I138 (o_0r0[1:1], op3_1_0[0:0], op3_1_0[1:1], op3_1_0[2:2]);
  BUFF I139 (o_0r1[1:1], op3_1_0[3:3]);
  C2 I140 (op3_2_0[0:0], termf_2[2:2], termf_1[2:2]);
  C2 I141 (op3_2_0[1:1], termf_2[2:2], termt_1[2:2]);
  C2 I142 (op3_2_0[2:2], termt_2[2:2], termf_1[2:2]);
  C2 I143 (op3_2_0[3:3], termt_2[2:2], termt_1[2:2]);
  OR3 I144 (o_0r0[2:2], op3_2_0[0:0], op3_2_0[1:1], op3_2_0[2:2]);
  BUFF I145 (o_0r1[2:2], op3_2_0[3:3]);
  C2 I146 (op3_3_0[0:0], termf_2[3:3], termf_1[3:3]);
  C2 I147 (op3_3_0[1:1], termf_2[3:3], termt_1[3:3]);
  C2 I148 (op3_3_0[2:2], termt_2[3:3], termf_1[3:3]);
  C2 I149 (op3_3_0[3:3], termt_2[3:3], termt_1[3:3]);
  OR3 I150 (o_0r0[3:3], op3_3_0[0:0], op3_3_0[1:1], op3_3_0[2:2]);
  BUFF I151 (o_0r1[3:3], op3_3_0[3:3]);
  C2 I152 (op3_4_0[0:0], termf_2[4:4], termf_1[4:4]);
  C2 I153 (op3_4_0[1:1], termf_2[4:4], termt_1[4:4]);
  C2 I154 (op3_4_0[2:2], termt_2[4:4], termf_1[4:4]);
  C2 I155 (op3_4_0[3:3], termt_2[4:4], termt_1[4:4]);
  OR3 I156 (o_0r0[4:4], op3_4_0[0:0], op3_4_0[1:1], op3_4_0[2:2]);
  BUFF I157 (o_0r1[4:4], op3_4_0[3:3]);
  C2 I158 (op3_5_0[0:0], termf_2[5:5], termf_1[5:5]);
  C2 I159 (op3_5_0[1:1], termf_2[5:5], termt_1[5:5]);
  C2 I160 (op3_5_0[2:2], termt_2[5:5], termf_1[5:5]);
  C2 I161 (op3_5_0[3:3], termt_2[5:5], termt_1[5:5]);
  OR3 I162 (o_0r0[5:5], op3_5_0[0:0], op3_5_0[1:1], op3_5_0[2:2]);
  BUFF I163 (o_0r1[5:5], op3_5_0[3:3]);
  C2 I164 (op3_6_0[0:0], termf_2[6:6], termf_1[6:6]);
  C2 I165 (op3_6_0[1:1], termf_2[6:6], termt_1[6:6]);
  C2 I166 (op3_6_0[2:2], termt_2[6:6], termf_1[6:6]);
  C2 I167 (op3_6_0[3:3], termt_2[6:6], termt_1[6:6]);
  OR3 I168 (o_0r0[6:6], op3_6_0[0:0], op3_6_0[1:1], op3_6_0[2:2]);
  BUFF I169 (o_0r1[6:6], op3_6_0[3:3]);
  C2 I170 (op3_7_0[0:0], termf_2[7:7], termf_1[7:7]);
  C2 I171 (op3_7_0[1:1], termf_2[7:7], termt_1[7:7]);
  C2 I172 (op3_7_0[2:2], termt_2[7:7], termf_1[7:7]);
  C2 I173 (op3_7_0[3:3], termt_2[7:7], termt_1[7:7]);
  OR3 I174 (o_0r0[7:7], op3_7_0[0:0], op3_7_0[1:1], op3_7_0[2:2]);
  BUFF I175 (o_0r1[7:7], op3_7_0[3:3]);
  C2 I176 (op3_8_0[0:0], termf_2[8:8], termf_1[8:8]);
  C2 I177 (op3_8_0[1:1], termf_2[8:8], termt_1[8:8]);
  C2 I178 (op3_8_0[2:2], termt_2[8:8], termf_1[8:8]);
  C2 I179 (op3_8_0[3:3], termt_2[8:8], termt_1[8:8]);
  OR3 I180 (o_0r0[8:8], op3_8_0[0:0], op3_8_0[1:1], op3_8_0[2:2]);
  BUFF I181 (o_0r1[8:8], op3_8_0[3:3]);
  C2 I182 (op3_9_0[0:0], termf_2[9:9], termf_1[9:9]);
  C2 I183 (op3_9_0[1:1], termf_2[9:9], termt_1[9:9]);
  C2 I184 (op3_9_0[2:2], termt_2[9:9], termf_1[9:9]);
  C2 I185 (op3_9_0[3:3], termt_2[9:9], termt_1[9:9]);
  OR3 I186 (o_0r0[9:9], op3_9_0[0:0], op3_9_0[1:1], op3_9_0[2:2]);
  BUFF I187 (o_0r1[9:9], op3_9_0[3:3]);
  C2 I188 (op3_10_0[0:0], termf_2[10:10], termf_1[10:10]);
  C2 I189 (op3_10_0[1:1], termf_2[10:10], termt_1[10:10]);
  C2 I190 (op3_10_0[2:2], termt_2[10:10], termf_1[10:10]);
  C2 I191 (op3_10_0[3:3], termt_2[10:10], termt_1[10:10]);
  OR3 I192 (o_0r0[10:10], op3_10_0[0:0], op3_10_0[1:1], op3_10_0[2:2]);
  BUFF I193 (o_0r1[10:10], op3_10_0[3:3]);
  C2 I194 (op3_11_0[0:0], termf_2[11:11], termf_1[11:11]);
  C2 I195 (op3_11_0[1:1], termf_2[11:11], termt_1[11:11]);
  C2 I196 (op3_11_0[2:2], termt_2[11:11], termf_1[11:11]);
  C2 I197 (op3_11_0[3:3], termt_2[11:11], termt_1[11:11]);
  OR3 I198 (o_0r0[11:11], op3_11_0[0:0], op3_11_0[1:1], op3_11_0[2:2]);
  BUFF I199 (o_0r1[11:11], op3_11_0[3:3]);
  C2 I200 (op3_12_0[0:0], termf_2[12:12], termf_1[12:12]);
  C2 I201 (op3_12_0[1:1], termf_2[12:12], termt_1[12:12]);
  C2 I202 (op3_12_0[2:2], termt_2[12:12], termf_1[12:12]);
  C2 I203 (op3_12_0[3:3], termt_2[12:12], termt_1[12:12]);
  OR3 I204 (o_0r0[12:12], op3_12_0[0:0], op3_12_0[1:1], op3_12_0[2:2]);
  BUFF I205 (o_0r1[12:12], op3_12_0[3:3]);
  C2 I206 (op3_13_0[0:0], termf_2[13:13], termf_1[13:13]);
  C2 I207 (op3_13_0[1:1], termf_2[13:13], termt_1[13:13]);
  C2 I208 (op3_13_0[2:2], termt_2[13:13], termf_1[13:13]);
  C2 I209 (op3_13_0[3:3], termt_2[13:13], termt_1[13:13]);
  OR3 I210 (o_0r0[13:13], op3_13_0[0:0], op3_13_0[1:1], op3_13_0[2:2]);
  BUFF I211 (o_0r1[13:13], op3_13_0[3:3]);
  C2 I212 (op3_14_0[0:0], termf_2[14:14], termf_1[14:14]);
  C2 I213 (op3_14_0[1:1], termf_2[14:14], termt_1[14:14]);
  C2 I214 (op3_14_0[2:2], termt_2[14:14], termf_1[14:14]);
  C2 I215 (op3_14_0[3:3], termt_2[14:14], termt_1[14:14]);
  OR3 I216 (o_0r0[14:14], op3_14_0[0:0], op3_14_0[1:1], op3_14_0[2:2]);
  BUFF I217 (o_0r1[14:14], op3_14_0[3:3]);
  C2 I218 (op3_15_0[0:0], termf_2[15:15], termf_1[15:15]);
  C2 I219 (op3_15_0[1:1], termf_2[15:15], termt_1[15:15]);
  C2 I220 (op3_15_0[2:2], termt_2[15:15], termf_1[15:15]);
  C2 I221 (op3_15_0[3:3], termt_2[15:15], termt_1[15:15]);
  OR3 I222 (o_0r0[15:15], op3_15_0[0:0], op3_15_0[1:1], op3_15_0[2:2]);
  BUFF I223 (o_0r1[15:15], op3_15_0[3:3]);
  C2 I224 (op3_16_0[0:0], termf_2[16:16], termf_1[16:16]);
  C2 I225 (op3_16_0[1:1], termf_2[16:16], termt_1[16:16]);
  C2 I226 (op3_16_0[2:2], termt_2[16:16], termf_1[16:16]);
  C2 I227 (op3_16_0[3:3], termt_2[16:16], termt_1[16:16]);
  OR3 I228 (o_0r0[16:16], op3_16_0[0:0], op3_16_0[1:1], op3_16_0[2:2]);
  BUFF I229 (o_0r1[16:16], op3_16_0[3:3]);
  C2 I230 (op3_17_0[0:0], termf_2[17:17], termf_1[17:17]);
  C2 I231 (op3_17_0[1:1], termf_2[17:17], termt_1[17:17]);
  C2 I232 (op3_17_0[2:2], termt_2[17:17], termf_1[17:17]);
  C2 I233 (op3_17_0[3:3], termt_2[17:17], termt_1[17:17]);
  OR3 I234 (o_0r0[17:17], op3_17_0[0:0], op3_17_0[1:1], op3_17_0[2:2]);
  BUFF I235 (o_0r1[17:17], op3_17_0[3:3]);
  C2 I236 (op3_18_0[0:0], termf_2[18:18], termf_1[18:18]);
  C2 I237 (op3_18_0[1:1], termf_2[18:18], termt_1[18:18]);
  C2 I238 (op3_18_0[2:2], termt_2[18:18], termf_1[18:18]);
  C2 I239 (op3_18_0[3:3], termt_2[18:18], termt_1[18:18]);
  OR3 I240 (o_0r0[18:18], op3_18_0[0:0], op3_18_0[1:1], op3_18_0[2:2]);
  BUFF I241 (o_0r1[18:18], op3_18_0[3:3]);
  C2 I242 (op3_19_0[0:0], termf_2[19:19], termf_1[19:19]);
  C2 I243 (op3_19_0[1:1], termf_2[19:19], termt_1[19:19]);
  C2 I244 (op3_19_0[2:2], termt_2[19:19], termf_1[19:19]);
  C2 I245 (op3_19_0[3:3], termt_2[19:19], termt_1[19:19]);
  OR3 I246 (o_0r0[19:19], op3_19_0[0:0], op3_19_0[1:1], op3_19_0[2:2]);
  BUFF I247 (o_0r1[19:19], op3_19_0[3:3]);
  C2 I248 (op3_20_0[0:0], termf_2[20:20], termf_1[20:20]);
  C2 I249 (op3_20_0[1:1], termf_2[20:20], termt_1[20:20]);
  C2 I250 (op3_20_0[2:2], termt_2[20:20], termf_1[20:20]);
  C2 I251 (op3_20_0[3:3], termt_2[20:20], termt_1[20:20]);
  OR3 I252 (o_0r0[20:20], op3_20_0[0:0], op3_20_0[1:1], op3_20_0[2:2]);
  BUFF I253 (o_0r1[20:20], op3_20_0[3:3]);
  C2 I254 (op3_21_0[0:0], termf_2[21:21], termf_1[21:21]);
  C2 I255 (op3_21_0[1:1], termf_2[21:21], termt_1[21:21]);
  C2 I256 (op3_21_0[2:2], termt_2[21:21], termf_1[21:21]);
  C2 I257 (op3_21_0[3:3], termt_2[21:21], termt_1[21:21]);
  OR3 I258 (o_0r0[21:21], op3_21_0[0:0], op3_21_0[1:1], op3_21_0[2:2]);
  BUFF I259 (o_0r1[21:21], op3_21_0[3:3]);
  C2 I260 (op3_22_0[0:0], termf_2[22:22], termf_1[22:22]);
  C2 I261 (op3_22_0[1:1], termf_2[22:22], termt_1[22:22]);
  C2 I262 (op3_22_0[2:2], termt_2[22:22], termf_1[22:22]);
  C2 I263 (op3_22_0[3:3], termt_2[22:22], termt_1[22:22]);
  OR3 I264 (o_0r0[22:22], op3_22_0[0:0], op3_22_0[1:1], op3_22_0[2:2]);
  BUFF I265 (o_0r1[22:22], op3_22_0[3:3]);
  C2 I266 (op3_23_0[0:0], termf_2[23:23], termf_1[23:23]);
  C2 I267 (op3_23_0[1:1], termf_2[23:23], termt_1[23:23]);
  C2 I268 (op3_23_0[2:2], termt_2[23:23], termf_1[23:23]);
  C2 I269 (op3_23_0[3:3], termt_2[23:23], termt_1[23:23]);
  OR3 I270 (o_0r0[23:23], op3_23_0[0:0], op3_23_0[1:1], op3_23_0[2:2]);
  BUFF I271 (o_0r1[23:23], op3_23_0[3:3]);
  C2 I272 (op3_24_0[0:0], termf_2[24:24], termf_1[24:24]);
  C2 I273 (op3_24_0[1:1], termf_2[24:24], termt_1[24:24]);
  C2 I274 (op3_24_0[2:2], termt_2[24:24], termf_1[24:24]);
  C2 I275 (op3_24_0[3:3], termt_2[24:24], termt_1[24:24]);
  OR3 I276 (o_0r0[24:24], op3_24_0[0:0], op3_24_0[1:1], op3_24_0[2:2]);
  BUFF I277 (o_0r1[24:24], op3_24_0[3:3]);
  C2 I278 (op3_25_0[0:0], termf_2[25:25], termf_1[25:25]);
  C2 I279 (op3_25_0[1:1], termf_2[25:25], termt_1[25:25]);
  C2 I280 (op3_25_0[2:2], termt_2[25:25], termf_1[25:25]);
  C2 I281 (op3_25_0[3:3], termt_2[25:25], termt_1[25:25]);
  OR3 I282 (o_0r0[25:25], op3_25_0[0:0], op3_25_0[1:1], op3_25_0[2:2]);
  BUFF I283 (o_0r1[25:25], op3_25_0[3:3]);
  C2 I284 (op3_26_0[0:0], termf_2[26:26], termf_1[26:26]);
  C2 I285 (op3_26_0[1:1], termf_2[26:26], termt_1[26:26]);
  C2 I286 (op3_26_0[2:2], termt_2[26:26], termf_1[26:26]);
  C2 I287 (op3_26_0[3:3], termt_2[26:26], termt_1[26:26]);
  OR3 I288 (o_0r0[26:26], op3_26_0[0:0], op3_26_0[1:1], op3_26_0[2:2]);
  BUFF I289 (o_0r1[26:26], op3_26_0[3:3]);
  C2 I290 (op3_27_0[0:0], termf_2[27:27], termf_1[27:27]);
  C2 I291 (op3_27_0[1:1], termf_2[27:27], termt_1[27:27]);
  C2 I292 (op3_27_0[2:2], termt_2[27:27], termf_1[27:27]);
  C2 I293 (op3_27_0[3:3], termt_2[27:27], termt_1[27:27]);
  OR3 I294 (o_0r0[27:27], op3_27_0[0:0], op3_27_0[1:1], op3_27_0[2:2]);
  BUFF I295 (o_0r1[27:27], op3_27_0[3:3]);
  C2 I296 (op3_28_0[0:0], termf_2[28:28], termf_1[28:28]);
  C2 I297 (op3_28_0[1:1], termf_2[28:28], termt_1[28:28]);
  C2 I298 (op3_28_0[2:2], termt_2[28:28], termf_1[28:28]);
  C2 I299 (op3_28_0[3:3], termt_2[28:28], termt_1[28:28]);
  OR3 I300 (o_0r0[28:28], op3_28_0[0:0], op3_28_0[1:1], op3_28_0[2:2]);
  BUFF I301 (o_0r1[28:28], op3_28_0[3:3]);
  C2 I302 (op3_29_0[0:0], termf_2[29:29], termf_1[29:29]);
  C2 I303 (op3_29_0[1:1], termf_2[29:29], termt_1[29:29]);
  C2 I304 (op3_29_0[2:2], termt_2[29:29], termf_1[29:29]);
  C2 I305 (op3_29_0[3:3], termt_2[29:29], termt_1[29:29]);
  OR3 I306 (o_0r0[29:29], op3_29_0[0:0], op3_29_0[1:1], op3_29_0[2:2]);
  BUFF I307 (o_0r1[29:29], op3_29_0[3:3]);
  C2 I308 (op3_30_0[0:0], termf_2[30:30], termf_1[30:30]);
  C2 I309 (op3_30_0[1:1], termf_2[30:30], termt_1[30:30]);
  C2 I310 (op3_30_0[2:2], termt_2[30:30], termf_1[30:30]);
  C2 I311 (op3_30_0[3:3], termt_2[30:30], termt_1[30:30]);
  OR3 I312 (o_0r0[30:30], op3_30_0[0:0], op3_30_0[1:1], op3_30_0[2:2]);
  BUFF I313 (o_0r1[30:30], op3_30_0[3:3]);
  C2 I314 (op3_31_0[0:0], termf_2[31:31], termf_1[31:31]);
  C2 I315 (op3_31_0[1:1], termf_2[31:31], termt_1[31:31]);
  C2 I316 (op3_31_0[2:2], termt_2[31:31], termf_1[31:31]);
  C2 I317 (op3_31_0[3:3], termt_2[31:31], termt_1[31:31]);
  OR3 I318 (o_0r0[31:31], op3_31_0[0:0], op3_31_0[1:1], op3_31_0[2:2]);
  BUFF I319 (o_0r1[31:31], op3_31_0[3:3]);
  BUFF I320 (i_0a, o_0a);
endmodule

// tko64m32_1api0w32b_2api32w32b_3ort1o0w32bt2o0w32b TeakO [
//     (1,TeakOAppend 1 [(0,0+:32)]),
//     (2,TeakOAppend 1 [(0,32+:32)]),
//     (3,TeakOp TeakOpOr [(1,0+:32),(2,0+:32)])] [One 64,One 32]
module tko64m32_1api0w32b_2api32w32b_3ort1o0w32bt2o0w32b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [63:0] i_0r0;
  input [63:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire [31:0] termf_1;
  wire [31:0] termf_2;
  wire [31:0] termt_1;
  wire [31:0] termt_2;
  wire [3:0] op3_0_0;
  wire [3:0] op3_1_0;
  wire [3:0] op3_2_0;
  wire [3:0] op3_3_0;
  wire [3:0] op3_4_0;
  wire [3:0] op3_5_0;
  wire [3:0] op3_6_0;
  wire [3:0] op3_7_0;
  wire [3:0] op3_8_0;
  wire [3:0] op3_9_0;
  wire [3:0] op3_10_0;
  wire [3:0] op3_11_0;
  wire [3:0] op3_12_0;
  wire [3:0] op3_13_0;
  wire [3:0] op3_14_0;
  wire [3:0] op3_15_0;
  wire [3:0] op3_16_0;
  wire [3:0] op3_17_0;
  wire [3:0] op3_18_0;
  wire [3:0] op3_19_0;
  wire [3:0] op3_20_0;
  wire [3:0] op3_21_0;
  wire [3:0] op3_22_0;
  wire [3:0] op3_23_0;
  wire [3:0] op3_24_0;
  wire [3:0] op3_25_0;
  wire [3:0] op3_26_0;
  wire [3:0] op3_27_0;
  wire [3:0] op3_28_0;
  wire [3:0] op3_29_0;
  wire [3:0] op3_30_0;
  wire [3:0] op3_31_0;
  BUFF I0 (termf_1[0:0], i_0r0[0:0]);
  BUFF I1 (termf_1[1:1], i_0r0[1:1]);
  BUFF I2 (termf_1[2:2], i_0r0[2:2]);
  BUFF I3 (termf_1[3:3], i_0r0[3:3]);
  BUFF I4 (termf_1[4:4], i_0r0[4:4]);
  BUFF I5 (termf_1[5:5], i_0r0[5:5]);
  BUFF I6 (termf_1[6:6], i_0r0[6:6]);
  BUFF I7 (termf_1[7:7], i_0r0[7:7]);
  BUFF I8 (termf_1[8:8], i_0r0[8:8]);
  BUFF I9 (termf_1[9:9], i_0r0[9:9]);
  BUFF I10 (termf_1[10:10], i_0r0[10:10]);
  BUFF I11 (termf_1[11:11], i_0r0[11:11]);
  BUFF I12 (termf_1[12:12], i_0r0[12:12]);
  BUFF I13 (termf_1[13:13], i_0r0[13:13]);
  BUFF I14 (termf_1[14:14], i_0r0[14:14]);
  BUFF I15 (termf_1[15:15], i_0r0[15:15]);
  BUFF I16 (termf_1[16:16], i_0r0[16:16]);
  BUFF I17 (termf_1[17:17], i_0r0[17:17]);
  BUFF I18 (termf_1[18:18], i_0r0[18:18]);
  BUFF I19 (termf_1[19:19], i_0r0[19:19]);
  BUFF I20 (termf_1[20:20], i_0r0[20:20]);
  BUFF I21 (termf_1[21:21], i_0r0[21:21]);
  BUFF I22 (termf_1[22:22], i_0r0[22:22]);
  BUFF I23 (termf_1[23:23], i_0r0[23:23]);
  BUFF I24 (termf_1[24:24], i_0r0[24:24]);
  BUFF I25 (termf_1[25:25], i_0r0[25:25]);
  BUFF I26 (termf_1[26:26], i_0r0[26:26]);
  BUFF I27 (termf_1[27:27], i_0r0[27:27]);
  BUFF I28 (termf_1[28:28], i_0r0[28:28]);
  BUFF I29 (termf_1[29:29], i_0r0[29:29]);
  BUFF I30 (termf_1[30:30], i_0r0[30:30]);
  BUFF I31 (termf_1[31:31], i_0r0[31:31]);
  BUFF I32 (termt_1[0:0], i_0r1[0:0]);
  BUFF I33 (termt_1[1:1], i_0r1[1:1]);
  BUFF I34 (termt_1[2:2], i_0r1[2:2]);
  BUFF I35 (termt_1[3:3], i_0r1[3:3]);
  BUFF I36 (termt_1[4:4], i_0r1[4:4]);
  BUFF I37 (termt_1[5:5], i_0r1[5:5]);
  BUFF I38 (termt_1[6:6], i_0r1[6:6]);
  BUFF I39 (termt_1[7:7], i_0r1[7:7]);
  BUFF I40 (termt_1[8:8], i_0r1[8:8]);
  BUFF I41 (termt_1[9:9], i_0r1[9:9]);
  BUFF I42 (termt_1[10:10], i_0r1[10:10]);
  BUFF I43 (termt_1[11:11], i_0r1[11:11]);
  BUFF I44 (termt_1[12:12], i_0r1[12:12]);
  BUFF I45 (termt_1[13:13], i_0r1[13:13]);
  BUFF I46 (termt_1[14:14], i_0r1[14:14]);
  BUFF I47 (termt_1[15:15], i_0r1[15:15]);
  BUFF I48 (termt_1[16:16], i_0r1[16:16]);
  BUFF I49 (termt_1[17:17], i_0r1[17:17]);
  BUFF I50 (termt_1[18:18], i_0r1[18:18]);
  BUFF I51 (termt_1[19:19], i_0r1[19:19]);
  BUFF I52 (termt_1[20:20], i_0r1[20:20]);
  BUFF I53 (termt_1[21:21], i_0r1[21:21]);
  BUFF I54 (termt_1[22:22], i_0r1[22:22]);
  BUFF I55 (termt_1[23:23], i_0r1[23:23]);
  BUFF I56 (termt_1[24:24], i_0r1[24:24]);
  BUFF I57 (termt_1[25:25], i_0r1[25:25]);
  BUFF I58 (termt_1[26:26], i_0r1[26:26]);
  BUFF I59 (termt_1[27:27], i_0r1[27:27]);
  BUFF I60 (termt_1[28:28], i_0r1[28:28]);
  BUFF I61 (termt_1[29:29], i_0r1[29:29]);
  BUFF I62 (termt_1[30:30], i_0r1[30:30]);
  BUFF I63 (termt_1[31:31], i_0r1[31:31]);
  BUFF I64 (termf_2[0:0], i_0r0[32:32]);
  BUFF I65 (termf_2[1:1], i_0r0[33:33]);
  BUFF I66 (termf_2[2:2], i_0r0[34:34]);
  BUFF I67 (termf_2[3:3], i_0r0[35:35]);
  BUFF I68 (termf_2[4:4], i_0r0[36:36]);
  BUFF I69 (termf_2[5:5], i_0r0[37:37]);
  BUFF I70 (termf_2[6:6], i_0r0[38:38]);
  BUFF I71 (termf_2[7:7], i_0r0[39:39]);
  BUFF I72 (termf_2[8:8], i_0r0[40:40]);
  BUFF I73 (termf_2[9:9], i_0r0[41:41]);
  BUFF I74 (termf_2[10:10], i_0r0[42:42]);
  BUFF I75 (termf_2[11:11], i_0r0[43:43]);
  BUFF I76 (termf_2[12:12], i_0r0[44:44]);
  BUFF I77 (termf_2[13:13], i_0r0[45:45]);
  BUFF I78 (termf_2[14:14], i_0r0[46:46]);
  BUFF I79 (termf_2[15:15], i_0r0[47:47]);
  BUFF I80 (termf_2[16:16], i_0r0[48:48]);
  BUFF I81 (termf_2[17:17], i_0r0[49:49]);
  BUFF I82 (termf_2[18:18], i_0r0[50:50]);
  BUFF I83 (termf_2[19:19], i_0r0[51:51]);
  BUFF I84 (termf_2[20:20], i_0r0[52:52]);
  BUFF I85 (termf_2[21:21], i_0r0[53:53]);
  BUFF I86 (termf_2[22:22], i_0r0[54:54]);
  BUFF I87 (termf_2[23:23], i_0r0[55:55]);
  BUFF I88 (termf_2[24:24], i_0r0[56:56]);
  BUFF I89 (termf_2[25:25], i_0r0[57:57]);
  BUFF I90 (termf_2[26:26], i_0r0[58:58]);
  BUFF I91 (termf_2[27:27], i_0r0[59:59]);
  BUFF I92 (termf_2[28:28], i_0r0[60:60]);
  BUFF I93 (termf_2[29:29], i_0r0[61:61]);
  BUFF I94 (termf_2[30:30], i_0r0[62:62]);
  BUFF I95 (termf_2[31:31], i_0r0[63:63]);
  BUFF I96 (termt_2[0:0], i_0r1[32:32]);
  BUFF I97 (termt_2[1:1], i_0r1[33:33]);
  BUFF I98 (termt_2[2:2], i_0r1[34:34]);
  BUFF I99 (termt_2[3:3], i_0r1[35:35]);
  BUFF I100 (termt_2[4:4], i_0r1[36:36]);
  BUFF I101 (termt_2[5:5], i_0r1[37:37]);
  BUFF I102 (termt_2[6:6], i_0r1[38:38]);
  BUFF I103 (termt_2[7:7], i_0r1[39:39]);
  BUFF I104 (termt_2[8:8], i_0r1[40:40]);
  BUFF I105 (termt_2[9:9], i_0r1[41:41]);
  BUFF I106 (termt_2[10:10], i_0r1[42:42]);
  BUFF I107 (termt_2[11:11], i_0r1[43:43]);
  BUFF I108 (termt_2[12:12], i_0r1[44:44]);
  BUFF I109 (termt_2[13:13], i_0r1[45:45]);
  BUFF I110 (termt_2[14:14], i_0r1[46:46]);
  BUFF I111 (termt_2[15:15], i_0r1[47:47]);
  BUFF I112 (termt_2[16:16], i_0r1[48:48]);
  BUFF I113 (termt_2[17:17], i_0r1[49:49]);
  BUFF I114 (termt_2[18:18], i_0r1[50:50]);
  BUFF I115 (termt_2[19:19], i_0r1[51:51]);
  BUFF I116 (termt_2[20:20], i_0r1[52:52]);
  BUFF I117 (termt_2[21:21], i_0r1[53:53]);
  BUFF I118 (termt_2[22:22], i_0r1[54:54]);
  BUFF I119 (termt_2[23:23], i_0r1[55:55]);
  BUFF I120 (termt_2[24:24], i_0r1[56:56]);
  BUFF I121 (termt_2[25:25], i_0r1[57:57]);
  BUFF I122 (termt_2[26:26], i_0r1[58:58]);
  BUFF I123 (termt_2[27:27], i_0r1[59:59]);
  BUFF I124 (termt_2[28:28], i_0r1[60:60]);
  BUFF I125 (termt_2[29:29], i_0r1[61:61]);
  BUFF I126 (termt_2[30:30], i_0r1[62:62]);
  BUFF I127 (termt_2[31:31], i_0r1[63:63]);
  C2 I128 (op3_0_0[0:0], termf_2[0:0], termf_1[0:0]);
  C2 I129 (op3_0_0[1:1], termf_2[0:0], termt_1[0:0]);
  C2 I130 (op3_0_0[2:2], termt_2[0:0], termf_1[0:0]);
  C2 I131 (op3_0_0[3:3], termt_2[0:0], termt_1[0:0]);
  BUFF I132 (o_0r0[0:0], op3_0_0[0:0]);
  OR3 I133 (o_0r1[0:0], op3_0_0[1:1], op3_0_0[2:2], op3_0_0[3:3]);
  C2 I134 (op3_1_0[0:0], termf_2[1:1], termf_1[1:1]);
  C2 I135 (op3_1_0[1:1], termf_2[1:1], termt_1[1:1]);
  C2 I136 (op3_1_0[2:2], termt_2[1:1], termf_1[1:1]);
  C2 I137 (op3_1_0[3:3], termt_2[1:1], termt_1[1:1]);
  BUFF I138 (o_0r0[1:1], op3_1_0[0:0]);
  OR3 I139 (o_0r1[1:1], op3_1_0[1:1], op3_1_0[2:2], op3_1_0[3:3]);
  C2 I140 (op3_2_0[0:0], termf_2[2:2], termf_1[2:2]);
  C2 I141 (op3_2_0[1:1], termf_2[2:2], termt_1[2:2]);
  C2 I142 (op3_2_0[2:2], termt_2[2:2], termf_1[2:2]);
  C2 I143 (op3_2_0[3:3], termt_2[2:2], termt_1[2:2]);
  BUFF I144 (o_0r0[2:2], op3_2_0[0:0]);
  OR3 I145 (o_0r1[2:2], op3_2_0[1:1], op3_2_0[2:2], op3_2_0[3:3]);
  C2 I146 (op3_3_0[0:0], termf_2[3:3], termf_1[3:3]);
  C2 I147 (op3_3_0[1:1], termf_2[3:3], termt_1[3:3]);
  C2 I148 (op3_3_0[2:2], termt_2[3:3], termf_1[3:3]);
  C2 I149 (op3_3_0[3:3], termt_2[3:3], termt_1[3:3]);
  BUFF I150 (o_0r0[3:3], op3_3_0[0:0]);
  OR3 I151 (o_0r1[3:3], op3_3_0[1:1], op3_3_0[2:2], op3_3_0[3:3]);
  C2 I152 (op3_4_0[0:0], termf_2[4:4], termf_1[4:4]);
  C2 I153 (op3_4_0[1:1], termf_2[4:4], termt_1[4:4]);
  C2 I154 (op3_4_0[2:2], termt_2[4:4], termf_1[4:4]);
  C2 I155 (op3_4_0[3:3], termt_2[4:4], termt_1[4:4]);
  BUFF I156 (o_0r0[4:4], op3_4_0[0:0]);
  OR3 I157 (o_0r1[4:4], op3_4_0[1:1], op3_4_0[2:2], op3_4_0[3:3]);
  C2 I158 (op3_5_0[0:0], termf_2[5:5], termf_1[5:5]);
  C2 I159 (op3_5_0[1:1], termf_2[5:5], termt_1[5:5]);
  C2 I160 (op3_5_0[2:2], termt_2[5:5], termf_1[5:5]);
  C2 I161 (op3_5_0[3:3], termt_2[5:5], termt_1[5:5]);
  BUFF I162 (o_0r0[5:5], op3_5_0[0:0]);
  OR3 I163 (o_0r1[5:5], op3_5_0[1:1], op3_5_0[2:2], op3_5_0[3:3]);
  C2 I164 (op3_6_0[0:0], termf_2[6:6], termf_1[6:6]);
  C2 I165 (op3_6_0[1:1], termf_2[6:6], termt_1[6:6]);
  C2 I166 (op3_6_0[2:2], termt_2[6:6], termf_1[6:6]);
  C2 I167 (op3_6_0[3:3], termt_2[6:6], termt_1[6:6]);
  BUFF I168 (o_0r0[6:6], op3_6_0[0:0]);
  OR3 I169 (o_0r1[6:6], op3_6_0[1:1], op3_6_0[2:2], op3_6_0[3:3]);
  C2 I170 (op3_7_0[0:0], termf_2[7:7], termf_1[7:7]);
  C2 I171 (op3_7_0[1:1], termf_2[7:7], termt_1[7:7]);
  C2 I172 (op3_7_0[2:2], termt_2[7:7], termf_1[7:7]);
  C2 I173 (op3_7_0[3:3], termt_2[7:7], termt_1[7:7]);
  BUFF I174 (o_0r0[7:7], op3_7_0[0:0]);
  OR3 I175 (o_0r1[7:7], op3_7_0[1:1], op3_7_0[2:2], op3_7_0[3:3]);
  C2 I176 (op3_8_0[0:0], termf_2[8:8], termf_1[8:8]);
  C2 I177 (op3_8_0[1:1], termf_2[8:8], termt_1[8:8]);
  C2 I178 (op3_8_0[2:2], termt_2[8:8], termf_1[8:8]);
  C2 I179 (op3_8_0[3:3], termt_2[8:8], termt_1[8:8]);
  BUFF I180 (o_0r0[8:8], op3_8_0[0:0]);
  OR3 I181 (o_0r1[8:8], op3_8_0[1:1], op3_8_0[2:2], op3_8_0[3:3]);
  C2 I182 (op3_9_0[0:0], termf_2[9:9], termf_1[9:9]);
  C2 I183 (op3_9_0[1:1], termf_2[9:9], termt_1[9:9]);
  C2 I184 (op3_9_0[2:2], termt_2[9:9], termf_1[9:9]);
  C2 I185 (op3_9_0[3:3], termt_2[9:9], termt_1[9:9]);
  BUFF I186 (o_0r0[9:9], op3_9_0[0:0]);
  OR3 I187 (o_0r1[9:9], op3_9_0[1:1], op3_9_0[2:2], op3_9_0[3:3]);
  C2 I188 (op3_10_0[0:0], termf_2[10:10], termf_1[10:10]);
  C2 I189 (op3_10_0[1:1], termf_2[10:10], termt_1[10:10]);
  C2 I190 (op3_10_0[2:2], termt_2[10:10], termf_1[10:10]);
  C2 I191 (op3_10_0[3:3], termt_2[10:10], termt_1[10:10]);
  BUFF I192 (o_0r0[10:10], op3_10_0[0:0]);
  OR3 I193 (o_0r1[10:10], op3_10_0[1:1], op3_10_0[2:2], op3_10_0[3:3]);
  C2 I194 (op3_11_0[0:0], termf_2[11:11], termf_1[11:11]);
  C2 I195 (op3_11_0[1:1], termf_2[11:11], termt_1[11:11]);
  C2 I196 (op3_11_0[2:2], termt_2[11:11], termf_1[11:11]);
  C2 I197 (op3_11_0[3:3], termt_2[11:11], termt_1[11:11]);
  BUFF I198 (o_0r0[11:11], op3_11_0[0:0]);
  OR3 I199 (o_0r1[11:11], op3_11_0[1:1], op3_11_0[2:2], op3_11_0[3:3]);
  C2 I200 (op3_12_0[0:0], termf_2[12:12], termf_1[12:12]);
  C2 I201 (op3_12_0[1:1], termf_2[12:12], termt_1[12:12]);
  C2 I202 (op3_12_0[2:2], termt_2[12:12], termf_1[12:12]);
  C2 I203 (op3_12_0[3:3], termt_2[12:12], termt_1[12:12]);
  BUFF I204 (o_0r0[12:12], op3_12_0[0:0]);
  OR3 I205 (o_0r1[12:12], op3_12_0[1:1], op3_12_0[2:2], op3_12_0[3:3]);
  C2 I206 (op3_13_0[0:0], termf_2[13:13], termf_1[13:13]);
  C2 I207 (op3_13_0[1:1], termf_2[13:13], termt_1[13:13]);
  C2 I208 (op3_13_0[2:2], termt_2[13:13], termf_1[13:13]);
  C2 I209 (op3_13_0[3:3], termt_2[13:13], termt_1[13:13]);
  BUFF I210 (o_0r0[13:13], op3_13_0[0:0]);
  OR3 I211 (o_0r1[13:13], op3_13_0[1:1], op3_13_0[2:2], op3_13_0[3:3]);
  C2 I212 (op3_14_0[0:0], termf_2[14:14], termf_1[14:14]);
  C2 I213 (op3_14_0[1:1], termf_2[14:14], termt_1[14:14]);
  C2 I214 (op3_14_0[2:2], termt_2[14:14], termf_1[14:14]);
  C2 I215 (op3_14_0[3:3], termt_2[14:14], termt_1[14:14]);
  BUFF I216 (o_0r0[14:14], op3_14_0[0:0]);
  OR3 I217 (o_0r1[14:14], op3_14_0[1:1], op3_14_0[2:2], op3_14_0[3:3]);
  C2 I218 (op3_15_0[0:0], termf_2[15:15], termf_1[15:15]);
  C2 I219 (op3_15_0[1:1], termf_2[15:15], termt_1[15:15]);
  C2 I220 (op3_15_0[2:2], termt_2[15:15], termf_1[15:15]);
  C2 I221 (op3_15_0[3:3], termt_2[15:15], termt_1[15:15]);
  BUFF I222 (o_0r0[15:15], op3_15_0[0:0]);
  OR3 I223 (o_0r1[15:15], op3_15_0[1:1], op3_15_0[2:2], op3_15_0[3:3]);
  C2 I224 (op3_16_0[0:0], termf_2[16:16], termf_1[16:16]);
  C2 I225 (op3_16_0[1:1], termf_2[16:16], termt_1[16:16]);
  C2 I226 (op3_16_0[2:2], termt_2[16:16], termf_1[16:16]);
  C2 I227 (op3_16_0[3:3], termt_2[16:16], termt_1[16:16]);
  BUFF I228 (o_0r0[16:16], op3_16_0[0:0]);
  OR3 I229 (o_0r1[16:16], op3_16_0[1:1], op3_16_0[2:2], op3_16_0[3:3]);
  C2 I230 (op3_17_0[0:0], termf_2[17:17], termf_1[17:17]);
  C2 I231 (op3_17_0[1:1], termf_2[17:17], termt_1[17:17]);
  C2 I232 (op3_17_0[2:2], termt_2[17:17], termf_1[17:17]);
  C2 I233 (op3_17_0[3:3], termt_2[17:17], termt_1[17:17]);
  BUFF I234 (o_0r0[17:17], op3_17_0[0:0]);
  OR3 I235 (o_0r1[17:17], op3_17_0[1:1], op3_17_0[2:2], op3_17_0[3:3]);
  C2 I236 (op3_18_0[0:0], termf_2[18:18], termf_1[18:18]);
  C2 I237 (op3_18_0[1:1], termf_2[18:18], termt_1[18:18]);
  C2 I238 (op3_18_0[2:2], termt_2[18:18], termf_1[18:18]);
  C2 I239 (op3_18_0[3:3], termt_2[18:18], termt_1[18:18]);
  BUFF I240 (o_0r0[18:18], op3_18_0[0:0]);
  OR3 I241 (o_0r1[18:18], op3_18_0[1:1], op3_18_0[2:2], op3_18_0[3:3]);
  C2 I242 (op3_19_0[0:0], termf_2[19:19], termf_1[19:19]);
  C2 I243 (op3_19_0[1:1], termf_2[19:19], termt_1[19:19]);
  C2 I244 (op3_19_0[2:2], termt_2[19:19], termf_1[19:19]);
  C2 I245 (op3_19_0[3:3], termt_2[19:19], termt_1[19:19]);
  BUFF I246 (o_0r0[19:19], op3_19_0[0:0]);
  OR3 I247 (o_0r1[19:19], op3_19_0[1:1], op3_19_0[2:2], op3_19_0[3:3]);
  C2 I248 (op3_20_0[0:0], termf_2[20:20], termf_1[20:20]);
  C2 I249 (op3_20_0[1:1], termf_2[20:20], termt_1[20:20]);
  C2 I250 (op3_20_0[2:2], termt_2[20:20], termf_1[20:20]);
  C2 I251 (op3_20_0[3:3], termt_2[20:20], termt_1[20:20]);
  BUFF I252 (o_0r0[20:20], op3_20_0[0:0]);
  OR3 I253 (o_0r1[20:20], op3_20_0[1:1], op3_20_0[2:2], op3_20_0[3:3]);
  C2 I254 (op3_21_0[0:0], termf_2[21:21], termf_1[21:21]);
  C2 I255 (op3_21_0[1:1], termf_2[21:21], termt_1[21:21]);
  C2 I256 (op3_21_0[2:2], termt_2[21:21], termf_1[21:21]);
  C2 I257 (op3_21_0[3:3], termt_2[21:21], termt_1[21:21]);
  BUFF I258 (o_0r0[21:21], op3_21_0[0:0]);
  OR3 I259 (o_0r1[21:21], op3_21_0[1:1], op3_21_0[2:2], op3_21_0[3:3]);
  C2 I260 (op3_22_0[0:0], termf_2[22:22], termf_1[22:22]);
  C2 I261 (op3_22_0[1:1], termf_2[22:22], termt_1[22:22]);
  C2 I262 (op3_22_0[2:2], termt_2[22:22], termf_1[22:22]);
  C2 I263 (op3_22_0[3:3], termt_2[22:22], termt_1[22:22]);
  BUFF I264 (o_0r0[22:22], op3_22_0[0:0]);
  OR3 I265 (o_0r1[22:22], op3_22_0[1:1], op3_22_0[2:2], op3_22_0[3:3]);
  C2 I266 (op3_23_0[0:0], termf_2[23:23], termf_1[23:23]);
  C2 I267 (op3_23_0[1:1], termf_2[23:23], termt_1[23:23]);
  C2 I268 (op3_23_0[2:2], termt_2[23:23], termf_1[23:23]);
  C2 I269 (op3_23_0[3:3], termt_2[23:23], termt_1[23:23]);
  BUFF I270 (o_0r0[23:23], op3_23_0[0:0]);
  OR3 I271 (o_0r1[23:23], op3_23_0[1:1], op3_23_0[2:2], op3_23_0[3:3]);
  C2 I272 (op3_24_0[0:0], termf_2[24:24], termf_1[24:24]);
  C2 I273 (op3_24_0[1:1], termf_2[24:24], termt_1[24:24]);
  C2 I274 (op3_24_0[2:2], termt_2[24:24], termf_1[24:24]);
  C2 I275 (op3_24_0[3:3], termt_2[24:24], termt_1[24:24]);
  BUFF I276 (o_0r0[24:24], op3_24_0[0:0]);
  OR3 I277 (o_0r1[24:24], op3_24_0[1:1], op3_24_0[2:2], op3_24_0[3:3]);
  C2 I278 (op3_25_0[0:0], termf_2[25:25], termf_1[25:25]);
  C2 I279 (op3_25_0[1:1], termf_2[25:25], termt_1[25:25]);
  C2 I280 (op3_25_0[2:2], termt_2[25:25], termf_1[25:25]);
  C2 I281 (op3_25_0[3:3], termt_2[25:25], termt_1[25:25]);
  BUFF I282 (o_0r0[25:25], op3_25_0[0:0]);
  OR3 I283 (o_0r1[25:25], op3_25_0[1:1], op3_25_0[2:2], op3_25_0[3:3]);
  C2 I284 (op3_26_0[0:0], termf_2[26:26], termf_1[26:26]);
  C2 I285 (op3_26_0[1:1], termf_2[26:26], termt_1[26:26]);
  C2 I286 (op3_26_0[2:2], termt_2[26:26], termf_1[26:26]);
  C2 I287 (op3_26_0[3:3], termt_2[26:26], termt_1[26:26]);
  BUFF I288 (o_0r0[26:26], op3_26_0[0:0]);
  OR3 I289 (o_0r1[26:26], op3_26_0[1:1], op3_26_0[2:2], op3_26_0[3:3]);
  C2 I290 (op3_27_0[0:0], termf_2[27:27], termf_1[27:27]);
  C2 I291 (op3_27_0[1:1], termf_2[27:27], termt_1[27:27]);
  C2 I292 (op3_27_0[2:2], termt_2[27:27], termf_1[27:27]);
  C2 I293 (op3_27_0[3:3], termt_2[27:27], termt_1[27:27]);
  BUFF I294 (o_0r0[27:27], op3_27_0[0:0]);
  OR3 I295 (o_0r1[27:27], op3_27_0[1:1], op3_27_0[2:2], op3_27_0[3:3]);
  C2 I296 (op3_28_0[0:0], termf_2[28:28], termf_1[28:28]);
  C2 I297 (op3_28_0[1:1], termf_2[28:28], termt_1[28:28]);
  C2 I298 (op3_28_0[2:2], termt_2[28:28], termf_1[28:28]);
  C2 I299 (op3_28_0[3:3], termt_2[28:28], termt_1[28:28]);
  BUFF I300 (o_0r0[28:28], op3_28_0[0:0]);
  OR3 I301 (o_0r1[28:28], op3_28_0[1:1], op3_28_0[2:2], op3_28_0[3:3]);
  C2 I302 (op3_29_0[0:0], termf_2[29:29], termf_1[29:29]);
  C2 I303 (op3_29_0[1:1], termf_2[29:29], termt_1[29:29]);
  C2 I304 (op3_29_0[2:2], termt_2[29:29], termf_1[29:29]);
  C2 I305 (op3_29_0[3:3], termt_2[29:29], termt_1[29:29]);
  BUFF I306 (o_0r0[29:29], op3_29_0[0:0]);
  OR3 I307 (o_0r1[29:29], op3_29_0[1:1], op3_29_0[2:2], op3_29_0[3:3]);
  C2 I308 (op3_30_0[0:0], termf_2[30:30], termf_1[30:30]);
  C2 I309 (op3_30_0[1:1], termf_2[30:30], termt_1[30:30]);
  C2 I310 (op3_30_0[2:2], termt_2[30:30], termf_1[30:30]);
  C2 I311 (op3_30_0[3:3], termt_2[30:30], termt_1[30:30]);
  BUFF I312 (o_0r0[30:30], op3_30_0[0:0]);
  OR3 I313 (o_0r1[30:30], op3_30_0[1:1], op3_30_0[2:2], op3_30_0[3:3]);
  C2 I314 (op3_31_0[0:0], termf_2[31:31], termf_1[31:31]);
  C2 I315 (op3_31_0[1:1], termf_2[31:31], termt_1[31:31]);
  C2 I316 (op3_31_0[2:2], termt_2[31:31], termf_1[31:31]);
  C2 I317 (op3_31_0[3:3], termt_2[31:31], termt_1[31:31]);
  BUFF I318 (o_0r0[31:31], op3_31_0[0:0]);
  OR3 I319 (o_0r1[31:31], op3_31_0[1:1], op3_31_0[2:2], op3_31_0[3:3]);
  BUFF I320 (i_0a, o_0a);
endmodule

// tko64m32_1api0w32b_2api32w32b_3xort1o0w32bt2o0w32b TeakO [
//     (1,TeakOAppend 1 [(0,0+:32)]),
//     (2,TeakOAppend 1 [(0,32+:32)]),
//     (3,TeakOp TeakOpXor [(1,0+:32),(2,0+:32)])] [One 64,One 32]
module tko64m32_1api0w32b_2api32w32b_3xort1o0w32bt2o0w32b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [63:0] i_0r0;
  input [63:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire [31:0] termf_1;
  wire [31:0] termf_2;
  wire [31:0] termt_1;
  wire [31:0] termt_2;
  wire [3:0] op3_0_0;
  wire [3:0] op3_1_0;
  wire [3:0] op3_2_0;
  wire [3:0] op3_3_0;
  wire [3:0] op3_4_0;
  wire [3:0] op3_5_0;
  wire [3:0] op3_6_0;
  wire [3:0] op3_7_0;
  wire [3:0] op3_8_0;
  wire [3:0] op3_9_0;
  wire [3:0] op3_10_0;
  wire [3:0] op3_11_0;
  wire [3:0] op3_12_0;
  wire [3:0] op3_13_0;
  wire [3:0] op3_14_0;
  wire [3:0] op3_15_0;
  wire [3:0] op3_16_0;
  wire [3:0] op3_17_0;
  wire [3:0] op3_18_0;
  wire [3:0] op3_19_0;
  wire [3:0] op3_20_0;
  wire [3:0] op3_21_0;
  wire [3:0] op3_22_0;
  wire [3:0] op3_23_0;
  wire [3:0] op3_24_0;
  wire [3:0] op3_25_0;
  wire [3:0] op3_26_0;
  wire [3:0] op3_27_0;
  wire [3:0] op3_28_0;
  wire [3:0] op3_29_0;
  wire [3:0] op3_30_0;
  wire [3:0] op3_31_0;
  BUFF I0 (termf_1[0:0], i_0r0[0:0]);
  BUFF I1 (termf_1[1:1], i_0r0[1:1]);
  BUFF I2 (termf_1[2:2], i_0r0[2:2]);
  BUFF I3 (termf_1[3:3], i_0r0[3:3]);
  BUFF I4 (termf_1[4:4], i_0r0[4:4]);
  BUFF I5 (termf_1[5:5], i_0r0[5:5]);
  BUFF I6 (termf_1[6:6], i_0r0[6:6]);
  BUFF I7 (termf_1[7:7], i_0r0[7:7]);
  BUFF I8 (termf_1[8:8], i_0r0[8:8]);
  BUFF I9 (termf_1[9:9], i_0r0[9:9]);
  BUFF I10 (termf_1[10:10], i_0r0[10:10]);
  BUFF I11 (termf_1[11:11], i_0r0[11:11]);
  BUFF I12 (termf_1[12:12], i_0r0[12:12]);
  BUFF I13 (termf_1[13:13], i_0r0[13:13]);
  BUFF I14 (termf_1[14:14], i_0r0[14:14]);
  BUFF I15 (termf_1[15:15], i_0r0[15:15]);
  BUFF I16 (termf_1[16:16], i_0r0[16:16]);
  BUFF I17 (termf_1[17:17], i_0r0[17:17]);
  BUFF I18 (termf_1[18:18], i_0r0[18:18]);
  BUFF I19 (termf_1[19:19], i_0r0[19:19]);
  BUFF I20 (termf_1[20:20], i_0r0[20:20]);
  BUFF I21 (termf_1[21:21], i_0r0[21:21]);
  BUFF I22 (termf_1[22:22], i_0r0[22:22]);
  BUFF I23 (termf_1[23:23], i_0r0[23:23]);
  BUFF I24 (termf_1[24:24], i_0r0[24:24]);
  BUFF I25 (termf_1[25:25], i_0r0[25:25]);
  BUFF I26 (termf_1[26:26], i_0r0[26:26]);
  BUFF I27 (termf_1[27:27], i_0r0[27:27]);
  BUFF I28 (termf_1[28:28], i_0r0[28:28]);
  BUFF I29 (termf_1[29:29], i_0r0[29:29]);
  BUFF I30 (termf_1[30:30], i_0r0[30:30]);
  BUFF I31 (termf_1[31:31], i_0r0[31:31]);
  BUFF I32 (termt_1[0:0], i_0r1[0:0]);
  BUFF I33 (termt_1[1:1], i_0r1[1:1]);
  BUFF I34 (termt_1[2:2], i_0r1[2:2]);
  BUFF I35 (termt_1[3:3], i_0r1[3:3]);
  BUFF I36 (termt_1[4:4], i_0r1[4:4]);
  BUFF I37 (termt_1[5:5], i_0r1[5:5]);
  BUFF I38 (termt_1[6:6], i_0r1[6:6]);
  BUFF I39 (termt_1[7:7], i_0r1[7:7]);
  BUFF I40 (termt_1[8:8], i_0r1[8:8]);
  BUFF I41 (termt_1[9:9], i_0r1[9:9]);
  BUFF I42 (termt_1[10:10], i_0r1[10:10]);
  BUFF I43 (termt_1[11:11], i_0r1[11:11]);
  BUFF I44 (termt_1[12:12], i_0r1[12:12]);
  BUFF I45 (termt_1[13:13], i_0r1[13:13]);
  BUFF I46 (termt_1[14:14], i_0r1[14:14]);
  BUFF I47 (termt_1[15:15], i_0r1[15:15]);
  BUFF I48 (termt_1[16:16], i_0r1[16:16]);
  BUFF I49 (termt_1[17:17], i_0r1[17:17]);
  BUFF I50 (termt_1[18:18], i_0r1[18:18]);
  BUFF I51 (termt_1[19:19], i_0r1[19:19]);
  BUFF I52 (termt_1[20:20], i_0r1[20:20]);
  BUFF I53 (termt_1[21:21], i_0r1[21:21]);
  BUFF I54 (termt_1[22:22], i_0r1[22:22]);
  BUFF I55 (termt_1[23:23], i_0r1[23:23]);
  BUFF I56 (termt_1[24:24], i_0r1[24:24]);
  BUFF I57 (termt_1[25:25], i_0r1[25:25]);
  BUFF I58 (termt_1[26:26], i_0r1[26:26]);
  BUFF I59 (termt_1[27:27], i_0r1[27:27]);
  BUFF I60 (termt_1[28:28], i_0r1[28:28]);
  BUFF I61 (termt_1[29:29], i_0r1[29:29]);
  BUFF I62 (termt_1[30:30], i_0r1[30:30]);
  BUFF I63 (termt_1[31:31], i_0r1[31:31]);
  BUFF I64 (termf_2[0:0], i_0r0[32:32]);
  BUFF I65 (termf_2[1:1], i_0r0[33:33]);
  BUFF I66 (termf_2[2:2], i_0r0[34:34]);
  BUFF I67 (termf_2[3:3], i_0r0[35:35]);
  BUFF I68 (termf_2[4:4], i_0r0[36:36]);
  BUFF I69 (termf_2[5:5], i_0r0[37:37]);
  BUFF I70 (termf_2[6:6], i_0r0[38:38]);
  BUFF I71 (termf_2[7:7], i_0r0[39:39]);
  BUFF I72 (termf_2[8:8], i_0r0[40:40]);
  BUFF I73 (termf_2[9:9], i_0r0[41:41]);
  BUFF I74 (termf_2[10:10], i_0r0[42:42]);
  BUFF I75 (termf_2[11:11], i_0r0[43:43]);
  BUFF I76 (termf_2[12:12], i_0r0[44:44]);
  BUFF I77 (termf_2[13:13], i_0r0[45:45]);
  BUFF I78 (termf_2[14:14], i_0r0[46:46]);
  BUFF I79 (termf_2[15:15], i_0r0[47:47]);
  BUFF I80 (termf_2[16:16], i_0r0[48:48]);
  BUFF I81 (termf_2[17:17], i_0r0[49:49]);
  BUFF I82 (termf_2[18:18], i_0r0[50:50]);
  BUFF I83 (termf_2[19:19], i_0r0[51:51]);
  BUFF I84 (termf_2[20:20], i_0r0[52:52]);
  BUFF I85 (termf_2[21:21], i_0r0[53:53]);
  BUFF I86 (termf_2[22:22], i_0r0[54:54]);
  BUFF I87 (termf_2[23:23], i_0r0[55:55]);
  BUFF I88 (termf_2[24:24], i_0r0[56:56]);
  BUFF I89 (termf_2[25:25], i_0r0[57:57]);
  BUFF I90 (termf_2[26:26], i_0r0[58:58]);
  BUFF I91 (termf_2[27:27], i_0r0[59:59]);
  BUFF I92 (termf_2[28:28], i_0r0[60:60]);
  BUFF I93 (termf_2[29:29], i_0r0[61:61]);
  BUFF I94 (termf_2[30:30], i_0r0[62:62]);
  BUFF I95 (termf_2[31:31], i_0r0[63:63]);
  BUFF I96 (termt_2[0:0], i_0r1[32:32]);
  BUFF I97 (termt_2[1:1], i_0r1[33:33]);
  BUFF I98 (termt_2[2:2], i_0r1[34:34]);
  BUFF I99 (termt_2[3:3], i_0r1[35:35]);
  BUFF I100 (termt_2[4:4], i_0r1[36:36]);
  BUFF I101 (termt_2[5:5], i_0r1[37:37]);
  BUFF I102 (termt_2[6:6], i_0r1[38:38]);
  BUFF I103 (termt_2[7:7], i_0r1[39:39]);
  BUFF I104 (termt_2[8:8], i_0r1[40:40]);
  BUFF I105 (termt_2[9:9], i_0r1[41:41]);
  BUFF I106 (termt_2[10:10], i_0r1[42:42]);
  BUFF I107 (termt_2[11:11], i_0r1[43:43]);
  BUFF I108 (termt_2[12:12], i_0r1[44:44]);
  BUFF I109 (termt_2[13:13], i_0r1[45:45]);
  BUFF I110 (termt_2[14:14], i_0r1[46:46]);
  BUFF I111 (termt_2[15:15], i_0r1[47:47]);
  BUFF I112 (termt_2[16:16], i_0r1[48:48]);
  BUFF I113 (termt_2[17:17], i_0r1[49:49]);
  BUFF I114 (termt_2[18:18], i_0r1[50:50]);
  BUFF I115 (termt_2[19:19], i_0r1[51:51]);
  BUFF I116 (termt_2[20:20], i_0r1[52:52]);
  BUFF I117 (termt_2[21:21], i_0r1[53:53]);
  BUFF I118 (termt_2[22:22], i_0r1[54:54]);
  BUFF I119 (termt_2[23:23], i_0r1[55:55]);
  BUFF I120 (termt_2[24:24], i_0r1[56:56]);
  BUFF I121 (termt_2[25:25], i_0r1[57:57]);
  BUFF I122 (termt_2[26:26], i_0r1[58:58]);
  BUFF I123 (termt_2[27:27], i_0r1[59:59]);
  BUFF I124 (termt_2[28:28], i_0r1[60:60]);
  BUFF I125 (termt_2[29:29], i_0r1[61:61]);
  BUFF I126 (termt_2[30:30], i_0r1[62:62]);
  BUFF I127 (termt_2[31:31], i_0r1[63:63]);
  C2 I128 (op3_0_0[0:0], termf_2[0:0], termf_1[0:0]);
  C2 I129 (op3_0_0[1:1], termf_2[0:0], termt_1[0:0]);
  C2 I130 (op3_0_0[2:2], termt_2[0:0], termf_1[0:0]);
  C2 I131 (op3_0_0[3:3], termt_2[0:0], termt_1[0:0]);
  OR2 I132 (o_0r0[0:0], op3_0_0[0:0], op3_0_0[3:3]);
  OR2 I133 (o_0r1[0:0], op3_0_0[1:1], op3_0_0[2:2]);
  C2 I134 (op3_1_0[0:0], termf_2[1:1], termf_1[1:1]);
  C2 I135 (op3_1_0[1:1], termf_2[1:1], termt_1[1:1]);
  C2 I136 (op3_1_0[2:2], termt_2[1:1], termf_1[1:1]);
  C2 I137 (op3_1_0[3:3], termt_2[1:1], termt_1[1:1]);
  OR2 I138 (o_0r0[1:1], op3_1_0[0:0], op3_1_0[3:3]);
  OR2 I139 (o_0r1[1:1], op3_1_0[1:1], op3_1_0[2:2]);
  C2 I140 (op3_2_0[0:0], termf_2[2:2], termf_1[2:2]);
  C2 I141 (op3_2_0[1:1], termf_2[2:2], termt_1[2:2]);
  C2 I142 (op3_2_0[2:2], termt_2[2:2], termf_1[2:2]);
  C2 I143 (op3_2_0[3:3], termt_2[2:2], termt_1[2:2]);
  OR2 I144 (o_0r0[2:2], op3_2_0[0:0], op3_2_0[3:3]);
  OR2 I145 (o_0r1[2:2], op3_2_0[1:1], op3_2_0[2:2]);
  C2 I146 (op3_3_0[0:0], termf_2[3:3], termf_1[3:3]);
  C2 I147 (op3_3_0[1:1], termf_2[3:3], termt_1[3:3]);
  C2 I148 (op3_3_0[2:2], termt_2[3:3], termf_1[3:3]);
  C2 I149 (op3_3_0[3:3], termt_2[3:3], termt_1[3:3]);
  OR2 I150 (o_0r0[3:3], op3_3_0[0:0], op3_3_0[3:3]);
  OR2 I151 (o_0r1[3:3], op3_3_0[1:1], op3_3_0[2:2]);
  C2 I152 (op3_4_0[0:0], termf_2[4:4], termf_1[4:4]);
  C2 I153 (op3_4_0[1:1], termf_2[4:4], termt_1[4:4]);
  C2 I154 (op3_4_0[2:2], termt_2[4:4], termf_1[4:4]);
  C2 I155 (op3_4_0[3:3], termt_2[4:4], termt_1[4:4]);
  OR2 I156 (o_0r0[4:4], op3_4_0[0:0], op3_4_0[3:3]);
  OR2 I157 (o_0r1[4:4], op3_4_0[1:1], op3_4_0[2:2]);
  C2 I158 (op3_5_0[0:0], termf_2[5:5], termf_1[5:5]);
  C2 I159 (op3_5_0[1:1], termf_2[5:5], termt_1[5:5]);
  C2 I160 (op3_5_0[2:2], termt_2[5:5], termf_1[5:5]);
  C2 I161 (op3_5_0[3:3], termt_2[5:5], termt_1[5:5]);
  OR2 I162 (o_0r0[5:5], op3_5_0[0:0], op3_5_0[3:3]);
  OR2 I163 (o_0r1[5:5], op3_5_0[1:1], op3_5_0[2:2]);
  C2 I164 (op3_6_0[0:0], termf_2[6:6], termf_1[6:6]);
  C2 I165 (op3_6_0[1:1], termf_2[6:6], termt_1[6:6]);
  C2 I166 (op3_6_0[2:2], termt_2[6:6], termf_1[6:6]);
  C2 I167 (op3_6_0[3:3], termt_2[6:6], termt_1[6:6]);
  OR2 I168 (o_0r0[6:6], op3_6_0[0:0], op3_6_0[3:3]);
  OR2 I169 (o_0r1[6:6], op3_6_0[1:1], op3_6_0[2:2]);
  C2 I170 (op3_7_0[0:0], termf_2[7:7], termf_1[7:7]);
  C2 I171 (op3_7_0[1:1], termf_2[7:7], termt_1[7:7]);
  C2 I172 (op3_7_0[2:2], termt_2[7:7], termf_1[7:7]);
  C2 I173 (op3_7_0[3:3], termt_2[7:7], termt_1[7:7]);
  OR2 I174 (o_0r0[7:7], op3_7_0[0:0], op3_7_0[3:3]);
  OR2 I175 (o_0r1[7:7], op3_7_0[1:1], op3_7_0[2:2]);
  C2 I176 (op3_8_0[0:0], termf_2[8:8], termf_1[8:8]);
  C2 I177 (op3_8_0[1:1], termf_2[8:8], termt_1[8:8]);
  C2 I178 (op3_8_0[2:2], termt_2[8:8], termf_1[8:8]);
  C2 I179 (op3_8_0[3:3], termt_2[8:8], termt_1[8:8]);
  OR2 I180 (o_0r0[8:8], op3_8_0[0:0], op3_8_0[3:3]);
  OR2 I181 (o_0r1[8:8], op3_8_0[1:1], op3_8_0[2:2]);
  C2 I182 (op3_9_0[0:0], termf_2[9:9], termf_1[9:9]);
  C2 I183 (op3_9_0[1:1], termf_2[9:9], termt_1[9:9]);
  C2 I184 (op3_9_0[2:2], termt_2[9:9], termf_1[9:9]);
  C2 I185 (op3_9_0[3:3], termt_2[9:9], termt_1[9:9]);
  OR2 I186 (o_0r0[9:9], op3_9_0[0:0], op3_9_0[3:3]);
  OR2 I187 (o_0r1[9:9], op3_9_0[1:1], op3_9_0[2:2]);
  C2 I188 (op3_10_0[0:0], termf_2[10:10], termf_1[10:10]);
  C2 I189 (op3_10_0[1:1], termf_2[10:10], termt_1[10:10]);
  C2 I190 (op3_10_0[2:2], termt_2[10:10], termf_1[10:10]);
  C2 I191 (op3_10_0[3:3], termt_2[10:10], termt_1[10:10]);
  OR2 I192 (o_0r0[10:10], op3_10_0[0:0], op3_10_0[3:3]);
  OR2 I193 (o_0r1[10:10], op3_10_0[1:1], op3_10_0[2:2]);
  C2 I194 (op3_11_0[0:0], termf_2[11:11], termf_1[11:11]);
  C2 I195 (op3_11_0[1:1], termf_2[11:11], termt_1[11:11]);
  C2 I196 (op3_11_0[2:2], termt_2[11:11], termf_1[11:11]);
  C2 I197 (op3_11_0[3:3], termt_2[11:11], termt_1[11:11]);
  OR2 I198 (o_0r0[11:11], op3_11_0[0:0], op3_11_0[3:3]);
  OR2 I199 (o_0r1[11:11], op3_11_0[1:1], op3_11_0[2:2]);
  C2 I200 (op3_12_0[0:0], termf_2[12:12], termf_1[12:12]);
  C2 I201 (op3_12_0[1:1], termf_2[12:12], termt_1[12:12]);
  C2 I202 (op3_12_0[2:2], termt_2[12:12], termf_1[12:12]);
  C2 I203 (op3_12_0[3:3], termt_2[12:12], termt_1[12:12]);
  OR2 I204 (o_0r0[12:12], op3_12_0[0:0], op3_12_0[3:3]);
  OR2 I205 (o_0r1[12:12], op3_12_0[1:1], op3_12_0[2:2]);
  C2 I206 (op3_13_0[0:0], termf_2[13:13], termf_1[13:13]);
  C2 I207 (op3_13_0[1:1], termf_2[13:13], termt_1[13:13]);
  C2 I208 (op3_13_0[2:2], termt_2[13:13], termf_1[13:13]);
  C2 I209 (op3_13_0[3:3], termt_2[13:13], termt_1[13:13]);
  OR2 I210 (o_0r0[13:13], op3_13_0[0:0], op3_13_0[3:3]);
  OR2 I211 (o_0r1[13:13], op3_13_0[1:1], op3_13_0[2:2]);
  C2 I212 (op3_14_0[0:0], termf_2[14:14], termf_1[14:14]);
  C2 I213 (op3_14_0[1:1], termf_2[14:14], termt_1[14:14]);
  C2 I214 (op3_14_0[2:2], termt_2[14:14], termf_1[14:14]);
  C2 I215 (op3_14_0[3:3], termt_2[14:14], termt_1[14:14]);
  OR2 I216 (o_0r0[14:14], op3_14_0[0:0], op3_14_0[3:3]);
  OR2 I217 (o_0r1[14:14], op3_14_0[1:1], op3_14_0[2:2]);
  C2 I218 (op3_15_0[0:0], termf_2[15:15], termf_1[15:15]);
  C2 I219 (op3_15_0[1:1], termf_2[15:15], termt_1[15:15]);
  C2 I220 (op3_15_0[2:2], termt_2[15:15], termf_1[15:15]);
  C2 I221 (op3_15_0[3:3], termt_2[15:15], termt_1[15:15]);
  OR2 I222 (o_0r0[15:15], op3_15_0[0:0], op3_15_0[3:3]);
  OR2 I223 (o_0r1[15:15], op3_15_0[1:1], op3_15_0[2:2]);
  C2 I224 (op3_16_0[0:0], termf_2[16:16], termf_1[16:16]);
  C2 I225 (op3_16_0[1:1], termf_2[16:16], termt_1[16:16]);
  C2 I226 (op3_16_0[2:2], termt_2[16:16], termf_1[16:16]);
  C2 I227 (op3_16_0[3:3], termt_2[16:16], termt_1[16:16]);
  OR2 I228 (o_0r0[16:16], op3_16_0[0:0], op3_16_0[3:3]);
  OR2 I229 (o_0r1[16:16], op3_16_0[1:1], op3_16_0[2:2]);
  C2 I230 (op3_17_0[0:0], termf_2[17:17], termf_1[17:17]);
  C2 I231 (op3_17_0[1:1], termf_2[17:17], termt_1[17:17]);
  C2 I232 (op3_17_0[2:2], termt_2[17:17], termf_1[17:17]);
  C2 I233 (op3_17_0[3:3], termt_2[17:17], termt_1[17:17]);
  OR2 I234 (o_0r0[17:17], op3_17_0[0:0], op3_17_0[3:3]);
  OR2 I235 (o_0r1[17:17], op3_17_0[1:1], op3_17_0[2:2]);
  C2 I236 (op3_18_0[0:0], termf_2[18:18], termf_1[18:18]);
  C2 I237 (op3_18_0[1:1], termf_2[18:18], termt_1[18:18]);
  C2 I238 (op3_18_0[2:2], termt_2[18:18], termf_1[18:18]);
  C2 I239 (op3_18_0[3:3], termt_2[18:18], termt_1[18:18]);
  OR2 I240 (o_0r0[18:18], op3_18_0[0:0], op3_18_0[3:3]);
  OR2 I241 (o_0r1[18:18], op3_18_0[1:1], op3_18_0[2:2]);
  C2 I242 (op3_19_0[0:0], termf_2[19:19], termf_1[19:19]);
  C2 I243 (op3_19_0[1:1], termf_2[19:19], termt_1[19:19]);
  C2 I244 (op3_19_0[2:2], termt_2[19:19], termf_1[19:19]);
  C2 I245 (op3_19_0[3:3], termt_2[19:19], termt_1[19:19]);
  OR2 I246 (o_0r0[19:19], op3_19_0[0:0], op3_19_0[3:3]);
  OR2 I247 (o_0r1[19:19], op3_19_0[1:1], op3_19_0[2:2]);
  C2 I248 (op3_20_0[0:0], termf_2[20:20], termf_1[20:20]);
  C2 I249 (op3_20_0[1:1], termf_2[20:20], termt_1[20:20]);
  C2 I250 (op3_20_0[2:2], termt_2[20:20], termf_1[20:20]);
  C2 I251 (op3_20_0[3:3], termt_2[20:20], termt_1[20:20]);
  OR2 I252 (o_0r0[20:20], op3_20_0[0:0], op3_20_0[3:3]);
  OR2 I253 (o_0r1[20:20], op3_20_0[1:1], op3_20_0[2:2]);
  C2 I254 (op3_21_0[0:0], termf_2[21:21], termf_1[21:21]);
  C2 I255 (op3_21_0[1:1], termf_2[21:21], termt_1[21:21]);
  C2 I256 (op3_21_0[2:2], termt_2[21:21], termf_1[21:21]);
  C2 I257 (op3_21_0[3:3], termt_2[21:21], termt_1[21:21]);
  OR2 I258 (o_0r0[21:21], op3_21_0[0:0], op3_21_0[3:3]);
  OR2 I259 (o_0r1[21:21], op3_21_0[1:1], op3_21_0[2:2]);
  C2 I260 (op3_22_0[0:0], termf_2[22:22], termf_1[22:22]);
  C2 I261 (op3_22_0[1:1], termf_2[22:22], termt_1[22:22]);
  C2 I262 (op3_22_0[2:2], termt_2[22:22], termf_1[22:22]);
  C2 I263 (op3_22_0[3:3], termt_2[22:22], termt_1[22:22]);
  OR2 I264 (o_0r0[22:22], op3_22_0[0:0], op3_22_0[3:3]);
  OR2 I265 (o_0r1[22:22], op3_22_0[1:1], op3_22_0[2:2]);
  C2 I266 (op3_23_0[0:0], termf_2[23:23], termf_1[23:23]);
  C2 I267 (op3_23_0[1:1], termf_2[23:23], termt_1[23:23]);
  C2 I268 (op3_23_0[2:2], termt_2[23:23], termf_1[23:23]);
  C2 I269 (op3_23_0[3:3], termt_2[23:23], termt_1[23:23]);
  OR2 I270 (o_0r0[23:23], op3_23_0[0:0], op3_23_0[3:3]);
  OR2 I271 (o_0r1[23:23], op3_23_0[1:1], op3_23_0[2:2]);
  C2 I272 (op3_24_0[0:0], termf_2[24:24], termf_1[24:24]);
  C2 I273 (op3_24_0[1:1], termf_2[24:24], termt_1[24:24]);
  C2 I274 (op3_24_0[2:2], termt_2[24:24], termf_1[24:24]);
  C2 I275 (op3_24_0[3:3], termt_2[24:24], termt_1[24:24]);
  OR2 I276 (o_0r0[24:24], op3_24_0[0:0], op3_24_0[3:3]);
  OR2 I277 (o_0r1[24:24], op3_24_0[1:1], op3_24_0[2:2]);
  C2 I278 (op3_25_0[0:0], termf_2[25:25], termf_1[25:25]);
  C2 I279 (op3_25_0[1:1], termf_2[25:25], termt_1[25:25]);
  C2 I280 (op3_25_0[2:2], termt_2[25:25], termf_1[25:25]);
  C2 I281 (op3_25_0[3:3], termt_2[25:25], termt_1[25:25]);
  OR2 I282 (o_0r0[25:25], op3_25_0[0:0], op3_25_0[3:3]);
  OR2 I283 (o_0r1[25:25], op3_25_0[1:1], op3_25_0[2:2]);
  C2 I284 (op3_26_0[0:0], termf_2[26:26], termf_1[26:26]);
  C2 I285 (op3_26_0[1:1], termf_2[26:26], termt_1[26:26]);
  C2 I286 (op3_26_0[2:2], termt_2[26:26], termf_1[26:26]);
  C2 I287 (op3_26_0[3:3], termt_2[26:26], termt_1[26:26]);
  OR2 I288 (o_0r0[26:26], op3_26_0[0:0], op3_26_0[3:3]);
  OR2 I289 (o_0r1[26:26], op3_26_0[1:1], op3_26_0[2:2]);
  C2 I290 (op3_27_0[0:0], termf_2[27:27], termf_1[27:27]);
  C2 I291 (op3_27_0[1:1], termf_2[27:27], termt_1[27:27]);
  C2 I292 (op3_27_0[2:2], termt_2[27:27], termf_1[27:27]);
  C2 I293 (op3_27_0[3:3], termt_2[27:27], termt_1[27:27]);
  OR2 I294 (o_0r0[27:27], op3_27_0[0:0], op3_27_0[3:3]);
  OR2 I295 (o_0r1[27:27], op3_27_0[1:1], op3_27_0[2:2]);
  C2 I296 (op3_28_0[0:0], termf_2[28:28], termf_1[28:28]);
  C2 I297 (op3_28_0[1:1], termf_2[28:28], termt_1[28:28]);
  C2 I298 (op3_28_0[2:2], termt_2[28:28], termf_1[28:28]);
  C2 I299 (op3_28_0[3:3], termt_2[28:28], termt_1[28:28]);
  OR2 I300 (o_0r0[28:28], op3_28_0[0:0], op3_28_0[3:3]);
  OR2 I301 (o_0r1[28:28], op3_28_0[1:1], op3_28_0[2:2]);
  C2 I302 (op3_29_0[0:0], termf_2[29:29], termf_1[29:29]);
  C2 I303 (op3_29_0[1:1], termf_2[29:29], termt_1[29:29]);
  C2 I304 (op3_29_0[2:2], termt_2[29:29], termf_1[29:29]);
  C2 I305 (op3_29_0[3:3], termt_2[29:29], termt_1[29:29]);
  OR2 I306 (o_0r0[29:29], op3_29_0[0:0], op3_29_0[3:3]);
  OR2 I307 (o_0r1[29:29], op3_29_0[1:1], op3_29_0[2:2]);
  C2 I308 (op3_30_0[0:0], termf_2[30:30], termf_1[30:30]);
  C2 I309 (op3_30_0[1:1], termf_2[30:30], termt_1[30:30]);
  C2 I310 (op3_30_0[2:2], termt_2[30:30], termf_1[30:30]);
  C2 I311 (op3_30_0[3:3], termt_2[30:30], termt_1[30:30]);
  OR2 I312 (o_0r0[30:30], op3_30_0[0:0], op3_30_0[3:3]);
  OR2 I313 (o_0r1[30:30], op3_30_0[1:1], op3_30_0[2:2]);
  C2 I314 (op3_31_0[0:0], termf_2[31:31], termf_1[31:31]);
  C2 I315 (op3_31_0[1:1], termf_2[31:31], termt_1[31:31]);
  C2 I316 (op3_31_0[2:2], termt_2[31:31], termf_1[31:31]);
  C2 I317 (op3_31_0[3:3], termt_2[31:31], termt_1[31:31]);
  OR2 I318 (o_0r0[31:31], op3_31_0[0:0], op3_31_0[3:3]);
  OR2 I319 (o_0r1[31:31], op3_31_0[1:1], op3_31_0[2:2]);
  BUFF I320 (i_0a, o_0a);
endmodule

// tkj2m1_1 TeakJ [Many [1,1],One 2]
module tkj2m1_1 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input i_1r0;
  input i_1r1;
  output i_1a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [1:0] joinf_0;
  wire [1:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0);
  BUFF I1 (joinf_0[1:1], i_1r0);
  BUFF I2 (joint_0[0:0], i_0r1);
  BUFF I3 (joint_0[1:1], i_1r1);
  OR2 I4 (dcomplete_0, i_1r0, i_1r1);
  BUFF I5 (icomplete_0, dcomplete_0);
  C2 I6 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I7 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I8 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I9 (o_0r1[1:1], joint_0[1:1]);
  BUFF I10 (i_0a, o_0a);
  BUFF I11 (i_1a, o_0a);
endmodule

// tks6_o0w6_4c20m9c30mac30mbc30mdc30mec30mfc30m20m21m22m23m28m2cm30m31m32m33m34m35m36m37m38m3co0w0_0m8
//   mcm10m14m18m1co0w0_1m5m11m15o0w0_2m6m12m16o0w0_3m7m13m17o0w0_25o0w0_26o0w0_27o0w0 TeakS (0+:6) [([Im
//   p 4 32,Imp 9 48,Imp 10 48,Imp 11 48,Imp 13 48,Imp 14 48,Imp 15 48,Imp 32 0,Imp 33 0,Imp 34 0,Imp 35 
//   0,Imp 40 0,Imp 44 0,Imp 48 0,Imp 49 0,Imp 50 0,Imp 51 0,Imp 52 0,Imp 53 0,Imp 54 0,Imp 55 0,Imp 56 0
//   ,Imp 60 0],0),([Imp 0 0,Imp 8 0,Imp 12 0,Imp 16 0,Imp 20 0,Imp 24 0,Imp 28 0],0),([Imp 1 0,Imp 5 0,I
//   mp 17 0,Imp 21 0],0),([Imp 2 0,Imp 6 0,Imp 18 0,Imp 22 0],0),([Imp 3 0,Imp 7 0,Imp 19 0,Imp 23 0],0)
//   ,([Imp 37 0],0),([Imp 38 0],0),([Imp 39 0],0)] [One 6,Many [0,0,0,0,0,0,0,0]]
module tks6_o0w6_4c20m9c30mac30mbc30mdc30mec30mfc30m20m21m22m23m28m2cm30m31m32m33m34m35m36m37m38m3co0w0_0m8mcm10m14m18m1co0w0_1m5m11m15o0w0_2m6m12m16o0w0_3m7m13m17o0w0_25o0w0_26o0w0_27o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, o_5r, o_5a, o_6r, o_6a, o_7r, o_7a, reset);
  input [5:0] i_0r0;
  input [5:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  output o_7r;
  input o_7a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire sel_4;
  wire sel_5;
  wire sel_6;
  wire sel_7;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire gsel_4;
  wire gsel_5;
  wire gsel_6;
  wire gsel_7;
  wire oack_0;
  wire [22:0] match0_0;
  wire [7:0] simp191_0;
  wire [2:0] simp192_0;
  wire [1:0] simp201_0;
  wire [1:0] simp211_0;
  wire [1:0] simp221_0;
  wire [1:0] simp231_0;
  wire [1:0] simp241_0;
  wire [1:0] simp251_0;
  wire [1:0] simp261_0;
  wire [1:0] simp271_0;
  wire [1:0] simp281_0;
  wire [1:0] simp291_0;
  wire [1:0] simp301_0;
  wire [1:0] simp311_0;
  wire [1:0] simp321_0;
  wire [1:0] simp331_0;
  wire [1:0] simp341_0;
  wire [1:0] simp351_0;
  wire [1:0] simp361_0;
  wire [1:0] simp371_0;
  wire [1:0] simp381_0;
  wire [1:0] simp391_0;
  wire [1:0] simp401_0;
  wire [1:0] simp411_0;
  wire [1:0] simp421_0;
  wire [6:0] match1_0;
  wire [2:0] simp441_0;
  wire [1:0] simp451_0;
  wire [1:0] simp461_0;
  wire [1:0] simp471_0;
  wire [1:0] simp481_0;
  wire [1:0] simp491_0;
  wire [1:0] simp501_0;
  wire [1:0] simp511_0;
  wire [3:0] match2_0;
  wire [1:0] simp531_0;
  wire [1:0] simp541_0;
  wire [1:0] simp551_0;
  wire [1:0] simp561_0;
  wire [1:0] simp571_0;
  wire [3:0] match3_0;
  wire [1:0] simp591_0;
  wire [1:0] simp601_0;
  wire [1:0] simp611_0;
  wire [1:0] simp621_0;
  wire [1:0] simp631_0;
  wire [3:0] match4_0;
  wire [1:0] simp651_0;
  wire [1:0] simp661_0;
  wire [1:0] simp671_0;
  wire [1:0] simp681_0;
  wire [1:0] simp691_0;
  wire match5_0;
  wire [1:0] simp721_0;
  wire match6_0;
  wire [1:0] simp751_0;
  wire match7_0;
  wire [1:0] simp781_0;
  wire [5:0] comp_0;
  wire [1:0] simp941_0;
  wire [2:0] simp1031_0;
  NOR3 I0 (simp191_0[0:0], match0_0[0:0], match0_0[1:1], match0_0[2:2]);
  NOR3 I1 (simp191_0[1:1], match0_0[3:3], match0_0[4:4], match0_0[5:5]);
  NOR3 I2 (simp191_0[2:2], match0_0[6:6], match0_0[7:7], match0_0[8:8]);
  NOR3 I3 (simp191_0[3:3], match0_0[9:9], match0_0[10:10], match0_0[11:11]);
  NOR3 I4 (simp191_0[4:4], match0_0[12:12], match0_0[13:13], match0_0[14:14]);
  NOR3 I5 (simp191_0[5:5], match0_0[15:15], match0_0[16:16], match0_0[17:17]);
  NOR3 I6 (simp191_0[6:6], match0_0[18:18], match0_0[19:19], match0_0[20:20]);
  NOR2 I7 (simp191_0[7:7], match0_0[21:21], match0_0[22:22]);
  NAND3 I8 (simp192_0[0:0], simp191_0[0:0], simp191_0[1:1], simp191_0[2:2]);
  NAND3 I9 (simp192_0[1:1], simp191_0[3:3], simp191_0[4:4], simp191_0[5:5]);
  NAND2 I10 (simp192_0[2:2], simp191_0[6:6], simp191_0[7:7]);
  OR3 I11 (sel_0, simp192_0[0:0], simp192_0[1:1], simp192_0[2:2]);
  C3 I12 (simp201_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C2 I13 (simp201_0[1:1], i_0r0[3:3], i_0r0[4:4]);
  C2 I14 (match0_0[0:0], simp201_0[0:0], simp201_0[1:1]);
  C3 I15 (simp211_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I16 (simp211_0[1:1], i_0r1[3:3]);
  C2 I17 (match0_0[1:1], simp211_0[0:0], simp211_0[1:1]);
  C3 I18 (simp221_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I19 (simp221_0[1:1], i_0r1[3:3]);
  C2 I20 (match0_0[2:2], simp221_0[0:0], simp221_0[1:1]);
  C3 I21 (simp231_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I22 (simp231_0[1:1], i_0r1[3:3]);
  C2 I23 (match0_0[3:3], simp231_0[0:0], simp231_0[1:1]);
  C3 I24 (simp241_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I25 (simp241_0[1:1], i_0r1[3:3]);
  C2 I26 (match0_0[4:4], simp241_0[0:0], simp241_0[1:1]);
  C3 I27 (simp251_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I28 (simp251_0[1:1], i_0r1[3:3]);
  C2 I29 (match0_0[5:5], simp251_0[0:0], simp251_0[1:1]);
  C3 I30 (simp261_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I31 (simp261_0[1:1], i_0r1[3:3]);
  C2 I32 (match0_0[6:6], simp261_0[0:0], simp261_0[1:1]);
  C3 I33 (simp271_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I34 (simp271_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I35 (match0_0[7:7], simp271_0[0:0], simp271_0[1:1]);
  C3 I36 (simp281_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I37 (simp281_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I38 (match0_0[8:8], simp281_0[0:0], simp281_0[1:1]);
  C3 I39 (simp291_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I40 (simp291_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I41 (match0_0[9:9], simp291_0[0:0], simp291_0[1:1]);
  C3 I42 (simp301_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I43 (simp301_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I44 (match0_0[10:10], simp301_0[0:0], simp301_0[1:1]);
  C3 I45 (simp311_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I46 (simp311_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I47 (match0_0[11:11], simp311_0[0:0], simp311_0[1:1]);
  C3 I48 (simp321_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I49 (simp321_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I50 (match0_0[12:12], simp321_0[0:0], simp321_0[1:1]);
  C3 I51 (simp331_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I52 (simp331_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I53 (match0_0[13:13], simp331_0[0:0], simp331_0[1:1]);
  C3 I54 (simp341_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I55 (simp341_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I56 (match0_0[14:14], simp341_0[0:0], simp341_0[1:1]);
  C3 I57 (simp351_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I58 (simp351_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I59 (match0_0[15:15], simp351_0[0:0], simp351_0[1:1]);
  C3 I60 (simp361_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I61 (simp361_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I62 (match0_0[16:16], simp361_0[0:0], simp361_0[1:1]);
  C3 I63 (simp371_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I64 (simp371_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I65 (match0_0[17:17], simp371_0[0:0], simp371_0[1:1]);
  C3 I66 (simp381_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I67 (simp381_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I68 (match0_0[18:18], simp381_0[0:0], simp381_0[1:1]);
  C3 I69 (simp391_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I70 (simp391_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I71 (match0_0[19:19], simp391_0[0:0], simp391_0[1:1]);
  C3 I72 (simp401_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I73 (simp401_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I74 (match0_0[20:20], simp401_0[0:0], simp401_0[1:1]);
  C3 I75 (simp411_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I76 (simp411_0[1:1], i_0r1[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I77 (match0_0[21:21], simp411_0[0:0], simp411_0[1:1]);
  C3 I78 (simp421_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I79 (simp421_0[1:1], i_0r1[3:3], i_0r1[4:4], i_0r1[5:5]);
  C2 I80 (match0_0[22:22], simp421_0[0:0], simp421_0[1:1]);
  NOR3 I81 (simp441_0[0:0], match1_0[0:0], match1_0[1:1], match1_0[2:2]);
  NOR3 I82 (simp441_0[1:1], match1_0[3:3], match1_0[4:4], match1_0[5:5]);
  INV I83 (simp441_0[2:2], match1_0[6:6]);
  NAND3 I84 (sel_1, simp441_0[0:0], simp441_0[1:1], simp441_0[2:2]);
  C3 I85 (simp451_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I86 (simp451_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I87 (match1_0[0:0], simp451_0[0:0], simp451_0[1:1]);
  C3 I88 (simp461_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I89 (simp461_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I90 (match1_0[1:1], simp461_0[0:0], simp461_0[1:1]);
  C3 I91 (simp471_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I92 (simp471_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I93 (match1_0[2:2], simp471_0[0:0], simp471_0[1:1]);
  C3 I94 (simp481_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I95 (simp481_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I96 (match1_0[3:3], simp481_0[0:0], simp481_0[1:1]);
  C3 I97 (simp491_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I98 (simp491_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I99 (match1_0[4:4], simp491_0[0:0], simp491_0[1:1]);
  C3 I100 (simp501_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I101 (simp501_0[1:1], i_0r1[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I102 (match1_0[5:5], simp501_0[0:0], simp501_0[1:1]);
  C3 I103 (simp511_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I104 (simp511_0[1:1], i_0r1[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I105 (match1_0[6:6], simp511_0[0:0], simp511_0[1:1]);
  NOR3 I106 (simp531_0[0:0], match2_0[0:0], match2_0[1:1], match2_0[2:2]);
  INV I107 (simp531_0[1:1], match2_0[3:3]);
  NAND2 I108 (sel_2, simp531_0[0:0], simp531_0[1:1]);
  C3 I109 (simp541_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I110 (simp541_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I111 (match2_0[0:0], simp541_0[0:0], simp541_0[1:1]);
  C3 I112 (simp551_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I113 (simp551_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I114 (match2_0[1:1], simp551_0[0:0], simp551_0[1:1]);
  C3 I115 (simp561_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I116 (simp561_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I117 (match2_0[2:2], simp561_0[0:0], simp561_0[1:1]);
  C3 I118 (simp571_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I119 (simp571_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I120 (match2_0[3:3], simp571_0[0:0], simp571_0[1:1]);
  NOR3 I121 (simp591_0[0:0], match3_0[0:0], match3_0[1:1], match3_0[2:2]);
  INV I122 (simp591_0[1:1], match3_0[3:3]);
  NAND2 I123 (sel_3, simp591_0[0:0], simp591_0[1:1]);
  C3 I124 (simp601_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I125 (simp601_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I126 (match3_0[0:0], simp601_0[0:0], simp601_0[1:1]);
  C3 I127 (simp611_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I128 (simp611_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I129 (match3_0[1:1], simp611_0[0:0], simp611_0[1:1]);
  C3 I130 (simp621_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I131 (simp621_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I132 (match3_0[2:2], simp621_0[0:0], simp621_0[1:1]);
  C3 I133 (simp631_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I134 (simp631_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I135 (match3_0[3:3], simp631_0[0:0], simp631_0[1:1]);
  NOR3 I136 (simp651_0[0:0], match4_0[0:0], match4_0[1:1], match4_0[2:2]);
  INV I137 (simp651_0[1:1], match4_0[3:3]);
  NAND2 I138 (sel_4, simp651_0[0:0], simp651_0[1:1]);
  C3 I139 (simp661_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I140 (simp661_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I141 (match4_0[0:0], simp661_0[0:0], simp661_0[1:1]);
  C3 I142 (simp671_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I143 (simp671_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I144 (match4_0[1:1], simp671_0[0:0], simp671_0[1:1]);
  C3 I145 (simp681_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I146 (simp681_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I147 (match4_0[2:2], simp681_0[0:0], simp681_0[1:1]);
  C3 I148 (simp691_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I149 (simp691_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I150 (match4_0[3:3], simp691_0[0:0], simp691_0[1:1]);
  BUFF I151 (sel_5, match5_0);
  C3 I152 (simp721_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I153 (simp721_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I154 (match5_0, simp721_0[0:0], simp721_0[1:1]);
  BUFF I155 (sel_6, match6_0);
  C3 I156 (simp751_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I157 (simp751_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I158 (match6_0, simp751_0[0:0], simp751_0[1:1]);
  BUFF I159 (sel_7, match7_0);
  C3 I160 (simp781_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I161 (simp781_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I162 (match7_0, simp781_0[0:0], simp781_0[1:1]);
  C2 I163 (gsel_0, sel_0, icomplete_0);
  C2 I164 (gsel_1, sel_1, icomplete_0);
  C2 I165 (gsel_2, sel_2, icomplete_0);
  C2 I166 (gsel_3, sel_3, icomplete_0);
  C2 I167 (gsel_4, sel_4, icomplete_0);
  C2 I168 (gsel_5, sel_5, icomplete_0);
  C2 I169 (gsel_6, sel_6, icomplete_0);
  C2 I170 (gsel_7, sel_7, icomplete_0);
  OR2 I171 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I172 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I173 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I174 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I175 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I176 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  C3 I177 (simp941_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I178 (simp941_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C2 I179 (icomplete_0, simp941_0[0:0], simp941_0[1:1]);
  BUFF I180 (o_0r, gsel_0);
  BUFF I181 (o_1r, gsel_1);
  BUFF I182 (o_2r, gsel_2);
  BUFF I183 (o_3r, gsel_3);
  BUFF I184 (o_4r, gsel_4);
  BUFF I185 (o_5r, gsel_5);
  BUFF I186 (o_6r, gsel_6);
  BUFF I187 (o_7r, gsel_7);
  NOR3 I188 (simp1031_0[0:0], o_0a, o_1a, o_2a);
  NOR3 I189 (simp1031_0[1:1], o_3a, o_4a, o_5a);
  NOR2 I190 (simp1031_0[2:2], o_6a, o_7a);
  NAND3 I191 (oack_0, simp1031_0[0:0], simp1031_0[1:1], simp1031_0[2:2]);
  C2 I192 (i_0a, oack_0, icomplete_0);
endmodule

// tkm8x0b TeakM [Many [0,0,0,0,0,0,0,0],One 0]
module tkm8x0b (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, i_3r, i_3a, i_4r, i_4a, i_5r, i_5a, i_6r, i_6a, i_7r, i_7a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  input i_4r;
  output i_4a;
  input i_5r;
  output i_5a;
  input i_6r;
  output i_6a;
  input i_7r;
  output i_7a;
  output o_0r;
  input o_0a;
  input reset;
  wire nchosen_0;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire choice_4;
  wire choice_5;
  wire choice_6;
  wire choice_7;
  wire [2:0] simp181_0;
  C2R I0 (choice_0, i_0r, nchosen_0, reset);
  C2R I1 (choice_1, i_1r, nchosen_0, reset);
  C2R I2 (choice_2, i_2r, nchosen_0, reset);
  C2R I3 (choice_3, i_3r, nchosen_0, reset);
  C2R I4 (choice_4, i_4r, nchosen_0, reset);
  C2R I5 (choice_5, i_5r, nchosen_0, reset);
  C2R I6 (choice_6, i_6r, nchosen_0, reset);
  C2R I7 (choice_7, i_7r, nchosen_0, reset);
  NOR2 I8 (nchosen_0, o_0r, o_0a);
  NOR3 I9 (simp181_0[0:0], choice_0, choice_1, choice_2);
  NOR3 I10 (simp181_0[1:1], choice_3, choice_4, choice_5);
  NOR2 I11 (simp181_0[2:2], choice_6, choice_7);
  NAND3 I12 (o_0r, simp181_0[0:0], simp181_0[1:1], simp181_0[2:2]);
  C2R I13 (i_0a, choice_0, o_0a, reset);
  C2R I14 (i_1a, choice_1, o_0a, reset);
  C2R I15 (i_2a, choice_2, o_0a, reset);
  C2R I16 (i_3a, choice_3, o_0a, reset);
  C2R I17 (i_4a, choice_4, o_0a, reset);
  C2R I18 (i_5a, choice_5, o_0a, reset);
  C2R I19 (i_6a, choice_6, o_0a, reset);
  C2R I20 (i_7a, choice_7, o_0a, reset);
endmodule

// tks6_o0w6_0c3cm1c38m2c38m3c38m5m6m7mdc30mec30mfc30m15c20m16c20m17c20o0w0_25m26m27o0w0 TeakS (0+:6) [
//   ([Imp 0 60,Imp 1 56,Imp 2 56,Imp 3 56,Imp 5 0,Imp 6 0,Imp 7 0,Imp 13 48,Imp 14 48,Imp 15 48,Imp 21 3
//   2,Imp 22 32,Imp 23 32],0),([Imp 37 0,Imp 38 0,Imp 39 0],0)] [One 6,Many [0,0]]
module tks6_o0w6_0c3cm1c38m2c38m3c38m5m6m7mdc30mec30mfc30m15c20m16c20m17c20o0w0_25m26m27o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, reset);
  input [5:0] i_0r0;
  input [5:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire [12:0] match0_0;
  wire [4:0] simp71_0;
  wire [1:0] simp72_0;
  wire [1:0] simp121_0;
  wire [1:0] simp131_0;
  wire [1:0] simp141_0;
  wire [1:0] simp151_0;
  wire [1:0] simp161_0;
  wire [1:0] simp171_0;
  wire [1:0] simp181_0;
  wire [1:0] simp191_0;
  wire [1:0] simp201_0;
  wire [2:0] match1_0;
  wire [1:0] simp231_0;
  wire [1:0] simp241_0;
  wire [1:0] simp251_0;
  wire [5:0] comp_0;
  wire [1:0] simp351_0;
  NOR3 I0 (simp71_0[0:0], match0_0[0:0], match0_0[1:1], match0_0[2:2]);
  NOR3 I1 (simp71_0[1:1], match0_0[3:3], match0_0[4:4], match0_0[5:5]);
  NOR3 I2 (simp71_0[2:2], match0_0[6:6], match0_0[7:7], match0_0[8:8]);
  NOR3 I3 (simp71_0[3:3], match0_0[9:9], match0_0[10:10], match0_0[11:11]);
  INV I4 (simp71_0[4:4], match0_0[12:12]);
  NAND3 I5 (simp72_0[0:0], simp71_0[0:0], simp71_0[1:1], simp71_0[2:2]);
  NAND2 I6 (simp72_0[1:1], simp71_0[3:3], simp71_0[4:4]);
  OR2 I7 (sel_0, simp72_0[0:0], simp72_0[1:1]);
  C2 I8 (match0_0[0:0], i_0r0[0:0], i_0r0[1:1]);
  C3 I9 (match0_0[1:1], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I10 (match0_0[2:2], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I11 (match0_0[3:3], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I12 (simp121_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I13 (simp121_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I14 (match0_0[4:4], simp121_0[0:0], simp121_0[1:1]);
  C3 I15 (simp131_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I16 (simp131_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I17 (match0_0[5:5], simp131_0[0:0], simp131_0[1:1]);
  C3 I18 (simp141_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I19 (simp141_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I20 (match0_0[6:6], simp141_0[0:0], simp141_0[1:1]);
  C3 I21 (simp151_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I22 (simp151_0[1:1], i_0r1[3:3]);
  C2 I23 (match0_0[7:7], simp151_0[0:0], simp151_0[1:1]);
  C3 I24 (simp161_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I25 (simp161_0[1:1], i_0r1[3:3]);
  C2 I26 (match0_0[8:8], simp161_0[0:0], simp161_0[1:1]);
  C3 I27 (simp171_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I28 (simp171_0[1:1], i_0r1[3:3]);
  C2 I29 (match0_0[9:9], simp171_0[0:0], simp171_0[1:1]);
  C3 I30 (simp181_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  C2 I31 (simp181_0[1:1], i_0r0[3:3], i_0r1[4:4]);
  C2 I32 (match0_0[10:10], simp181_0[0:0], simp181_0[1:1]);
  C3 I33 (simp191_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  C2 I34 (simp191_0[1:1], i_0r0[3:3], i_0r1[4:4]);
  C2 I35 (match0_0[11:11], simp191_0[0:0], simp191_0[1:1]);
  C3 I36 (simp201_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  C2 I37 (simp201_0[1:1], i_0r0[3:3], i_0r1[4:4]);
  C2 I38 (match0_0[12:12], simp201_0[0:0], simp201_0[1:1]);
  OR3 I39 (sel_1, match1_0[0:0], match1_0[1:1], match1_0[2:2]);
  C3 I40 (simp231_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I41 (simp231_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I42 (match1_0[0:0], simp231_0[0:0], simp231_0[1:1]);
  C3 I43 (simp241_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I44 (simp241_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I45 (match1_0[1:1], simp241_0[0:0], simp241_0[1:1]);
  C3 I46 (simp251_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  C3 I47 (simp251_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I48 (match1_0[2:2], simp251_0[0:0], simp251_0[1:1]);
  C2 I49 (gsel_0, sel_0, icomplete_0);
  C2 I50 (gsel_1, sel_1, icomplete_0);
  OR2 I51 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I52 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I53 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I54 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I55 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I56 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  C3 I57 (simp351_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I58 (simp351_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C2 I59 (icomplete_0, simp351_0[0:0], simp351_0[1:1]);
  BUFF I60 (o_0r, gsel_0);
  BUFF I61 (o_1r, gsel_1);
  OR2 I62 (oack_0, o_0a, o_1a);
  C2 I63 (i_0a, oack_0, icomplete_0);
endmodule

// tkvaddResult33_wo0w33_ro0w33 TeakV "addResult" 33 [] [0] [0] [Many [33],Many [0],Many [0],Many [33]]
module tkvaddResult33_wo0w33_ro0w33 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [32:0] wg_0r0;
  input [32:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [32:0] rd_0r0;
  output [32:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [32:0] wf_0;
  wire [32:0] wt_0;
  wire [32:0] df_0;
  wire [32:0] dt_0;
  wire wc_0;
  wire [32:0] wacks_0;
  wire [32:0] wenr_0;
  wire [32:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [32:0] drlgf_0;
  wire [32:0] drlgt_0;
  wire [32:0] comp0_0;
  wire [10:0] simp2451_0;
  wire [3:0] simp2452_0;
  wire [1:0] simp2453_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [32:0] conwgit_0;
  wire [32:0] conwgif_0;
  wire conwig_0;
  wire [11:0] simp4191_0;
  wire [3:0] simp4192_0;
  wire [1:0] simp4193_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (wen_0[32:32], wenr_0[32:32], nreset_0);
  AND2 I34 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I35 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I36 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I37 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I38 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I39 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I40 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I41 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I42 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I43 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I44 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I45 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I46 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I47 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I48 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I49 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I50 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I51 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I52 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I53 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I54 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I55 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I56 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I57 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I58 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I59 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I60 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I61 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I62 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I63 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I64 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I65 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I66 (drlgf_0[32:32], wf_0[32:32], wen_0[32:32]);
  AND2 I67 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I68 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I69 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I70 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I71 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I72 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I73 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I74 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I75 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I76 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I77 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I78 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I79 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I80 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I81 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I82 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I83 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I84 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I85 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I86 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I87 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I88 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I89 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I90 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I91 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I92 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I93 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I94 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I95 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I96 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I97 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I98 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  AND2 I99 (drlgt_0[32:32], wt_0[32:32], wen_0[32:32]);
  NOR2 I100 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I101 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I102 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I103 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I104 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I105 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I106 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I107 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I108 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I109 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I110 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I111 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I112 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I113 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I114 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I115 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I116 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I117 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I118 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I119 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I120 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I121 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I122 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I123 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I124 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I125 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I126 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I127 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I128 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I129 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I130 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I131 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR2 I132 (df_0[32:32], dt_0[32:32], drlgt_0[32:32]);
  NOR3 I133 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I134 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I135 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I136 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I137 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I138 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I139 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I140 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I141 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I142 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I143 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I144 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I145 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I146 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I147 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I148 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I149 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I150 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I151 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I152 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I153 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I154 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I155 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I156 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I157 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I158 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I159 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I160 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I161 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I162 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I163 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I164 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  NOR3 I165 (dt_0[32:32], df_0[32:32], drlgf_0[32:32], reset);
  AO22 I166 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I167 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I168 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I169 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I170 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I171 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I172 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I173 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I174 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I175 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I176 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I177 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I178 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I179 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I180 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I181 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I182 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I183 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I184 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I185 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I186 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I187 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I188 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I189 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I190 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I191 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I192 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I193 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I194 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I195 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I196 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I197 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  AO22 I198 (wacks_0[32:32], drlgf_0[32:32], df_0[32:32], drlgt_0[32:32], dt_0[32:32]);
  OR2 I199 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I200 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I201 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I202 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I203 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I204 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I205 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I206 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I207 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I208 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I209 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I210 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I211 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I212 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I213 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I214 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I215 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I216 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I217 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I218 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I219 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I220 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I221 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I222 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I223 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I224 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I225 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I226 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I227 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I228 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I229 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I230 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  OR2 I231 (comp0_0[32:32], wg_0r0[32:32], wg_0r1[32:32]);
  C3 I232 (simp2451_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I233 (simp2451_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I234 (simp2451_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I235 (simp2451_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I236 (simp2451_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I237 (simp2451_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I238 (simp2451_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I239 (simp2451_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I240 (simp2451_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I241 (simp2451_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C3 I242 (simp2451_0[10:10], comp0_0[30:30], comp0_0[31:31], comp0_0[32:32]);
  C3 I243 (simp2452_0[0:0], simp2451_0[0:0], simp2451_0[1:1], simp2451_0[2:2]);
  C3 I244 (simp2452_0[1:1], simp2451_0[3:3], simp2451_0[4:4], simp2451_0[5:5]);
  C3 I245 (simp2452_0[2:2], simp2451_0[6:6], simp2451_0[7:7], simp2451_0[8:8]);
  C2 I246 (simp2452_0[3:3], simp2451_0[9:9], simp2451_0[10:10]);
  C3 I247 (simp2453_0[0:0], simp2452_0[0:0], simp2452_0[1:1], simp2452_0[2:2]);
  BUFF I248 (simp2453_0[1:1], simp2452_0[3:3]);
  C2 I249 (wc_0, simp2453_0[0:0], simp2453_0[1:1]);
  AND2 I250 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I251 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I252 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I253 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I254 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I255 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I256 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I257 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I258 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I259 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I260 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I261 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I262 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I263 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I264 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I265 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I266 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I267 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I268 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I269 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I270 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I271 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I272 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I273 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I274 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I275 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I276 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I277 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I278 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I279 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I280 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I281 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I282 (conwgif_0[32:32], wg_0r0[32:32], conwig_0);
  AND2 I283 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I284 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I285 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I286 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I287 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I288 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I289 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I290 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I291 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I292 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I293 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I294 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I295 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I296 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I297 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I298 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I299 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I300 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I301 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I302 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I303 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I304 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I305 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I306 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I307 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I308 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I309 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I310 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I311 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I312 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I313 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I314 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  AND2 I315 (conwgit_0[32:32], wg_0r1[32:32], conwig_0);
  BUFF I316 (conwigc_0, wc_0);
  AO22 I317 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I318 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I319 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I320 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I321 (wenr_0[0:0], wc_0);
  BUFF I322 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I323 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I324 (wenr_0[1:1], wc_0);
  BUFF I325 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I326 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I327 (wenr_0[2:2], wc_0);
  BUFF I328 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I329 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I330 (wenr_0[3:3], wc_0);
  BUFF I331 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I332 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I333 (wenr_0[4:4], wc_0);
  BUFF I334 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I335 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I336 (wenr_0[5:5], wc_0);
  BUFF I337 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I338 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I339 (wenr_0[6:6], wc_0);
  BUFF I340 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I341 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I342 (wenr_0[7:7], wc_0);
  BUFF I343 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I344 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I345 (wenr_0[8:8], wc_0);
  BUFF I346 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I347 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I348 (wenr_0[9:9], wc_0);
  BUFF I349 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I350 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I351 (wenr_0[10:10], wc_0);
  BUFF I352 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I353 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I354 (wenr_0[11:11], wc_0);
  BUFF I355 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I356 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I357 (wenr_0[12:12], wc_0);
  BUFF I358 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I359 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I360 (wenr_0[13:13], wc_0);
  BUFF I361 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I362 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I363 (wenr_0[14:14], wc_0);
  BUFF I364 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I365 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I366 (wenr_0[15:15], wc_0);
  BUFF I367 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I368 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I369 (wenr_0[16:16], wc_0);
  BUFF I370 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I371 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I372 (wenr_0[17:17], wc_0);
  BUFF I373 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I374 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I375 (wenr_0[18:18], wc_0);
  BUFF I376 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I377 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I378 (wenr_0[19:19], wc_0);
  BUFF I379 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I380 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I381 (wenr_0[20:20], wc_0);
  BUFF I382 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I383 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I384 (wenr_0[21:21], wc_0);
  BUFF I385 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I386 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I387 (wenr_0[22:22], wc_0);
  BUFF I388 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I389 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I390 (wenr_0[23:23], wc_0);
  BUFF I391 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I392 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I393 (wenr_0[24:24], wc_0);
  BUFF I394 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I395 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I396 (wenr_0[25:25], wc_0);
  BUFF I397 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I398 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I399 (wenr_0[26:26], wc_0);
  BUFF I400 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I401 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I402 (wenr_0[27:27], wc_0);
  BUFF I403 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I404 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I405 (wenr_0[28:28], wc_0);
  BUFF I406 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I407 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I408 (wenr_0[29:29], wc_0);
  BUFF I409 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I410 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I411 (wenr_0[30:30], wc_0);
  BUFF I412 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I413 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I414 (wenr_0[31:31], wc_0);
  BUFF I415 (wf_0[32:32], conwgif_0[32:32]);
  BUFF I416 (wt_0[32:32], conwgit_0[32:32]);
  BUFF I417 (wenr_0[32:32], wc_0);
  C3 I418 (simp4191_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I419 (simp4191_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I420 (simp4191_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I421 (simp4191_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I422 (simp4191_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I423 (simp4191_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I424 (simp4191_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I425 (simp4191_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I426 (simp4191_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I427 (simp4191_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I428 (simp4191_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  BUFF I429 (simp4191_0[11:11], wacks_0[32:32]);
  C3 I430 (simp4192_0[0:0], simp4191_0[0:0], simp4191_0[1:1], simp4191_0[2:2]);
  C3 I431 (simp4192_0[1:1], simp4191_0[3:3], simp4191_0[4:4], simp4191_0[5:5]);
  C3 I432 (simp4192_0[2:2], simp4191_0[6:6], simp4191_0[7:7], simp4191_0[8:8]);
  C3 I433 (simp4192_0[3:3], simp4191_0[9:9], simp4191_0[10:10], simp4191_0[11:11]);
  C3 I434 (simp4193_0[0:0], simp4192_0[0:0], simp4192_0[1:1], simp4192_0[2:2]);
  BUFF I435 (simp4193_0[1:1], simp4192_0[3:3]);
  C2 I436 (wd_0r, simp4193_0[0:0], simp4193_0[1:1]);
  AND2 I437 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I438 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I439 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I440 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I441 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I442 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I443 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I444 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I445 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I446 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I447 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I448 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I449 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I450 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I451 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I452 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I453 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I454 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I455 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I456 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I457 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I458 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I459 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I460 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I461 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I462 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I463 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I464 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I465 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I466 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I467 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I468 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I469 (rd_0r0[32:32], df_0[32:32], rg_0r);
  AND2 I470 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I471 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I472 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I473 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I474 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I475 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I476 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I477 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I478 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I479 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I480 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I481 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I482 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I483 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I484 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I485 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I486 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I487 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I488 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I489 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I490 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I491 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I492 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I493 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I494 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I495 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I496 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I497 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I498 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I499 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I500 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I501 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I502 (rd_0r1[32:32], dt_0[32:32], rg_0r);
  OR2 I503 (anyread_0, rg_0r, rg_0a);
  BUFF I504 (wg_0a, wd_0a);
  BUFF I505 (rg_0a, rd_0a);
endmodule

// tkj33m0_33 TeakJ [Many [0,33],One 33]
module tkj33m0_33 (i_0r, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  input [32:0] i_1r0;
  input [32:0] i_1r1;
  output i_1a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [32:0] joinf_0;
  wire [32:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_1r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_1r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_1r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_1r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_1r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_1r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_1r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_1r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_1r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_1r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_1r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_1r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_1r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_1r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_1r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_1r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_1r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_1r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_1r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_1r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_1r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_1r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_1r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_1r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_1r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_1r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_1r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_1r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_1r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_1r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_1r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_1r0[31:31]);
  BUFF I32 (joinf_0[32:32], i_1r0[32:32]);
  BUFF I33 (joint_0[0:0], i_1r1[0:0]);
  BUFF I34 (joint_0[1:1], i_1r1[1:1]);
  BUFF I35 (joint_0[2:2], i_1r1[2:2]);
  BUFF I36 (joint_0[3:3], i_1r1[3:3]);
  BUFF I37 (joint_0[4:4], i_1r1[4:4]);
  BUFF I38 (joint_0[5:5], i_1r1[5:5]);
  BUFF I39 (joint_0[6:6], i_1r1[6:6]);
  BUFF I40 (joint_0[7:7], i_1r1[7:7]);
  BUFF I41 (joint_0[8:8], i_1r1[8:8]);
  BUFF I42 (joint_0[9:9], i_1r1[9:9]);
  BUFF I43 (joint_0[10:10], i_1r1[10:10]);
  BUFF I44 (joint_0[11:11], i_1r1[11:11]);
  BUFF I45 (joint_0[12:12], i_1r1[12:12]);
  BUFF I46 (joint_0[13:13], i_1r1[13:13]);
  BUFF I47 (joint_0[14:14], i_1r1[14:14]);
  BUFF I48 (joint_0[15:15], i_1r1[15:15]);
  BUFF I49 (joint_0[16:16], i_1r1[16:16]);
  BUFF I50 (joint_0[17:17], i_1r1[17:17]);
  BUFF I51 (joint_0[18:18], i_1r1[18:18]);
  BUFF I52 (joint_0[19:19], i_1r1[19:19]);
  BUFF I53 (joint_0[20:20], i_1r1[20:20]);
  BUFF I54 (joint_0[21:21], i_1r1[21:21]);
  BUFF I55 (joint_0[22:22], i_1r1[22:22]);
  BUFF I56 (joint_0[23:23], i_1r1[23:23]);
  BUFF I57 (joint_0[24:24], i_1r1[24:24]);
  BUFF I58 (joint_0[25:25], i_1r1[25:25]);
  BUFF I59 (joint_0[26:26], i_1r1[26:26]);
  BUFF I60 (joint_0[27:27], i_1r1[27:27]);
  BUFF I61 (joint_0[28:28], i_1r1[28:28]);
  BUFF I62 (joint_0[29:29], i_1r1[29:29]);
  BUFF I63 (joint_0[30:30], i_1r1[30:30]);
  BUFF I64 (joint_0[31:31], i_1r1[31:31]);
  BUFF I65 (joint_0[32:32], i_1r1[32:32]);
  BUFF I66 (icomplete_0, i_0r);
  C2 I67 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I68 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I69 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I70 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I71 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I72 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I73 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I74 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I75 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I76 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I77 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I78 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I79 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I80 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I81 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I82 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I83 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I84 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I85 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I86 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I87 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I88 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I89 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I90 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I91 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I92 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I93 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I94 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I95 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I96 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I97 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I98 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I99 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I100 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I101 (o_0r1[1:1], joint_0[1:1]);
  BUFF I102 (o_0r1[2:2], joint_0[2:2]);
  BUFF I103 (o_0r1[3:3], joint_0[3:3]);
  BUFF I104 (o_0r1[4:4], joint_0[4:4]);
  BUFF I105 (o_0r1[5:5], joint_0[5:5]);
  BUFF I106 (o_0r1[6:6], joint_0[6:6]);
  BUFF I107 (o_0r1[7:7], joint_0[7:7]);
  BUFF I108 (o_0r1[8:8], joint_0[8:8]);
  BUFF I109 (o_0r1[9:9], joint_0[9:9]);
  BUFF I110 (o_0r1[10:10], joint_0[10:10]);
  BUFF I111 (o_0r1[11:11], joint_0[11:11]);
  BUFF I112 (o_0r1[12:12], joint_0[12:12]);
  BUFF I113 (o_0r1[13:13], joint_0[13:13]);
  BUFF I114 (o_0r1[14:14], joint_0[14:14]);
  BUFF I115 (o_0r1[15:15], joint_0[15:15]);
  BUFF I116 (o_0r1[16:16], joint_0[16:16]);
  BUFF I117 (o_0r1[17:17], joint_0[17:17]);
  BUFF I118 (o_0r1[18:18], joint_0[18:18]);
  BUFF I119 (o_0r1[19:19], joint_0[19:19]);
  BUFF I120 (o_0r1[20:20], joint_0[20:20]);
  BUFF I121 (o_0r1[21:21], joint_0[21:21]);
  BUFF I122 (o_0r1[22:22], joint_0[22:22]);
  BUFF I123 (o_0r1[23:23], joint_0[23:23]);
  BUFF I124 (o_0r1[24:24], joint_0[24:24]);
  BUFF I125 (o_0r1[25:25], joint_0[25:25]);
  BUFF I126 (o_0r1[26:26], joint_0[26:26]);
  BUFF I127 (o_0r1[27:27], joint_0[27:27]);
  BUFF I128 (o_0r1[28:28], joint_0[28:28]);
  BUFF I129 (o_0r1[29:29], joint_0[29:29]);
  BUFF I130 (o_0r1[30:30], joint_0[30:30]);
  BUFF I131 (o_0r1[31:31], joint_0[31:31]);
  BUFF I132 (o_0r1[32:32], joint_0[32:32]);
  BUFF I133 (i_0a, o_0a);
  BUFF I134 (i_1a, o_0a);
endmodule

// tkvlogicResult32_wo0w32_ro0w32 TeakV "logicResult" 32 [] [0] [0] [Many [32],Many [0],Many [0],Many [
//   32]]
module tkvlogicResult32_wo0w32_ro0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I457 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I458 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I459 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I460 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I461 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I462 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I463 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I464 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I465 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I466 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I467 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I468 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I469 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I470 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I471 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I472 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I473 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I474 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I475 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I476 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I477 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I478 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I479 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I480 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I481 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I482 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I483 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I484 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I485 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I486 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I487 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  OR2 I488 (anyread_0, rg_0r, rg_0a);
  BUFF I489 (wg_0a, wd_0a);
  BUFF I490 (rg_0a, rd_0a);
endmodule

// tkj32m0_32 TeakJ [Many [0,32],One 32]
module tkj32m0_32 (i_0r, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [31:0] joinf_0;
  wire [31:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_1r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_1r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_1r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_1r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_1r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_1r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_1r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_1r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_1r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_1r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_1r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_1r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_1r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_1r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_1r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_1r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_1r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_1r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_1r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_1r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_1r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_1r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_1r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_1r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_1r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_1r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_1r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_1r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_1r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_1r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_1r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_1r0[31:31]);
  BUFF I32 (joint_0[0:0], i_1r1[0:0]);
  BUFF I33 (joint_0[1:1], i_1r1[1:1]);
  BUFF I34 (joint_0[2:2], i_1r1[2:2]);
  BUFF I35 (joint_0[3:3], i_1r1[3:3]);
  BUFF I36 (joint_0[4:4], i_1r1[4:4]);
  BUFF I37 (joint_0[5:5], i_1r1[5:5]);
  BUFF I38 (joint_0[6:6], i_1r1[6:6]);
  BUFF I39 (joint_0[7:7], i_1r1[7:7]);
  BUFF I40 (joint_0[8:8], i_1r1[8:8]);
  BUFF I41 (joint_0[9:9], i_1r1[9:9]);
  BUFF I42 (joint_0[10:10], i_1r1[10:10]);
  BUFF I43 (joint_0[11:11], i_1r1[11:11]);
  BUFF I44 (joint_0[12:12], i_1r1[12:12]);
  BUFF I45 (joint_0[13:13], i_1r1[13:13]);
  BUFF I46 (joint_0[14:14], i_1r1[14:14]);
  BUFF I47 (joint_0[15:15], i_1r1[15:15]);
  BUFF I48 (joint_0[16:16], i_1r1[16:16]);
  BUFF I49 (joint_0[17:17], i_1r1[17:17]);
  BUFF I50 (joint_0[18:18], i_1r1[18:18]);
  BUFF I51 (joint_0[19:19], i_1r1[19:19]);
  BUFF I52 (joint_0[20:20], i_1r1[20:20]);
  BUFF I53 (joint_0[21:21], i_1r1[21:21]);
  BUFF I54 (joint_0[22:22], i_1r1[22:22]);
  BUFF I55 (joint_0[23:23], i_1r1[23:23]);
  BUFF I56 (joint_0[24:24], i_1r1[24:24]);
  BUFF I57 (joint_0[25:25], i_1r1[25:25]);
  BUFF I58 (joint_0[26:26], i_1r1[26:26]);
  BUFF I59 (joint_0[27:27], i_1r1[27:27]);
  BUFF I60 (joint_0[28:28], i_1r1[28:28]);
  BUFF I61 (joint_0[29:29], i_1r1[29:29]);
  BUFF I62 (joint_0[30:30], i_1r1[30:30]);
  BUFF I63 (joint_0[31:31], i_1r1[31:31]);
  BUFF I64 (icomplete_0, i_0r);
  C2 I65 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I66 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I67 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I68 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I69 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I70 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I71 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I72 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I73 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I74 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I75 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I76 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I77 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I78 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I79 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I80 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I81 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I82 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I83 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I84 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I85 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I86 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I87 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I88 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I89 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I90 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I91 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I92 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I93 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I94 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I95 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I96 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I97 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I98 (o_0r1[1:1], joint_0[1:1]);
  BUFF I99 (o_0r1[2:2], joint_0[2:2]);
  BUFF I100 (o_0r1[3:3], joint_0[3:3]);
  BUFF I101 (o_0r1[4:4], joint_0[4:4]);
  BUFF I102 (o_0r1[5:5], joint_0[5:5]);
  BUFF I103 (o_0r1[6:6], joint_0[6:6]);
  BUFF I104 (o_0r1[7:7], joint_0[7:7]);
  BUFF I105 (o_0r1[8:8], joint_0[8:8]);
  BUFF I106 (o_0r1[9:9], joint_0[9:9]);
  BUFF I107 (o_0r1[10:10], joint_0[10:10]);
  BUFF I108 (o_0r1[11:11], joint_0[11:11]);
  BUFF I109 (o_0r1[12:12], joint_0[12:12]);
  BUFF I110 (o_0r1[13:13], joint_0[13:13]);
  BUFF I111 (o_0r1[14:14], joint_0[14:14]);
  BUFF I112 (o_0r1[15:15], joint_0[15:15]);
  BUFF I113 (o_0r1[16:16], joint_0[16:16]);
  BUFF I114 (o_0r1[17:17], joint_0[17:17]);
  BUFF I115 (o_0r1[18:18], joint_0[18:18]);
  BUFF I116 (o_0r1[19:19], joint_0[19:19]);
  BUFF I117 (o_0r1[20:20], joint_0[20:20]);
  BUFF I118 (o_0r1[21:21], joint_0[21:21]);
  BUFF I119 (o_0r1[22:22], joint_0[22:22]);
  BUFF I120 (o_0r1[23:23], joint_0[23:23]);
  BUFF I121 (o_0r1[24:24], joint_0[24:24]);
  BUFF I122 (o_0r1[25:25], joint_0[25:25]);
  BUFF I123 (o_0r1[26:26], joint_0[26:26]);
  BUFF I124 (o_0r1[27:27], joint_0[27:27]);
  BUFF I125 (o_0r1[28:28], joint_0[28:28]);
  BUFF I126 (o_0r1[29:29], joint_0[29:29]);
  BUFF I127 (o_0r1[30:30], joint_0[30:30]);
  BUFF I128 (o_0r1[31:31], joint_0[31:31]);
  BUFF I129 (i_0a, o_0a);
  BUFF I130 (i_1a, o_0a);
endmodule

// tkvshiftResult32_wo0w32_ro0w32 TeakV "shiftResult" 32 [] [0] [0] [Many [32],Many [0],Many [0],Many [
//   32]]
module tkvshiftResult32_wo0w32_ro0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I457 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I458 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I459 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I460 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I461 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I462 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I463 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I464 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I465 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I466 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I467 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I468 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I469 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I470 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I471 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I472 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I473 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I474 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I475 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I476 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I477 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I478 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I479 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I480 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I481 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I482 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I483 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I484 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I485 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I486 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I487 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  OR2 I488 (anyread_0, rg_0r, rg_0a);
  BUFF I489 (wg_0a, wd_0a);
  BUFF I490 (rg_0a, rd_0a);
endmodule

// tko33m1_1api0w32b_2api32w1b_3nm31b0_4apt2o0w1bt3o0w31b_5eqt1o0w32bt4o0w32b TeakO [
//     (1,TeakOAppend 1 [(0,0+:32)]),
//     (2,TeakOAppend 1 [(0,32+:1)]),
//     (3,TeakOConstant 31 0),
//     (4,TeakOAppend 1 [(2,0+:1),(3,0+:31)]),
//     (5,TeakOp TeakOpEqual [(1,0+:32),(4,0+:32)])] [One 33,One 1]
module tko33m1_1api0w32b_2api32w1b_3nm31b0_4apt2o0w1bt3o0w31b_5eqt1o0w32bt4o0w32b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [32:0] i_0r0;
  input [32:0] i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [32:0] gocomp_0;
  wire [10:0] simp351_0;
  wire [3:0] simp352_0;
  wire [1:0] simp353_0;
  wire [31:0] termf_1;
  wire termf_2;
  wire [30:0] termf_3;
  wire [31:0] termf_4;
  wire [31:0] termt_1;
  wire termt_2;
  wire [30:0] termt_3;
  wire [31:0] termt_4;
  wire [31:0] xf5_0;
  wire [31:0] xt5_0;
  wire [3:0] op5_0_0;
  wire [3:0] op5_1_0;
  wire [3:0] op5_2_0;
  wire [3:0] op5_3_0;
  wire [3:0] op5_4_0;
  wire [3:0] op5_5_0;
  wire [3:0] op5_6_0;
  wire [3:0] op5_7_0;
  wire [3:0] op5_8_0;
  wire [3:0] op5_9_0;
  wire [3:0] op5_10_0;
  wire [3:0] op5_11_0;
  wire [3:0] op5_12_0;
  wire [3:0] op5_13_0;
  wire [3:0] op5_14_0;
  wire [3:0] op5_15_0;
  wire [3:0] op5_16_0;
  wire [3:0] op5_17_0;
  wire [3:0] op5_18_0;
  wire [3:0] op5_19_0;
  wire [3:0] op5_20_0;
  wire [3:0] op5_21_0;
  wire [3:0] op5_22_0;
  wire [3:0] op5_23_0;
  wire [3:0] op5_24_0;
  wire [3:0] op5_25_0;
  wire [3:0] op5_26_0;
  wire [3:0] op5_27_0;
  wire [3:0] op5_28_0;
  wire [3:0] op5_29_0;
  wire [3:0] op5_30_0;
  wire [3:0] op5_31_0;
  wire [15:0] c5o_0;
  wire [15:0] c5o_1;
  wire [7:0] c5ro_0;
  wire [7:0] c5ro_1;
  wire [3:0] c5rro_0;
  wire [3:0] c5rro_1;
  wire [1:0] c5rrro_0;
  wire [1:0] c5rrro_1;
  wire [3:0] c5rrrr0_0;
  wire [3:0] c5rrr0_0;
  wire [3:0] c5rrr1_0;
  wire [3:0] c5rr0_0;
  wire [3:0] c5rr1_0;
  wire [3:0] c5rr2_0;
  wire [3:0] c5rr3_0;
  wire [3:0] c5r0_0;
  wire [3:0] c5r1_0;
  wire [3:0] c5r2_0;
  wire [3:0] c5r3_0;
  wire [3:0] c5r4_0;
  wire [3:0] c5r5_0;
  wire [3:0] c5r6_0;
  wire [3:0] c5r7_0;
  wire [3:0] c50_0;
  wire [3:0] c51_0;
  wire [3:0] c52_0;
  wire [3:0] c53_0;
  wire [3:0] c54_0;
  wire [3:0] c55_0;
  wire [3:0] c56_0;
  wire [3:0] c57_0;
  wire [3:0] c58_0;
  wire [3:0] c59_0;
  wire [3:0] c510_0;
  wire [3:0] c511_0;
  wire [3:0] c512_0;
  wire [3:0] c513_0;
  wire [3:0] c514_0;
  wire [3:0] c515_0;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I30 (gocomp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I31 (gocomp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I32 (gocomp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  C3 I33 (simp351_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  C3 I34 (simp351_0[1:1], gocomp_0[3:3], gocomp_0[4:4], gocomp_0[5:5]);
  C3 I35 (simp351_0[2:2], gocomp_0[6:6], gocomp_0[7:7], gocomp_0[8:8]);
  C3 I36 (simp351_0[3:3], gocomp_0[9:9], gocomp_0[10:10], gocomp_0[11:11]);
  C3 I37 (simp351_0[4:4], gocomp_0[12:12], gocomp_0[13:13], gocomp_0[14:14]);
  C3 I38 (simp351_0[5:5], gocomp_0[15:15], gocomp_0[16:16], gocomp_0[17:17]);
  C3 I39 (simp351_0[6:6], gocomp_0[18:18], gocomp_0[19:19], gocomp_0[20:20]);
  C3 I40 (simp351_0[7:7], gocomp_0[21:21], gocomp_0[22:22], gocomp_0[23:23]);
  C3 I41 (simp351_0[8:8], gocomp_0[24:24], gocomp_0[25:25], gocomp_0[26:26]);
  C3 I42 (simp351_0[9:9], gocomp_0[27:27], gocomp_0[28:28], gocomp_0[29:29]);
  C3 I43 (simp351_0[10:10], gocomp_0[30:30], gocomp_0[31:31], gocomp_0[32:32]);
  C3 I44 (simp352_0[0:0], simp351_0[0:0], simp351_0[1:1], simp351_0[2:2]);
  C3 I45 (simp352_0[1:1], simp351_0[3:3], simp351_0[4:4], simp351_0[5:5]);
  C3 I46 (simp352_0[2:2], simp351_0[6:6], simp351_0[7:7], simp351_0[8:8]);
  C2 I47 (simp352_0[3:3], simp351_0[9:9], simp351_0[10:10]);
  C3 I48 (simp353_0[0:0], simp352_0[0:0], simp352_0[1:1], simp352_0[2:2]);
  BUFF I49 (simp353_0[1:1], simp352_0[3:3]);
  C2 I50 (go_0, simp353_0[0:0], simp353_0[1:1]);
  BUFF I51 (termf_1[0:0], i_0r0[0:0]);
  BUFF I52 (termf_1[1:1], i_0r0[1:1]);
  BUFF I53 (termf_1[2:2], i_0r0[2:2]);
  BUFF I54 (termf_1[3:3], i_0r0[3:3]);
  BUFF I55 (termf_1[4:4], i_0r0[4:4]);
  BUFF I56 (termf_1[5:5], i_0r0[5:5]);
  BUFF I57 (termf_1[6:6], i_0r0[6:6]);
  BUFF I58 (termf_1[7:7], i_0r0[7:7]);
  BUFF I59 (termf_1[8:8], i_0r0[8:8]);
  BUFF I60 (termf_1[9:9], i_0r0[9:9]);
  BUFF I61 (termf_1[10:10], i_0r0[10:10]);
  BUFF I62 (termf_1[11:11], i_0r0[11:11]);
  BUFF I63 (termf_1[12:12], i_0r0[12:12]);
  BUFF I64 (termf_1[13:13], i_0r0[13:13]);
  BUFF I65 (termf_1[14:14], i_0r0[14:14]);
  BUFF I66 (termf_1[15:15], i_0r0[15:15]);
  BUFF I67 (termf_1[16:16], i_0r0[16:16]);
  BUFF I68 (termf_1[17:17], i_0r0[17:17]);
  BUFF I69 (termf_1[18:18], i_0r0[18:18]);
  BUFF I70 (termf_1[19:19], i_0r0[19:19]);
  BUFF I71 (termf_1[20:20], i_0r0[20:20]);
  BUFF I72 (termf_1[21:21], i_0r0[21:21]);
  BUFF I73 (termf_1[22:22], i_0r0[22:22]);
  BUFF I74 (termf_1[23:23], i_0r0[23:23]);
  BUFF I75 (termf_1[24:24], i_0r0[24:24]);
  BUFF I76 (termf_1[25:25], i_0r0[25:25]);
  BUFF I77 (termf_1[26:26], i_0r0[26:26]);
  BUFF I78 (termf_1[27:27], i_0r0[27:27]);
  BUFF I79 (termf_1[28:28], i_0r0[28:28]);
  BUFF I80 (termf_1[29:29], i_0r0[29:29]);
  BUFF I81 (termf_1[30:30], i_0r0[30:30]);
  BUFF I82 (termf_1[31:31], i_0r0[31:31]);
  BUFF I83 (termt_1[0:0], i_0r1[0:0]);
  BUFF I84 (termt_1[1:1], i_0r1[1:1]);
  BUFF I85 (termt_1[2:2], i_0r1[2:2]);
  BUFF I86 (termt_1[3:3], i_0r1[3:3]);
  BUFF I87 (termt_1[4:4], i_0r1[4:4]);
  BUFF I88 (termt_1[5:5], i_0r1[5:5]);
  BUFF I89 (termt_1[6:6], i_0r1[6:6]);
  BUFF I90 (termt_1[7:7], i_0r1[7:7]);
  BUFF I91 (termt_1[8:8], i_0r1[8:8]);
  BUFF I92 (termt_1[9:9], i_0r1[9:9]);
  BUFF I93 (termt_1[10:10], i_0r1[10:10]);
  BUFF I94 (termt_1[11:11], i_0r1[11:11]);
  BUFF I95 (termt_1[12:12], i_0r1[12:12]);
  BUFF I96 (termt_1[13:13], i_0r1[13:13]);
  BUFF I97 (termt_1[14:14], i_0r1[14:14]);
  BUFF I98 (termt_1[15:15], i_0r1[15:15]);
  BUFF I99 (termt_1[16:16], i_0r1[16:16]);
  BUFF I100 (termt_1[17:17], i_0r1[17:17]);
  BUFF I101 (termt_1[18:18], i_0r1[18:18]);
  BUFF I102 (termt_1[19:19], i_0r1[19:19]);
  BUFF I103 (termt_1[20:20], i_0r1[20:20]);
  BUFF I104 (termt_1[21:21], i_0r1[21:21]);
  BUFF I105 (termt_1[22:22], i_0r1[22:22]);
  BUFF I106 (termt_1[23:23], i_0r1[23:23]);
  BUFF I107 (termt_1[24:24], i_0r1[24:24]);
  BUFF I108 (termt_1[25:25], i_0r1[25:25]);
  BUFF I109 (termt_1[26:26], i_0r1[26:26]);
  BUFF I110 (termt_1[27:27], i_0r1[27:27]);
  BUFF I111 (termt_1[28:28], i_0r1[28:28]);
  BUFF I112 (termt_1[29:29], i_0r1[29:29]);
  BUFF I113 (termt_1[30:30], i_0r1[30:30]);
  BUFF I114 (termt_1[31:31], i_0r1[31:31]);
  BUFF I115 (termf_2, i_0r0[32:32]);
  BUFF I116 (termt_2, i_0r1[32:32]);
  BUFF I117 (termf_3[0:0], go_0);
  BUFF I118 (termf_3[1:1], go_0);
  BUFF I119 (termf_3[2:2], go_0);
  BUFF I120 (termf_3[3:3], go_0);
  BUFF I121 (termf_3[4:4], go_0);
  BUFF I122 (termf_3[5:5], go_0);
  BUFF I123 (termf_3[6:6], go_0);
  BUFF I124 (termf_3[7:7], go_0);
  BUFF I125 (termf_3[8:8], go_0);
  BUFF I126 (termf_3[9:9], go_0);
  BUFF I127 (termf_3[10:10], go_0);
  BUFF I128 (termf_3[11:11], go_0);
  BUFF I129 (termf_3[12:12], go_0);
  BUFF I130 (termf_3[13:13], go_0);
  BUFF I131 (termf_3[14:14], go_0);
  BUFF I132 (termf_3[15:15], go_0);
  BUFF I133 (termf_3[16:16], go_0);
  BUFF I134 (termf_3[17:17], go_0);
  BUFF I135 (termf_3[18:18], go_0);
  BUFF I136 (termf_3[19:19], go_0);
  BUFF I137 (termf_3[20:20], go_0);
  BUFF I138 (termf_3[21:21], go_0);
  BUFF I139 (termf_3[22:22], go_0);
  BUFF I140 (termf_3[23:23], go_0);
  BUFF I141 (termf_3[24:24], go_0);
  BUFF I142 (termf_3[25:25], go_0);
  BUFF I143 (termf_3[26:26], go_0);
  BUFF I144 (termf_3[27:27], go_0);
  BUFF I145 (termf_3[28:28], go_0);
  BUFF I146 (termf_3[29:29], go_0);
  BUFF I147 (termf_3[30:30], go_0);
  GND I148 (termt_3[0:0]);
  GND I149 (termt_3[1:1]);
  GND I150 (termt_3[2:2]);
  GND I151 (termt_3[3:3]);
  GND I152 (termt_3[4:4]);
  GND I153 (termt_3[5:5]);
  GND I154 (termt_3[6:6]);
  GND I155 (termt_3[7:7]);
  GND I156 (termt_3[8:8]);
  GND I157 (termt_3[9:9]);
  GND I158 (termt_3[10:10]);
  GND I159 (termt_3[11:11]);
  GND I160 (termt_3[12:12]);
  GND I161 (termt_3[13:13]);
  GND I162 (termt_3[14:14]);
  GND I163 (termt_3[15:15]);
  GND I164 (termt_3[16:16]);
  GND I165 (termt_3[17:17]);
  GND I166 (termt_3[18:18]);
  GND I167 (termt_3[19:19]);
  GND I168 (termt_3[20:20]);
  GND I169 (termt_3[21:21]);
  GND I170 (termt_3[22:22]);
  GND I171 (termt_3[23:23]);
  GND I172 (termt_3[24:24]);
  GND I173 (termt_3[25:25]);
  GND I174 (termt_3[26:26]);
  GND I175 (termt_3[27:27]);
  GND I176 (termt_3[28:28]);
  GND I177 (termt_3[29:29]);
  GND I178 (termt_3[30:30]);
  BUFF I179 (termf_4[0:0], termf_2);
  BUFF I180 (termf_4[1:1], termf_3[0:0]);
  BUFF I181 (termf_4[2:2], termf_3[1:1]);
  BUFF I182 (termf_4[3:3], termf_3[2:2]);
  BUFF I183 (termf_4[4:4], termf_3[3:3]);
  BUFF I184 (termf_4[5:5], termf_3[4:4]);
  BUFF I185 (termf_4[6:6], termf_3[5:5]);
  BUFF I186 (termf_4[7:7], termf_3[6:6]);
  BUFF I187 (termf_4[8:8], termf_3[7:7]);
  BUFF I188 (termf_4[9:9], termf_3[8:8]);
  BUFF I189 (termf_4[10:10], termf_3[9:9]);
  BUFF I190 (termf_4[11:11], termf_3[10:10]);
  BUFF I191 (termf_4[12:12], termf_3[11:11]);
  BUFF I192 (termf_4[13:13], termf_3[12:12]);
  BUFF I193 (termf_4[14:14], termf_3[13:13]);
  BUFF I194 (termf_4[15:15], termf_3[14:14]);
  BUFF I195 (termf_4[16:16], termf_3[15:15]);
  BUFF I196 (termf_4[17:17], termf_3[16:16]);
  BUFF I197 (termf_4[18:18], termf_3[17:17]);
  BUFF I198 (termf_4[19:19], termf_3[18:18]);
  BUFF I199 (termf_4[20:20], termf_3[19:19]);
  BUFF I200 (termf_4[21:21], termf_3[20:20]);
  BUFF I201 (termf_4[22:22], termf_3[21:21]);
  BUFF I202 (termf_4[23:23], termf_3[22:22]);
  BUFF I203 (termf_4[24:24], termf_3[23:23]);
  BUFF I204 (termf_4[25:25], termf_3[24:24]);
  BUFF I205 (termf_4[26:26], termf_3[25:25]);
  BUFF I206 (termf_4[27:27], termf_3[26:26]);
  BUFF I207 (termf_4[28:28], termf_3[27:27]);
  BUFF I208 (termf_4[29:29], termf_3[28:28]);
  BUFF I209 (termf_4[30:30], termf_3[29:29]);
  BUFF I210 (termf_4[31:31], termf_3[30:30]);
  BUFF I211 (termt_4[0:0], termt_2);
  BUFF I212 (termt_4[1:1], termt_3[0:0]);
  BUFF I213 (termt_4[2:2], termt_3[1:1]);
  BUFF I214 (termt_4[3:3], termt_3[2:2]);
  BUFF I215 (termt_4[4:4], termt_3[3:3]);
  BUFF I216 (termt_4[5:5], termt_3[4:4]);
  BUFF I217 (termt_4[6:6], termt_3[5:5]);
  BUFF I218 (termt_4[7:7], termt_3[6:6]);
  BUFF I219 (termt_4[8:8], termt_3[7:7]);
  BUFF I220 (termt_4[9:9], termt_3[8:8]);
  BUFF I221 (termt_4[10:10], termt_3[9:9]);
  BUFF I222 (termt_4[11:11], termt_3[10:10]);
  BUFF I223 (termt_4[12:12], termt_3[11:11]);
  BUFF I224 (termt_4[13:13], termt_3[12:12]);
  BUFF I225 (termt_4[14:14], termt_3[13:13]);
  BUFF I226 (termt_4[15:15], termt_3[14:14]);
  BUFF I227 (termt_4[16:16], termt_3[15:15]);
  BUFF I228 (termt_4[17:17], termt_3[16:16]);
  BUFF I229 (termt_4[18:18], termt_3[17:17]);
  BUFF I230 (termt_4[19:19], termt_3[18:18]);
  BUFF I231 (termt_4[20:20], termt_3[19:19]);
  BUFF I232 (termt_4[21:21], termt_3[20:20]);
  BUFF I233 (termt_4[22:22], termt_3[21:21]);
  BUFF I234 (termt_4[23:23], termt_3[22:22]);
  BUFF I235 (termt_4[24:24], termt_3[23:23]);
  BUFF I236 (termt_4[25:25], termt_3[24:24]);
  BUFF I237 (termt_4[26:26], termt_3[25:25]);
  BUFF I238 (termt_4[27:27], termt_3[26:26]);
  BUFF I239 (termt_4[28:28], termt_3[27:27]);
  BUFF I240 (termt_4[29:29], termt_3[28:28]);
  BUFF I241 (termt_4[30:30], termt_3[29:29]);
  BUFF I242 (termt_4[31:31], termt_3[30:30]);
  C2 I243 (op5_0_0[0:0], termf_4[0:0], termf_1[0:0]);
  C2 I244 (op5_0_0[1:1], termf_4[0:0], termt_1[0:0]);
  C2 I245 (op5_0_0[2:2], termt_4[0:0], termf_1[0:0]);
  C2 I246 (op5_0_0[3:3], termt_4[0:0], termt_1[0:0]);
  OR2 I247 (xf5_0[0:0], op5_0_0[1:1], op5_0_0[2:2]);
  OR2 I248 (xt5_0[0:0], op5_0_0[0:0], op5_0_0[3:3]);
  C2 I249 (op5_1_0[0:0], termf_4[1:1], termf_1[1:1]);
  C2 I250 (op5_1_0[1:1], termf_4[1:1], termt_1[1:1]);
  C2 I251 (op5_1_0[2:2], termt_4[1:1], termf_1[1:1]);
  C2 I252 (op5_1_0[3:3], termt_4[1:1], termt_1[1:1]);
  OR2 I253 (xf5_0[1:1], op5_1_0[1:1], op5_1_0[2:2]);
  OR2 I254 (xt5_0[1:1], op5_1_0[0:0], op5_1_0[3:3]);
  C2 I255 (op5_2_0[0:0], termf_4[2:2], termf_1[2:2]);
  C2 I256 (op5_2_0[1:1], termf_4[2:2], termt_1[2:2]);
  C2 I257 (op5_2_0[2:2], termt_4[2:2], termf_1[2:2]);
  C2 I258 (op5_2_0[3:3], termt_4[2:2], termt_1[2:2]);
  OR2 I259 (xf5_0[2:2], op5_2_0[1:1], op5_2_0[2:2]);
  OR2 I260 (xt5_0[2:2], op5_2_0[0:0], op5_2_0[3:3]);
  C2 I261 (op5_3_0[0:0], termf_4[3:3], termf_1[3:3]);
  C2 I262 (op5_3_0[1:1], termf_4[3:3], termt_1[3:3]);
  C2 I263 (op5_3_0[2:2], termt_4[3:3], termf_1[3:3]);
  C2 I264 (op5_3_0[3:3], termt_4[3:3], termt_1[3:3]);
  OR2 I265 (xf5_0[3:3], op5_3_0[1:1], op5_3_0[2:2]);
  OR2 I266 (xt5_0[3:3], op5_3_0[0:0], op5_3_0[3:3]);
  C2 I267 (op5_4_0[0:0], termf_4[4:4], termf_1[4:4]);
  C2 I268 (op5_4_0[1:1], termf_4[4:4], termt_1[4:4]);
  C2 I269 (op5_4_0[2:2], termt_4[4:4], termf_1[4:4]);
  C2 I270 (op5_4_0[3:3], termt_4[4:4], termt_1[4:4]);
  OR2 I271 (xf5_0[4:4], op5_4_0[1:1], op5_4_0[2:2]);
  OR2 I272 (xt5_0[4:4], op5_4_0[0:0], op5_4_0[3:3]);
  C2 I273 (op5_5_0[0:0], termf_4[5:5], termf_1[5:5]);
  C2 I274 (op5_5_0[1:1], termf_4[5:5], termt_1[5:5]);
  C2 I275 (op5_5_0[2:2], termt_4[5:5], termf_1[5:5]);
  C2 I276 (op5_5_0[3:3], termt_4[5:5], termt_1[5:5]);
  OR2 I277 (xf5_0[5:5], op5_5_0[1:1], op5_5_0[2:2]);
  OR2 I278 (xt5_0[5:5], op5_5_0[0:0], op5_5_0[3:3]);
  C2 I279 (op5_6_0[0:0], termf_4[6:6], termf_1[6:6]);
  C2 I280 (op5_6_0[1:1], termf_4[6:6], termt_1[6:6]);
  C2 I281 (op5_6_0[2:2], termt_4[6:6], termf_1[6:6]);
  C2 I282 (op5_6_0[3:3], termt_4[6:6], termt_1[6:6]);
  OR2 I283 (xf5_0[6:6], op5_6_0[1:1], op5_6_0[2:2]);
  OR2 I284 (xt5_0[6:6], op5_6_0[0:0], op5_6_0[3:3]);
  C2 I285 (op5_7_0[0:0], termf_4[7:7], termf_1[7:7]);
  C2 I286 (op5_7_0[1:1], termf_4[7:7], termt_1[7:7]);
  C2 I287 (op5_7_0[2:2], termt_4[7:7], termf_1[7:7]);
  C2 I288 (op5_7_0[3:3], termt_4[7:7], termt_1[7:7]);
  OR2 I289 (xf5_0[7:7], op5_7_0[1:1], op5_7_0[2:2]);
  OR2 I290 (xt5_0[7:7], op5_7_0[0:0], op5_7_0[3:3]);
  C2 I291 (op5_8_0[0:0], termf_4[8:8], termf_1[8:8]);
  C2 I292 (op5_8_0[1:1], termf_4[8:8], termt_1[8:8]);
  C2 I293 (op5_8_0[2:2], termt_4[8:8], termf_1[8:8]);
  C2 I294 (op5_8_0[3:3], termt_4[8:8], termt_1[8:8]);
  OR2 I295 (xf5_0[8:8], op5_8_0[1:1], op5_8_0[2:2]);
  OR2 I296 (xt5_0[8:8], op5_8_0[0:0], op5_8_0[3:3]);
  C2 I297 (op5_9_0[0:0], termf_4[9:9], termf_1[9:9]);
  C2 I298 (op5_9_0[1:1], termf_4[9:9], termt_1[9:9]);
  C2 I299 (op5_9_0[2:2], termt_4[9:9], termf_1[9:9]);
  C2 I300 (op5_9_0[3:3], termt_4[9:9], termt_1[9:9]);
  OR2 I301 (xf5_0[9:9], op5_9_0[1:1], op5_9_0[2:2]);
  OR2 I302 (xt5_0[9:9], op5_9_0[0:0], op5_9_0[3:3]);
  C2 I303 (op5_10_0[0:0], termf_4[10:10], termf_1[10:10]);
  C2 I304 (op5_10_0[1:1], termf_4[10:10], termt_1[10:10]);
  C2 I305 (op5_10_0[2:2], termt_4[10:10], termf_1[10:10]);
  C2 I306 (op5_10_0[3:3], termt_4[10:10], termt_1[10:10]);
  OR2 I307 (xf5_0[10:10], op5_10_0[1:1], op5_10_0[2:2]);
  OR2 I308 (xt5_0[10:10], op5_10_0[0:0], op5_10_0[3:3]);
  C2 I309 (op5_11_0[0:0], termf_4[11:11], termf_1[11:11]);
  C2 I310 (op5_11_0[1:1], termf_4[11:11], termt_1[11:11]);
  C2 I311 (op5_11_0[2:2], termt_4[11:11], termf_1[11:11]);
  C2 I312 (op5_11_0[3:3], termt_4[11:11], termt_1[11:11]);
  OR2 I313 (xf5_0[11:11], op5_11_0[1:1], op5_11_0[2:2]);
  OR2 I314 (xt5_0[11:11], op5_11_0[0:0], op5_11_0[3:3]);
  C2 I315 (op5_12_0[0:0], termf_4[12:12], termf_1[12:12]);
  C2 I316 (op5_12_0[1:1], termf_4[12:12], termt_1[12:12]);
  C2 I317 (op5_12_0[2:2], termt_4[12:12], termf_1[12:12]);
  C2 I318 (op5_12_0[3:3], termt_4[12:12], termt_1[12:12]);
  OR2 I319 (xf5_0[12:12], op5_12_0[1:1], op5_12_0[2:2]);
  OR2 I320 (xt5_0[12:12], op5_12_0[0:0], op5_12_0[3:3]);
  C2 I321 (op5_13_0[0:0], termf_4[13:13], termf_1[13:13]);
  C2 I322 (op5_13_0[1:1], termf_4[13:13], termt_1[13:13]);
  C2 I323 (op5_13_0[2:2], termt_4[13:13], termf_1[13:13]);
  C2 I324 (op5_13_0[3:3], termt_4[13:13], termt_1[13:13]);
  OR2 I325 (xf5_0[13:13], op5_13_0[1:1], op5_13_0[2:2]);
  OR2 I326 (xt5_0[13:13], op5_13_0[0:0], op5_13_0[3:3]);
  C2 I327 (op5_14_0[0:0], termf_4[14:14], termf_1[14:14]);
  C2 I328 (op5_14_0[1:1], termf_4[14:14], termt_1[14:14]);
  C2 I329 (op5_14_0[2:2], termt_4[14:14], termf_1[14:14]);
  C2 I330 (op5_14_0[3:3], termt_4[14:14], termt_1[14:14]);
  OR2 I331 (xf5_0[14:14], op5_14_0[1:1], op5_14_0[2:2]);
  OR2 I332 (xt5_0[14:14], op5_14_0[0:0], op5_14_0[3:3]);
  C2 I333 (op5_15_0[0:0], termf_4[15:15], termf_1[15:15]);
  C2 I334 (op5_15_0[1:1], termf_4[15:15], termt_1[15:15]);
  C2 I335 (op5_15_0[2:2], termt_4[15:15], termf_1[15:15]);
  C2 I336 (op5_15_0[3:3], termt_4[15:15], termt_1[15:15]);
  OR2 I337 (xf5_0[15:15], op5_15_0[1:1], op5_15_0[2:2]);
  OR2 I338 (xt5_0[15:15], op5_15_0[0:0], op5_15_0[3:3]);
  C2 I339 (op5_16_0[0:0], termf_4[16:16], termf_1[16:16]);
  C2 I340 (op5_16_0[1:1], termf_4[16:16], termt_1[16:16]);
  C2 I341 (op5_16_0[2:2], termt_4[16:16], termf_1[16:16]);
  C2 I342 (op5_16_0[3:3], termt_4[16:16], termt_1[16:16]);
  OR2 I343 (xf5_0[16:16], op5_16_0[1:1], op5_16_0[2:2]);
  OR2 I344 (xt5_0[16:16], op5_16_0[0:0], op5_16_0[3:3]);
  C2 I345 (op5_17_0[0:0], termf_4[17:17], termf_1[17:17]);
  C2 I346 (op5_17_0[1:1], termf_4[17:17], termt_1[17:17]);
  C2 I347 (op5_17_0[2:2], termt_4[17:17], termf_1[17:17]);
  C2 I348 (op5_17_0[3:3], termt_4[17:17], termt_1[17:17]);
  OR2 I349 (xf5_0[17:17], op5_17_0[1:1], op5_17_0[2:2]);
  OR2 I350 (xt5_0[17:17], op5_17_0[0:0], op5_17_0[3:3]);
  C2 I351 (op5_18_0[0:0], termf_4[18:18], termf_1[18:18]);
  C2 I352 (op5_18_0[1:1], termf_4[18:18], termt_1[18:18]);
  C2 I353 (op5_18_0[2:2], termt_4[18:18], termf_1[18:18]);
  C2 I354 (op5_18_0[3:3], termt_4[18:18], termt_1[18:18]);
  OR2 I355 (xf5_0[18:18], op5_18_0[1:1], op5_18_0[2:2]);
  OR2 I356 (xt5_0[18:18], op5_18_0[0:0], op5_18_0[3:3]);
  C2 I357 (op5_19_0[0:0], termf_4[19:19], termf_1[19:19]);
  C2 I358 (op5_19_0[1:1], termf_4[19:19], termt_1[19:19]);
  C2 I359 (op5_19_0[2:2], termt_4[19:19], termf_1[19:19]);
  C2 I360 (op5_19_0[3:3], termt_4[19:19], termt_1[19:19]);
  OR2 I361 (xf5_0[19:19], op5_19_0[1:1], op5_19_0[2:2]);
  OR2 I362 (xt5_0[19:19], op5_19_0[0:0], op5_19_0[3:3]);
  C2 I363 (op5_20_0[0:0], termf_4[20:20], termf_1[20:20]);
  C2 I364 (op5_20_0[1:1], termf_4[20:20], termt_1[20:20]);
  C2 I365 (op5_20_0[2:2], termt_4[20:20], termf_1[20:20]);
  C2 I366 (op5_20_0[3:3], termt_4[20:20], termt_1[20:20]);
  OR2 I367 (xf5_0[20:20], op5_20_0[1:1], op5_20_0[2:2]);
  OR2 I368 (xt5_0[20:20], op5_20_0[0:0], op5_20_0[3:3]);
  C2 I369 (op5_21_0[0:0], termf_4[21:21], termf_1[21:21]);
  C2 I370 (op5_21_0[1:1], termf_4[21:21], termt_1[21:21]);
  C2 I371 (op5_21_0[2:2], termt_4[21:21], termf_1[21:21]);
  C2 I372 (op5_21_0[3:3], termt_4[21:21], termt_1[21:21]);
  OR2 I373 (xf5_0[21:21], op5_21_0[1:1], op5_21_0[2:2]);
  OR2 I374 (xt5_0[21:21], op5_21_0[0:0], op5_21_0[3:3]);
  C2 I375 (op5_22_0[0:0], termf_4[22:22], termf_1[22:22]);
  C2 I376 (op5_22_0[1:1], termf_4[22:22], termt_1[22:22]);
  C2 I377 (op5_22_0[2:2], termt_4[22:22], termf_1[22:22]);
  C2 I378 (op5_22_0[3:3], termt_4[22:22], termt_1[22:22]);
  OR2 I379 (xf5_0[22:22], op5_22_0[1:1], op5_22_0[2:2]);
  OR2 I380 (xt5_0[22:22], op5_22_0[0:0], op5_22_0[3:3]);
  C2 I381 (op5_23_0[0:0], termf_4[23:23], termf_1[23:23]);
  C2 I382 (op5_23_0[1:1], termf_4[23:23], termt_1[23:23]);
  C2 I383 (op5_23_0[2:2], termt_4[23:23], termf_1[23:23]);
  C2 I384 (op5_23_0[3:3], termt_4[23:23], termt_1[23:23]);
  OR2 I385 (xf5_0[23:23], op5_23_0[1:1], op5_23_0[2:2]);
  OR2 I386 (xt5_0[23:23], op5_23_0[0:0], op5_23_0[3:3]);
  C2 I387 (op5_24_0[0:0], termf_4[24:24], termf_1[24:24]);
  C2 I388 (op5_24_0[1:1], termf_4[24:24], termt_1[24:24]);
  C2 I389 (op5_24_0[2:2], termt_4[24:24], termf_1[24:24]);
  C2 I390 (op5_24_0[3:3], termt_4[24:24], termt_1[24:24]);
  OR2 I391 (xf5_0[24:24], op5_24_0[1:1], op5_24_0[2:2]);
  OR2 I392 (xt5_0[24:24], op5_24_0[0:0], op5_24_0[3:3]);
  C2 I393 (op5_25_0[0:0], termf_4[25:25], termf_1[25:25]);
  C2 I394 (op5_25_0[1:1], termf_4[25:25], termt_1[25:25]);
  C2 I395 (op5_25_0[2:2], termt_4[25:25], termf_1[25:25]);
  C2 I396 (op5_25_0[3:3], termt_4[25:25], termt_1[25:25]);
  OR2 I397 (xf5_0[25:25], op5_25_0[1:1], op5_25_0[2:2]);
  OR2 I398 (xt5_0[25:25], op5_25_0[0:0], op5_25_0[3:3]);
  C2 I399 (op5_26_0[0:0], termf_4[26:26], termf_1[26:26]);
  C2 I400 (op5_26_0[1:1], termf_4[26:26], termt_1[26:26]);
  C2 I401 (op5_26_0[2:2], termt_4[26:26], termf_1[26:26]);
  C2 I402 (op5_26_0[3:3], termt_4[26:26], termt_1[26:26]);
  OR2 I403 (xf5_0[26:26], op5_26_0[1:1], op5_26_0[2:2]);
  OR2 I404 (xt5_0[26:26], op5_26_0[0:0], op5_26_0[3:3]);
  C2 I405 (op5_27_0[0:0], termf_4[27:27], termf_1[27:27]);
  C2 I406 (op5_27_0[1:1], termf_4[27:27], termt_1[27:27]);
  C2 I407 (op5_27_0[2:2], termt_4[27:27], termf_1[27:27]);
  C2 I408 (op5_27_0[3:3], termt_4[27:27], termt_1[27:27]);
  OR2 I409 (xf5_0[27:27], op5_27_0[1:1], op5_27_0[2:2]);
  OR2 I410 (xt5_0[27:27], op5_27_0[0:0], op5_27_0[3:3]);
  C2 I411 (op5_28_0[0:0], termf_4[28:28], termf_1[28:28]);
  C2 I412 (op5_28_0[1:1], termf_4[28:28], termt_1[28:28]);
  C2 I413 (op5_28_0[2:2], termt_4[28:28], termf_1[28:28]);
  C2 I414 (op5_28_0[3:3], termt_4[28:28], termt_1[28:28]);
  OR2 I415 (xf5_0[28:28], op5_28_0[1:1], op5_28_0[2:2]);
  OR2 I416 (xt5_0[28:28], op5_28_0[0:0], op5_28_0[3:3]);
  C2 I417 (op5_29_0[0:0], termf_4[29:29], termf_1[29:29]);
  C2 I418 (op5_29_0[1:1], termf_4[29:29], termt_1[29:29]);
  C2 I419 (op5_29_0[2:2], termt_4[29:29], termf_1[29:29]);
  C2 I420 (op5_29_0[3:3], termt_4[29:29], termt_1[29:29]);
  OR2 I421 (xf5_0[29:29], op5_29_0[1:1], op5_29_0[2:2]);
  OR2 I422 (xt5_0[29:29], op5_29_0[0:0], op5_29_0[3:3]);
  C2 I423 (op5_30_0[0:0], termf_4[30:30], termf_1[30:30]);
  C2 I424 (op5_30_0[1:1], termf_4[30:30], termt_1[30:30]);
  C2 I425 (op5_30_0[2:2], termt_4[30:30], termf_1[30:30]);
  C2 I426 (op5_30_0[3:3], termt_4[30:30], termt_1[30:30]);
  OR2 I427 (xf5_0[30:30], op5_30_0[1:1], op5_30_0[2:2]);
  OR2 I428 (xt5_0[30:30], op5_30_0[0:0], op5_30_0[3:3]);
  C2 I429 (op5_31_0[0:0], termf_4[31:31], termf_1[31:31]);
  C2 I430 (op5_31_0[1:1], termf_4[31:31], termt_1[31:31]);
  C2 I431 (op5_31_0[2:2], termt_4[31:31], termf_1[31:31]);
  C2 I432 (op5_31_0[3:3], termt_4[31:31], termt_1[31:31]);
  OR2 I433 (xf5_0[31:31], op5_31_0[1:1], op5_31_0[2:2]);
  OR2 I434 (xt5_0[31:31], op5_31_0[0:0], op5_31_0[3:3]);
  C2 I435 (c5rrrr0_0[0:0], c5rrro_0[1:1], c5rrro_0[0:0]);
  C2 I436 (c5rrrr0_0[1:1], c5rrro_0[1:1], c5rrro_1[0:0]);
  C2 I437 (c5rrrr0_0[2:2], c5rrro_1[1:1], c5rrro_0[0:0]);
  C2 I438 (c5rrrr0_0[3:3], c5rrro_1[1:1], c5rrro_1[0:0]);
  OR3 I439 (o_0r0, c5rrrr0_0[0:0], c5rrrr0_0[1:1], c5rrrr0_0[2:2]);
  BUFF I440 (o_0r1, c5rrrr0_0[3:3]);
  C2 I441 (c5rrr0_0[0:0], c5rro_0[1:1], c5rro_0[0:0]);
  C2 I442 (c5rrr0_0[1:1], c5rro_0[1:1], c5rro_1[0:0]);
  C2 I443 (c5rrr0_0[2:2], c5rro_1[1:1], c5rro_0[0:0]);
  C2 I444 (c5rrr0_0[3:3], c5rro_1[1:1], c5rro_1[0:0]);
  OR3 I445 (c5rrro_0[0:0], c5rrr0_0[0:0], c5rrr0_0[1:1], c5rrr0_0[2:2]);
  BUFF I446 (c5rrro_1[0:0], c5rrr0_0[3:3]);
  C2 I447 (c5rrr1_0[0:0], c5rro_0[3:3], c5rro_0[2:2]);
  C2 I448 (c5rrr1_0[1:1], c5rro_0[3:3], c5rro_1[2:2]);
  C2 I449 (c5rrr1_0[2:2], c5rro_1[3:3], c5rro_0[2:2]);
  C2 I450 (c5rrr1_0[3:3], c5rro_1[3:3], c5rro_1[2:2]);
  OR3 I451 (c5rrro_0[1:1], c5rrr1_0[0:0], c5rrr1_0[1:1], c5rrr1_0[2:2]);
  BUFF I452 (c5rrro_1[1:1], c5rrr1_0[3:3]);
  C2 I453 (c5rr0_0[0:0], c5ro_0[1:1], c5ro_0[0:0]);
  C2 I454 (c5rr0_0[1:1], c5ro_0[1:1], c5ro_1[0:0]);
  C2 I455 (c5rr0_0[2:2], c5ro_1[1:1], c5ro_0[0:0]);
  C2 I456 (c5rr0_0[3:3], c5ro_1[1:1], c5ro_1[0:0]);
  OR3 I457 (c5rro_0[0:0], c5rr0_0[0:0], c5rr0_0[1:1], c5rr0_0[2:2]);
  BUFF I458 (c5rro_1[0:0], c5rr0_0[3:3]);
  C2 I459 (c5rr1_0[0:0], c5ro_0[3:3], c5ro_0[2:2]);
  C2 I460 (c5rr1_0[1:1], c5ro_0[3:3], c5ro_1[2:2]);
  C2 I461 (c5rr1_0[2:2], c5ro_1[3:3], c5ro_0[2:2]);
  C2 I462 (c5rr1_0[3:3], c5ro_1[3:3], c5ro_1[2:2]);
  OR3 I463 (c5rro_0[1:1], c5rr1_0[0:0], c5rr1_0[1:1], c5rr1_0[2:2]);
  BUFF I464 (c5rro_1[1:1], c5rr1_0[3:3]);
  C2 I465 (c5rr2_0[0:0], c5ro_0[5:5], c5ro_0[4:4]);
  C2 I466 (c5rr2_0[1:1], c5ro_0[5:5], c5ro_1[4:4]);
  C2 I467 (c5rr2_0[2:2], c5ro_1[5:5], c5ro_0[4:4]);
  C2 I468 (c5rr2_0[3:3], c5ro_1[5:5], c5ro_1[4:4]);
  OR3 I469 (c5rro_0[2:2], c5rr2_0[0:0], c5rr2_0[1:1], c5rr2_0[2:2]);
  BUFF I470 (c5rro_1[2:2], c5rr2_0[3:3]);
  C2 I471 (c5rr3_0[0:0], c5ro_0[7:7], c5ro_0[6:6]);
  C2 I472 (c5rr3_0[1:1], c5ro_0[7:7], c5ro_1[6:6]);
  C2 I473 (c5rr3_0[2:2], c5ro_1[7:7], c5ro_0[6:6]);
  C2 I474 (c5rr3_0[3:3], c5ro_1[7:7], c5ro_1[6:6]);
  OR3 I475 (c5rro_0[3:3], c5rr3_0[0:0], c5rr3_0[1:1], c5rr3_0[2:2]);
  BUFF I476 (c5rro_1[3:3], c5rr3_0[3:3]);
  C2 I477 (c5r0_0[0:0], c5o_0[1:1], c5o_0[0:0]);
  C2 I478 (c5r0_0[1:1], c5o_0[1:1], c5o_1[0:0]);
  C2 I479 (c5r0_0[2:2], c5o_1[1:1], c5o_0[0:0]);
  C2 I480 (c5r0_0[3:3], c5o_1[1:1], c5o_1[0:0]);
  OR3 I481 (c5ro_0[0:0], c5r0_0[0:0], c5r0_0[1:1], c5r0_0[2:2]);
  BUFF I482 (c5ro_1[0:0], c5r0_0[3:3]);
  C2 I483 (c5r1_0[0:0], c5o_0[3:3], c5o_0[2:2]);
  C2 I484 (c5r1_0[1:1], c5o_0[3:3], c5o_1[2:2]);
  C2 I485 (c5r1_0[2:2], c5o_1[3:3], c5o_0[2:2]);
  C2 I486 (c5r1_0[3:3], c5o_1[3:3], c5o_1[2:2]);
  OR3 I487 (c5ro_0[1:1], c5r1_0[0:0], c5r1_0[1:1], c5r1_0[2:2]);
  BUFF I488 (c5ro_1[1:1], c5r1_0[3:3]);
  C2 I489 (c5r2_0[0:0], c5o_0[5:5], c5o_0[4:4]);
  C2 I490 (c5r2_0[1:1], c5o_0[5:5], c5o_1[4:4]);
  C2 I491 (c5r2_0[2:2], c5o_1[5:5], c5o_0[4:4]);
  C2 I492 (c5r2_0[3:3], c5o_1[5:5], c5o_1[4:4]);
  OR3 I493 (c5ro_0[2:2], c5r2_0[0:0], c5r2_0[1:1], c5r2_0[2:2]);
  BUFF I494 (c5ro_1[2:2], c5r2_0[3:3]);
  C2 I495 (c5r3_0[0:0], c5o_0[7:7], c5o_0[6:6]);
  C2 I496 (c5r3_0[1:1], c5o_0[7:7], c5o_1[6:6]);
  C2 I497 (c5r3_0[2:2], c5o_1[7:7], c5o_0[6:6]);
  C2 I498 (c5r3_0[3:3], c5o_1[7:7], c5o_1[6:6]);
  OR3 I499 (c5ro_0[3:3], c5r3_0[0:0], c5r3_0[1:1], c5r3_0[2:2]);
  BUFF I500 (c5ro_1[3:3], c5r3_0[3:3]);
  C2 I501 (c5r4_0[0:0], c5o_0[9:9], c5o_0[8:8]);
  C2 I502 (c5r4_0[1:1], c5o_0[9:9], c5o_1[8:8]);
  C2 I503 (c5r4_0[2:2], c5o_1[9:9], c5o_0[8:8]);
  C2 I504 (c5r4_0[3:3], c5o_1[9:9], c5o_1[8:8]);
  OR3 I505 (c5ro_0[4:4], c5r4_0[0:0], c5r4_0[1:1], c5r4_0[2:2]);
  BUFF I506 (c5ro_1[4:4], c5r4_0[3:3]);
  C2 I507 (c5r5_0[0:0], c5o_0[11:11], c5o_0[10:10]);
  C2 I508 (c5r5_0[1:1], c5o_0[11:11], c5o_1[10:10]);
  C2 I509 (c5r5_0[2:2], c5o_1[11:11], c5o_0[10:10]);
  C2 I510 (c5r5_0[3:3], c5o_1[11:11], c5o_1[10:10]);
  OR3 I511 (c5ro_0[5:5], c5r5_0[0:0], c5r5_0[1:1], c5r5_0[2:2]);
  BUFF I512 (c5ro_1[5:5], c5r5_0[3:3]);
  C2 I513 (c5r6_0[0:0], c5o_0[13:13], c5o_0[12:12]);
  C2 I514 (c5r6_0[1:1], c5o_0[13:13], c5o_1[12:12]);
  C2 I515 (c5r6_0[2:2], c5o_1[13:13], c5o_0[12:12]);
  C2 I516 (c5r6_0[3:3], c5o_1[13:13], c5o_1[12:12]);
  OR3 I517 (c5ro_0[6:6], c5r6_0[0:0], c5r6_0[1:1], c5r6_0[2:2]);
  BUFF I518 (c5ro_1[6:6], c5r6_0[3:3]);
  C2 I519 (c5r7_0[0:0], c5o_0[15:15], c5o_0[14:14]);
  C2 I520 (c5r7_0[1:1], c5o_0[15:15], c5o_1[14:14]);
  C2 I521 (c5r7_0[2:2], c5o_1[15:15], c5o_0[14:14]);
  C2 I522 (c5r7_0[3:3], c5o_1[15:15], c5o_1[14:14]);
  OR3 I523 (c5ro_0[7:7], c5r7_0[0:0], c5r7_0[1:1], c5r7_0[2:2]);
  BUFF I524 (c5ro_1[7:7], c5r7_0[3:3]);
  C2 I525 (c50_0[0:0], xf5_0[1:1], xf5_0[0:0]);
  C2 I526 (c50_0[1:1], xf5_0[1:1], xt5_0[0:0]);
  C2 I527 (c50_0[2:2], xt5_0[1:1], xf5_0[0:0]);
  C2 I528 (c50_0[3:3], xt5_0[1:1], xt5_0[0:0]);
  OR3 I529 (c5o_0[0:0], c50_0[0:0], c50_0[1:1], c50_0[2:2]);
  BUFF I530 (c5o_1[0:0], c50_0[3:3]);
  C2 I531 (c51_0[0:0], xf5_0[3:3], xf5_0[2:2]);
  C2 I532 (c51_0[1:1], xf5_0[3:3], xt5_0[2:2]);
  C2 I533 (c51_0[2:2], xt5_0[3:3], xf5_0[2:2]);
  C2 I534 (c51_0[3:3], xt5_0[3:3], xt5_0[2:2]);
  OR3 I535 (c5o_0[1:1], c51_0[0:0], c51_0[1:1], c51_0[2:2]);
  BUFF I536 (c5o_1[1:1], c51_0[3:3]);
  C2 I537 (c52_0[0:0], xf5_0[5:5], xf5_0[4:4]);
  C2 I538 (c52_0[1:1], xf5_0[5:5], xt5_0[4:4]);
  C2 I539 (c52_0[2:2], xt5_0[5:5], xf5_0[4:4]);
  C2 I540 (c52_0[3:3], xt5_0[5:5], xt5_0[4:4]);
  OR3 I541 (c5o_0[2:2], c52_0[0:0], c52_0[1:1], c52_0[2:2]);
  BUFF I542 (c5o_1[2:2], c52_0[3:3]);
  C2 I543 (c53_0[0:0], xf5_0[7:7], xf5_0[6:6]);
  C2 I544 (c53_0[1:1], xf5_0[7:7], xt5_0[6:6]);
  C2 I545 (c53_0[2:2], xt5_0[7:7], xf5_0[6:6]);
  C2 I546 (c53_0[3:3], xt5_0[7:7], xt5_0[6:6]);
  OR3 I547 (c5o_0[3:3], c53_0[0:0], c53_0[1:1], c53_0[2:2]);
  BUFF I548 (c5o_1[3:3], c53_0[3:3]);
  C2 I549 (c54_0[0:0], xf5_0[9:9], xf5_0[8:8]);
  C2 I550 (c54_0[1:1], xf5_0[9:9], xt5_0[8:8]);
  C2 I551 (c54_0[2:2], xt5_0[9:9], xf5_0[8:8]);
  C2 I552 (c54_0[3:3], xt5_0[9:9], xt5_0[8:8]);
  OR3 I553 (c5o_0[4:4], c54_0[0:0], c54_0[1:1], c54_0[2:2]);
  BUFF I554 (c5o_1[4:4], c54_0[3:3]);
  C2 I555 (c55_0[0:0], xf5_0[11:11], xf5_0[10:10]);
  C2 I556 (c55_0[1:1], xf5_0[11:11], xt5_0[10:10]);
  C2 I557 (c55_0[2:2], xt5_0[11:11], xf5_0[10:10]);
  C2 I558 (c55_0[3:3], xt5_0[11:11], xt5_0[10:10]);
  OR3 I559 (c5o_0[5:5], c55_0[0:0], c55_0[1:1], c55_0[2:2]);
  BUFF I560 (c5o_1[5:5], c55_0[3:3]);
  C2 I561 (c56_0[0:0], xf5_0[13:13], xf5_0[12:12]);
  C2 I562 (c56_0[1:1], xf5_0[13:13], xt5_0[12:12]);
  C2 I563 (c56_0[2:2], xt5_0[13:13], xf5_0[12:12]);
  C2 I564 (c56_0[3:3], xt5_0[13:13], xt5_0[12:12]);
  OR3 I565 (c5o_0[6:6], c56_0[0:0], c56_0[1:1], c56_0[2:2]);
  BUFF I566 (c5o_1[6:6], c56_0[3:3]);
  C2 I567 (c57_0[0:0], xf5_0[15:15], xf5_0[14:14]);
  C2 I568 (c57_0[1:1], xf5_0[15:15], xt5_0[14:14]);
  C2 I569 (c57_0[2:2], xt5_0[15:15], xf5_0[14:14]);
  C2 I570 (c57_0[3:3], xt5_0[15:15], xt5_0[14:14]);
  OR3 I571 (c5o_0[7:7], c57_0[0:0], c57_0[1:1], c57_0[2:2]);
  BUFF I572 (c5o_1[7:7], c57_0[3:3]);
  C2 I573 (c58_0[0:0], xf5_0[17:17], xf5_0[16:16]);
  C2 I574 (c58_0[1:1], xf5_0[17:17], xt5_0[16:16]);
  C2 I575 (c58_0[2:2], xt5_0[17:17], xf5_0[16:16]);
  C2 I576 (c58_0[3:3], xt5_0[17:17], xt5_0[16:16]);
  OR3 I577 (c5o_0[8:8], c58_0[0:0], c58_0[1:1], c58_0[2:2]);
  BUFF I578 (c5o_1[8:8], c58_0[3:3]);
  C2 I579 (c59_0[0:0], xf5_0[19:19], xf5_0[18:18]);
  C2 I580 (c59_0[1:1], xf5_0[19:19], xt5_0[18:18]);
  C2 I581 (c59_0[2:2], xt5_0[19:19], xf5_0[18:18]);
  C2 I582 (c59_0[3:3], xt5_0[19:19], xt5_0[18:18]);
  OR3 I583 (c5o_0[9:9], c59_0[0:0], c59_0[1:1], c59_0[2:2]);
  BUFF I584 (c5o_1[9:9], c59_0[3:3]);
  C2 I585 (c510_0[0:0], xf5_0[21:21], xf5_0[20:20]);
  C2 I586 (c510_0[1:1], xf5_0[21:21], xt5_0[20:20]);
  C2 I587 (c510_0[2:2], xt5_0[21:21], xf5_0[20:20]);
  C2 I588 (c510_0[3:3], xt5_0[21:21], xt5_0[20:20]);
  OR3 I589 (c5o_0[10:10], c510_0[0:0], c510_0[1:1], c510_0[2:2]);
  BUFF I590 (c5o_1[10:10], c510_0[3:3]);
  C2 I591 (c511_0[0:0], xf5_0[23:23], xf5_0[22:22]);
  C2 I592 (c511_0[1:1], xf5_0[23:23], xt5_0[22:22]);
  C2 I593 (c511_0[2:2], xt5_0[23:23], xf5_0[22:22]);
  C2 I594 (c511_0[3:3], xt5_0[23:23], xt5_0[22:22]);
  OR3 I595 (c5o_0[11:11], c511_0[0:0], c511_0[1:1], c511_0[2:2]);
  BUFF I596 (c5o_1[11:11], c511_0[3:3]);
  C2 I597 (c512_0[0:0], xf5_0[25:25], xf5_0[24:24]);
  C2 I598 (c512_0[1:1], xf5_0[25:25], xt5_0[24:24]);
  C2 I599 (c512_0[2:2], xt5_0[25:25], xf5_0[24:24]);
  C2 I600 (c512_0[3:3], xt5_0[25:25], xt5_0[24:24]);
  OR3 I601 (c5o_0[12:12], c512_0[0:0], c512_0[1:1], c512_0[2:2]);
  BUFF I602 (c5o_1[12:12], c512_0[3:3]);
  C2 I603 (c513_0[0:0], xf5_0[27:27], xf5_0[26:26]);
  C2 I604 (c513_0[1:1], xf5_0[27:27], xt5_0[26:26]);
  C2 I605 (c513_0[2:2], xt5_0[27:27], xf5_0[26:26]);
  C2 I606 (c513_0[3:3], xt5_0[27:27], xt5_0[26:26]);
  OR3 I607 (c5o_0[13:13], c513_0[0:0], c513_0[1:1], c513_0[2:2]);
  BUFF I608 (c5o_1[13:13], c513_0[3:3]);
  C2 I609 (c514_0[0:0], xf5_0[29:29], xf5_0[28:28]);
  C2 I610 (c514_0[1:1], xf5_0[29:29], xt5_0[28:28]);
  C2 I611 (c514_0[2:2], xt5_0[29:29], xf5_0[28:28]);
  C2 I612 (c514_0[3:3], xt5_0[29:29], xt5_0[28:28]);
  OR3 I613 (c5o_0[14:14], c514_0[0:0], c514_0[1:1], c514_0[2:2]);
  BUFF I614 (c5o_1[14:14], c514_0[3:3]);
  C2 I615 (c515_0[0:0], xf5_0[31:31], xf5_0[30:30]);
  C2 I616 (c515_0[1:1], xf5_0[31:31], xt5_0[30:30]);
  C2 I617 (c515_0[2:2], xt5_0[31:31], xf5_0[30:30]);
  C2 I618 (c515_0[3:3], xt5_0[31:31], xt5_0[30:30]);
  OR3 I619 (c5o_0[15:15], c515_0[0:0], c515_0[1:1], c515_0[2:2]);
  BUFF I620 (c5o_1[15:15], c515_0[3:3]);
  BUFF I621 (i_0a, o_0a);
endmodule

// tko2m1_1api0w1b_2api1w1b_3xort1o0w1bt2o0w1b TeakO [
//     (1,TeakOAppend 1 [(0,0+:1)]),
//     (2,TeakOAppend 1 [(0,1+:1)]),
//     (3,TeakOp TeakOpXor [(1,0+:1),(2,0+:1)])] [One 2,One 1]
module tko2m1_1api0w1b_2api1w1b_3xort1o0w1bt2o0w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire termf_1;
  wire termf_2;
  wire termt_1;
  wire termt_2;
  wire [3:0] op3_0_0;
  BUFF I0 (termf_1, i_0r0[0:0]);
  BUFF I1 (termt_1, i_0r1[0:0]);
  BUFF I2 (termf_2, i_0r0[1:1]);
  BUFF I3 (termt_2, i_0r1[1:1]);
  C2 I4 (op3_0_0[0:0], termf_2, termf_1);
  C2 I5 (op3_0_0[1:1], termf_2, termt_1);
  C2 I6 (op3_0_0[2:2], termt_2, termf_1);
  C2 I7 (op3_0_0[3:3], termt_2, termt_1);
  OR2 I8 (o_0r0, op3_0_0[0:0], op3_0_0[3:3]);
  OR2 I9 (o_0r1, op3_0_0[1:1], op3_0_0[2:2]);
  BUFF I10 (i_0a, o_0a);
endmodule

// tko0m6_1nm6b4 TeakO [
//     (1,TeakOConstant 6 4)] [One 0,One 6]
module tko0m6_1nm6b4 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [5:0] o_0r0;
  output [5:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[2:2], i_0r);
  GND I1 (o_0r0[2:2]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  BUFF I6 (o_0r0[5:5], i_0r);
  GND I7 (o_0r1[0:0]);
  GND I8 (o_0r1[1:1]);
  GND I9 (o_0r1[3:3]);
  GND I10 (o_0r1[4:4]);
  GND I11 (o_0r1[5:5]);
  BUFF I12 (i_0a, o_0a);
endmodule

// tkj12m6_6 TeakJ [Many [6,6],One 12]
module tkj12m6_6 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [5:0] i_0r0;
  input [5:0] i_0r1;
  output i_0a;
  input [5:0] i_1r0;
  input [5:0] i_1r1;
  output i_1a;
  output [11:0] o_0r0;
  output [11:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [11:0] joinf_0;
  wire [11:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_1r0[0:0]);
  BUFF I7 (joinf_0[7:7], i_1r0[1:1]);
  BUFF I8 (joinf_0[8:8], i_1r0[2:2]);
  BUFF I9 (joinf_0[9:9], i_1r0[3:3]);
  BUFF I10 (joinf_0[10:10], i_1r0[4:4]);
  BUFF I11 (joinf_0[11:11], i_1r0[5:5]);
  BUFF I12 (joint_0[0:0], i_0r1[0:0]);
  BUFF I13 (joint_0[1:1], i_0r1[1:1]);
  BUFF I14 (joint_0[2:2], i_0r1[2:2]);
  BUFF I15 (joint_0[3:3], i_0r1[3:3]);
  BUFF I16 (joint_0[4:4], i_0r1[4:4]);
  BUFF I17 (joint_0[5:5], i_0r1[5:5]);
  BUFF I18 (joint_0[6:6], i_1r1[0:0]);
  BUFF I19 (joint_0[7:7], i_1r1[1:1]);
  BUFF I20 (joint_0[8:8], i_1r1[2:2]);
  BUFF I21 (joint_0[9:9], i_1r1[3:3]);
  BUFF I22 (joint_0[10:10], i_1r1[4:4]);
  BUFF I23 (joint_0[11:11], i_1r1[5:5]);
  OR2 I24 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I25 (icomplete_0, dcomplete_0);
  C2 I26 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I27 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I28 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I29 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I30 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I31 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I32 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I33 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I34 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I35 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I36 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I37 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I38 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I39 (o_0r1[1:1], joint_0[1:1]);
  BUFF I40 (o_0r1[2:2], joint_0[2:2]);
  BUFF I41 (o_0r1[3:3], joint_0[3:3]);
  BUFF I42 (o_0r1[4:4], joint_0[4:4]);
  BUFF I43 (o_0r1[5:5], joint_0[5:5]);
  BUFF I44 (o_0r1[6:6], joint_0[6:6]);
  BUFF I45 (o_0r1[7:7], joint_0[7:7]);
  BUFF I46 (o_0r1[8:8], joint_0[8:8]);
  BUFF I47 (o_0r1[9:9], joint_0[9:9]);
  BUFF I48 (o_0r1[10:10], joint_0[10:10]);
  BUFF I49 (o_0r1[11:11], joint_0[11:11]);
  BUFF I50 (i_0a, o_0a);
  BUFF I51 (i_1a, o_0a);
endmodule

// tko12m1_1api0w6b_2api6w6b_3eqt1o0w6bt2o0w6b TeakO [
//     (1,TeakOAppend 1 [(0,0+:6)]),
//     (2,TeakOAppend 1 [(0,6+:6)]),
//     (3,TeakOp TeakOpEqual [(1,0+:6),(2,0+:6)])] [One 12,One 1]
module tko12m1_1api0w6b_2api6w6b_3eqt1o0w6bt2o0w6b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [11:0] i_0r0;
  input [11:0] i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire [5:0] termf_1;
  wire [5:0] termf_2;
  wire [5:0] termt_1;
  wire [5:0] termt_2;
  wire [5:0] xf3_0;
  wire [5:0] xt3_0;
  wire [3:0] op3_0_0;
  wire [3:0] op3_1_0;
  wire [3:0] op3_2_0;
  wire [3:0] op3_3_0;
  wire [3:0] op3_4_0;
  wire [3:0] op3_5_0;
  wire [2:0] c3o_0;
  wire [2:0] c3o_1;
  wire [1:0] c3ro_0;
  wire [1:0] c3ro_1;
  wire [3:0] c3rr0_0;
  wire [3:0] c3r0_0;
  wire [3:0] c30_0;
  wire [3:0] c31_0;
  wire [3:0] c32_0;
  BUFF I0 (termf_1[0:0], i_0r0[0:0]);
  BUFF I1 (termf_1[1:1], i_0r0[1:1]);
  BUFF I2 (termf_1[2:2], i_0r0[2:2]);
  BUFF I3 (termf_1[3:3], i_0r0[3:3]);
  BUFF I4 (termf_1[4:4], i_0r0[4:4]);
  BUFF I5 (termf_1[5:5], i_0r0[5:5]);
  BUFF I6 (termt_1[0:0], i_0r1[0:0]);
  BUFF I7 (termt_1[1:1], i_0r1[1:1]);
  BUFF I8 (termt_1[2:2], i_0r1[2:2]);
  BUFF I9 (termt_1[3:3], i_0r1[3:3]);
  BUFF I10 (termt_1[4:4], i_0r1[4:4]);
  BUFF I11 (termt_1[5:5], i_0r1[5:5]);
  BUFF I12 (termf_2[0:0], i_0r0[6:6]);
  BUFF I13 (termf_2[1:1], i_0r0[7:7]);
  BUFF I14 (termf_2[2:2], i_0r0[8:8]);
  BUFF I15 (termf_2[3:3], i_0r0[9:9]);
  BUFF I16 (termf_2[4:4], i_0r0[10:10]);
  BUFF I17 (termf_2[5:5], i_0r0[11:11]);
  BUFF I18 (termt_2[0:0], i_0r1[6:6]);
  BUFF I19 (termt_2[1:1], i_0r1[7:7]);
  BUFF I20 (termt_2[2:2], i_0r1[8:8]);
  BUFF I21 (termt_2[3:3], i_0r1[9:9]);
  BUFF I22 (termt_2[4:4], i_0r1[10:10]);
  BUFF I23 (termt_2[5:5], i_0r1[11:11]);
  C2 I24 (op3_0_0[0:0], termf_2[0:0], termf_1[0:0]);
  C2 I25 (op3_0_0[1:1], termf_2[0:0], termt_1[0:0]);
  C2 I26 (op3_0_0[2:2], termt_2[0:0], termf_1[0:0]);
  C2 I27 (op3_0_0[3:3], termt_2[0:0], termt_1[0:0]);
  OR2 I28 (xf3_0[0:0], op3_0_0[1:1], op3_0_0[2:2]);
  OR2 I29 (xt3_0[0:0], op3_0_0[0:0], op3_0_0[3:3]);
  C2 I30 (op3_1_0[0:0], termf_2[1:1], termf_1[1:1]);
  C2 I31 (op3_1_0[1:1], termf_2[1:1], termt_1[1:1]);
  C2 I32 (op3_1_0[2:2], termt_2[1:1], termf_1[1:1]);
  C2 I33 (op3_1_0[3:3], termt_2[1:1], termt_1[1:1]);
  OR2 I34 (xf3_0[1:1], op3_1_0[1:1], op3_1_0[2:2]);
  OR2 I35 (xt3_0[1:1], op3_1_0[0:0], op3_1_0[3:3]);
  C2 I36 (op3_2_0[0:0], termf_2[2:2], termf_1[2:2]);
  C2 I37 (op3_2_0[1:1], termf_2[2:2], termt_1[2:2]);
  C2 I38 (op3_2_0[2:2], termt_2[2:2], termf_1[2:2]);
  C2 I39 (op3_2_0[3:3], termt_2[2:2], termt_1[2:2]);
  OR2 I40 (xf3_0[2:2], op3_2_0[1:1], op3_2_0[2:2]);
  OR2 I41 (xt3_0[2:2], op3_2_0[0:0], op3_2_0[3:3]);
  C2 I42 (op3_3_0[0:0], termf_2[3:3], termf_1[3:3]);
  C2 I43 (op3_3_0[1:1], termf_2[3:3], termt_1[3:3]);
  C2 I44 (op3_3_0[2:2], termt_2[3:3], termf_1[3:3]);
  C2 I45 (op3_3_0[3:3], termt_2[3:3], termt_1[3:3]);
  OR2 I46 (xf3_0[3:3], op3_3_0[1:1], op3_3_0[2:2]);
  OR2 I47 (xt3_0[3:3], op3_3_0[0:0], op3_3_0[3:3]);
  C2 I48 (op3_4_0[0:0], termf_2[4:4], termf_1[4:4]);
  C2 I49 (op3_4_0[1:1], termf_2[4:4], termt_1[4:4]);
  C2 I50 (op3_4_0[2:2], termt_2[4:4], termf_1[4:4]);
  C2 I51 (op3_4_0[3:3], termt_2[4:4], termt_1[4:4]);
  OR2 I52 (xf3_0[4:4], op3_4_0[1:1], op3_4_0[2:2]);
  OR2 I53 (xt3_0[4:4], op3_4_0[0:0], op3_4_0[3:3]);
  C2 I54 (op3_5_0[0:0], termf_2[5:5], termf_1[5:5]);
  C2 I55 (op3_5_0[1:1], termf_2[5:5], termt_1[5:5]);
  C2 I56 (op3_5_0[2:2], termt_2[5:5], termf_1[5:5]);
  C2 I57 (op3_5_0[3:3], termt_2[5:5], termt_1[5:5]);
  OR2 I58 (xf3_0[5:5], op3_5_0[1:1], op3_5_0[2:2]);
  OR2 I59 (xt3_0[5:5], op3_5_0[0:0], op3_5_0[3:3]);
  C2 I60 (c3rr0_0[0:0], c3ro_0[1:1], c3ro_0[0:0]);
  C2 I61 (c3rr0_0[1:1], c3ro_0[1:1], c3ro_1[0:0]);
  C2 I62 (c3rr0_0[2:2], c3ro_1[1:1], c3ro_0[0:0]);
  C2 I63 (c3rr0_0[3:3], c3ro_1[1:1], c3ro_1[0:0]);
  OR3 I64 (o_0r0, c3rr0_0[0:0], c3rr0_0[1:1], c3rr0_0[2:2]);
  BUFF I65 (o_0r1, c3rr0_0[3:3]);
  BUFF I66 (c3ro_0[1:1], c3o_0[2:2]);
  BUFF I67 (c3ro_1[1:1], c3o_1[2:2]);
  C2 I68 (c3r0_0[0:0], c3o_0[1:1], c3o_0[0:0]);
  C2 I69 (c3r0_0[1:1], c3o_0[1:1], c3o_1[0:0]);
  C2 I70 (c3r0_0[2:2], c3o_1[1:1], c3o_0[0:0]);
  C2 I71 (c3r0_0[3:3], c3o_1[1:1], c3o_1[0:0]);
  OR3 I72 (c3ro_0[0:0], c3r0_0[0:0], c3r0_0[1:1], c3r0_0[2:2]);
  BUFF I73 (c3ro_1[0:0], c3r0_0[3:3]);
  C2 I74 (c30_0[0:0], xf3_0[1:1], xf3_0[0:0]);
  C2 I75 (c30_0[1:1], xf3_0[1:1], xt3_0[0:0]);
  C2 I76 (c30_0[2:2], xt3_0[1:1], xf3_0[0:0]);
  C2 I77 (c30_0[3:3], xt3_0[1:1], xt3_0[0:0]);
  OR3 I78 (c3o_0[0:0], c30_0[0:0], c30_0[1:1], c30_0[2:2]);
  BUFF I79 (c3o_1[0:0], c30_0[3:3]);
  C2 I80 (c31_0[0:0], xf3_0[3:3], xf3_0[2:2]);
  C2 I81 (c31_0[1:1], xf3_0[3:3], xt3_0[2:2]);
  C2 I82 (c31_0[2:2], xt3_0[3:3], xf3_0[2:2]);
  C2 I83 (c31_0[3:3], xt3_0[3:3], xt3_0[2:2]);
  OR3 I84 (c3o_0[1:1], c31_0[0:0], c31_0[1:1], c31_0[2:2]);
  BUFF I85 (c3o_1[1:1], c31_0[3:3]);
  C2 I86 (c32_0[0:0], xf3_0[5:5], xf3_0[4:4]);
  C2 I87 (c32_0[1:1], xf3_0[5:5], xt3_0[4:4]);
  C2 I88 (c32_0[2:2], xt3_0[5:5], xf3_0[4:4]);
  C2 I89 (c32_0[3:3], xt3_0[5:5], xt3_0[4:4]);
  OR3 I90 (c3o_0[2:2], c32_0[0:0], c32_0[1:1], c32_0[2:2]);
  BUFF I91 (c3o_1[2:2], c32_0[3:3]);
  BUFF I92 (i_0a, o_0a);
endmodule

// tko2m1_1api0w1b_2api1w1b_3net1o0w1bt2o0w1b TeakO [
//     (1,TeakOAppend 1 [(0,0+:1)]),
//     (2,TeakOAppend 1 [(0,1+:1)]),
//     (3,TeakOp TeakOpNotEqual [(1,0+:1),(2,0+:1)])] [One 2,One 1]
module tko2m1_1api0w1b_2api1w1b_3net1o0w1bt2o0w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire termf_1;
  wire termf_2;
  wire termt_1;
  wire termt_2;
  wire xf3_0;
  wire xt3_0;
  wire [3:0] op3_0_0;
  BUFF I0 (termf_1, i_0r0[0:0]);
  BUFF I1 (termt_1, i_0r1[0:0]);
  BUFF I2 (termf_2, i_0r0[1:1]);
  BUFF I3 (termt_2, i_0r1[1:1]);
  C2 I4 (op3_0_0[0:0], termf_2, termf_1);
  C2 I5 (op3_0_0[1:1], termf_2, termt_1);
  C2 I6 (op3_0_0[2:2], termt_2, termf_1);
  C2 I7 (op3_0_0[3:3], termt_2, termt_1);
  OR2 I8 (xf3_0, op3_0_0[1:1], op3_0_0[2:2]);
  OR2 I9 (xt3_0, op3_0_0[0:0], op3_0_0[3:3]);
  BUFF I10 (o_0r1, xf3_0);
  BUFF I11 (o_0r0, xt3_0);
  BUFF I12 (i_0a, o_0a);
endmodule

// tkj4m1_1_1_1 TeakJ [Many [1,1,1,1],One 4]
module tkj4m1_1_1_1 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input i_1r0;
  input i_1r1;
  output i_1a;
  input i_2r0;
  input i_2r1;
  output i_2a;
  input i_3r0;
  input i_3r1;
  output i_3a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [3:0] joinf_0;
  wire [3:0] joint_0;
  wire dcomplete_0;
  wire dcomplete_1;
  wire dcomplete_2;
  BUFF I0 (joinf_0[0:0], i_0r0);
  BUFF I1 (joinf_0[1:1], i_1r0);
  BUFF I2 (joinf_0[2:2], i_2r0);
  BUFF I3 (joinf_0[3:3], i_3r0);
  BUFF I4 (joint_0[0:0], i_0r1);
  BUFF I5 (joint_0[1:1], i_1r1);
  BUFF I6 (joint_0[2:2], i_2r1);
  BUFF I7 (joint_0[3:3], i_3r1);
  OR2 I8 (dcomplete_0, i_1r0, i_1r1);
  OR2 I9 (dcomplete_1, i_2r0, i_2r1);
  OR2 I10 (dcomplete_2, i_3r0, i_3r1);
  C3 I11 (icomplete_0, dcomplete_0, dcomplete_1, dcomplete_2);
  C2 I12 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I13 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I14 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I15 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I16 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I17 (o_0r1[1:1], joint_0[1:1]);
  BUFF I18 (o_0r1[2:2], joint_0[2:2]);
  BUFF I19 (o_0r1[3:3], joint_0[3:3]);
  BUFF I20 (i_0a, o_0a);
  BUFF I21 (i_1a, o_0a);
  BUFF I22 (i_2a, o_0a);
  BUFF I23 (i_3a, o_0a);
endmodule

// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 TeakF [0,0,0,0,0,0,0,0,0,0] [One 0,Many [0,0,
//   0,0,0,0,0,0,0,0]]
module tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, o_5r, o_5a, o_6r, o_6a, o_7r, o_7a, o_8r, o_8a, o_9r, o_9a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  output o_7r;
  input o_7a;
  output o_8r;
  input o_8a;
  output o_9r;
  input o_9a;
  input reset;
  wire [3:0] simp11_0;
  wire [1:0] simp12_0;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  BUFF I2 (o_2r, i_0r);
  BUFF I3 (o_3r, i_0r);
  BUFF I4 (o_4r, i_0r);
  BUFF I5 (o_5r, i_0r);
  BUFF I6 (o_6r, i_0r);
  BUFF I7 (o_7r, i_0r);
  BUFF I8 (o_8r, i_0r);
  BUFF I9 (o_9r, i_0r);
  C3 I10 (simp11_0[0:0], o_0a, o_1a, o_2a);
  C3 I11 (simp11_0[1:1], o_3a, o_4a, o_5a);
  C3 I12 (simp11_0[2:2], o_6a, o_7a, o_8a);
  BUFF I13 (simp11_0[3:3], o_9a);
  C3 I14 (simp12_0[0:0], simp11_0[0:0], simp11_0[1:1], simp11_0[2:2]);
  BUFF I15 (simp12_0[1:1], simp11_0[3:3]);
  C2 I16 (i_0a, simp12_0[0:0], simp12_0[1:1]);
endmodule

// tkvmergedResult33_wo0w33_ro0w32o0w32o31w1o32w1o31w1o32w1 TeakV "mergedResult" 33 [] [0] [0,0,31,32,3
//   1,32] [Many [33],Many [0],Many [0,0,0,0,0,0],Many [32,32,1,1,1,1]]
module tkvmergedResult33_wo0w33_ro0w32o0w32o31w1o32w1o31w1o32w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rg_5r, rg_5a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, rd_5r0, rd_5r1, rd_5a, reset);
  input [32:0] wg_0r0;
  input [32:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  input rg_5r;
  output rg_5a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output rd_2r0;
  output rd_2r1;
  input rd_2a;
  output rd_3r0;
  output rd_3r1;
  input rd_3a;
  output rd_4r0;
  output rd_4r1;
  input rd_4a;
  output rd_5r0;
  output rd_5r1;
  input rd_5a;
  input reset;
  wire [32:0] wf_0;
  wire [32:0] wt_0;
  wire [32:0] df_0;
  wire [32:0] dt_0;
  wire wc_0;
  wire [32:0] wacks_0;
  wire [32:0] wenr_0;
  wire [32:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [32:0] drlgf_0;
  wire [32:0] drlgt_0;
  wire [32:0] comp0_0;
  wire [10:0] simp2451_0;
  wire [3:0] simp2452_0;
  wire [1:0] simp2453_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [32:0] conwgit_0;
  wire [32:0] conwgif_0;
  wire conwig_0;
  wire [11:0] simp4191_0;
  wire [3:0] simp4192_0;
  wire [1:0] simp4193_0;
  wire [3:0] simp5561_0;
  wire [1:0] simp5562_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (wen_0[32:32], wenr_0[32:32], nreset_0);
  AND2 I34 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I35 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I36 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I37 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I38 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I39 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I40 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I41 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I42 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I43 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I44 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I45 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I46 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I47 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I48 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I49 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I50 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I51 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I52 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I53 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I54 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I55 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I56 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I57 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I58 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I59 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I60 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I61 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I62 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I63 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I64 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I65 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I66 (drlgf_0[32:32], wf_0[32:32], wen_0[32:32]);
  AND2 I67 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I68 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I69 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I70 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I71 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I72 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I73 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I74 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I75 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I76 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I77 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I78 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I79 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I80 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I81 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I82 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I83 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I84 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I85 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I86 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I87 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I88 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I89 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I90 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I91 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I92 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I93 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I94 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I95 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I96 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I97 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I98 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  AND2 I99 (drlgt_0[32:32], wt_0[32:32], wen_0[32:32]);
  NOR2 I100 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I101 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I102 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I103 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I104 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I105 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I106 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I107 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I108 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I109 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I110 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I111 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I112 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I113 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I114 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I115 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I116 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I117 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I118 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I119 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I120 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I121 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I122 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I123 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I124 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I125 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I126 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I127 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I128 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I129 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I130 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I131 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR2 I132 (df_0[32:32], dt_0[32:32], drlgt_0[32:32]);
  NOR3 I133 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I134 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I135 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I136 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I137 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I138 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I139 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I140 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I141 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I142 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I143 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I144 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I145 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I146 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I147 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I148 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I149 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I150 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I151 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I152 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I153 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I154 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I155 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I156 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I157 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I158 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I159 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I160 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I161 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I162 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I163 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I164 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  NOR3 I165 (dt_0[32:32], df_0[32:32], drlgf_0[32:32], reset);
  AO22 I166 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I167 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I168 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I169 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I170 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I171 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I172 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I173 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I174 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I175 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I176 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I177 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I178 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I179 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I180 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I181 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I182 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I183 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I184 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I185 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I186 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I187 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I188 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I189 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I190 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I191 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I192 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I193 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I194 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I195 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I196 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I197 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  AO22 I198 (wacks_0[32:32], drlgf_0[32:32], df_0[32:32], drlgt_0[32:32], dt_0[32:32]);
  OR2 I199 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I200 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I201 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I202 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I203 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I204 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I205 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I206 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I207 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I208 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I209 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I210 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I211 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I212 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I213 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I214 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I215 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I216 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I217 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I218 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I219 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I220 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I221 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I222 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I223 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I224 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I225 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I226 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I227 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I228 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I229 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I230 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  OR2 I231 (comp0_0[32:32], wg_0r0[32:32], wg_0r1[32:32]);
  C3 I232 (simp2451_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I233 (simp2451_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I234 (simp2451_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I235 (simp2451_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I236 (simp2451_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I237 (simp2451_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I238 (simp2451_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I239 (simp2451_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I240 (simp2451_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I241 (simp2451_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C3 I242 (simp2451_0[10:10], comp0_0[30:30], comp0_0[31:31], comp0_0[32:32]);
  C3 I243 (simp2452_0[0:0], simp2451_0[0:0], simp2451_0[1:1], simp2451_0[2:2]);
  C3 I244 (simp2452_0[1:1], simp2451_0[3:3], simp2451_0[4:4], simp2451_0[5:5]);
  C3 I245 (simp2452_0[2:2], simp2451_0[6:6], simp2451_0[7:7], simp2451_0[8:8]);
  C2 I246 (simp2452_0[3:3], simp2451_0[9:9], simp2451_0[10:10]);
  C3 I247 (simp2453_0[0:0], simp2452_0[0:0], simp2452_0[1:1], simp2452_0[2:2]);
  BUFF I248 (simp2453_0[1:1], simp2452_0[3:3]);
  C2 I249 (wc_0, simp2453_0[0:0], simp2453_0[1:1]);
  AND2 I250 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I251 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I252 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I253 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I254 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I255 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I256 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I257 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I258 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I259 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I260 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I261 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I262 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I263 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I264 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I265 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I266 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I267 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I268 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I269 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I270 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I271 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I272 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I273 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I274 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I275 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I276 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I277 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I278 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I279 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I280 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I281 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I282 (conwgif_0[32:32], wg_0r0[32:32], conwig_0);
  AND2 I283 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I284 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I285 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I286 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I287 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I288 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I289 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I290 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I291 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I292 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I293 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I294 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I295 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I296 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I297 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I298 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I299 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I300 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I301 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I302 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I303 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I304 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I305 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I306 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I307 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I308 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I309 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I310 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I311 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I312 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I313 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I314 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  AND2 I315 (conwgit_0[32:32], wg_0r1[32:32], conwig_0);
  BUFF I316 (conwigc_0, wc_0);
  AO22 I317 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I318 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I319 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I320 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I321 (wenr_0[0:0], wc_0);
  BUFF I322 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I323 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I324 (wenr_0[1:1], wc_0);
  BUFF I325 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I326 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I327 (wenr_0[2:2], wc_0);
  BUFF I328 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I329 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I330 (wenr_0[3:3], wc_0);
  BUFF I331 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I332 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I333 (wenr_0[4:4], wc_0);
  BUFF I334 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I335 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I336 (wenr_0[5:5], wc_0);
  BUFF I337 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I338 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I339 (wenr_0[6:6], wc_0);
  BUFF I340 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I341 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I342 (wenr_0[7:7], wc_0);
  BUFF I343 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I344 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I345 (wenr_0[8:8], wc_0);
  BUFF I346 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I347 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I348 (wenr_0[9:9], wc_0);
  BUFF I349 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I350 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I351 (wenr_0[10:10], wc_0);
  BUFF I352 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I353 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I354 (wenr_0[11:11], wc_0);
  BUFF I355 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I356 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I357 (wenr_0[12:12], wc_0);
  BUFF I358 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I359 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I360 (wenr_0[13:13], wc_0);
  BUFF I361 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I362 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I363 (wenr_0[14:14], wc_0);
  BUFF I364 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I365 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I366 (wenr_0[15:15], wc_0);
  BUFF I367 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I368 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I369 (wenr_0[16:16], wc_0);
  BUFF I370 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I371 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I372 (wenr_0[17:17], wc_0);
  BUFF I373 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I374 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I375 (wenr_0[18:18], wc_0);
  BUFF I376 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I377 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I378 (wenr_0[19:19], wc_0);
  BUFF I379 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I380 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I381 (wenr_0[20:20], wc_0);
  BUFF I382 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I383 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I384 (wenr_0[21:21], wc_0);
  BUFF I385 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I386 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I387 (wenr_0[22:22], wc_0);
  BUFF I388 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I389 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I390 (wenr_0[23:23], wc_0);
  BUFF I391 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I392 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I393 (wenr_0[24:24], wc_0);
  BUFF I394 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I395 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I396 (wenr_0[25:25], wc_0);
  BUFF I397 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I398 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I399 (wenr_0[26:26], wc_0);
  BUFF I400 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I401 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I402 (wenr_0[27:27], wc_0);
  BUFF I403 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I404 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I405 (wenr_0[28:28], wc_0);
  BUFF I406 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I407 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I408 (wenr_0[29:29], wc_0);
  BUFF I409 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I410 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I411 (wenr_0[30:30], wc_0);
  BUFF I412 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I413 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I414 (wenr_0[31:31], wc_0);
  BUFF I415 (wf_0[32:32], conwgif_0[32:32]);
  BUFF I416 (wt_0[32:32], conwgit_0[32:32]);
  BUFF I417 (wenr_0[32:32], wc_0);
  C3 I418 (simp4191_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I419 (simp4191_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I420 (simp4191_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I421 (simp4191_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I422 (simp4191_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I423 (simp4191_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I424 (simp4191_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I425 (simp4191_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I426 (simp4191_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I427 (simp4191_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I428 (simp4191_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  BUFF I429 (simp4191_0[11:11], wacks_0[32:32]);
  C3 I430 (simp4192_0[0:0], simp4191_0[0:0], simp4191_0[1:1], simp4191_0[2:2]);
  C3 I431 (simp4192_0[1:1], simp4191_0[3:3], simp4191_0[4:4], simp4191_0[5:5]);
  C3 I432 (simp4192_0[2:2], simp4191_0[6:6], simp4191_0[7:7], simp4191_0[8:8]);
  C3 I433 (simp4192_0[3:3], simp4191_0[9:9], simp4191_0[10:10], simp4191_0[11:11]);
  C3 I434 (simp4193_0[0:0], simp4192_0[0:0], simp4192_0[1:1], simp4192_0[2:2]);
  BUFF I435 (simp4193_0[1:1], simp4192_0[3:3]);
  C2 I436 (wd_0r, simp4193_0[0:0], simp4193_0[1:1]);
  AND2 I437 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I438 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I439 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I440 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I441 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I442 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I443 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I444 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I445 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I446 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I447 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I448 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I449 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I450 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I451 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I452 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I453 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I454 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I455 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I456 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I457 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I458 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I459 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I460 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I461 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I462 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I463 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I464 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I465 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I466 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I467 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I468 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I469 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I470 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I471 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I472 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I473 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I474 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I475 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I476 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I477 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I478 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I479 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I480 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I481 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I482 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I483 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I484 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I485 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I486 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I487 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I488 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I489 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I490 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I491 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I492 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I493 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I494 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I495 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I496 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I497 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I498 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I499 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I500 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I501 (rd_2r0, df_0[31:31], rg_2r);
  AND2 I502 (rd_3r0, df_0[32:32], rg_3r);
  AND2 I503 (rd_4r0, df_0[31:31], rg_4r);
  AND2 I504 (rd_5r0, df_0[32:32], rg_5r);
  AND2 I505 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I506 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I507 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I508 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I509 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I510 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I511 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I512 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I513 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I514 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I515 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I516 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I517 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I518 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I519 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I520 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I521 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I522 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I523 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I524 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I525 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I526 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I527 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I528 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I529 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I530 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I531 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I532 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I533 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I534 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I535 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I536 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I537 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I538 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I539 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I540 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I541 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I542 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I543 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I544 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I545 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I546 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I547 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I548 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I549 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I550 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I551 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I552 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I553 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I554 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I555 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I556 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I557 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I558 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I559 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I560 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I561 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I562 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I563 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I564 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I565 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I566 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I567 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I568 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I569 (rd_2r1, dt_0[31:31], rg_2r);
  AND2 I570 (rd_3r1, dt_0[32:32], rg_3r);
  AND2 I571 (rd_4r1, dt_0[31:31], rg_4r);
  AND2 I572 (rd_5r1, dt_0[32:32], rg_5r);
  NOR3 I573 (simp5561_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I574 (simp5561_0[1:1], rg_3r, rg_4r, rg_5r);
  NOR3 I575 (simp5561_0[2:2], rg_0a, rg_1a, rg_2a);
  NOR3 I576 (simp5561_0[3:3], rg_3a, rg_4a, rg_5a);
  NAND3 I577 (simp5562_0[0:0], simp5561_0[0:0], simp5561_0[1:1], simp5561_0[2:2]);
  INV I578 (simp5562_0[1:1], simp5561_0[3:3]);
  OR2 I579 (anyread_0, simp5562_0[0:0], simp5562_0[1:1]);
  BUFF I580 (wg_0a, wd_0a);
  BUFF I581 (rg_0a, rd_0a);
  BUFF I582 (rg_1a, rd_1a);
  BUFF I583 (rg_2a, rd_2a);
  BUFF I584 (rg_3a, rd_3a);
  BUFF I585 (rg_4a, rd_4a);
  BUFF I586 (rg_5a, rd_5a);
endmodule

// tkm3x33b TeakM [Many [33,33,33],One 33]
module tkm3x33b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, o_0r0, o_0r1, o_0a, reset);
  input [32:0] i_0r0;
  input [32:0] i_0r1;
  output i_0a;
  input [32:0] i_1r0;
  input [32:0] i_1r1;
  output i_1a;
  input [32:0] i_2r0;
  input [32:0] i_2r1;
  output i_2a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  wire [32:0] gfint_0;
  wire [32:0] gfint_1;
  wire [32:0] gfint_2;
  wire [32:0] gtint_0;
  wire [32:0] gtint_1;
  wire [32:0] gtint_2;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire nchosen_0;
  wire [32:0] comp0_0;
  wire [10:0] simp3121_0;
  wire [3:0] simp3122_0;
  wire [1:0] simp3123_0;
  wire [32:0] comp1_0;
  wire [10:0] simp3471_0;
  wire [3:0] simp3472_0;
  wire [1:0] simp3473_0;
  wire [32:0] comp2_0;
  wire [10:0] simp3821_0;
  wire [3:0] simp3822_0;
  wire [1:0] simp3823_0;
  OR3 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  OR3 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  OR3 I2 (o_0r0[2:2], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  OR3 I3 (o_0r0[3:3], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  OR3 I4 (o_0r0[4:4], gfint_0[4:4], gfint_1[4:4], gfint_2[4:4]);
  OR3 I5 (o_0r0[5:5], gfint_0[5:5], gfint_1[5:5], gfint_2[5:5]);
  OR3 I6 (o_0r0[6:6], gfint_0[6:6], gfint_1[6:6], gfint_2[6:6]);
  OR3 I7 (o_0r0[7:7], gfint_0[7:7], gfint_1[7:7], gfint_2[7:7]);
  OR3 I8 (o_0r0[8:8], gfint_0[8:8], gfint_1[8:8], gfint_2[8:8]);
  OR3 I9 (o_0r0[9:9], gfint_0[9:9], gfint_1[9:9], gfint_2[9:9]);
  OR3 I10 (o_0r0[10:10], gfint_0[10:10], gfint_1[10:10], gfint_2[10:10]);
  OR3 I11 (o_0r0[11:11], gfint_0[11:11], gfint_1[11:11], gfint_2[11:11]);
  OR3 I12 (o_0r0[12:12], gfint_0[12:12], gfint_1[12:12], gfint_2[12:12]);
  OR3 I13 (o_0r0[13:13], gfint_0[13:13], gfint_1[13:13], gfint_2[13:13]);
  OR3 I14 (o_0r0[14:14], gfint_0[14:14], gfint_1[14:14], gfint_2[14:14]);
  OR3 I15 (o_0r0[15:15], gfint_0[15:15], gfint_1[15:15], gfint_2[15:15]);
  OR3 I16 (o_0r0[16:16], gfint_0[16:16], gfint_1[16:16], gfint_2[16:16]);
  OR3 I17 (o_0r0[17:17], gfint_0[17:17], gfint_1[17:17], gfint_2[17:17]);
  OR3 I18 (o_0r0[18:18], gfint_0[18:18], gfint_1[18:18], gfint_2[18:18]);
  OR3 I19 (o_0r0[19:19], gfint_0[19:19], gfint_1[19:19], gfint_2[19:19]);
  OR3 I20 (o_0r0[20:20], gfint_0[20:20], gfint_1[20:20], gfint_2[20:20]);
  OR3 I21 (o_0r0[21:21], gfint_0[21:21], gfint_1[21:21], gfint_2[21:21]);
  OR3 I22 (o_0r0[22:22], gfint_0[22:22], gfint_1[22:22], gfint_2[22:22]);
  OR3 I23 (o_0r0[23:23], gfint_0[23:23], gfint_1[23:23], gfint_2[23:23]);
  OR3 I24 (o_0r0[24:24], gfint_0[24:24], gfint_1[24:24], gfint_2[24:24]);
  OR3 I25 (o_0r0[25:25], gfint_0[25:25], gfint_1[25:25], gfint_2[25:25]);
  OR3 I26 (o_0r0[26:26], gfint_0[26:26], gfint_1[26:26], gfint_2[26:26]);
  OR3 I27 (o_0r0[27:27], gfint_0[27:27], gfint_1[27:27], gfint_2[27:27]);
  OR3 I28 (o_0r0[28:28], gfint_0[28:28], gfint_1[28:28], gfint_2[28:28]);
  OR3 I29 (o_0r0[29:29], gfint_0[29:29], gfint_1[29:29], gfint_2[29:29]);
  OR3 I30 (o_0r0[30:30], gfint_0[30:30], gfint_1[30:30], gfint_2[30:30]);
  OR3 I31 (o_0r0[31:31], gfint_0[31:31], gfint_1[31:31], gfint_2[31:31]);
  OR3 I32 (o_0r0[32:32], gfint_0[32:32], gfint_1[32:32], gfint_2[32:32]);
  OR3 I33 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  OR3 I34 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  OR3 I35 (o_0r1[2:2], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  OR3 I36 (o_0r1[3:3], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  OR3 I37 (o_0r1[4:4], gtint_0[4:4], gtint_1[4:4], gtint_2[4:4]);
  OR3 I38 (o_0r1[5:5], gtint_0[5:5], gtint_1[5:5], gtint_2[5:5]);
  OR3 I39 (o_0r1[6:6], gtint_0[6:6], gtint_1[6:6], gtint_2[6:6]);
  OR3 I40 (o_0r1[7:7], gtint_0[7:7], gtint_1[7:7], gtint_2[7:7]);
  OR3 I41 (o_0r1[8:8], gtint_0[8:8], gtint_1[8:8], gtint_2[8:8]);
  OR3 I42 (o_0r1[9:9], gtint_0[9:9], gtint_1[9:9], gtint_2[9:9]);
  OR3 I43 (o_0r1[10:10], gtint_0[10:10], gtint_1[10:10], gtint_2[10:10]);
  OR3 I44 (o_0r1[11:11], gtint_0[11:11], gtint_1[11:11], gtint_2[11:11]);
  OR3 I45 (o_0r1[12:12], gtint_0[12:12], gtint_1[12:12], gtint_2[12:12]);
  OR3 I46 (o_0r1[13:13], gtint_0[13:13], gtint_1[13:13], gtint_2[13:13]);
  OR3 I47 (o_0r1[14:14], gtint_0[14:14], gtint_1[14:14], gtint_2[14:14]);
  OR3 I48 (o_0r1[15:15], gtint_0[15:15], gtint_1[15:15], gtint_2[15:15]);
  OR3 I49 (o_0r1[16:16], gtint_0[16:16], gtint_1[16:16], gtint_2[16:16]);
  OR3 I50 (o_0r1[17:17], gtint_0[17:17], gtint_1[17:17], gtint_2[17:17]);
  OR3 I51 (o_0r1[18:18], gtint_0[18:18], gtint_1[18:18], gtint_2[18:18]);
  OR3 I52 (o_0r1[19:19], gtint_0[19:19], gtint_1[19:19], gtint_2[19:19]);
  OR3 I53 (o_0r1[20:20], gtint_0[20:20], gtint_1[20:20], gtint_2[20:20]);
  OR3 I54 (o_0r1[21:21], gtint_0[21:21], gtint_1[21:21], gtint_2[21:21]);
  OR3 I55 (o_0r1[22:22], gtint_0[22:22], gtint_1[22:22], gtint_2[22:22]);
  OR3 I56 (o_0r1[23:23], gtint_0[23:23], gtint_1[23:23], gtint_2[23:23]);
  OR3 I57 (o_0r1[24:24], gtint_0[24:24], gtint_1[24:24], gtint_2[24:24]);
  OR3 I58 (o_0r1[25:25], gtint_0[25:25], gtint_1[25:25], gtint_2[25:25]);
  OR3 I59 (o_0r1[26:26], gtint_0[26:26], gtint_1[26:26], gtint_2[26:26]);
  OR3 I60 (o_0r1[27:27], gtint_0[27:27], gtint_1[27:27], gtint_2[27:27]);
  OR3 I61 (o_0r1[28:28], gtint_0[28:28], gtint_1[28:28], gtint_2[28:28]);
  OR3 I62 (o_0r1[29:29], gtint_0[29:29], gtint_1[29:29], gtint_2[29:29]);
  OR3 I63 (o_0r1[30:30], gtint_0[30:30], gtint_1[30:30], gtint_2[30:30]);
  OR3 I64 (o_0r1[31:31], gtint_0[31:31], gtint_1[31:31], gtint_2[31:31]);
  OR3 I65 (o_0r1[32:32], gtint_0[32:32], gtint_1[32:32], gtint_2[32:32]);
  AND2 I66 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I67 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I68 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I69 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I70 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I71 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I72 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I73 (gtint_0[7:7], choice_0, i_0r1[7:7]);
  AND2 I74 (gtint_0[8:8], choice_0, i_0r1[8:8]);
  AND2 I75 (gtint_0[9:9], choice_0, i_0r1[9:9]);
  AND2 I76 (gtint_0[10:10], choice_0, i_0r1[10:10]);
  AND2 I77 (gtint_0[11:11], choice_0, i_0r1[11:11]);
  AND2 I78 (gtint_0[12:12], choice_0, i_0r1[12:12]);
  AND2 I79 (gtint_0[13:13], choice_0, i_0r1[13:13]);
  AND2 I80 (gtint_0[14:14], choice_0, i_0r1[14:14]);
  AND2 I81 (gtint_0[15:15], choice_0, i_0r1[15:15]);
  AND2 I82 (gtint_0[16:16], choice_0, i_0r1[16:16]);
  AND2 I83 (gtint_0[17:17], choice_0, i_0r1[17:17]);
  AND2 I84 (gtint_0[18:18], choice_0, i_0r1[18:18]);
  AND2 I85 (gtint_0[19:19], choice_0, i_0r1[19:19]);
  AND2 I86 (gtint_0[20:20], choice_0, i_0r1[20:20]);
  AND2 I87 (gtint_0[21:21], choice_0, i_0r1[21:21]);
  AND2 I88 (gtint_0[22:22], choice_0, i_0r1[22:22]);
  AND2 I89 (gtint_0[23:23], choice_0, i_0r1[23:23]);
  AND2 I90 (gtint_0[24:24], choice_0, i_0r1[24:24]);
  AND2 I91 (gtint_0[25:25], choice_0, i_0r1[25:25]);
  AND2 I92 (gtint_0[26:26], choice_0, i_0r1[26:26]);
  AND2 I93 (gtint_0[27:27], choice_0, i_0r1[27:27]);
  AND2 I94 (gtint_0[28:28], choice_0, i_0r1[28:28]);
  AND2 I95 (gtint_0[29:29], choice_0, i_0r1[29:29]);
  AND2 I96 (gtint_0[30:30], choice_0, i_0r1[30:30]);
  AND2 I97 (gtint_0[31:31], choice_0, i_0r1[31:31]);
  AND2 I98 (gtint_0[32:32], choice_0, i_0r1[32:32]);
  AND2 I99 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I100 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I101 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I102 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I103 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I104 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I105 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I106 (gtint_1[7:7], choice_1, i_1r1[7:7]);
  AND2 I107 (gtint_1[8:8], choice_1, i_1r1[8:8]);
  AND2 I108 (gtint_1[9:9], choice_1, i_1r1[9:9]);
  AND2 I109 (gtint_1[10:10], choice_1, i_1r1[10:10]);
  AND2 I110 (gtint_1[11:11], choice_1, i_1r1[11:11]);
  AND2 I111 (gtint_1[12:12], choice_1, i_1r1[12:12]);
  AND2 I112 (gtint_1[13:13], choice_1, i_1r1[13:13]);
  AND2 I113 (gtint_1[14:14], choice_1, i_1r1[14:14]);
  AND2 I114 (gtint_1[15:15], choice_1, i_1r1[15:15]);
  AND2 I115 (gtint_1[16:16], choice_1, i_1r1[16:16]);
  AND2 I116 (gtint_1[17:17], choice_1, i_1r1[17:17]);
  AND2 I117 (gtint_1[18:18], choice_1, i_1r1[18:18]);
  AND2 I118 (gtint_1[19:19], choice_1, i_1r1[19:19]);
  AND2 I119 (gtint_1[20:20], choice_1, i_1r1[20:20]);
  AND2 I120 (gtint_1[21:21], choice_1, i_1r1[21:21]);
  AND2 I121 (gtint_1[22:22], choice_1, i_1r1[22:22]);
  AND2 I122 (gtint_1[23:23], choice_1, i_1r1[23:23]);
  AND2 I123 (gtint_1[24:24], choice_1, i_1r1[24:24]);
  AND2 I124 (gtint_1[25:25], choice_1, i_1r1[25:25]);
  AND2 I125 (gtint_1[26:26], choice_1, i_1r1[26:26]);
  AND2 I126 (gtint_1[27:27], choice_1, i_1r1[27:27]);
  AND2 I127 (gtint_1[28:28], choice_1, i_1r1[28:28]);
  AND2 I128 (gtint_1[29:29], choice_1, i_1r1[29:29]);
  AND2 I129 (gtint_1[30:30], choice_1, i_1r1[30:30]);
  AND2 I130 (gtint_1[31:31], choice_1, i_1r1[31:31]);
  AND2 I131 (gtint_1[32:32], choice_1, i_1r1[32:32]);
  AND2 I132 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I133 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I134 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I135 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AND2 I136 (gtint_2[4:4], choice_2, i_2r1[4:4]);
  AND2 I137 (gtint_2[5:5], choice_2, i_2r1[5:5]);
  AND2 I138 (gtint_2[6:6], choice_2, i_2r1[6:6]);
  AND2 I139 (gtint_2[7:7], choice_2, i_2r1[7:7]);
  AND2 I140 (gtint_2[8:8], choice_2, i_2r1[8:8]);
  AND2 I141 (gtint_2[9:9], choice_2, i_2r1[9:9]);
  AND2 I142 (gtint_2[10:10], choice_2, i_2r1[10:10]);
  AND2 I143 (gtint_2[11:11], choice_2, i_2r1[11:11]);
  AND2 I144 (gtint_2[12:12], choice_2, i_2r1[12:12]);
  AND2 I145 (gtint_2[13:13], choice_2, i_2r1[13:13]);
  AND2 I146 (gtint_2[14:14], choice_2, i_2r1[14:14]);
  AND2 I147 (gtint_2[15:15], choice_2, i_2r1[15:15]);
  AND2 I148 (gtint_2[16:16], choice_2, i_2r1[16:16]);
  AND2 I149 (gtint_2[17:17], choice_2, i_2r1[17:17]);
  AND2 I150 (gtint_2[18:18], choice_2, i_2r1[18:18]);
  AND2 I151 (gtint_2[19:19], choice_2, i_2r1[19:19]);
  AND2 I152 (gtint_2[20:20], choice_2, i_2r1[20:20]);
  AND2 I153 (gtint_2[21:21], choice_2, i_2r1[21:21]);
  AND2 I154 (gtint_2[22:22], choice_2, i_2r1[22:22]);
  AND2 I155 (gtint_2[23:23], choice_2, i_2r1[23:23]);
  AND2 I156 (gtint_2[24:24], choice_2, i_2r1[24:24]);
  AND2 I157 (gtint_2[25:25], choice_2, i_2r1[25:25]);
  AND2 I158 (gtint_2[26:26], choice_2, i_2r1[26:26]);
  AND2 I159 (gtint_2[27:27], choice_2, i_2r1[27:27]);
  AND2 I160 (gtint_2[28:28], choice_2, i_2r1[28:28]);
  AND2 I161 (gtint_2[29:29], choice_2, i_2r1[29:29]);
  AND2 I162 (gtint_2[30:30], choice_2, i_2r1[30:30]);
  AND2 I163 (gtint_2[31:31], choice_2, i_2r1[31:31]);
  AND2 I164 (gtint_2[32:32], choice_2, i_2r1[32:32]);
  AND2 I165 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I166 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I167 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I168 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I169 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I170 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I171 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I172 (gfint_0[7:7], choice_0, i_0r0[7:7]);
  AND2 I173 (gfint_0[8:8], choice_0, i_0r0[8:8]);
  AND2 I174 (gfint_0[9:9], choice_0, i_0r0[9:9]);
  AND2 I175 (gfint_0[10:10], choice_0, i_0r0[10:10]);
  AND2 I176 (gfint_0[11:11], choice_0, i_0r0[11:11]);
  AND2 I177 (gfint_0[12:12], choice_0, i_0r0[12:12]);
  AND2 I178 (gfint_0[13:13], choice_0, i_0r0[13:13]);
  AND2 I179 (gfint_0[14:14], choice_0, i_0r0[14:14]);
  AND2 I180 (gfint_0[15:15], choice_0, i_0r0[15:15]);
  AND2 I181 (gfint_0[16:16], choice_0, i_0r0[16:16]);
  AND2 I182 (gfint_0[17:17], choice_0, i_0r0[17:17]);
  AND2 I183 (gfint_0[18:18], choice_0, i_0r0[18:18]);
  AND2 I184 (gfint_0[19:19], choice_0, i_0r0[19:19]);
  AND2 I185 (gfint_0[20:20], choice_0, i_0r0[20:20]);
  AND2 I186 (gfint_0[21:21], choice_0, i_0r0[21:21]);
  AND2 I187 (gfint_0[22:22], choice_0, i_0r0[22:22]);
  AND2 I188 (gfint_0[23:23], choice_0, i_0r0[23:23]);
  AND2 I189 (gfint_0[24:24], choice_0, i_0r0[24:24]);
  AND2 I190 (gfint_0[25:25], choice_0, i_0r0[25:25]);
  AND2 I191 (gfint_0[26:26], choice_0, i_0r0[26:26]);
  AND2 I192 (gfint_0[27:27], choice_0, i_0r0[27:27]);
  AND2 I193 (gfint_0[28:28], choice_0, i_0r0[28:28]);
  AND2 I194 (gfint_0[29:29], choice_0, i_0r0[29:29]);
  AND2 I195 (gfint_0[30:30], choice_0, i_0r0[30:30]);
  AND2 I196 (gfint_0[31:31], choice_0, i_0r0[31:31]);
  AND2 I197 (gfint_0[32:32], choice_0, i_0r0[32:32]);
  AND2 I198 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I199 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I200 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I201 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I202 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I203 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I204 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I205 (gfint_1[7:7], choice_1, i_1r0[7:7]);
  AND2 I206 (gfint_1[8:8], choice_1, i_1r0[8:8]);
  AND2 I207 (gfint_1[9:9], choice_1, i_1r0[9:9]);
  AND2 I208 (gfint_1[10:10], choice_1, i_1r0[10:10]);
  AND2 I209 (gfint_1[11:11], choice_1, i_1r0[11:11]);
  AND2 I210 (gfint_1[12:12], choice_1, i_1r0[12:12]);
  AND2 I211 (gfint_1[13:13], choice_1, i_1r0[13:13]);
  AND2 I212 (gfint_1[14:14], choice_1, i_1r0[14:14]);
  AND2 I213 (gfint_1[15:15], choice_1, i_1r0[15:15]);
  AND2 I214 (gfint_1[16:16], choice_1, i_1r0[16:16]);
  AND2 I215 (gfint_1[17:17], choice_1, i_1r0[17:17]);
  AND2 I216 (gfint_1[18:18], choice_1, i_1r0[18:18]);
  AND2 I217 (gfint_1[19:19], choice_1, i_1r0[19:19]);
  AND2 I218 (gfint_1[20:20], choice_1, i_1r0[20:20]);
  AND2 I219 (gfint_1[21:21], choice_1, i_1r0[21:21]);
  AND2 I220 (gfint_1[22:22], choice_1, i_1r0[22:22]);
  AND2 I221 (gfint_1[23:23], choice_1, i_1r0[23:23]);
  AND2 I222 (gfint_1[24:24], choice_1, i_1r0[24:24]);
  AND2 I223 (gfint_1[25:25], choice_1, i_1r0[25:25]);
  AND2 I224 (gfint_1[26:26], choice_1, i_1r0[26:26]);
  AND2 I225 (gfint_1[27:27], choice_1, i_1r0[27:27]);
  AND2 I226 (gfint_1[28:28], choice_1, i_1r0[28:28]);
  AND2 I227 (gfint_1[29:29], choice_1, i_1r0[29:29]);
  AND2 I228 (gfint_1[30:30], choice_1, i_1r0[30:30]);
  AND2 I229 (gfint_1[31:31], choice_1, i_1r0[31:31]);
  AND2 I230 (gfint_1[32:32], choice_1, i_1r0[32:32]);
  AND2 I231 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I232 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I233 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I234 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AND2 I235 (gfint_2[4:4], choice_2, i_2r0[4:4]);
  AND2 I236 (gfint_2[5:5], choice_2, i_2r0[5:5]);
  AND2 I237 (gfint_2[6:6], choice_2, i_2r0[6:6]);
  AND2 I238 (gfint_2[7:7], choice_2, i_2r0[7:7]);
  AND2 I239 (gfint_2[8:8], choice_2, i_2r0[8:8]);
  AND2 I240 (gfint_2[9:9], choice_2, i_2r0[9:9]);
  AND2 I241 (gfint_2[10:10], choice_2, i_2r0[10:10]);
  AND2 I242 (gfint_2[11:11], choice_2, i_2r0[11:11]);
  AND2 I243 (gfint_2[12:12], choice_2, i_2r0[12:12]);
  AND2 I244 (gfint_2[13:13], choice_2, i_2r0[13:13]);
  AND2 I245 (gfint_2[14:14], choice_2, i_2r0[14:14]);
  AND2 I246 (gfint_2[15:15], choice_2, i_2r0[15:15]);
  AND2 I247 (gfint_2[16:16], choice_2, i_2r0[16:16]);
  AND2 I248 (gfint_2[17:17], choice_2, i_2r0[17:17]);
  AND2 I249 (gfint_2[18:18], choice_2, i_2r0[18:18]);
  AND2 I250 (gfint_2[19:19], choice_2, i_2r0[19:19]);
  AND2 I251 (gfint_2[20:20], choice_2, i_2r0[20:20]);
  AND2 I252 (gfint_2[21:21], choice_2, i_2r0[21:21]);
  AND2 I253 (gfint_2[22:22], choice_2, i_2r0[22:22]);
  AND2 I254 (gfint_2[23:23], choice_2, i_2r0[23:23]);
  AND2 I255 (gfint_2[24:24], choice_2, i_2r0[24:24]);
  AND2 I256 (gfint_2[25:25], choice_2, i_2r0[25:25]);
  AND2 I257 (gfint_2[26:26], choice_2, i_2r0[26:26]);
  AND2 I258 (gfint_2[27:27], choice_2, i_2r0[27:27]);
  AND2 I259 (gfint_2[28:28], choice_2, i_2r0[28:28]);
  AND2 I260 (gfint_2[29:29], choice_2, i_2r0[29:29]);
  AND2 I261 (gfint_2[30:30], choice_2, i_2r0[30:30]);
  AND2 I262 (gfint_2[31:31], choice_2, i_2r0[31:31]);
  AND2 I263 (gfint_2[32:32], choice_2, i_2r0[32:32]);
  OR2 I264 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I265 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I266 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I267 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I268 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I269 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I270 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I271 (comp0_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I272 (comp0_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I273 (comp0_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I274 (comp0_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I275 (comp0_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I276 (comp0_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I277 (comp0_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I278 (comp0_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I279 (comp0_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I280 (comp0_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I281 (comp0_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I282 (comp0_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I283 (comp0_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I284 (comp0_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I285 (comp0_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I286 (comp0_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I287 (comp0_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I288 (comp0_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I289 (comp0_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I290 (comp0_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I291 (comp0_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I292 (comp0_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I293 (comp0_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I294 (comp0_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I295 (comp0_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I296 (comp0_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  C3 I297 (simp3121_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I298 (simp3121_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I299 (simp3121_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I300 (simp3121_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I301 (simp3121_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I302 (simp3121_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I303 (simp3121_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I304 (simp3121_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I305 (simp3121_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I306 (simp3121_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C3 I307 (simp3121_0[10:10], comp0_0[30:30], comp0_0[31:31], comp0_0[32:32]);
  C3 I308 (simp3122_0[0:0], simp3121_0[0:0], simp3121_0[1:1], simp3121_0[2:2]);
  C3 I309 (simp3122_0[1:1], simp3121_0[3:3], simp3121_0[4:4], simp3121_0[5:5]);
  C3 I310 (simp3122_0[2:2], simp3121_0[6:6], simp3121_0[7:7], simp3121_0[8:8]);
  C2 I311 (simp3122_0[3:3], simp3121_0[9:9], simp3121_0[10:10]);
  C3 I312 (simp3123_0[0:0], simp3122_0[0:0], simp3122_0[1:1], simp3122_0[2:2]);
  BUFF I313 (simp3123_0[1:1], simp3122_0[3:3]);
  C2 I314 (icomp_0, simp3123_0[0:0], simp3123_0[1:1]);
  OR2 I315 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I316 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I317 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I318 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I319 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I320 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I321 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  OR2 I322 (comp1_0[7:7], i_1r0[7:7], i_1r1[7:7]);
  OR2 I323 (comp1_0[8:8], i_1r0[8:8], i_1r1[8:8]);
  OR2 I324 (comp1_0[9:9], i_1r0[9:9], i_1r1[9:9]);
  OR2 I325 (comp1_0[10:10], i_1r0[10:10], i_1r1[10:10]);
  OR2 I326 (comp1_0[11:11], i_1r0[11:11], i_1r1[11:11]);
  OR2 I327 (comp1_0[12:12], i_1r0[12:12], i_1r1[12:12]);
  OR2 I328 (comp1_0[13:13], i_1r0[13:13], i_1r1[13:13]);
  OR2 I329 (comp1_0[14:14], i_1r0[14:14], i_1r1[14:14]);
  OR2 I330 (comp1_0[15:15], i_1r0[15:15], i_1r1[15:15]);
  OR2 I331 (comp1_0[16:16], i_1r0[16:16], i_1r1[16:16]);
  OR2 I332 (comp1_0[17:17], i_1r0[17:17], i_1r1[17:17]);
  OR2 I333 (comp1_0[18:18], i_1r0[18:18], i_1r1[18:18]);
  OR2 I334 (comp1_0[19:19], i_1r0[19:19], i_1r1[19:19]);
  OR2 I335 (comp1_0[20:20], i_1r0[20:20], i_1r1[20:20]);
  OR2 I336 (comp1_0[21:21], i_1r0[21:21], i_1r1[21:21]);
  OR2 I337 (comp1_0[22:22], i_1r0[22:22], i_1r1[22:22]);
  OR2 I338 (comp1_0[23:23], i_1r0[23:23], i_1r1[23:23]);
  OR2 I339 (comp1_0[24:24], i_1r0[24:24], i_1r1[24:24]);
  OR2 I340 (comp1_0[25:25], i_1r0[25:25], i_1r1[25:25]);
  OR2 I341 (comp1_0[26:26], i_1r0[26:26], i_1r1[26:26]);
  OR2 I342 (comp1_0[27:27], i_1r0[27:27], i_1r1[27:27]);
  OR2 I343 (comp1_0[28:28], i_1r0[28:28], i_1r1[28:28]);
  OR2 I344 (comp1_0[29:29], i_1r0[29:29], i_1r1[29:29]);
  OR2 I345 (comp1_0[30:30], i_1r0[30:30], i_1r1[30:30]);
  OR2 I346 (comp1_0[31:31], i_1r0[31:31], i_1r1[31:31]);
  OR2 I347 (comp1_0[32:32], i_1r0[32:32], i_1r1[32:32]);
  C3 I348 (simp3471_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I349 (simp3471_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  C3 I350 (simp3471_0[2:2], comp1_0[6:6], comp1_0[7:7], comp1_0[8:8]);
  C3 I351 (simp3471_0[3:3], comp1_0[9:9], comp1_0[10:10], comp1_0[11:11]);
  C3 I352 (simp3471_0[4:4], comp1_0[12:12], comp1_0[13:13], comp1_0[14:14]);
  C3 I353 (simp3471_0[5:5], comp1_0[15:15], comp1_0[16:16], comp1_0[17:17]);
  C3 I354 (simp3471_0[6:6], comp1_0[18:18], comp1_0[19:19], comp1_0[20:20]);
  C3 I355 (simp3471_0[7:7], comp1_0[21:21], comp1_0[22:22], comp1_0[23:23]);
  C3 I356 (simp3471_0[8:8], comp1_0[24:24], comp1_0[25:25], comp1_0[26:26]);
  C3 I357 (simp3471_0[9:9], comp1_0[27:27], comp1_0[28:28], comp1_0[29:29]);
  C3 I358 (simp3471_0[10:10], comp1_0[30:30], comp1_0[31:31], comp1_0[32:32]);
  C3 I359 (simp3472_0[0:0], simp3471_0[0:0], simp3471_0[1:1], simp3471_0[2:2]);
  C3 I360 (simp3472_0[1:1], simp3471_0[3:3], simp3471_0[4:4], simp3471_0[5:5]);
  C3 I361 (simp3472_0[2:2], simp3471_0[6:6], simp3471_0[7:7], simp3471_0[8:8]);
  C2 I362 (simp3472_0[3:3], simp3471_0[9:9], simp3471_0[10:10]);
  C3 I363 (simp3473_0[0:0], simp3472_0[0:0], simp3472_0[1:1], simp3472_0[2:2]);
  BUFF I364 (simp3473_0[1:1], simp3472_0[3:3]);
  C2 I365 (icomp_1, simp3473_0[0:0], simp3473_0[1:1]);
  OR2 I366 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I367 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I368 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2 I369 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  OR2 I370 (comp2_0[4:4], i_2r0[4:4], i_2r1[4:4]);
  OR2 I371 (comp2_0[5:5], i_2r0[5:5], i_2r1[5:5]);
  OR2 I372 (comp2_0[6:6], i_2r0[6:6], i_2r1[6:6]);
  OR2 I373 (comp2_0[7:7], i_2r0[7:7], i_2r1[7:7]);
  OR2 I374 (comp2_0[8:8], i_2r0[8:8], i_2r1[8:8]);
  OR2 I375 (comp2_0[9:9], i_2r0[9:9], i_2r1[9:9]);
  OR2 I376 (comp2_0[10:10], i_2r0[10:10], i_2r1[10:10]);
  OR2 I377 (comp2_0[11:11], i_2r0[11:11], i_2r1[11:11]);
  OR2 I378 (comp2_0[12:12], i_2r0[12:12], i_2r1[12:12]);
  OR2 I379 (comp2_0[13:13], i_2r0[13:13], i_2r1[13:13]);
  OR2 I380 (comp2_0[14:14], i_2r0[14:14], i_2r1[14:14]);
  OR2 I381 (comp2_0[15:15], i_2r0[15:15], i_2r1[15:15]);
  OR2 I382 (comp2_0[16:16], i_2r0[16:16], i_2r1[16:16]);
  OR2 I383 (comp2_0[17:17], i_2r0[17:17], i_2r1[17:17]);
  OR2 I384 (comp2_0[18:18], i_2r0[18:18], i_2r1[18:18]);
  OR2 I385 (comp2_0[19:19], i_2r0[19:19], i_2r1[19:19]);
  OR2 I386 (comp2_0[20:20], i_2r0[20:20], i_2r1[20:20]);
  OR2 I387 (comp2_0[21:21], i_2r0[21:21], i_2r1[21:21]);
  OR2 I388 (comp2_0[22:22], i_2r0[22:22], i_2r1[22:22]);
  OR2 I389 (comp2_0[23:23], i_2r0[23:23], i_2r1[23:23]);
  OR2 I390 (comp2_0[24:24], i_2r0[24:24], i_2r1[24:24]);
  OR2 I391 (comp2_0[25:25], i_2r0[25:25], i_2r1[25:25]);
  OR2 I392 (comp2_0[26:26], i_2r0[26:26], i_2r1[26:26]);
  OR2 I393 (comp2_0[27:27], i_2r0[27:27], i_2r1[27:27]);
  OR2 I394 (comp2_0[28:28], i_2r0[28:28], i_2r1[28:28]);
  OR2 I395 (comp2_0[29:29], i_2r0[29:29], i_2r1[29:29]);
  OR2 I396 (comp2_0[30:30], i_2r0[30:30], i_2r1[30:30]);
  OR2 I397 (comp2_0[31:31], i_2r0[31:31], i_2r1[31:31]);
  OR2 I398 (comp2_0[32:32], i_2r0[32:32], i_2r1[32:32]);
  C3 I399 (simp3821_0[0:0], comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C3 I400 (simp3821_0[1:1], comp2_0[3:3], comp2_0[4:4], comp2_0[5:5]);
  C3 I401 (simp3821_0[2:2], comp2_0[6:6], comp2_0[7:7], comp2_0[8:8]);
  C3 I402 (simp3821_0[3:3], comp2_0[9:9], comp2_0[10:10], comp2_0[11:11]);
  C3 I403 (simp3821_0[4:4], comp2_0[12:12], comp2_0[13:13], comp2_0[14:14]);
  C3 I404 (simp3821_0[5:5], comp2_0[15:15], comp2_0[16:16], comp2_0[17:17]);
  C3 I405 (simp3821_0[6:6], comp2_0[18:18], comp2_0[19:19], comp2_0[20:20]);
  C3 I406 (simp3821_0[7:7], comp2_0[21:21], comp2_0[22:22], comp2_0[23:23]);
  C3 I407 (simp3821_0[8:8], comp2_0[24:24], comp2_0[25:25], comp2_0[26:26]);
  C3 I408 (simp3821_0[9:9], comp2_0[27:27], comp2_0[28:28], comp2_0[29:29]);
  C3 I409 (simp3821_0[10:10], comp2_0[30:30], comp2_0[31:31], comp2_0[32:32]);
  C3 I410 (simp3822_0[0:0], simp3821_0[0:0], simp3821_0[1:1], simp3821_0[2:2]);
  C3 I411 (simp3822_0[1:1], simp3821_0[3:3], simp3821_0[4:4], simp3821_0[5:5]);
  C3 I412 (simp3822_0[2:2], simp3821_0[6:6], simp3821_0[7:7], simp3821_0[8:8]);
  C2 I413 (simp3822_0[3:3], simp3821_0[9:9], simp3821_0[10:10]);
  C3 I414 (simp3823_0[0:0], simp3822_0[0:0], simp3822_0[1:1], simp3822_0[2:2]);
  BUFF I415 (simp3823_0[1:1], simp3822_0[3:3]);
  C2 I416 (icomp_2, simp3823_0[0:0], simp3823_0[1:1]);
  C2R I417 (choice_0, icomp_0, nchosen_0, reset);
  C2R I418 (choice_1, icomp_1, nchosen_0, reset);
  C2R I419 (choice_2, icomp_2, nchosen_0, reset);
  OR3 I420 (anychoice_0, choice_0, choice_1, choice_2);
  NOR2 I421 (nchosen_0, anychoice_0, o_0a);
  C2R I422 (i_0a, choice_0, o_0a, reset);
  C2R I423 (i_1a, choice_1, o_0a, reset);
  C2R I424 (i_2a, choice_2, o_0a, reset);
endmodule

// tkj33m33_0 TeakJ [Many [33,0],One 33]
module tkj33m33_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [32:0] i_0r0;
  input [32:0] i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [32:0] joinf_0;
  wire [32:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joinf_0[32:32], i_0r0[32:32]);
  BUFF I33 (joint_0[0:0], i_0r1[0:0]);
  BUFF I34 (joint_0[1:1], i_0r1[1:1]);
  BUFF I35 (joint_0[2:2], i_0r1[2:2]);
  BUFF I36 (joint_0[3:3], i_0r1[3:3]);
  BUFF I37 (joint_0[4:4], i_0r1[4:4]);
  BUFF I38 (joint_0[5:5], i_0r1[5:5]);
  BUFF I39 (joint_0[6:6], i_0r1[6:6]);
  BUFF I40 (joint_0[7:7], i_0r1[7:7]);
  BUFF I41 (joint_0[8:8], i_0r1[8:8]);
  BUFF I42 (joint_0[9:9], i_0r1[9:9]);
  BUFF I43 (joint_0[10:10], i_0r1[10:10]);
  BUFF I44 (joint_0[11:11], i_0r1[11:11]);
  BUFF I45 (joint_0[12:12], i_0r1[12:12]);
  BUFF I46 (joint_0[13:13], i_0r1[13:13]);
  BUFF I47 (joint_0[14:14], i_0r1[14:14]);
  BUFF I48 (joint_0[15:15], i_0r1[15:15]);
  BUFF I49 (joint_0[16:16], i_0r1[16:16]);
  BUFF I50 (joint_0[17:17], i_0r1[17:17]);
  BUFF I51 (joint_0[18:18], i_0r1[18:18]);
  BUFF I52 (joint_0[19:19], i_0r1[19:19]);
  BUFF I53 (joint_0[20:20], i_0r1[20:20]);
  BUFF I54 (joint_0[21:21], i_0r1[21:21]);
  BUFF I55 (joint_0[22:22], i_0r1[22:22]);
  BUFF I56 (joint_0[23:23], i_0r1[23:23]);
  BUFF I57 (joint_0[24:24], i_0r1[24:24]);
  BUFF I58 (joint_0[25:25], i_0r1[25:25]);
  BUFF I59 (joint_0[26:26], i_0r1[26:26]);
  BUFF I60 (joint_0[27:27], i_0r1[27:27]);
  BUFF I61 (joint_0[28:28], i_0r1[28:28]);
  BUFF I62 (joint_0[29:29], i_0r1[29:29]);
  BUFF I63 (joint_0[30:30], i_0r1[30:30]);
  BUFF I64 (joint_0[31:31], i_0r1[31:31]);
  BUFF I65 (joint_0[32:32], i_0r1[32:32]);
  BUFF I66 (icomplete_0, i_1r);
  C2 I67 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I68 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I69 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I70 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I71 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I72 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I73 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I74 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I75 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I76 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I77 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I78 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I79 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I80 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I81 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I82 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I83 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I84 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I85 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I86 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I87 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I88 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I89 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I90 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I91 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I92 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I93 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I94 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I95 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I96 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I97 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I98 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I99 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I100 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I101 (o_0r1[1:1], joint_0[1:1]);
  BUFF I102 (o_0r1[2:2], joint_0[2:2]);
  BUFF I103 (o_0r1[3:3], joint_0[3:3]);
  BUFF I104 (o_0r1[4:4], joint_0[4:4]);
  BUFF I105 (o_0r1[5:5], joint_0[5:5]);
  BUFF I106 (o_0r1[6:6], joint_0[6:6]);
  BUFF I107 (o_0r1[7:7], joint_0[7:7]);
  BUFF I108 (o_0r1[8:8], joint_0[8:8]);
  BUFF I109 (o_0r1[9:9], joint_0[9:9]);
  BUFF I110 (o_0r1[10:10], joint_0[10:10]);
  BUFF I111 (o_0r1[11:11], joint_0[11:11]);
  BUFF I112 (o_0r1[12:12], joint_0[12:12]);
  BUFF I113 (o_0r1[13:13], joint_0[13:13]);
  BUFF I114 (o_0r1[14:14], joint_0[14:14]);
  BUFF I115 (o_0r1[15:15], joint_0[15:15]);
  BUFF I116 (o_0r1[16:16], joint_0[16:16]);
  BUFF I117 (o_0r1[17:17], joint_0[17:17]);
  BUFF I118 (o_0r1[18:18], joint_0[18:18]);
  BUFF I119 (o_0r1[19:19], joint_0[19:19]);
  BUFF I120 (o_0r1[20:20], joint_0[20:20]);
  BUFF I121 (o_0r1[21:21], joint_0[21:21]);
  BUFF I122 (o_0r1[22:22], joint_0[22:22]);
  BUFF I123 (o_0r1[23:23], joint_0[23:23]);
  BUFF I124 (o_0r1[24:24], joint_0[24:24]);
  BUFF I125 (o_0r1[25:25], joint_0[25:25]);
  BUFF I126 (o_0r1[26:26], joint_0[26:26]);
  BUFF I127 (o_0r1[27:27], joint_0[27:27]);
  BUFF I128 (o_0r1[28:28], joint_0[28:28]);
  BUFF I129 (o_0r1[29:29], joint_0[29:29]);
  BUFF I130 (o_0r1[30:30], joint_0[30:30]);
  BUFF I131 (o_0r1[31:31], joint_0[31:31]);
  BUFF I132 (o_0r1[32:32], joint_0[32:32]);
  BUFF I133 (i_0a, o_0a);
  BUFF I134 (i_1a, o_0a);
endmodule

// tkvpostRhs32_wo0w32_ro0w32o31w1o0w5o31w1 TeakV "postRhs" 32 [] [0] [0,31,0,31] [Many [32],Many [0],M
//   any [0,0,0,0],Many [32,1,5,1]]
module tkvpostRhs32_wo0w32_ro0w32o31w1o0w5o31w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output rd_1r0;
  output rd_1r1;
  input rd_1a;
  output [4:0] rd_2r0;
  output [4:0] rd_2r1;
  input rd_2a;
  output rd_3r0;
  output rd_3r1;
  input rd_3a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [2:0] simp4861_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0, df_0[31:31], rg_1r);
  AND2 I457 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I458 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I459 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I460 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I461 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I462 (rd_3r0, df_0[31:31], rg_3r);
  AND2 I463 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I464 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I465 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I466 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I467 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I468 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I469 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I470 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I471 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I472 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I473 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I474 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I475 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I476 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I477 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I478 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I479 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I480 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I481 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I482 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I483 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I484 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I485 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I486 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I487 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I488 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I489 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I490 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I491 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I492 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I493 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I494 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I495 (rd_1r1, dt_0[31:31], rg_1r);
  AND2 I496 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I497 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I498 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I499 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I500 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I501 (rd_3r1, dt_0[31:31], rg_3r);
  NOR3 I502 (simp4861_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I503 (simp4861_0[1:1], rg_3r, rg_0a, rg_1a);
  NOR2 I504 (simp4861_0[2:2], rg_2a, rg_3a);
  NAND3 I505 (anyread_0, simp4861_0[0:0], simp4861_0[1:1], simp4861_0[2:2]);
  BUFF I506 (wg_0a, wd_0a);
  BUFF I507 (rg_0a, rd_0a);
  BUFF I508 (rg_1a, rd_1a);
  BUFF I509 (rg_2a, rd_2a);
  BUFF I510 (rg_3a, rd_3a);
endmodule

// tkvaddCarryIn1_wo0w1_ro0w1o0w1 TeakV "addCarryIn" 1 [] [0] [0,0] [Many [1],Many [0],Many [0,0],Many 
//   [1,1]]
module tkvaddCarryIn1_wo0w1_ro0w1o0w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, reset);
  input wg_0r0;
  input wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  output rd_1r0;
  output rd_1r1;
  input rd_1a;
  input reset;
  wire wf_0;
  wire wt_0;
  wire df_0;
  wire dt_0;
  wire wc_0;
  wire wacks_0;
  wire wenr_0;
  wire wen_0;
  wire anyread_0;
  wire nreset_0;
  wire drlgf_0;
  wire drlgt_0;
  wire comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire conwgit_0;
  wire conwgif_0;
  wire conwig_0;
  wire [1:0] simp401_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0, wenr_0, nreset_0);
  AND2 I2 (drlgf_0, wf_0, wen_0);
  AND2 I3 (drlgt_0, wt_0, wen_0);
  NOR2 I4 (df_0, dt_0, drlgt_0);
  NOR3 I5 (dt_0, df_0, drlgf_0, reset);
  AO22 I6 (wacks_0, drlgf_0, df_0, drlgt_0, dt_0);
  OR2 I7 (comp0_0, wg_0r0, wg_0r1);
  BUFF I8 (wc_0, comp0_0);
  AND2 I9 (conwgif_0, wg_0r0, conwig_0);
  AND2 I10 (conwgit_0, wg_0r1, conwig_0);
  BUFF I11 (conwigc_0, wc_0);
  AO22 I12 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I13 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I14 (wf_0, conwgif_0);
  BUFF I15 (wt_0, conwgit_0);
  BUFF I16 (wenr_0, wc_0);
  C2 I17 (wd_0r, conwig_0, wacks_0);
  AND2 I18 (rd_0r0, df_0, rg_0r);
  AND2 I19 (rd_1r0, df_0, rg_1r);
  AND2 I20 (rd_0r1, dt_0, rg_0r);
  AND2 I21 (rd_1r1, dt_0, rg_1r);
  NOR3 I22 (simp401_0[0:0], rg_0r, rg_1r, rg_0a);
  INV I23 (simp401_0[1:1], rg_1a);
  NAND2 I24 (anyread_0, simp401_0[0:0], simp401_0[1:1]);
  BUFF I25 (wg_0a, wd_0a);
  BUFF I26 (rg_0a, rd_0a);
  BUFF I27 (rg_1a, rd_1a);
endmodule

// tkvop7_wo0w7_ro0w6o0w6o6w1o6w1o0w6o0w6o0w6 TeakV "op" 7 [] [0] [0,0,6,6,0,0,0] [Many [7],Many [0],Ma
//   ny [0,0,0,0,0,0,0],Many [6,6,1,1,6,6,6]]
module tkvop7_wo0w7_ro0w6o0w6o6w1o6w1o0w6o0w6o0w6 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rg_5r, rg_5a, rg_6r, rg_6a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, rd_5r0, rd_5r1, rd_5a, rd_6r0, rd_6r1, rd_6a, reset);
  input [6:0] wg_0r0;
  input [6:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  input rg_5r;
  output rg_5a;
  input rg_6r;
  output rg_6a;
  output [5:0] rd_0r0;
  output [5:0] rd_0r1;
  input rd_0a;
  output [5:0] rd_1r0;
  output [5:0] rd_1r1;
  input rd_1a;
  output rd_2r0;
  output rd_2r1;
  input rd_2a;
  output rd_3r0;
  output rd_3r1;
  input rd_3a;
  output [5:0] rd_4r0;
  output [5:0] rd_4r1;
  input rd_4a;
  output [5:0] rd_5r0;
  output [5:0] rd_5r1;
  input rd_5a;
  output [5:0] rd_6r0;
  output [5:0] rd_6r1;
  input rd_6a;
  input reset;
  wire [6:0] wf_0;
  wire [6:0] wt_0;
  wire [6:0] df_0;
  wire [6:0] dt_0;
  wire wc_0;
  wire [6:0] wacks_0;
  wire [6:0] wenr_0;
  wire [6:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [6:0] drlgf_0;
  wire [6:0] drlgt_0;
  wire [6:0] comp0_0;
  wire [2:0] simp631_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [6:0] conwgit_0;
  wire [6:0] conwgif_0;
  wire conwig_0;
  wire [2:0] simp1071_0;
  wire [4:0] simp1721_0;
  wire [1:0] simp1722_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I9 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I10 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I11 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I12 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I13 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I14 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I15 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I16 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I17 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I18 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I19 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I20 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I21 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  NOR2 I22 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I23 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I24 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I25 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I26 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I27 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I28 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR3 I29 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I30 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I31 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I32 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I33 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I34 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I35 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  AO22 I36 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I37 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I38 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I39 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I40 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I41 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I42 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  OR2 I43 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I44 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I45 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I46 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I47 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I48 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I49 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  C3 I50 (simp631_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I51 (simp631_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  BUFF I52 (simp631_0[2:2], comp0_0[6:6]);
  C3 I53 (wc_0, simp631_0[0:0], simp631_0[1:1], simp631_0[2:2]);
  AND2 I54 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I55 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I56 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I57 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I58 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I59 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I60 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I61 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I62 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I63 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I64 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I65 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I66 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I67 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  BUFF I68 (conwigc_0, wc_0);
  AO22 I69 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I70 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I71 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I72 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I73 (wenr_0[0:0], wc_0);
  BUFF I74 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I75 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I76 (wenr_0[1:1], wc_0);
  BUFF I77 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I78 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I79 (wenr_0[2:2], wc_0);
  BUFF I80 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I81 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I82 (wenr_0[3:3], wc_0);
  BUFF I83 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I84 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I85 (wenr_0[4:4], wc_0);
  BUFF I86 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I87 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I88 (wenr_0[5:5], wc_0);
  BUFF I89 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I90 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I91 (wenr_0[6:6], wc_0);
  C3 I92 (simp1071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I93 (simp1071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C2 I94 (simp1071_0[2:2], wacks_0[5:5], wacks_0[6:6]);
  C3 I95 (wd_0r, simp1071_0[0:0], simp1071_0[1:1], simp1071_0[2:2]);
  AND2 I96 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I97 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I98 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I99 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I100 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I101 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I102 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I103 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I104 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I105 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I106 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I107 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I108 (rd_2r0, df_0[6:6], rg_2r);
  AND2 I109 (rd_3r0, df_0[6:6], rg_3r);
  AND2 I110 (rd_4r0[0:0], df_0[0:0], rg_4r);
  AND2 I111 (rd_4r0[1:1], df_0[1:1], rg_4r);
  AND2 I112 (rd_4r0[2:2], df_0[2:2], rg_4r);
  AND2 I113 (rd_4r0[3:3], df_0[3:3], rg_4r);
  AND2 I114 (rd_4r0[4:4], df_0[4:4], rg_4r);
  AND2 I115 (rd_4r0[5:5], df_0[5:5], rg_4r);
  AND2 I116 (rd_5r0[0:0], df_0[0:0], rg_5r);
  AND2 I117 (rd_5r0[1:1], df_0[1:1], rg_5r);
  AND2 I118 (rd_5r0[2:2], df_0[2:2], rg_5r);
  AND2 I119 (rd_5r0[3:3], df_0[3:3], rg_5r);
  AND2 I120 (rd_5r0[4:4], df_0[4:4], rg_5r);
  AND2 I121 (rd_5r0[5:5], df_0[5:5], rg_5r);
  AND2 I122 (rd_6r0[0:0], df_0[0:0], rg_6r);
  AND2 I123 (rd_6r0[1:1], df_0[1:1], rg_6r);
  AND2 I124 (rd_6r0[2:2], df_0[2:2], rg_6r);
  AND2 I125 (rd_6r0[3:3], df_0[3:3], rg_6r);
  AND2 I126 (rd_6r0[4:4], df_0[4:4], rg_6r);
  AND2 I127 (rd_6r0[5:5], df_0[5:5], rg_6r);
  AND2 I128 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I129 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I130 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I131 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I132 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I133 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I134 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I135 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I136 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I137 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I138 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I139 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I140 (rd_2r1, dt_0[6:6], rg_2r);
  AND2 I141 (rd_3r1, dt_0[6:6], rg_3r);
  AND2 I142 (rd_4r1[0:0], dt_0[0:0], rg_4r);
  AND2 I143 (rd_4r1[1:1], dt_0[1:1], rg_4r);
  AND2 I144 (rd_4r1[2:2], dt_0[2:2], rg_4r);
  AND2 I145 (rd_4r1[3:3], dt_0[3:3], rg_4r);
  AND2 I146 (rd_4r1[4:4], dt_0[4:4], rg_4r);
  AND2 I147 (rd_4r1[5:5], dt_0[5:5], rg_4r);
  AND2 I148 (rd_5r1[0:0], dt_0[0:0], rg_5r);
  AND2 I149 (rd_5r1[1:1], dt_0[1:1], rg_5r);
  AND2 I150 (rd_5r1[2:2], dt_0[2:2], rg_5r);
  AND2 I151 (rd_5r1[3:3], dt_0[3:3], rg_5r);
  AND2 I152 (rd_5r1[4:4], dt_0[4:4], rg_5r);
  AND2 I153 (rd_5r1[5:5], dt_0[5:5], rg_5r);
  AND2 I154 (rd_6r1[0:0], dt_0[0:0], rg_6r);
  AND2 I155 (rd_6r1[1:1], dt_0[1:1], rg_6r);
  AND2 I156 (rd_6r1[2:2], dt_0[2:2], rg_6r);
  AND2 I157 (rd_6r1[3:3], dt_0[3:3], rg_6r);
  AND2 I158 (rd_6r1[4:4], dt_0[4:4], rg_6r);
  AND2 I159 (rd_6r1[5:5], dt_0[5:5], rg_6r);
  NOR3 I160 (simp1721_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I161 (simp1721_0[1:1], rg_3r, rg_4r, rg_5r);
  NOR3 I162 (simp1721_0[2:2], rg_6r, rg_0a, rg_1a);
  NOR3 I163 (simp1721_0[3:3], rg_2a, rg_3a, rg_4a);
  NOR2 I164 (simp1721_0[4:4], rg_5a, rg_6a);
  NAND3 I165 (simp1722_0[0:0], simp1721_0[0:0], simp1721_0[1:1], simp1721_0[2:2]);
  NAND2 I166 (simp1722_0[1:1], simp1721_0[3:3], simp1721_0[4:4]);
  OR2 I167 (anyread_0, simp1722_0[0:0], simp1722_0[1:1]);
  BUFF I168 (wg_0a, wd_0a);
  BUFF I169 (rg_0a, rd_0a);
  BUFF I170 (rg_1a, rd_1a);
  BUFF I171 (rg_2a, rd_2a);
  BUFF I172 (rg_3a, rd_3a);
  BUFF I173 (rg_4a, rd_4a);
  BUFF I174 (rg_5a, rd_5a);
  BUFF I175 (rg_6a, rd_6a);
endmodule

// tkvlhs32_wo0w32_ro0w32o0w32o0w32o0w32o0w32o31w1 TeakV "lhs" 32 [] [0] [0,0,0,0,0,31] [Many [32],Many
//    [0],Many [0,0,0,0,0,0],Many [32,32,32,32,32,1]]
module tkvlhs32_wo0w32_ro0w32o0w32o0w32o0w32o0w32o31w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rg_5r, rg_5a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, rd_5r0, rd_5r1, rd_5a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  input rg_5r;
  output rg_5a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  output [31:0] rd_3r0;
  output [31:0] rd_3r1;
  input rd_3a;
  output [31:0] rd_4r0;
  output [31:0] rd_4r1;
  input rd_4a;
  output rd_5r0;
  output rd_5r1;
  input rd_5a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [3:0] simp7301_0;
  wire [1:0] simp7302_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_3r0[0:0], df_0[0:0], rg_3r);
  AND2 I521 (rd_3r0[1:1], df_0[1:1], rg_3r);
  AND2 I522 (rd_3r0[2:2], df_0[2:2], rg_3r);
  AND2 I523 (rd_3r0[3:3], df_0[3:3], rg_3r);
  AND2 I524 (rd_3r0[4:4], df_0[4:4], rg_3r);
  AND2 I525 (rd_3r0[5:5], df_0[5:5], rg_3r);
  AND2 I526 (rd_3r0[6:6], df_0[6:6], rg_3r);
  AND2 I527 (rd_3r0[7:7], df_0[7:7], rg_3r);
  AND2 I528 (rd_3r0[8:8], df_0[8:8], rg_3r);
  AND2 I529 (rd_3r0[9:9], df_0[9:9], rg_3r);
  AND2 I530 (rd_3r0[10:10], df_0[10:10], rg_3r);
  AND2 I531 (rd_3r0[11:11], df_0[11:11], rg_3r);
  AND2 I532 (rd_3r0[12:12], df_0[12:12], rg_3r);
  AND2 I533 (rd_3r0[13:13], df_0[13:13], rg_3r);
  AND2 I534 (rd_3r0[14:14], df_0[14:14], rg_3r);
  AND2 I535 (rd_3r0[15:15], df_0[15:15], rg_3r);
  AND2 I536 (rd_3r0[16:16], df_0[16:16], rg_3r);
  AND2 I537 (rd_3r0[17:17], df_0[17:17], rg_3r);
  AND2 I538 (rd_3r0[18:18], df_0[18:18], rg_3r);
  AND2 I539 (rd_3r0[19:19], df_0[19:19], rg_3r);
  AND2 I540 (rd_3r0[20:20], df_0[20:20], rg_3r);
  AND2 I541 (rd_3r0[21:21], df_0[21:21], rg_3r);
  AND2 I542 (rd_3r0[22:22], df_0[22:22], rg_3r);
  AND2 I543 (rd_3r0[23:23], df_0[23:23], rg_3r);
  AND2 I544 (rd_3r0[24:24], df_0[24:24], rg_3r);
  AND2 I545 (rd_3r0[25:25], df_0[25:25], rg_3r);
  AND2 I546 (rd_3r0[26:26], df_0[26:26], rg_3r);
  AND2 I547 (rd_3r0[27:27], df_0[27:27], rg_3r);
  AND2 I548 (rd_3r0[28:28], df_0[28:28], rg_3r);
  AND2 I549 (rd_3r0[29:29], df_0[29:29], rg_3r);
  AND2 I550 (rd_3r0[30:30], df_0[30:30], rg_3r);
  AND2 I551 (rd_3r0[31:31], df_0[31:31], rg_3r);
  AND2 I552 (rd_4r0[0:0], df_0[0:0], rg_4r);
  AND2 I553 (rd_4r0[1:1], df_0[1:1], rg_4r);
  AND2 I554 (rd_4r0[2:2], df_0[2:2], rg_4r);
  AND2 I555 (rd_4r0[3:3], df_0[3:3], rg_4r);
  AND2 I556 (rd_4r0[4:4], df_0[4:4], rg_4r);
  AND2 I557 (rd_4r0[5:5], df_0[5:5], rg_4r);
  AND2 I558 (rd_4r0[6:6], df_0[6:6], rg_4r);
  AND2 I559 (rd_4r0[7:7], df_0[7:7], rg_4r);
  AND2 I560 (rd_4r0[8:8], df_0[8:8], rg_4r);
  AND2 I561 (rd_4r0[9:9], df_0[9:9], rg_4r);
  AND2 I562 (rd_4r0[10:10], df_0[10:10], rg_4r);
  AND2 I563 (rd_4r0[11:11], df_0[11:11], rg_4r);
  AND2 I564 (rd_4r0[12:12], df_0[12:12], rg_4r);
  AND2 I565 (rd_4r0[13:13], df_0[13:13], rg_4r);
  AND2 I566 (rd_4r0[14:14], df_0[14:14], rg_4r);
  AND2 I567 (rd_4r0[15:15], df_0[15:15], rg_4r);
  AND2 I568 (rd_4r0[16:16], df_0[16:16], rg_4r);
  AND2 I569 (rd_4r0[17:17], df_0[17:17], rg_4r);
  AND2 I570 (rd_4r0[18:18], df_0[18:18], rg_4r);
  AND2 I571 (rd_4r0[19:19], df_0[19:19], rg_4r);
  AND2 I572 (rd_4r0[20:20], df_0[20:20], rg_4r);
  AND2 I573 (rd_4r0[21:21], df_0[21:21], rg_4r);
  AND2 I574 (rd_4r0[22:22], df_0[22:22], rg_4r);
  AND2 I575 (rd_4r0[23:23], df_0[23:23], rg_4r);
  AND2 I576 (rd_4r0[24:24], df_0[24:24], rg_4r);
  AND2 I577 (rd_4r0[25:25], df_0[25:25], rg_4r);
  AND2 I578 (rd_4r0[26:26], df_0[26:26], rg_4r);
  AND2 I579 (rd_4r0[27:27], df_0[27:27], rg_4r);
  AND2 I580 (rd_4r0[28:28], df_0[28:28], rg_4r);
  AND2 I581 (rd_4r0[29:29], df_0[29:29], rg_4r);
  AND2 I582 (rd_4r0[30:30], df_0[30:30], rg_4r);
  AND2 I583 (rd_4r0[31:31], df_0[31:31], rg_4r);
  AND2 I584 (rd_5r0, df_0[31:31], rg_5r);
  AND2 I585 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I586 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I587 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I588 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I589 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I590 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I591 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I592 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I593 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I594 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I595 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I596 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I597 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I598 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I599 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I600 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I601 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I602 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I603 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I604 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I605 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I606 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I607 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I608 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I609 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I610 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I611 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I612 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I613 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I614 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I615 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I616 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I617 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I618 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I619 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I620 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I621 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I622 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I623 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I624 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I625 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I626 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I627 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I628 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I629 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I630 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I631 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I632 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I633 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I634 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I635 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I636 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I637 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I638 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I639 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I640 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I641 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I642 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I643 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I644 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I645 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I646 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I647 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I648 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I649 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I650 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I651 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I652 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I653 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I654 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I655 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I656 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I657 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I658 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I659 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I660 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I661 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I662 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I663 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I664 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I665 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I666 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I667 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I668 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I669 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I670 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I671 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I672 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I673 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I674 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I675 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I676 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I677 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I678 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I679 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I680 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  AND2 I681 (rd_3r1[0:0], dt_0[0:0], rg_3r);
  AND2 I682 (rd_3r1[1:1], dt_0[1:1], rg_3r);
  AND2 I683 (rd_3r1[2:2], dt_0[2:2], rg_3r);
  AND2 I684 (rd_3r1[3:3], dt_0[3:3], rg_3r);
  AND2 I685 (rd_3r1[4:4], dt_0[4:4], rg_3r);
  AND2 I686 (rd_3r1[5:5], dt_0[5:5], rg_3r);
  AND2 I687 (rd_3r1[6:6], dt_0[6:6], rg_3r);
  AND2 I688 (rd_3r1[7:7], dt_0[7:7], rg_3r);
  AND2 I689 (rd_3r1[8:8], dt_0[8:8], rg_3r);
  AND2 I690 (rd_3r1[9:9], dt_0[9:9], rg_3r);
  AND2 I691 (rd_3r1[10:10], dt_0[10:10], rg_3r);
  AND2 I692 (rd_3r1[11:11], dt_0[11:11], rg_3r);
  AND2 I693 (rd_3r1[12:12], dt_0[12:12], rg_3r);
  AND2 I694 (rd_3r1[13:13], dt_0[13:13], rg_3r);
  AND2 I695 (rd_3r1[14:14], dt_0[14:14], rg_3r);
  AND2 I696 (rd_3r1[15:15], dt_0[15:15], rg_3r);
  AND2 I697 (rd_3r1[16:16], dt_0[16:16], rg_3r);
  AND2 I698 (rd_3r1[17:17], dt_0[17:17], rg_3r);
  AND2 I699 (rd_3r1[18:18], dt_0[18:18], rg_3r);
  AND2 I700 (rd_3r1[19:19], dt_0[19:19], rg_3r);
  AND2 I701 (rd_3r1[20:20], dt_0[20:20], rg_3r);
  AND2 I702 (rd_3r1[21:21], dt_0[21:21], rg_3r);
  AND2 I703 (rd_3r1[22:22], dt_0[22:22], rg_3r);
  AND2 I704 (rd_3r1[23:23], dt_0[23:23], rg_3r);
  AND2 I705 (rd_3r1[24:24], dt_0[24:24], rg_3r);
  AND2 I706 (rd_3r1[25:25], dt_0[25:25], rg_3r);
  AND2 I707 (rd_3r1[26:26], dt_0[26:26], rg_3r);
  AND2 I708 (rd_3r1[27:27], dt_0[27:27], rg_3r);
  AND2 I709 (rd_3r1[28:28], dt_0[28:28], rg_3r);
  AND2 I710 (rd_3r1[29:29], dt_0[29:29], rg_3r);
  AND2 I711 (rd_3r1[30:30], dt_0[30:30], rg_3r);
  AND2 I712 (rd_3r1[31:31], dt_0[31:31], rg_3r);
  AND2 I713 (rd_4r1[0:0], dt_0[0:0], rg_4r);
  AND2 I714 (rd_4r1[1:1], dt_0[1:1], rg_4r);
  AND2 I715 (rd_4r1[2:2], dt_0[2:2], rg_4r);
  AND2 I716 (rd_4r1[3:3], dt_0[3:3], rg_4r);
  AND2 I717 (rd_4r1[4:4], dt_0[4:4], rg_4r);
  AND2 I718 (rd_4r1[5:5], dt_0[5:5], rg_4r);
  AND2 I719 (rd_4r1[6:6], dt_0[6:6], rg_4r);
  AND2 I720 (rd_4r1[7:7], dt_0[7:7], rg_4r);
  AND2 I721 (rd_4r1[8:8], dt_0[8:8], rg_4r);
  AND2 I722 (rd_4r1[9:9], dt_0[9:9], rg_4r);
  AND2 I723 (rd_4r1[10:10], dt_0[10:10], rg_4r);
  AND2 I724 (rd_4r1[11:11], dt_0[11:11], rg_4r);
  AND2 I725 (rd_4r1[12:12], dt_0[12:12], rg_4r);
  AND2 I726 (rd_4r1[13:13], dt_0[13:13], rg_4r);
  AND2 I727 (rd_4r1[14:14], dt_0[14:14], rg_4r);
  AND2 I728 (rd_4r1[15:15], dt_0[15:15], rg_4r);
  AND2 I729 (rd_4r1[16:16], dt_0[16:16], rg_4r);
  AND2 I730 (rd_4r1[17:17], dt_0[17:17], rg_4r);
  AND2 I731 (rd_4r1[18:18], dt_0[18:18], rg_4r);
  AND2 I732 (rd_4r1[19:19], dt_0[19:19], rg_4r);
  AND2 I733 (rd_4r1[20:20], dt_0[20:20], rg_4r);
  AND2 I734 (rd_4r1[21:21], dt_0[21:21], rg_4r);
  AND2 I735 (rd_4r1[22:22], dt_0[22:22], rg_4r);
  AND2 I736 (rd_4r1[23:23], dt_0[23:23], rg_4r);
  AND2 I737 (rd_4r1[24:24], dt_0[24:24], rg_4r);
  AND2 I738 (rd_4r1[25:25], dt_0[25:25], rg_4r);
  AND2 I739 (rd_4r1[26:26], dt_0[26:26], rg_4r);
  AND2 I740 (rd_4r1[27:27], dt_0[27:27], rg_4r);
  AND2 I741 (rd_4r1[28:28], dt_0[28:28], rg_4r);
  AND2 I742 (rd_4r1[29:29], dt_0[29:29], rg_4r);
  AND2 I743 (rd_4r1[30:30], dt_0[30:30], rg_4r);
  AND2 I744 (rd_4r1[31:31], dt_0[31:31], rg_4r);
  AND2 I745 (rd_5r1, dt_0[31:31], rg_5r);
  NOR3 I746 (simp7301_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I747 (simp7301_0[1:1], rg_3r, rg_4r, rg_5r);
  NOR3 I748 (simp7301_0[2:2], rg_0a, rg_1a, rg_2a);
  NOR3 I749 (simp7301_0[3:3], rg_3a, rg_4a, rg_5a);
  NAND3 I750 (simp7302_0[0:0], simp7301_0[0:0], simp7301_0[1:1], simp7301_0[2:2]);
  INV I751 (simp7302_0[1:1], simp7301_0[3:3]);
  OR2 I752 (anyread_0, simp7302_0[0:0], simp7302_0[1:1]);
  BUFF I753 (wg_0a, wd_0a);
  BUFF I754 (rg_0a, rd_0a);
  BUFF I755 (rg_1a, rd_1a);
  BUFF I756 (rg_2a, rd_2a);
  BUFF I757 (rg_3a, rd_3a);
  BUFF I758 (rg_4a, rd_4a);
  BUFF I759 (rg_5a, rd_5a);
endmodule

// tkvrhs32_wo0w32_ro0w32o0w32o0w32o0w32o0w32 TeakV "rhs" 32 [] [0] [0,0,0,0,0] [Many [32],Many [0],Man
//   y [0,0,0,0,0],Many [32,32,32,32,32]]
module tkvrhs32_wo0w32_ro0w32o0w32o0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  output [31:0] rd_3r0;
  output [31:0] rd_3r1;
  input rd_3a;
  output [31:0] rd_4r0;
  output [31:0] rd_4r1;
  input rd_4a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [3:0] simp7281_0;
  wire [1:0] simp7282_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_3r0[0:0], df_0[0:0], rg_3r);
  AND2 I521 (rd_3r0[1:1], df_0[1:1], rg_3r);
  AND2 I522 (rd_3r0[2:2], df_0[2:2], rg_3r);
  AND2 I523 (rd_3r0[3:3], df_0[3:3], rg_3r);
  AND2 I524 (rd_3r0[4:4], df_0[4:4], rg_3r);
  AND2 I525 (rd_3r0[5:5], df_0[5:5], rg_3r);
  AND2 I526 (rd_3r0[6:6], df_0[6:6], rg_3r);
  AND2 I527 (rd_3r0[7:7], df_0[7:7], rg_3r);
  AND2 I528 (rd_3r0[8:8], df_0[8:8], rg_3r);
  AND2 I529 (rd_3r0[9:9], df_0[9:9], rg_3r);
  AND2 I530 (rd_3r0[10:10], df_0[10:10], rg_3r);
  AND2 I531 (rd_3r0[11:11], df_0[11:11], rg_3r);
  AND2 I532 (rd_3r0[12:12], df_0[12:12], rg_3r);
  AND2 I533 (rd_3r0[13:13], df_0[13:13], rg_3r);
  AND2 I534 (rd_3r0[14:14], df_0[14:14], rg_3r);
  AND2 I535 (rd_3r0[15:15], df_0[15:15], rg_3r);
  AND2 I536 (rd_3r0[16:16], df_0[16:16], rg_3r);
  AND2 I537 (rd_3r0[17:17], df_0[17:17], rg_3r);
  AND2 I538 (rd_3r0[18:18], df_0[18:18], rg_3r);
  AND2 I539 (rd_3r0[19:19], df_0[19:19], rg_3r);
  AND2 I540 (rd_3r0[20:20], df_0[20:20], rg_3r);
  AND2 I541 (rd_3r0[21:21], df_0[21:21], rg_3r);
  AND2 I542 (rd_3r0[22:22], df_0[22:22], rg_3r);
  AND2 I543 (rd_3r0[23:23], df_0[23:23], rg_3r);
  AND2 I544 (rd_3r0[24:24], df_0[24:24], rg_3r);
  AND2 I545 (rd_3r0[25:25], df_0[25:25], rg_3r);
  AND2 I546 (rd_3r0[26:26], df_0[26:26], rg_3r);
  AND2 I547 (rd_3r0[27:27], df_0[27:27], rg_3r);
  AND2 I548 (rd_3r0[28:28], df_0[28:28], rg_3r);
  AND2 I549 (rd_3r0[29:29], df_0[29:29], rg_3r);
  AND2 I550 (rd_3r0[30:30], df_0[30:30], rg_3r);
  AND2 I551 (rd_3r0[31:31], df_0[31:31], rg_3r);
  AND2 I552 (rd_4r0[0:0], df_0[0:0], rg_4r);
  AND2 I553 (rd_4r0[1:1], df_0[1:1], rg_4r);
  AND2 I554 (rd_4r0[2:2], df_0[2:2], rg_4r);
  AND2 I555 (rd_4r0[3:3], df_0[3:3], rg_4r);
  AND2 I556 (rd_4r0[4:4], df_0[4:4], rg_4r);
  AND2 I557 (rd_4r0[5:5], df_0[5:5], rg_4r);
  AND2 I558 (rd_4r0[6:6], df_0[6:6], rg_4r);
  AND2 I559 (rd_4r0[7:7], df_0[7:7], rg_4r);
  AND2 I560 (rd_4r0[8:8], df_0[8:8], rg_4r);
  AND2 I561 (rd_4r0[9:9], df_0[9:9], rg_4r);
  AND2 I562 (rd_4r0[10:10], df_0[10:10], rg_4r);
  AND2 I563 (rd_4r0[11:11], df_0[11:11], rg_4r);
  AND2 I564 (rd_4r0[12:12], df_0[12:12], rg_4r);
  AND2 I565 (rd_4r0[13:13], df_0[13:13], rg_4r);
  AND2 I566 (rd_4r0[14:14], df_0[14:14], rg_4r);
  AND2 I567 (rd_4r0[15:15], df_0[15:15], rg_4r);
  AND2 I568 (rd_4r0[16:16], df_0[16:16], rg_4r);
  AND2 I569 (rd_4r0[17:17], df_0[17:17], rg_4r);
  AND2 I570 (rd_4r0[18:18], df_0[18:18], rg_4r);
  AND2 I571 (rd_4r0[19:19], df_0[19:19], rg_4r);
  AND2 I572 (rd_4r0[20:20], df_0[20:20], rg_4r);
  AND2 I573 (rd_4r0[21:21], df_0[21:21], rg_4r);
  AND2 I574 (rd_4r0[22:22], df_0[22:22], rg_4r);
  AND2 I575 (rd_4r0[23:23], df_0[23:23], rg_4r);
  AND2 I576 (rd_4r0[24:24], df_0[24:24], rg_4r);
  AND2 I577 (rd_4r0[25:25], df_0[25:25], rg_4r);
  AND2 I578 (rd_4r0[26:26], df_0[26:26], rg_4r);
  AND2 I579 (rd_4r0[27:27], df_0[27:27], rg_4r);
  AND2 I580 (rd_4r0[28:28], df_0[28:28], rg_4r);
  AND2 I581 (rd_4r0[29:29], df_0[29:29], rg_4r);
  AND2 I582 (rd_4r0[30:30], df_0[30:30], rg_4r);
  AND2 I583 (rd_4r0[31:31], df_0[31:31], rg_4r);
  AND2 I584 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I585 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I586 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I587 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I588 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I589 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I590 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I591 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I592 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I593 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I594 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I595 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I596 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I597 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I598 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I599 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I600 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I601 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I602 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I603 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I604 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I605 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I606 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I607 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I608 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I609 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I610 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I611 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I612 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I613 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I614 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I615 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I616 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I617 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I618 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I619 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I620 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I621 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I622 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I623 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I624 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I625 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I626 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I627 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I628 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I629 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I630 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I631 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I632 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I633 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I634 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I635 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I636 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I637 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I638 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I639 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I640 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I641 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I642 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I643 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I644 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I645 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I646 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I647 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I648 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I649 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I650 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I651 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I652 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I653 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I654 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I655 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I656 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I657 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I658 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I659 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I660 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I661 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I662 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I663 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I664 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I665 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I666 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I667 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I668 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I669 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I670 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I671 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I672 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I673 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I674 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I675 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I676 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I677 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I678 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I679 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  AND2 I680 (rd_3r1[0:0], dt_0[0:0], rg_3r);
  AND2 I681 (rd_3r1[1:1], dt_0[1:1], rg_3r);
  AND2 I682 (rd_3r1[2:2], dt_0[2:2], rg_3r);
  AND2 I683 (rd_3r1[3:3], dt_0[3:3], rg_3r);
  AND2 I684 (rd_3r1[4:4], dt_0[4:4], rg_3r);
  AND2 I685 (rd_3r1[5:5], dt_0[5:5], rg_3r);
  AND2 I686 (rd_3r1[6:6], dt_0[6:6], rg_3r);
  AND2 I687 (rd_3r1[7:7], dt_0[7:7], rg_3r);
  AND2 I688 (rd_3r1[8:8], dt_0[8:8], rg_3r);
  AND2 I689 (rd_3r1[9:9], dt_0[9:9], rg_3r);
  AND2 I690 (rd_3r1[10:10], dt_0[10:10], rg_3r);
  AND2 I691 (rd_3r1[11:11], dt_0[11:11], rg_3r);
  AND2 I692 (rd_3r1[12:12], dt_0[12:12], rg_3r);
  AND2 I693 (rd_3r1[13:13], dt_0[13:13], rg_3r);
  AND2 I694 (rd_3r1[14:14], dt_0[14:14], rg_3r);
  AND2 I695 (rd_3r1[15:15], dt_0[15:15], rg_3r);
  AND2 I696 (rd_3r1[16:16], dt_0[16:16], rg_3r);
  AND2 I697 (rd_3r1[17:17], dt_0[17:17], rg_3r);
  AND2 I698 (rd_3r1[18:18], dt_0[18:18], rg_3r);
  AND2 I699 (rd_3r1[19:19], dt_0[19:19], rg_3r);
  AND2 I700 (rd_3r1[20:20], dt_0[20:20], rg_3r);
  AND2 I701 (rd_3r1[21:21], dt_0[21:21], rg_3r);
  AND2 I702 (rd_3r1[22:22], dt_0[22:22], rg_3r);
  AND2 I703 (rd_3r1[23:23], dt_0[23:23], rg_3r);
  AND2 I704 (rd_3r1[24:24], dt_0[24:24], rg_3r);
  AND2 I705 (rd_3r1[25:25], dt_0[25:25], rg_3r);
  AND2 I706 (rd_3r1[26:26], dt_0[26:26], rg_3r);
  AND2 I707 (rd_3r1[27:27], dt_0[27:27], rg_3r);
  AND2 I708 (rd_3r1[28:28], dt_0[28:28], rg_3r);
  AND2 I709 (rd_3r1[29:29], dt_0[29:29], rg_3r);
  AND2 I710 (rd_3r1[30:30], dt_0[30:30], rg_3r);
  AND2 I711 (rd_3r1[31:31], dt_0[31:31], rg_3r);
  AND2 I712 (rd_4r1[0:0], dt_0[0:0], rg_4r);
  AND2 I713 (rd_4r1[1:1], dt_0[1:1], rg_4r);
  AND2 I714 (rd_4r1[2:2], dt_0[2:2], rg_4r);
  AND2 I715 (rd_4r1[3:3], dt_0[3:3], rg_4r);
  AND2 I716 (rd_4r1[4:4], dt_0[4:4], rg_4r);
  AND2 I717 (rd_4r1[5:5], dt_0[5:5], rg_4r);
  AND2 I718 (rd_4r1[6:6], dt_0[6:6], rg_4r);
  AND2 I719 (rd_4r1[7:7], dt_0[7:7], rg_4r);
  AND2 I720 (rd_4r1[8:8], dt_0[8:8], rg_4r);
  AND2 I721 (rd_4r1[9:9], dt_0[9:9], rg_4r);
  AND2 I722 (rd_4r1[10:10], dt_0[10:10], rg_4r);
  AND2 I723 (rd_4r1[11:11], dt_0[11:11], rg_4r);
  AND2 I724 (rd_4r1[12:12], dt_0[12:12], rg_4r);
  AND2 I725 (rd_4r1[13:13], dt_0[13:13], rg_4r);
  AND2 I726 (rd_4r1[14:14], dt_0[14:14], rg_4r);
  AND2 I727 (rd_4r1[15:15], dt_0[15:15], rg_4r);
  AND2 I728 (rd_4r1[16:16], dt_0[16:16], rg_4r);
  AND2 I729 (rd_4r1[17:17], dt_0[17:17], rg_4r);
  AND2 I730 (rd_4r1[18:18], dt_0[18:18], rg_4r);
  AND2 I731 (rd_4r1[19:19], dt_0[19:19], rg_4r);
  AND2 I732 (rd_4r1[20:20], dt_0[20:20], rg_4r);
  AND2 I733 (rd_4r1[21:21], dt_0[21:21], rg_4r);
  AND2 I734 (rd_4r1[22:22], dt_0[22:22], rg_4r);
  AND2 I735 (rd_4r1[23:23], dt_0[23:23], rg_4r);
  AND2 I736 (rd_4r1[24:24], dt_0[24:24], rg_4r);
  AND2 I737 (rd_4r1[25:25], dt_0[25:25], rg_4r);
  AND2 I738 (rd_4r1[26:26], dt_0[26:26], rg_4r);
  AND2 I739 (rd_4r1[27:27], dt_0[27:27], rg_4r);
  AND2 I740 (rd_4r1[28:28], dt_0[28:28], rg_4r);
  AND2 I741 (rd_4r1[29:29], dt_0[29:29], rg_4r);
  AND2 I742 (rd_4r1[30:30], dt_0[30:30], rg_4r);
  AND2 I743 (rd_4r1[31:31], dt_0[31:31], rg_4r);
  NOR3 I744 (simp7281_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I745 (simp7281_0[1:1], rg_3r, rg_4r, rg_0a);
  NOR3 I746 (simp7281_0[2:2], rg_1a, rg_2a, rg_3a);
  INV I747 (simp7281_0[3:3], rg_4a);
  NAND3 I748 (simp7282_0[0:0], simp7281_0[0:0], simp7281_0[1:1], simp7281_0[2:2]);
  INV I749 (simp7282_0[1:1], simp7281_0[3:3]);
  OR2 I750 (anyread_0, simp7282_0[0:0], simp7282_0[1:1]);
  BUFF I751 (wg_0a, wd_0a);
  BUFF I752 (rg_0a, rd_0a);
  BUFF I753 (rg_1a, rd_1a);
  BUFF I754 (rg_2a, rd_2a);
  BUFF I755 (rg_3a, rd_3a);
  BUFF I756 (rg_4a, rd_4a);
endmodule

// tkf5mo0w0_o0w5 TeakF [0,0] [One 5,Many [0,5]]
module tkf5mo0w0_o0w5 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [4:0] i_0r0;
  input [4:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [4:0] o_1r0;
  output [4:0] o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_1r0[0:0], i_0r0[0:0]);
  BUFF I3 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I4 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I5 (o_1r0[3:3], i_0r0[3:3]);
  BUFF I6 (o_1r0[4:4], i_0r0[4:4]);
  BUFF I7 (o_1r1[0:0], i_0r1[0:0]);
  BUFF I8 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I9 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I10 (o_1r1[3:3], i_0r1[3:3]);
  BUFF I11 (o_1r1[4:4], i_0r1[4:4]);
  BUFF I12 (o_0r, icomplete_0);
  C3 I13 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tkf2mo0w0_o0w2 TeakF [0,0] [One 2,Many [0,2]]
module tkf2mo0w0_o0w2 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [1:0] o_1r0;
  output [1:0] o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_1r0[0:0], i_0r0[0:0]);
  BUFF I3 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I4 (o_1r1[0:0], i_0r1[0:0]);
  BUFF I5 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I6 (o_0r, icomplete_0);
  C3 I7 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tkm3x2b TeakM [Many [2,2,2],One 2]
module tkm3x2b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, o_0r0, o_0r1, o_0a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  input [1:0] i_1r0;
  input [1:0] i_1r1;
  output i_1a;
  input [1:0] i_2r0;
  input [1:0] i_2r1;
  output i_2a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  wire [1:0] gfint_0;
  wire [1:0] gfint_1;
  wire [1:0] gfint_2;
  wire [1:0] gtint_0;
  wire [1:0] gtint_1;
  wire [1:0] gtint_2;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire nchosen_0;
  wire [1:0] comp0_0;
  wire [1:0] comp1_0;
  wire [1:0] comp2_0;
  OR3 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  OR3 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  OR3 I2 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  OR3 I3 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  AND2 I4 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I5 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I6 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I7 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I8 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I9 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I10 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I11 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I12 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I13 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I14 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I15 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  OR2 I16 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I17 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  C2 I18 (icomp_0, comp0_0[0:0], comp0_0[1:1]);
  OR2 I19 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I20 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  C2 I21 (icomp_1, comp1_0[0:0], comp1_0[1:1]);
  OR2 I22 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I23 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  C2 I24 (icomp_2, comp2_0[0:0], comp2_0[1:1]);
  C2R I25 (choice_0, icomp_0, nchosen_0, reset);
  C2R I26 (choice_1, icomp_1, nchosen_0, reset);
  C2R I27 (choice_2, icomp_2, nchosen_0, reset);
  OR3 I28 (anychoice_0, choice_0, choice_1, choice_2);
  NOR2 I29 (nchosen_0, anychoice_0, o_0a);
  C2R I30 (i_0a, choice_0, o_0a, reset);
  C2R I31 (i_1a, choice_1, o_0a, reset);
  C2R I32 (i_2a, choice_2, o_0a, reset);
endmodule

// tkm4x1b TeakM [Many [1,1,1,1],One 1]
module tkm4x1b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input i_1r0;
  input i_1r1;
  output i_1a;
  input i_2r0;
  input i_2r1;
  output i_2a;
  input i_3r0;
  input i_3r1;
  output i_3a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire gfint_0;
  wire gfint_1;
  wire gfint_2;
  wire gfint_3;
  wire gtint_0;
  wire gtint_1;
  wire gtint_2;
  wire gtint_3;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire icomp_3;
  wire nchosen_0;
  wire [1:0] simp181_0;
  wire [1:0] simp191_0;
  wire comp0_0;
  wire comp1_0;
  wire comp2_0;
  wire comp3_0;
  wire [1:0] simp441_0;
  NOR3 I0 (simp181_0[0:0], gfint_0, gfint_1, gfint_2);
  INV I1 (simp181_0[1:1], gfint_3);
  NAND2 I2 (o_0r0, simp181_0[0:0], simp181_0[1:1]);
  NOR3 I3 (simp191_0[0:0], gtint_0, gtint_1, gtint_2);
  INV I4 (simp191_0[1:1], gtint_3);
  NAND2 I5 (o_0r1, simp191_0[0:0], simp191_0[1:1]);
  AND2 I6 (gtint_0, choice_0, i_0r1);
  AND2 I7 (gtint_1, choice_1, i_1r1);
  AND2 I8 (gtint_2, choice_2, i_2r1);
  AND2 I9 (gtint_3, choice_3, i_3r1);
  AND2 I10 (gfint_0, choice_0, i_0r0);
  AND2 I11 (gfint_1, choice_1, i_1r0);
  AND2 I12 (gfint_2, choice_2, i_2r0);
  AND2 I13 (gfint_3, choice_3, i_3r0);
  OR2 I14 (comp0_0, i_0r0, i_0r1);
  BUFF I15 (icomp_0, comp0_0);
  OR2 I16 (comp1_0, i_1r0, i_1r1);
  BUFF I17 (icomp_1, comp1_0);
  OR2 I18 (comp2_0, i_2r0, i_2r1);
  BUFF I19 (icomp_2, comp2_0);
  OR2 I20 (comp3_0, i_3r0, i_3r1);
  BUFF I21 (icomp_3, comp3_0);
  C2R I22 (choice_0, icomp_0, nchosen_0, reset);
  C2R I23 (choice_1, icomp_1, nchosen_0, reset);
  C2R I24 (choice_2, icomp_2, nchosen_0, reset);
  C2R I25 (choice_3, icomp_3, nchosen_0, reset);
  NOR3 I26 (simp441_0[0:0], choice_0, choice_1, choice_2);
  INV I27 (simp441_0[1:1], choice_3);
  NAND2 I28 (anychoice_0, simp441_0[0:0], simp441_0[1:1]);
  NOR2 I29 (nchosen_0, anychoice_0, o_0a);
  C2R I30 (i_0a, choice_0, o_0a, reset);
  C2R I31 (i_1a, choice_1, o_0a, reset);
  C2R I32 (i_2a, choice_2, o_0a, reset);
  C2R I33 (i_3a, choice_3, o_0a, reset);
endmodule

// tkm2x32b TeakM [Many [32,32],One 32]
module tkm2x32b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire [31:0] gfint_0;
  wire [31:0] gfint_1;
  wire [31:0] gtint_0;
  wire [31:0] gtint_1;
  wire choice_0;
  wire choice_1;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire nchosen_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2351_0;
  wire [3:0] simp2352_0;
  wire [1:0] simp2353_0;
  wire [31:0] comp1_0;
  wire [10:0] simp2691_0;
  wire [3:0] simp2692_0;
  wire [1:0] simp2693_0;
  OR2 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0]);
  OR2 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1]);
  OR2 I2 (o_0r0[2:2], gfint_0[2:2], gfint_1[2:2]);
  OR2 I3 (o_0r0[3:3], gfint_0[3:3], gfint_1[3:3]);
  OR2 I4 (o_0r0[4:4], gfint_0[4:4], gfint_1[4:4]);
  OR2 I5 (o_0r0[5:5], gfint_0[5:5], gfint_1[5:5]);
  OR2 I6 (o_0r0[6:6], gfint_0[6:6], gfint_1[6:6]);
  OR2 I7 (o_0r0[7:7], gfint_0[7:7], gfint_1[7:7]);
  OR2 I8 (o_0r0[8:8], gfint_0[8:8], gfint_1[8:8]);
  OR2 I9 (o_0r0[9:9], gfint_0[9:9], gfint_1[9:9]);
  OR2 I10 (o_0r0[10:10], gfint_0[10:10], gfint_1[10:10]);
  OR2 I11 (o_0r0[11:11], gfint_0[11:11], gfint_1[11:11]);
  OR2 I12 (o_0r0[12:12], gfint_0[12:12], gfint_1[12:12]);
  OR2 I13 (o_0r0[13:13], gfint_0[13:13], gfint_1[13:13]);
  OR2 I14 (o_0r0[14:14], gfint_0[14:14], gfint_1[14:14]);
  OR2 I15 (o_0r0[15:15], gfint_0[15:15], gfint_1[15:15]);
  OR2 I16 (o_0r0[16:16], gfint_0[16:16], gfint_1[16:16]);
  OR2 I17 (o_0r0[17:17], gfint_0[17:17], gfint_1[17:17]);
  OR2 I18 (o_0r0[18:18], gfint_0[18:18], gfint_1[18:18]);
  OR2 I19 (o_0r0[19:19], gfint_0[19:19], gfint_1[19:19]);
  OR2 I20 (o_0r0[20:20], gfint_0[20:20], gfint_1[20:20]);
  OR2 I21 (o_0r0[21:21], gfint_0[21:21], gfint_1[21:21]);
  OR2 I22 (o_0r0[22:22], gfint_0[22:22], gfint_1[22:22]);
  OR2 I23 (o_0r0[23:23], gfint_0[23:23], gfint_1[23:23]);
  OR2 I24 (o_0r0[24:24], gfint_0[24:24], gfint_1[24:24]);
  OR2 I25 (o_0r0[25:25], gfint_0[25:25], gfint_1[25:25]);
  OR2 I26 (o_0r0[26:26], gfint_0[26:26], gfint_1[26:26]);
  OR2 I27 (o_0r0[27:27], gfint_0[27:27], gfint_1[27:27]);
  OR2 I28 (o_0r0[28:28], gfint_0[28:28], gfint_1[28:28]);
  OR2 I29 (o_0r0[29:29], gfint_0[29:29], gfint_1[29:29]);
  OR2 I30 (o_0r0[30:30], gfint_0[30:30], gfint_1[30:30]);
  OR2 I31 (o_0r0[31:31], gfint_0[31:31], gfint_1[31:31]);
  OR2 I32 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0]);
  OR2 I33 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1]);
  OR2 I34 (o_0r1[2:2], gtint_0[2:2], gtint_1[2:2]);
  OR2 I35 (o_0r1[3:3], gtint_0[3:3], gtint_1[3:3]);
  OR2 I36 (o_0r1[4:4], gtint_0[4:4], gtint_1[4:4]);
  OR2 I37 (o_0r1[5:5], gtint_0[5:5], gtint_1[5:5]);
  OR2 I38 (o_0r1[6:6], gtint_0[6:6], gtint_1[6:6]);
  OR2 I39 (o_0r1[7:7], gtint_0[7:7], gtint_1[7:7]);
  OR2 I40 (o_0r1[8:8], gtint_0[8:8], gtint_1[8:8]);
  OR2 I41 (o_0r1[9:9], gtint_0[9:9], gtint_1[9:9]);
  OR2 I42 (o_0r1[10:10], gtint_0[10:10], gtint_1[10:10]);
  OR2 I43 (o_0r1[11:11], gtint_0[11:11], gtint_1[11:11]);
  OR2 I44 (o_0r1[12:12], gtint_0[12:12], gtint_1[12:12]);
  OR2 I45 (o_0r1[13:13], gtint_0[13:13], gtint_1[13:13]);
  OR2 I46 (o_0r1[14:14], gtint_0[14:14], gtint_1[14:14]);
  OR2 I47 (o_0r1[15:15], gtint_0[15:15], gtint_1[15:15]);
  OR2 I48 (o_0r1[16:16], gtint_0[16:16], gtint_1[16:16]);
  OR2 I49 (o_0r1[17:17], gtint_0[17:17], gtint_1[17:17]);
  OR2 I50 (o_0r1[18:18], gtint_0[18:18], gtint_1[18:18]);
  OR2 I51 (o_0r1[19:19], gtint_0[19:19], gtint_1[19:19]);
  OR2 I52 (o_0r1[20:20], gtint_0[20:20], gtint_1[20:20]);
  OR2 I53 (o_0r1[21:21], gtint_0[21:21], gtint_1[21:21]);
  OR2 I54 (o_0r1[22:22], gtint_0[22:22], gtint_1[22:22]);
  OR2 I55 (o_0r1[23:23], gtint_0[23:23], gtint_1[23:23]);
  OR2 I56 (o_0r1[24:24], gtint_0[24:24], gtint_1[24:24]);
  OR2 I57 (o_0r1[25:25], gtint_0[25:25], gtint_1[25:25]);
  OR2 I58 (o_0r1[26:26], gtint_0[26:26], gtint_1[26:26]);
  OR2 I59 (o_0r1[27:27], gtint_0[27:27], gtint_1[27:27]);
  OR2 I60 (o_0r1[28:28], gtint_0[28:28], gtint_1[28:28]);
  OR2 I61 (o_0r1[29:29], gtint_0[29:29], gtint_1[29:29]);
  OR2 I62 (o_0r1[30:30], gtint_0[30:30], gtint_1[30:30]);
  OR2 I63 (o_0r1[31:31], gtint_0[31:31], gtint_1[31:31]);
  AND2 I64 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I65 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I66 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I67 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I68 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I69 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I70 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I71 (gtint_0[7:7], choice_0, i_0r1[7:7]);
  AND2 I72 (gtint_0[8:8], choice_0, i_0r1[8:8]);
  AND2 I73 (gtint_0[9:9], choice_0, i_0r1[9:9]);
  AND2 I74 (gtint_0[10:10], choice_0, i_0r1[10:10]);
  AND2 I75 (gtint_0[11:11], choice_0, i_0r1[11:11]);
  AND2 I76 (gtint_0[12:12], choice_0, i_0r1[12:12]);
  AND2 I77 (gtint_0[13:13], choice_0, i_0r1[13:13]);
  AND2 I78 (gtint_0[14:14], choice_0, i_0r1[14:14]);
  AND2 I79 (gtint_0[15:15], choice_0, i_0r1[15:15]);
  AND2 I80 (gtint_0[16:16], choice_0, i_0r1[16:16]);
  AND2 I81 (gtint_0[17:17], choice_0, i_0r1[17:17]);
  AND2 I82 (gtint_0[18:18], choice_0, i_0r1[18:18]);
  AND2 I83 (gtint_0[19:19], choice_0, i_0r1[19:19]);
  AND2 I84 (gtint_0[20:20], choice_0, i_0r1[20:20]);
  AND2 I85 (gtint_0[21:21], choice_0, i_0r1[21:21]);
  AND2 I86 (gtint_0[22:22], choice_0, i_0r1[22:22]);
  AND2 I87 (gtint_0[23:23], choice_0, i_0r1[23:23]);
  AND2 I88 (gtint_0[24:24], choice_0, i_0r1[24:24]);
  AND2 I89 (gtint_0[25:25], choice_0, i_0r1[25:25]);
  AND2 I90 (gtint_0[26:26], choice_0, i_0r1[26:26]);
  AND2 I91 (gtint_0[27:27], choice_0, i_0r1[27:27]);
  AND2 I92 (gtint_0[28:28], choice_0, i_0r1[28:28]);
  AND2 I93 (gtint_0[29:29], choice_0, i_0r1[29:29]);
  AND2 I94 (gtint_0[30:30], choice_0, i_0r1[30:30]);
  AND2 I95 (gtint_0[31:31], choice_0, i_0r1[31:31]);
  AND2 I96 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I97 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I98 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I99 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I100 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I101 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I102 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I103 (gtint_1[7:7], choice_1, i_1r1[7:7]);
  AND2 I104 (gtint_1[8:8], choice_1, i_1r1[8:8]);
  AND2 I105 (gtint_1[9:9], choice_1, i_1r1[9:9]);
  AND2 I106 (gtint_1[10:10], choice_1, i_1r1[10:10]);
  AND2 I107 (gtint_1[11:11], choice_1, i_1r1[11:11]);
  AND2 I108 (gtint_1[12:12], choice_1, i_1r1[12:12]);
  AND2 I109 (gtint_1[13:13], choice_1, i_1r1[13:13]);
  AND2 I110 (gtint_1[14:14], choice_1, i_1r1[14:14]);
  AND2 I111 (gtint_1[15:15], choice_1, i_1r1[15:15]);
  AND2 I112 (gtint_1[16:16], choice_1, i_1r1[16:16]);
  AND2 I113 (gtint_1[17:17], choice_1, i_1r1[17:17]);
  AND2 I114 (gtint_1[18:18], choice_1, i_1r1[18:18]);
  AND2 I115 (gtint_1[19:19], choice_1, i_1r1[19:19]);
  AND2 I116 (gtint_1[20:20], choice_1, i_1r1[20:20]);
  AND2 I117 (gtint_1[21:21], choice_1, i_1r1[21:21]);
  AND2 I118 (gtint_1[22:22], choice_1, i_1r1[22:22]);
  AND2 I119 (gtint_1[23:23], choice_1, i_1r1[23:23]);
  AND2 I120 (gtint_1[24:24], choice_1, i_1r1[24:24]);
  AND2 I121 (gtint_1[25:25], choice_1, i_1r1[25:25]);
  AND2 I122 (gtint_1[26:26], choice_1, i_1r1[26:26]);
  AND2 I123 (gtint_1[27:27], choice_1, i_1r1[27:27]);
  AND2 I124 (gtint_1[28:28], choice_1, i_1r1[28:28]);
  AND2 I125 (gtint_1[29:29], choice_1, i_1r1[29:29]);
  AND2 I126 (gtint_1[30:30], choice_1, i_1r1[30:30]);
  AND2 I127 (gtint_1[31:31], choice_1, i_1r1[31:31]);
  AND2 I128 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I129 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I130 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I131 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I132 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I133 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I134 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I135 (gfint_0[7:7], choice_0, i_0r0[7:7]);
  AND2 I136 (gfint_0[8:8], choice_0, i_0r0[8:8]);
  AND2 I137 (gfint_0[9:9], choice_0, i_0r0[9:9]);
  AND2 I138 (gfint_0[10:10], choice_0, i_0r0[10:10]);
  AND2 I139 (gfint_0[11:11], choice_0, i_0r0[11:11]);
  AND2 I140 (gfint_0[12:12], choice_0, i_0r0[12:12]);
  AND2 I141 (gfint_0[13:13], choice_0, i_0r0[13:13]);
  AND2 I142 (gfint_0[14:14], choice_0, i_0r0[14:14]);
  AND2 I143 (gfint_0[15:15], choice_0, i_0r0[15:15]);
  AND2 I144 (gfint_0[16:16], choice_0, i_0r0[16:16]);
  AND2 I145 (gfint_0[17:17], choice_0, i_0r0[17:17]);
  AND2 I146 (gfint_0[18:18], choice_0, i_0r0[18:18]);
  AND2 I147 (gfint_0[19:19], choice_0, i_0r0[19:19]);
  AND2 I148 (gfint_0[20:20], choice_0, i_0r0[20:20]);
  AND2 I149 (gfint_0[21:21], choice_0, i_0r0[21:21]);
  AND2 I150 (gfint_0[22:22], choice_0, i_0r0[22:22]);
  AND2 I151 (gfint_0[23:23], choice_0, i_0r0[23:23]);
  AND2 I152 (gfint_0[24:24], choice_0, i_0r0[24:24]);
  AND2 I153 (gfint_0[25:25], choice_0, i_0r0[25:25]);
  AND2 I154 (gfint_0[26:26], choice_0, i_0r0[26:26]);
  AND2 I155 (gfint_0[27:27], choice_0, i_0r0[27:27]);
  AND2 I156 (gfint_0[28:28], choice_0, i_0r0[28:28]);
  AND2 I157 (gfint_0[29:29], choice_0, i_0r0[29:29]);
  AND2 I158 (gfint_0[30:30], choice_0, i_0r0[30:30]);
  AND2 I159 (gfint_0[31:31], choice_0, i_0r0[31:31]);
  AND2 I160 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I161 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I162 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I163 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I164 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I165 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I166 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I167 (gfint_1[7:7], choice_1, i_1r0[7:7]);
  AND2 I168 (gfint_1[8:8], choice_1, i_1r0[8:8]);
  AND2 I169 (gfint_1[9:9], choice_1, i_1r0[9:9]);
  AND2 I170 (gfint_1[10:10], choice_1, i_1r0[10:10]);
  AND2 I171 (gfint_1[11:11], choice_1, i_1r0[11:11]);
  AND2 I172 (gfint_1[12:12], choice_1, i_1r0[12:12]);
  AND2 I173 (gfint_1[13:13], choice_1, i_1r0[13:13]);
  AND2 I174 (gfint_1[14:14], choice_1, i_1r0[14:14]);
  AND2 I175 (gfint_1[15:15], choice_1, i_1r0[15:15]);
  AND2 I176 (gfint_1[16:16], choice_1, i_1r0[16:16]);
  AND2 I177 (gfint_1[17:17], choice_1, i_1r0[17:17]);
  AND2 I178 (gfint_1[18:18], choice_1, i_1r0[18:18]);
  AND2 I179 (gfint_1[19:19], choice_1, i_1r0[19:19]);
  AND2 I180 (gfint_1[20:20], choice_1, i_1r0[20:20]);
  AND2 I181 (gfint_1[21:21], choice_1, i_1r0[21:21]);
  AND2 I182 (gfint_1[22:22], choice_1, i_1r0[22:22]);
  AND2 I183 (gfint_1[23:23], choice_1, i_1r0[23:23]);
  AND2 I184 (gfint_1[24:24], choice_1, i_1r0[24:24]);
  AND2 I185 (gfint_1[25:25], choice_1, i_1r0[25:25]);
  AND2 I186 (gfint_1[26:26], choice_1, i_1r0[26:26]);
  AND2 I187 (gfint_1[27:27], choice_1, i_1r0[27:27]);
  AND2 I188 (gfint_1[28:28], choice_1, i_1r0[28:28]);
  AND2 I189 (gfint_1[29:29], choice_1, i_1r0[29:29]);
  AND2 I190 (gfint_1[30:30], choice_1, i_1r0[30:30]);
  AND2 I191 (gfint_1[31:31], choice_1, i_1r0[31:31]);
  OR2 I192 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I193 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I194 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I195 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I196 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I197 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I198 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I199 (comp0_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I200 (comp0_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I201 (comp0_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I202 (comp0_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I203 (comp0_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I204 (comp0_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I205 (comp0_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I206 (comp0_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I207 (comp0_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I208 (comp0_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I209 (comp0_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I210 (comp0_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I211 (comp0_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I212 (comp0_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I213 (comp0_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I214 (comp0_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I215 (comp0_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I216 (comp0_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I217 (comp0_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I218 (comp0_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I219 (comp0_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I220 (comp0_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I221 (comp0_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I222 (comp0_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I223 (comp0_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  C3 I224 (simp2351_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I225 (simp2351_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I226 (simp2351_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I227 (simp2351_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I228 (simp2351_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I229 (simp2351_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I230 (simp2351_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I231 (simp2351_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I232 (simp2351_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I233 (simp2351_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I234 (simp2351_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I235 (simp2352_0[0:0], simp2351_0[0:0], simp2351_0[1:1], simp2351_0[2:2]);
  C3 I236 (simp2352_0[1:1], simp2351_0[3:3], simp2351_0[4:4], simp2351_0[5:5]);
  C3 I237 (simp2352_0[2:2], simp2351_0[6:6], simp2351_0[7:7], simp2351_0[8:8]);
  C2 I238 (simp2352_0[3:3], simp2351_0[9:9], simp2351_0[10:10]);
  C3 I239 (simp2353_0[0:0], simp2352_0[0:0], simp2352_0[1:1], simp2352_0[2:2]);
  BUFF I240 (simp2353_0[1:1], simp2352_0[3:3]);
  C2 I241 (icomp_0, simp2353_0[0:0], simp2353_0[1:1]);
  OR2 I242 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I243 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I244 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I245 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I246 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I247 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I248 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  OR2 I249 (comp1_0[7:7], i_1r0[7:7], i_1r1[7:7]);
  OR2 I250 (comp1_0[8:8], i_1r0[8:8], i_1r1[8:8]);
  OR2 I251 (comp1_0[9:9], i_1r0[9:9], i_1r1[9:9]);
  OR2 I252 (comp1_0[10:10], i_1r0[10:10], i_1r1[10:10]);
  OR2 I253 (comp1_0[11:11], i_1r0[11:11], i_1r1[11:11]);
  OR2 I254 (comp1_0[12:12], i_1r0[12:12], i_1r1[12:12]);
  OR2 I255 (comp1_0[13:13], i_1r0[13:13], i_1r1[13:13]);
  OR2 I256 (comp1_0[14:14], i_1r0[14:14], i_1r1[14:14]);
  OR2 I257 (comp1_0[15:15], i_1r0[15:15], i_1r1[15:15]);
  OR2 I258 (comp1_0[16:16], i_1r0[16:16], i_1r1[16:16]);
  OR2 I259 (comp1_0[17:17], i_1r0[17:17], i_1r1[17:17]);
  OR2 I260 (comp1_0[18:18], i_1r0[18:18], i_1r1[18:18]);
  OR2 I261 (comp1_0[19:19], i_1r0[19:19], i_1r1[19:19]);
  OR2 I262 (comp1_0[20:20], i_1r0[20:20], i_1r1[20:20]);
  OR2 I263 (comp1_0[21:21], i_1r0[21:21], i_1r1[21:21]);
  OR2 I264 (comp1_0[22:22], i_1r0[22:22], i_1r1[22:22]);
  OR2 I265 (comp1_0[23:23], i_1r0[23:23], i_1r1[23:23]);
  OR2 I266 (comp1_0[24:24], i_1r0[24:24], i_1r1[24:24]);
  OR2 I267 (comp1_0[25:25], i_1r0[25:25], i_1r1[25:25]);
  OR2 I268 (comp1_0[26:26], i_1r0[26:26], i_1r1[26:26]);
  OR2 I269 (comp1_0[27:27], i_1r0[27:27], i_1r1[27:27]);
  OR2 I270 (comp1_0[28:28], i_1r0[28:28], i_1r1[28:28]);
  OR2 I271 (comp1_0[29:29], i_1r0[29:29], i_1r1[29:29]);
  OR2 I272 (comp1_0[30:30], i_1r0[30:30], i_1r1[30:30]);
  OR2 I273 (comp1_0[31:31], i_1r0[31:31], i_1r1[31:31]);
  C3 I274 (simp2691_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I275 (simp2691_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  C3 I276 (simp2691_0[2:2], comp1_0[6:6], comp1_0[7:7], comp1_0[8:8]);
  C3 I277 (simp2691_0[3:3], comp1_0[9:9], comp1_0[10:10], comp1_0[11:11]);
  C3 I278 (simp2691_0[4:4], comp1_0[12:12], comp1_0[13:13], comp1_0[14:14]);
  C3 I279 (simp2691_0[5:5], comp1_0[15:15], comp1_0[16:16], comp1_0[17:17]);
  C3 I280 (simp2691_0[6:6], comp1_0[18:18], comp1_0[19:19], comp1_0[20:20]);
  C3 I281 (simp2691_0[7:7], comp1_0[21:21], comp1_0[22:22], comp1_0[23:23]);
  C3 I282 (simp2691_0[8:8], comp1_0[24:24], comp1_0[25:25], comp1_0[26:26]);
  C3 I283 (simp2691_0[9:9], comp1_0[27:27], comp1_0[28:28], comp1_0[29:29]);
  C2 I284 (simp2691_0[10:10], comp1_0[30:30], comp1_0[31:31]);
  C3 I285 (simp2692_0[0:0], simp2691_0[0:0], simp2691_0[1:1], simp2691_0[2:2]);
  C3 I286 (simp2692_0[1:1], simp2691_0[3:3], simp2691_0[4:4], simp2691_0[5:5]);
  C3 I287 (simp2692_0[2:2], simp2691_0[6:6], simp2691_0[7:7], simp2691_0[8:8]);
  C2 I288 (simp2692_0[3:3], simp2691_0[9:9], simp2691_0[10:10]);
  C3 I289 (simp2693_0[0:0], simp2692_0[0:0], simp2692_0[1:1], simp2692_0[2:2]);
  BUFF I290 (simp2693_0[1:1], simp2692_0[3:3]);
  C2 I291 (icomp_1, simp2693_0[0:0], simp2693_0[1:1]);
  C2R I292 (choice_0, icomp_0, nchosen_0, reset);
  C2R I293 (choice_1, icomp_1, nchosen_0, reset);
  OR2 I294 (anychoice_0, choice_0, choice_1);
  NOR2 I295 (nchosen_0, anychoice_0, o_0a);
  C2R I296 (i_0a, choice_0, o_0a, reset);
  C2R I297 (i_1a, choice_1, o_0a, reset);
endmodule

// tkj7m7_0 TeakJ [Many [7,0],One 7]
module tkj7m7_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [6:0] i_0r0;
  input [6:0] i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  output [6:0] o_0r0;
  output [6:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [6:0] joinf_0;
  wire [6:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joint_0[0:0], i_0r1[0:0]);
  BUFF I8 (joint_0[1:1], i_0r1[1:1]);
  BUFF I9 (joint_0[2:2], i_0r1[2:2]);
  BUFF I10 (joint_0[3:3], i_0r1[3:3]);
  BUFF I11 (joint_0[4:4], i_0r1[4:4]);
  BUFF I12 (joint_0[5:5], i_0r1[5:5]);
  BUFF I13 (joint_0[6:6], i_0r1[6:6]);
  BUFF I14 (icomplete_0, i_1r);
  C2 I15 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I16 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I17 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I18 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I19 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I20 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I21 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I22 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I23 (o_0r1[1:1], joint_0[1:1]);
  BUFF I24 (o_0r1[2:2], joint_0[2:2]);
  BUFF I25 (o_0r1[3:3], joint_0[3:3]);
  BUFF I26 (o_0r1[4:4], joint_0[4:4]);
  BUFF I27 (o_0r1[5:5], joint_0[5:5]);
  BUFF I28 (o_0r1[6:6], joint_0[6:6]);
  BUFF I29 (i_0a, o_0a);
  BUFF I30 (i_1a, o_0a);
endmodule

// tks3_o0w3_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0 TeakS (0+:3) [([Imp 1 0],0),([Imp 2 0],0),([Imp 
//   3 0],0),([Imp 4 0],0),([Imp 5 0],0),([Imp 6 0],0),([Imp 7 0],0)] [One 3,Many [0,0,0,0,0,0,0]]
module tks3_o0w3_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, o_5r, o_5a, o_6r, o_6a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire sel_4;
  wire sel_5;
  wire sel_6;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire gsel_4;
  wire gsel_5;
  wire gsel_6;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire match2_0;
  wire match3_0;
  wire match4_0;
  wire match5_0;
  wire match6_0;
  wire [2:0] comp_0;
  wire [2:0] simp561_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (match0_0, i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I2 (sel_1, match1_0);
  C3 I3 (match1_0, i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I4 (sel_2, match2_0);
  C3 I5 (match2_0, i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I6 (sel_3, match3_0);
  C3 I7 (match3_0, i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I8 (sel_4, match4_0);
  C3 I9 (match4_0, i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I10 (sel_5, match5_0);
  C3 I11 (match5_0, i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I12 (sel_6, match6_0);
  C3 I13 (match6_0, i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  C2 I14 (gsel_0, sel_0, icomplete_0);
  C2 I15 (gsel_1, sel_1, icomplete_0);
  C2 I16 (gsel_2, sel_2, icomplete_0);
  C2 I17 (gsel_3, sel_3, icomplete_0);
  C2 I18 (gsel_4, sel_4, icomplete_0);
  C2 I19 (gsel_5, sel_5, icomplete_0);
  C2 I20 (gsel_6, sel_6, icomplete_0);
  OR2 I21 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I22 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I23 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I24 (icomplete_0, comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  BUFF I25 (o_0r, gsel_0);
  BUFF I26 (o_1r, gsel_1);
  BUFF I27 (o_2r, gsel_2);
  BUFF I28 (o_3r, gsel_3);
  BUFF I29 (o_4r, gsel_4);
  BUFF I30 (o_5r, gsel_5);
  BUFF I31 (o_6r, gsel_6);
  NOR3 I32 (simp561_0[0:0], o_0a, o_1a, o_2a);
  NOR3 I33 (simp561_0[1:1], o_3a, o_4a, o_5a);
  INV I34 (simp561_0[2:2], o_6a);
  NAND3 I35 (oack_0, simp561_0[0:0], simp561_0[1:1], simp561_0[2:2]);
  C2 I36 (i_0a, oack_0, icomplete_0);
endmodule

// tkm7x32b TeakM [Many [32,32,32,32,32,32,32],One 32]
module tkm7x32b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, i_4r0, i_4r1, i_4a, i_5r0, i_5r1, i_5a, i_6r0, i_6r1, i_6a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  input [31:0] i_2r0;
  input [31:0] i_2r1;
  output i_2a;
  input [31:0] i_3r0;
  input [31:0] i_3r1;
  output i_3a;
  input [31:0] i_4r0;
  input [31:0] i_4r1;
  output i_4a;
  input [31:0] i_5r0;
  input [31:0] i_5r1;
  output i_5a;
  input [31:0] i_6r0;
  input [31:0] i_6r1;
  output i_6a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire [31:0] gfint_0;
  wire [31:0] gfint_1;
  wire [31:0] gfint_2;
  wire [31:0] gfint_3;
  wire [31:0] gfint_4;
  wire [31:0] gfint_5;
  wire [31:0] gfint_6;
  wire [31:0] gtint_0;
  wire [31:0] gtint_1;
  wire [31:0] gtint_2;
  wire [31:0] gtint_3;
  wire [31:0] gtint_4;
  wire [31:0] gtint_5;
  wire [31:0] gtint_6;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire choice_4;
  wire choice_5;
  wire choice_6;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire icomp_3;
  wire icomp_4;
  wire icomp_5;
  wire icomp_6;
  wire nchosen_0;
  wire [2:0] simp301_0;
  wire [2:0] simp311_0;
  wire [2:0] simp321_0;
  wire [2:0] simp331_0;
  wire [2:0] simp341_0;
  wire [2:0] simp351_0;
  wire [2:0] simp361_0;
  wire [2:0] simp371_0;
  wire [2:0] simp381_0;
  wire [2:0] simp391_0;
  wire [2:0] simp401_0;
  wire [2:0] simp411_0;
  wire [2:0] simp421_0;
  wire [2:0] simp431_0;
  wire [2:0] simp441_0;
  wire [2:0] simp451_0;
  wire [2:0] simp461_0;
  wire [2:0] simp471_0;
  wire [2:0] simp481_0;
  wire [2:0] simp491_0;
  wire [2:0] simp501_0;
  wire [2:0] simp511_0;
  wire [2:0] simp521_0;
  wire [2:0] simp531_0;
  wire [2:0] simp541_0;
  wire [2:0] simp551_0;
  wire [2:0] simp561_0;
  wire [2:0] simp571_0;
  wire [2:0] simp581_0;
  wire [2:0] simp591_0;
  wire [2:0] simp601_0;
  wire [2:0] simp611_0;
  wire [2:0] simp621_0;
  wire [2:0] simp631_0;
  wire [2:0] simp641_0;
  wire [2:0] simp651_0;
  wire [2:0] simp661_0;
  wire [2:0] simp671_0;
  wire [2:0] simp681_0;
  wire [2:0] simp691_0;
  wire [2:0] simp701_0;
  wire [2:0] simp711_0;
  wire [2:0] simp721_0;
  wire [2:0] simp731_0;
  wire [2:0] simp741_0;
  wire [2:0] simp751_0;
  wire [2:0] simp761_0;
  wire [2:0] simp771_0;
  wire [2:0] simp781_0;
  wire [2:0] simp791_0;
  wire [2:0] simp801_0;
  wire [2:0] simp811_0;
  wire [2:0] simp821_0;
  wire [2:0] simp831_0;
  wire [2:0] simp841_0;
  wire [2:0] simp851_0;
  wire [2:0] simp861_0;
  wire [2:0] simp871_0;
  wire [2:0] simp881_0;
  wire [2:0] simp891_0;
  wire [2:0] simp901_0;
  wire [2:0] simp911_0;
  wire [2:0] simp921_0;
  wire [2:0] simp931_0;
  wire [31:0] comp0_0;
  wire [10:0] simp5751_0;
  wire [3:0] simp5752_0;
  wire [1:0] simp5753_0;
  wire [31:0] comp1_0;
  wire [10:0] simp6091_0;
  wire [3:0] simp6092_0;
  wire [1:0] simp6093_0;
  wire [31:0] comp2_0;
  wire [10:0] simp6431_0;
  wire [3:0] simp6432_0;
  wire [1:0] simp6433_0;
  wire [31:0] comp3_0;
  wire [10:0] simp6771_0;
  wire [3:0] simp6772_0;
  wire [1:0] simp6773_0;
  wire [31:0] comp4_0;
  wire [10:0] simp7111_0;
  wire [3:0] simp7112_0;
  wire [1:0] simp7113_0;
  wire [31:0] comp5_0;
  wire [10:0] simp7451_0;
  wire [3:0] simp7452_0;
  wire [1:0] simp7453_0;
  wire [31:0] comp6_0;
  wire [10:0] simp7791_0;
  wire [3:0] simp7792_0;
  wire [1:0] simp7793_0;
  wire [2:0] simp7871_0;
  NOR3 I0 (simp301_0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  NOR3 I1 (simp301_0[1:1], gfint_3[0:0], gfint_4[0:0], gfint_5[0:0]);
  INV I2 (simp301_0[2:2], gfint_6[0:0]);
  NAND3 I3 (o_0r0[0:0], simp301_0[0:0], simp301_0[1:1], simp301_0[2:2]);
  NOR3 I4 (simp311_0[0:0], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  NOR3 I5 (simp311_0[1:1], gfint_3[1:1], gfint_4[1:1], gfint_5[1:1]);
  INV I6 (simp311_0[2:2], gfint_6[1:1]);
  NAND3 I7 (o_0r0[1:1], simp311_0[0:0], simp311_0[1:1], simp311_0[2:2]);
  NOR3 I8 (simp321_0[0:0], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  NOR3 I9 (simp321_0[1:1], gfint_3[2:2], gfint_4[2:2], gfint_5[2:2]);
  INV I10 (simp321_0[2:2], gfint_6[2:2]);
  NAND3 I11 (o_0r0[2:2], simp321_0[0:0], simp321_0[1:1], simp321_0[2:2]);
  NOR3 I12 (simp331_0[0:0], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  NOR3 I13 (simp331_0[1:1], gfint_3[3:3], gfint_4[3:3], gfint_5[3:3]);
  INV I14 (simp331_0[2:2], gfint_6[3:3]);
  NAND3 I15 (o_0r0[3:3], simp331_0[0:0], simp331_0[1:1], simp331_0[2:2]);
  NOR3 I16 (simp341_0[0:0], gfint_0[4:4], gfint_1[4:4], gfint_2[4:4]);
  NOR3 I17 (simp341_0[1:1], gfint_3[4:4], gfint_4[4:4], gfint_5[4:4]);
  INV I18 (simp341_0[2:2], gfint_6[4:4]);
  NAND3 I19 (o_0r0[4:4], simp341_0[0:0], simp341_0[1:1], simp341_0[2:2]);
  NOR3 I20 (simp351_0[0:0], gfint_0[5:5], gfint_1[5:5], gfint_2[5:5]);
  NOR3 I21 (simp351_0[1:1], gfint_3[5:5], gfint_4[5:5], gfint_5[5:5]);
  INV I22 (simp351_0[2:2], gfint_6[5:5]);
  NAND3 I23 (o_0r0[5:5], simp351_0[0:0], simp351_0[1:1], simp351_0[2:2]);
  NOR3 I24 (simp361_0[0:0], gfint_0[6:6], gfint_1[6:6], gfint_2[6:6]);
  NOR3 I25 (simp361_0[1:1], gfint_3[6:6], gfint_4[6:6], gfint_5[6:6]);
  INV I26 (simp361_0[2:2], gfint_6[6:6]);
  NAND3 I27 (o_0r0[6:6], simp361_0[0:0], simp361_0[1:1], simp361_0[2:2]);
  NOR3 I28 (simp371_0[0:0], gfint_0[7:7], gfint_1[7:7], gfint_2[7:7]);
  NOR3 I29 (simp371_0[1:1], gfint_3[7:7], gfint_4[7:7], gfint_5[7:7]);
  INV I30 (simp371_0[2:2], gfint_6[7:7]);
  NAND3 I31 (o_0r0[7:7], simp371_0[0:0], simp371_0[1:1], simp371_0[2:2]);
  NOR3 I32 (simp381_0[0:0], gfint_0[8:8], gfint_1[8:8], gfint_2[8:8]);
  NOR3 I33 (simp381_0[1:1], gfint_3[8:8], gfint_4[8:8], gfint_5[8:8]);
  INV I34 (simp381_0[2:2], gfint_6[8:8]);
  NAND3 I35 (o_0r0[8:8], simp381_0[0:0], simp381_0[1:1], simp381_0[2:2]);
  NOR3 I36 (simp391_0[0:0], gfint_0[9:9], gfint_1[9:9], gfint_2[9:9]);
  NOR3 I37 (simp391_0[1:1], gfint_3[9:9], gfint_4[9:9], gfint_5[9:9]);
  INV I38 (simp391_0[2:2], gfint_6[9:9]);
  NAND3 I39 (o_0r0[9:9], simp391_0[0:0], simp391_0[1:1], simp391_0[2:2]);
  NOR3 I40 (simp401_0[0:0], gfint_0[10:10], gfint_1[10:10], gfint_2[10:10]);
  NOR3 I41 (simp401_0[1:1], gfint_3[10:10], gfint_4[10:10], gfint_5[10:10]);
  INV I42 (simp401_0[2:2], gfint_6[10:10]);
  NAND3 I43 (o_0r0[10:10], simp401_0[0:0], simp401_0[1:1], simp401_0[2:2]);
  NOR3 I44 (simp411_0[0:0], gfint_0[11:11], gfint_1[11:11], gfint_2[11:11]);
  NOR3 I45 (simp411_0[1:1], gfint_3[11:11], gfint_4[11:11], gfint_5[11:11]);
  INV I46 (simp411_0[2:2], gfint_6[11:11]);
  NAND3 I47 (o_0r0[11:11], simp411_0[0:0], simp411_0[1:1], simp411_0[2:2]);
  NOR3 I48 (simp421_0[0:0], gfint_0[12:12], gfint_1[12:12], gfint_2[12:12]);
  NOR3 I49 (simp421_0[1:1], gfint_3[12:12], gfint_4[12:12], gfint_5[12:12]);
  INV I50 (simp421_0[2:2], gfint_6[12:12]);
  NAND3 I51 (o_0r0[12:12], simp421_0[0:0], simp421_0[1:1], simp421_0[2:2]);
  NOR3 I52 (simp431_0[0:0], gfint_0[13:13], gfint_1[13:13], gfint_2[13:13]);
  NOR3 I53 (simp431_0[1:1], gfint_3[13:13], gfint_4[13:13], gfint_5[13:13]);
  INV I54 (simp431_0[2:2], gfint_6[13:13]);
  NAND3 I55 (o_0r0[13:13], simp431_0[0:0], simp431_0[1:1], simp431_0[2:2]);
  NOR3 I56 (simp441_0[0:0], gfint_0[14:14], gfint_1[14:14], gfint_2[14:14]);
  NOR3 I57 (simp441_0[1:1], gfint_3[14:14], gfint_4[14:14], gfint_5[14:14]);
  INV I58 (simp441_0[2:2], gfint_6[14:14]);
  NAND3 I59 (o_0r0[14:14], simp441_0[0:0], simp441_0[1:1], simp441_0[2:2]);
  NOR3 I60 (simp451_0[0:0], gfint_0[15:15], gfint_1[15:15], gfint_2[15:15]);
  NOR3 I61 (simp451_0[1:1], gfint_3[15:15], gfint_4[15:15], gfint_5[15:15]);
  INV I62 (simp451_0[2:2], gfint_6[15:15]);
  NAND3 I63 (o_0r0[15:15], simp451_0[0:0], simp451_0[1:1], simp451_0[2:2]);
  NOR3 I64 (simp461_0[0:0], gfint_0[16:16], gfint_1[16:16], gfint_2[16:16]);
  NOR3 I65 (simp461_0[1:1], gfint_3[16:16], gfint_4[16:16], gfint_5[16:16]);
  INV I66 (simp461_0[2:2], gfint_6[16:16]);
  NAND3 I67 (o_0r0[16:16], simp461_0[0:0], simp461_0[1:1], simp461_0[2:2]);
  NOR3 I68 (simp471_0[0:0], gfint_0[17:17], gfint_1[17:17], gfint_2[17:17]);
  NOR3 I69 (simp471_0[1:1], gfint_3[17:17], gfint_4[17:17], gfint_5[17:17]);
  INV I70 (simp471_0[2:2], gfint_6[17:17]);
  NAND3 I71 (o_0r0[17:17], simp471_0[0:0], simp471_0[1:1], simp471_0[2:2]);
  NOR3 I72 (simp481_0[0:0], gfint_0[18:18], gfint_1[18:18], gfint_2[18:18]);
  NOR3 I73 (simp481_0[1:1], gfint_3[18:18], gfint_4[18:18], gfint_5[18:18]);
  INV I74 (simp481_0[2:2], gfint_6[18:18]);
  NAND3 I75 (o_0r0[18:18], simp481_0[0:0], simp481_0[1:1], simp481_0[2:2]);
  NOR3 I76 (simp491_0[0:0], gfint_0[19:19], gfint_1[19:19], gfint_2[19:19]);
  NOR3 I77 (simp491_0[1:1], gfint_3[19:19], gfint_4[19:19], gfint_5[19:19]);
  INV I78 (simp491_0[2:2], gfint_6[19:19]);
  NAND3 I79 (o_0r0[19:19], simp491_0[0:0], simp491_0[1:1], simp491_0[2:2]);
  NOR3 I80 (simp501_0[0:0], gfint_0[20:20], gfint_1[20:20], gfint_2[20:20]);
  NOR3 I81 (simp501_0[1:1], gfint_3[20:20], gfint_4[20:20], gfint_5[20:20]);
  INV I82 (simp501_0[2:2], gfint_6[20:20]);
  NAND3 I83 (o_0r0[20:20], simp501_0[0:0], simp501_0[1:1], simp501_0[2:2]);
  NOR3 I84 (simp511_0[0:0], gfint_0[21:21], gfint_1[21:21], gfint_2[21:21]);
  NOR3 I85 (simp511_0[1:1], gfint_3[21:21], gfint_4[21:21], gfint_5[21:21]);
  INV I86 (simp511_0[2:2], gfint_6[21:21]);
  NAND3 I87 (o_0r0[21:21], simp511_0[0:0], simp511_0[1:1], simp511_0[2:2]);
  NOR3 I88 (simp521_0[0:0], gfint_0[22:22], gfint_1[22:22], gfint_2[22:22]);
  NOR3 I89 (simp521_0[1:1], gfint_3[22:22], gfint_4[22:22], gfint_5[22:22]);
  INV I90 (simp521_0[2:2], gfint_6[22:22]);
  NAND3 I91 (o_0r0[22:22], simp521_0[0:0], simp521_0[1:1], simp521_0[2:2]);
  NOR3 I92 (simp531_0[0:0], gfint_0[23:23], gfint_1[23:23], gfint_2[23:23]);
  NOR3 I93 (simp531_0[1:1], gfint_3[23:23], gfint_4[23:23], gfint_5[23:23]);
  INV I94 (simp531_0[2:2], gfint_6[23:23]);
  NAND3 I95 (o_0r0[23:23], simp531_0[0:0], simp531_0[1:1], simp531_0[2:2]);
  NOR3 I96 (simp541_0[0:0], gfint_0[24:24], gfint_1[24:24], gfint_2[24:24]);
  NOR3 I97 (simp541_0[1:1], gfint_3[24:24], gfint_4[24:24], gfint_5[24:24]);
  INV I98 (simp541_0[2:2], gfint_6[24:24]);
  NAND3 I99 (o_0r0[24:24], simp541_0[0:0], simp541_0[1:1], simp541_0[2:2]);
  NOR3 I100 (simp551_0[0:0], gfint_0[25:25], gfint_1[25:25], gfint_2[25:25]);
  NOR3 I101 (simp551_0[1:1], gfint_3[25:25], gfint_4[25:25], gfint_5[25:25]);
  INV I102 (simp551_0[2:2], gfint_6[25:25]);
  NAND3 I103 (o_0r0[25:25], simp551_0[0:0], simp551_0[1:1], simp551_0[2:2]);
  NOR3 I104 (simp561_0[0:0], gfint_0[26:26], gfint_1[26:26], gfint_2[26:26]);
  NOR3 I105 (simp561_0[1:1], gfint_3[26:26], gfint_4[26:26], gfint_5[26:26]);
  INV I106 (simp561_0[2:2], gfint_6[26:26]);
  NAND3 I107 (o_0r0[26:26], simp561_0[0:0], simp561_0[1:1], simp561_0[2:2]);
  NOR3 I108 (simp571_0[0:0], gfint_0[27:27], gfint_1[27:27], gfint_2[27:27]);
  NOR3 I109 (simp571_0[1:1], gfint_3[27:27], gfint_4[27:27], gfint_5[27:27]);
  INV I110 (simp571_0[2:2], gfint_6[27:27]);
  NAND3 I111 (o_0r0[27:27], simp571_0[0:0], simp571_0[1:1], simp571_0[2:2]);
  NOR3 I112 (simp581_0[0:0], gfint_0[28:28], gfint_1[28:28], gfint_2[28:28]);
  NOR3 I113 (simp581_0[1:1], gfint_3[28:28], gfint_4[28:28], gfint_5[28:28]);
  INV I114 (simp581_0[2:2], gfint_6[28:28]);
  NAND3 I115 (o_0r0[28:28], simp581_0[0:0], simp581_0[1:1], simp581_0[2:2]);
  NOR3 I116 (simp591_0[0:0], gfint_0[29:29], gfint_1[29:29], gfint_2[29:29]);
  NOR3 I117 (simp591_0[1:1], gfint_3[29:29], gfint_4[29:29], gfint_5[29:29]);
  INV I118 (simp591_0[2:2], gfint_6[29:29]);
  NAND3 I119 (o_0r0[29:29], simp591_0[0:0], simp591_0[1:1], simp591_0[2:2]);
  NOR3 I120 (simp601_0[0:0], gfint_0[30:30], gfint_1[30:30], gfint_2[30:30]);
  NOR3 I121 (simp601_0[1:1], gfint_3[30:30], gfint_4[30:30], gfint_5[30:30]);
  INV I122 (simp601_0[2:2], gfint_6[30:30]);
  NAND3 I123 (o_0r0[30:30], simp601_0[0:0], simp601_0[1:1], simp601_0[2:2]);
  NOR3 I124 (simp611_0[0:0], gfint_0[31:31], gfint_1[31:31], gfint_2[31:31]);
  NOR3 I125 (simp611_0[1:1], gfint_3[31:31], gfint_4[31:31], gfint_5[31:31]);
  INV I126 (simp611_0[2:2], gfint_6[31:31]);
  NAND3 I127 (o_0r0[31:31], simp611_0[0:0], simp611_0[1:1], simp611_0[2:2]);
  NOR3 I128 (simp621_0[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  NOR3 I129 (simp621_0[1:1], gtint_3[0:0], gtint_4[0:0], gtint_5[0:0]);
  INV I130 (simp621_0[2:2], gtint_6[0:0]);
  NAND3 I131 (o_0r1[0:0], simp621_0[0:0], simp621_0[1:1], simp621_0[2:2]);
  NOR3 I132 (simp631_0[0:0], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  NOR3 I133 (simp631_0[1:1], gtint_3[1:1], gtint_4[1:1], gtint_5[1:1]);
  INV I134 (simp631_0[2:2], gtint_6[1:1]);
  NAND3 I135 (o_0r1[1:1], simp631_0[0:0], simp631_0[1:1], simp631_0[2:2]);
  NOR3 I136 (simp641_0[0:0], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  NOR3 I137 (simp641_0[1:1], gtint_3[2:2], gtint_4[2:2], gtint_5[2:2]);
  INV I138 (simp641_0[2:2], gtint_6[2:2]);
  NAND3 I139 (o_0r1[2:2], simp641_0[0:0], simp641_0[1:1], simp641_0[2:2]);
  NOR3 I140 (simp651_0[0:0], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  NOR3 I141 (simp651_0[1:1], gtint_3[3:3], gtint_4[3:3], gtint_5[3:3]);
  INV I142 (simp651_0[2:2], gtint_6[3:3]);
  NAND3 I143 (o_0r1[3:3], simp651_0[0:0], simp651_0[1:1], simp651_0[2:2]);
  NOR3 I144 (simp661_0[0:0], gtint_0[4:4], gtint_1[4:4], gtint_2[4:4]);
  NOR3 I145 (simp661_0[1:1], gtint_3[4:4], gtint_4[4:4], gtint_5[4:4]);
  INV I146 (simp661_0[2:2], gtint_6[4:4]);
  NAND3 I147 (o_0r1[4:4], simp661_0[0:0], simp661_0[1:1], simp661_0[2:2]);
  NOR3 I148 (simp671_0[0:0], gtint_0[5:5], gtint_1[5:5], gtint_2[5:5]);
  NOR3 I149 (simp671_0[1:1], gtint_3[5:5], gtint_4[5:5], gtint_5[5:5]);
  INV I150 (simp671_0[2:2], gtint_6[5:5]);
  NAND3 I151 (o_0r1[5:5], simp671_0[0:0], simp671_0[1:1], simp671_0[2:2]);
  NOR3 I152 (simp681_0[0:0], gtint_0[6:6], gtint_1[6:6], gtint_2[6:6]);
  NOR3 I153 (simp681_0[1:1], gtint_3[6:6], gtint_4[6:6], gtint_5[6:6]);
  INV I154 (simp681_0[2:2], gtint_6[6:6]);
  NAND3 I155 (o_0r1[6:6], simp681_0[0:0], simp681_0[1:1], simp681_0[2:2]);
  NOR3 I156 (simp691_0[0:0], gtint_0[7:7], gtint_1[7:7], gtint_2[7:7]);
  NOR3 I157 (simp691_0[1:1], gtint_3[7:7], gtint_4[7:7], gtint_5[7:7]);
  INV I158 (simp691_0[2:2], gtint_6[7:7]);
  NAND3 I159 (o_0r1[7:7], simp691_0[0:0], simp691_0[1:1], simp691_0[2:2]);
  NOR3 I160 (simp701_0[0:0], gtint_0[8:8], gtint_1[8:8], gtint_2[8:8]);
  NOR3 I161 (simp701_0[1:1], gtint_3[8:8], gtint_4[8:8], gtint_5[8:8]);
  INV I162 (simp701_0[2:2], gtint_6[8:8]);
  NAND3 I163 (o_0r1[8:8], simp701_0[0:0], simp701_0[1:1], simp701_0[2:2]);
  NOR3 I164 (simp711_0[0:0], gtint_0[9:9], gtint_1[9:9], gtint_2[9:9]);
  NOR3 I165 (simp711_0[1:1], gtint_3[9:9], gtint_4[9:9], gtint_5[9:9]);
  INV I166 (simp711_0[2:2], gtint_6[9:9]);
  NAND3 I167 (o_0r1[9:9], simp711_0[0:0], simp711_0[1:1], simp711_0[2:2]);
  NOR3 I168 (simp721_0[0:0], gtint_0[10:10], gtint_1[10:10], gtint_2[10:10]);
  NOR3 I169 (simp721_0[1:1], gtint_3[10:10], gtint_4[10:10], gtint_5[10:10]);
  INV I170 (simp721_0[2:2], gtint_6[10:10]);
  NAND3 I171 (o_0r1[10:10], simp721_0[0:0], simp721_0[1:1], simp721_0[2:2]);
  NOR3 I172 (simp731_0[0:0], gtint_0[11:11], gtint_1[11:11], gtint_2[11:11]);
  NOR3 I173 (simp731_0[1:1], gtint_3[11:11], gtint_4[11:11], gtint_5[11:11]);
  INV I174 (simp731_0[2:2], gtint_6[11:11]);
  NAND3 I175 (o_0r1[11:11], simp731_0[0:0], simp731_0[1:1], simp731_0[2:2]);
  NOR3 I176 (simp741_0[0:0], gtint_0[12:12], gtint_1[12:12], gtint_2[12:12]);
  NOR3 I177 (simp741_0[1:1], gtint_3[12:12], gtint_4[12:12], gtint_5[12:12]);
  INV I178 (simp741_0[2:2], gtint_6[12:12]);
  NAND3 I179 (o_0r1[12:12], simp741_0[0:0], simp741_0[1:1], simp741_0[2:2]);
  NOR3 I180 (simp751_0[0:0], gtint_0[13:13], gtint_1[13:13], gtint_2[13:13]);
  NOR3 I181 (simp751_0[1:1], gtint_3[13:13], gtint_4[13:13], gtint_5[13:13]);
  INV I182 (simp751_0[2:2], gtint_6[13:13]);
  NAND3 I183 (o_0r1[13:13], simp751_0[0:0], simp751_0[1:1], simp751_0[2:2]);
  NOR3 I184 (simp761_0[0:0], gtint_0[14:14], gtint_1[14:14], gtint_2[14:14]);
  NOR3 I185 (simp761_0[1:1], gtint_3[14:14], gtint_4[14:14], gtint_5[14:14]);
  INV I186 (simp761_0[2:2], gtint_6[14:14]);
  NAND3 I187 (o_0r1[14:14], simp761_0[0:0], simp761_0[1:1], simp761_0[2:2]);
  NOR3 I188 (simp771_0[0:0], gtint_0[15:15], gtint_1[15:15], gtint_2[15:15]);
  NOR3 I189 (simp771_0[1:1], gtint_3[15:15], gtint_4[15:15], gtint_5[15:15]);
  INV I190 (simp771_0[2:2], gtint_6[15:15]);
  NAND3 I191 (o_0r1[15:15], simp771_0[0:0], simp771_0[1:1], simp771_0[2:2]);
  NOR3 I192 (simp781_0[0:0], gtint_0[16:16], gtint_1[16:16], gtint_2[16:16]);
  NOR3 I193 (simp781_0[1:1], gtint_3[16:16], gtint_4[16:16], gtint_5[16:16]);
  INV I194 (simp781_0[2:2], gtint_6[16:16]);
  NAND3 I195 (o_0r1[16:16], simp781_0[0:0], simp781_0[1:1], simp781_0[2:2]);
  NOR3 I196 (simp791_0[0:0], gtint_0[17:17], gtint_1[17:17], gtint_2[17:17]);
  NOR3 I197 (simp791_0[1:1], gtint_3[17:17], gtint_4[17:17], gtint_5[17:17]);
  INV I198 (simp791_0[2:2], gtint_6[17:17]);
  NAND3 I199 (o_0r1[17:17], simp791_0[0:0], simp791_0[1:1], simp791_0[2:2]);
  NOR3 I200 (simp801_0[0:0], gtint_0[18:18], gtint_1[18:18], gtint_2[18:18]);
  NOR3 I201 (simp801_0[1:1], gtint_3[18:18], gtint_4[18:18], gtint_5[18:18]);
  INV I202 (simp801_0[2:2], gtint_6[18:18]);
  NAND3 I203 (o_0r1[18:18], simp801_0[0:0], simp801_0[1:1], simp801_0[2:2]);
  NOR3 I204 (simp811_0[0:0], gtint_0[19:19], gtint_1[19:19], gtint_2[19:19]);
  NOR3 I205 (simp811_0[1:1], gtint_3[19:19], gtint_4[19:19], gtint_5[19:19]);
  INV I206 (simp811_0[2:2], gtint_6[19:19]);
  NAND3 I207 (o_0r1[19:19], simp811_0[0:0], simp811_0[1:1], simp811_0[2:2]);
  NOR3 I208 (simp821_0[0:0], gtint_0[20:20], gtint_1[20:20], gtint_2[20:20]);
  NOR3 I209 (simp821_0[1:1], gtint_3[20:20], gtint_4[20:20], gtint_5[20:20]);
  INV I210 (simp821_0[2:2], gtint_6[20:20]);
  NAND3 I211 (o_0r1[20:20], simp821_0[0:0], simp821_0[1:1], simp821_0[2:2]);
  NOR3 I212 (simp831_0[0:0], gtint_0[21:21], gtint_1[21:21], gtint_2[21:21]);
  NOR3 I213 (simp831_0[1:1], gtint_3[21:21], gtint_4[21:21], gtint_5[21:21]);
  INV I214 (simp831_0[2:2], gtint_6[21:21]);
  NAND3 I215 (o_0r1[21:21], simp831_0[0:0], simp831_0[1:1], simp831_0[2:2]);
  NOR3 I216 (simp841_0[0:0], gtint_0[22:22], gtint_1[22:22], gtint_2[22:22]);
  NOR3 I217 (simp841_0[1:1], gtint_3[22:22], gtint_4[22:22], gtint_5[22:22]);
  INV I218 (simp841_0[2:2], gtint_6[22:22]);
  NAND3 I219 (o_0r1[22:22], simp841_0[0:0], simp841_0[1:1], simp841_0[2:2]);
  NOR3 I220 (simp851_0[0:0], gtint_0[23:23], gtint_1[23:23], gtint_2[23:23]);
  NOR3 I221 (simp851_0[1:1], gtint_3[23:23], gtint_4[23:23], gtint_5[23:23]);
  INV I222 (simp851_0[2:2], gtint_6[23:23]);
  NAND3 I223 (o_0r1[23:23], simp851_0[0:0], simp851_0[1:1], simp851_0[2:2]);
  NOR3 I224 (simp861_0[0:0], gtint_0[24:24], gtint_1[24:24], gtint_2[24:24]);
  NOR3 I225 (simp861_0[1:1], gtint_3[24:24], gtint_4[24:24], gtint_5[24:24]);
  INV I226 (simp861_0[2:2], gtint_6[24:24]);
  NAND3 I227 (o_0r1[24:24], simp861_0[0:0], simp861_0[1:1], simp861_0[2:2]);
  NOR3 I228 (simp871_0[0:0], gtint_0[25:25], gtint_1[25:25], gtint_2[25:25]);
  NOR3 I229 (simp871_0[1:1], gtint_3[25:25], gtint_4[25:25], gtint_5[25:25]);
  INV I230 (simp871_0[2:2], gtint_6[25:25]);
  NAND3 I231 (o_0r1[25:25], simp871_0[0:0], simp871_0[1:1], simp871_0[2:2]);
  NOR3 I232 (simp881_0[0:0], gtint_0[26:26], gtint_1[26:26], gtint_2[26:26]);
  NOR3 I233 (simp881_0[1:1], gtint_3[26:26], gtint_4[26:26], gtint_5[26:26]);
  INV I234 (simp881_0[2:2], gtint_6[26:26]);
  NAND3 I235 (o_0r1[26:26], simp881_0[0:0], simp881_0[1:1], simp881_0[2:2]);
  NOR3 I236 (simp891_0[0:0], gtint_0[27:27], gtint_1[27:27], gtint_2[27:27]);
  NOR3 I237 (simp891_0[1:1], gtint_3[27:27], gtint_4[27:27], gtint_5[27:27]);
  INV I238 (simp891_0[2:2], gtint_6[27:27]);
  NAND3 I239 (o_0r1[27:27], simp891_0[0:0], simp891_0[1:1], simp891_0[2:2]);
  NOR3 I240 (simp901_0[0:0], gtint_0[28:28], gtint_1[28:28], gtint_2[28:28]);
  NOR3 I241 (simp901_0[1:1], gtint_3[28:28], gtint_4[28:28], gtint_5[28:28]);
  INV I242 (simp901_0[2:2], gtint_6[28:28]);
  NAND3 I243 (o_0r1[28:28], simp901_0[0:0], simp901_0[1:1], simp901_0[2:2]);
  NOR3 I244 (simp911_0[0:0], gtint_0[29:29], gtint_1[29:29], gtint_2[29:29]);
  NOR3 I245 (simp911_0[1:1], gtint_3[29:29], gtint_4[29:29], gtint_5[29:29]);
  INV I246 (simp911_0[2:2], gtint_6[29:29]);
  NAND3 I247 (o_0r1[29:29], simp911_0[0:0], simp911_0[1:1], simp911_0[2:2]);
  NOR3 I248 (simp921_0[0:0], gtint_0[30:30], gtint_1[30:30], gtint_2[30:30]);
  NOR3 I249 (simp921_0[1:1], gtint_3[30:30], gtint_4[30:30], gtint_5[30:30]);
  INV I250 (simp921_0[2:2], gtint_6[30:30]);
  NAND3 I251 (o_0r1[30:30], simp921_0[0:0], simp921_0[1:1], simp921_0[2:2]);
  NOR3 I252 (simp931_0[0:0], gtint_0[31:31], gtint_1[31:31], gtint_2[31:31]);
  NOR3 I253 (simp931_0[1:1], gtint_3[31:31], gtint_4[31:31], gtint_5[31:31]);
  INV I254 (simp931_0[2:2], gtint_6[31:31]);
  NAND3 I255 (o_0r1[31:31], simp931_0[0:0], simp931_0[1:1], simp931_0[2:2]);
  AND2 I256 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I257 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I258 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I259 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I260 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I261 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I262 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I263 (gtint_0[7:7], choice_0, i_0r1[7:7]);
  AND2 I264 (gtint_0[8:8], choice_0, i_0r1[8:8]);
  AND2 I265 (gtint_0[9:9], choice_0, i_0r1[9:9]);
  AND2 I266 (gtint_0[10:10], choice_0, i_0r1[10:10]);
  AND2 I267 (gtint_0[11:11], choice_0, i_0r1[11:11]);
  AND2 I268 (gtint_0[12:12], choice_0, i_0r1[12:12]);
  AND2 I269 (gtint_0[13:13], choice_0, i_0r1[13:13]);
  AND2 I270 (gtint_0[14:14], choice_0, i_0r1[14:14]);
  AND2 I271 (gtint_0[15:15], choice_0, i_0r1[15:15]);
  AND2 I272 (gtint_0[16:16], choice_0, i_0r1[16:16]);
  AND2 I273 (gtint_0[17:17], choice_0, i_0r1[17:17]);
  AND2 I274 (gtint_0[18:18], choice_0, i_0r1[18:18]);
  AND2 I275 (gtint_0[19:19], choice_0, i_0r1[19:19]);
  AND2 I276 (gtint_0[20:20], choice_0, i_0r1[20:20]);
  AND2 I277 (gtint_0[21:21], choice_0, i_0r1[21:21]);
  AND2 I278 (gtint_0[22:22], choice_0, i_0r1[22:22]);
  AND2 I279 (gtint_0[23:23], choice_0, i_0r1[23:23]);
  AND2 I280 (gtint_0[24:24], choice_0, i_0r1[24:24]);
  AND2 I281 (gtint_0[25:25], choice_0, i_0r1[25:25]);
  AND2 I282 (gtint_0[26:26], choice_0, i_0r1[26:26]);
  AND2 I283 (gtint_0[27:27], choice_0, i_0r1[27:27]);
  AND2 I284 (gtint_0[28:28], choice_0, i_0r1[28:28]);
  AND2 I285 (gtint_0[29:29], choice_0, i_0r1[29:29]);
  AND2 I286 (gtint_0[30:30], choice_0, i_0r1[30:30]);
  AND2 I287 (gtint_0[31:31], choice_0, i_0r1[31:31]);
  AND2 I288 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I289 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I290 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I291 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I292 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I293 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I294 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I295 (gtint_1[7:7], choice_1, i_1r1[7:7]);
  AND2 I296 (gtint_1[8:8], choice_1, i_1r1[8:8]);
  AND2 I297 (gtint_1[9:9], choice_1, i_1r1[9:9]);
  AND2 I298 (gtint_1[10:10], choice_1, i_1r1[10:10]);
  AND2 I299 (gtint_1[11:11], choice_1, i_1r1[11:11]);
  AND2 I300 (gtint_1[12:12], choice_1, i_1r1[12:12]);
  AND2 I301 (gtint_1[13:13], choice_1, i_1r1[13:13]);
  AND2 I302 (gtint_1[14:14], choice_1, i_1r1[14:14]);
  AND2 I303 (gtint_1[15:15], choice_1, i_1r1[15:15]);
  AND2 I304 (gtint_1[16:16], choice_1, i_1r1[16:16]);
  AND2 I305 (gtint_1[17:17], choice_1, i_1r1[17:17]);
  AND2 I306 (gtint_1[18:18], choice_1, i_1r1[18:18]);
  AND2 I307 (gtint_1[19:19], choice_1, i_1r1[19:19]);
  AND2 I308 (gtint_1[20:20], choice_1, i_1r1[20:20]);
  AND2 I309 (gtint_1[21:21], choice_1, i_1r1[21:21]);
  AND2 I310 (gtint_1[22:22], choice_1, i_1r1[22:22]);
  AND2 I311 (gtint_1[23:23], choice_1, i_1r1[23:23]);
  AND2 I312 (gtint_1[24:24], choice_1, i_1r1[24:24]);
  AND2 I313 (gtint_1[25:25], choice_1, i_1r1[25:25]);
  AND2 I314 (gtint_1[26:26], choice_1, i_1r1[26:26]);
  AND2 I315 (gtint_1[27:27], choice_1, i_1r1[27:27]);
  AND2 I316 (gtint_1[28:28], choice_1, i_1r1[28:28]);
  AND2 I317 (gtint_1[29:29], choice_1, i_1r1[29:29]);
  AND2 I318 (gtint_1[30:30], choice_1, i_1r1[30:30]);
  AND2 I319 (gtint_1[31:31], choice_1, i_1r1[31:31]);
  AND2 I320 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I321 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I322 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I323 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AND2 I324 (gtint_2[4:4], choice_2, i_2r1[4:4]);
  AND2 I325 (gtint_2[5:5], choice_2, i_2r1[5:5]);
  AND2 I326 (gtint_2[6:6], choice_2, i_2r1[6:6]);
  AND2 I327 (gtint_2[7:7], choice_2, i_2r1[7:7]);
  AND2 I328 (gtint_2[8:8], choice_2, i_2r1[8:8]);
  AND2 I329 (gtint_2[9:9], choice_2, i_2r1[9:9]);
  AND2 I330 (gtint_2[10:10], choice_2, i_2r1[10:10]);
  AND2 I331 (gtint_2[11:11], choice_2, i_2r1[11:11]);
  AND2 I332 (gtint_2[12:12], choice_2, i_2r1[12:12]);
  AND2 I333 (gtint_2[13:13], choice_2, i_2r1[13:13]);
  AND2 I334 (gtint_2[14:14], choice_2, i_2r1[14:14]);
  AND2 I335 (gtint_2[15:15], choice_2, i_2r1[15:15]);
  AND2 I336 (gtint_2[16:16], choice_2, i_2r1[16:16]);
  AND2 I337 (gtint_2[17:17], choice_2, i_2r1[17:17]);
  AND2 I338 (gtint_2[18:18], choice_2, i_2r1[18:18]);
  AND2 I339 (gtint_2[19:19], choice_2, i_2r1[19:19]);
  AND2 I340 (gtint_2[20:20], choice_2, i_2r1[20:20]);
  AND2 I341 (gtint_2[21:21], choice_2, i_2r1[21:21]);
  AND2 I342 (gtint_2[22:22], choice_2, i_2r1[22:22]);
  AND2 I343 (gtint_2[23:23], choice_2, i_2r1[23:23]);
  AND2 I344 (gtint_2[24:24], choice_2, i_2r1[24:24]);
  AND2 I345 (gtint_2[25:25], choice_2, i_2r1[25:25]);
  AND2 I346 (gtint_2[26:26], choice_2, i_2r1[26:26]);
  AND2 I347 (gtint_2[27:27], choice_2, i_2r1[27:27]);
  AND2 I348 (gtint_2[28:28], choice_2, i_2r1[28:28]);
  AND2 I349 (gtint_2[29:29], choice_2, i_2r1[29:29]);
  AND2 I350 (gtint_2[30:30], choice_2, i_2r1[30:30]);
  AND2 I351 (gtint_2[31:31], choice_2, i_2r1[31:31]);
  AND2 I352 (gtint_3[0:0], choice_3, i_3r1[0:0]);
  AND2 I353 (gtint_3[1:1], choice_3, i_3r1[1:1]);
  AND2 I354 (gtint_3[2:2], choice_3, i_3r1[2:2]);
  AND2 I355 (gtint_3[3:3], choice_3, i_3r1[3:3]);
  AND2 I356 (gtint_3[4:4], choice_3, i_3r1[4:4]);
  AND2 I357 (gtint_3[5:5], choice_3, i_3r1[5:5]);
  AND2 I358 (gtint_3[6:6], choice_3, i_3r1[6:6]);
  AND2 I359 (gtint_3[7:7], choice_3, i_3r1[7:7]);
  AND2 I360 (gtint_3[8:8], choice_3, i_3r1[8:8]);
  AND2 I361 (gtint_3[9:9], choice_3, i_3r1[9:9]);
  AND2 I362 (gtint_3[10:10], choice_3, i_3r1[10:10]);
  AND2 I363 (gtint_3[11:11], choice_3, i_3r1[11:11]);
  AND2 I364 (gtint_3[12:12], choice_3, i_3r1[12:12]);
  AND2 I365 (gtint_3[13:13], choice_3, i_3r1[13:13]);
  AND2 I366 (gtint_3[14:14], choice_3, i_3r1[14:14]);
  AND2 I367 (gtint_3[15:15], choice_3, i_3r1[15:15]);
  AND2 I368 (gtint_3[16:16], choice_3, i_3r1[16:16]);
  AND2 I369 (gtint_3[17:17], choice_3, i_3r1[17:17]);
  AND2 I370 (gtint_3[18:18], choice_3, i_3r1[18:18]);
  AND2 I371 (gtint_3[19:19], choice_3, i_3r1[19:19]);
  AND2 I372 (gtint_3[20:20], choice_3, i_3r1[20:20]);
  AND2 I373 (gtint_3[21:21], choice_3, i_3r1[21:21]);
  AND2 I374 (gtint_3[22:22], choice_3, i_3r1[22:22]);
  AND2 I375 (gtint_3[23:23], choice_3, i_3r1[23:23]);
  AND2 I376 (gtint_3[24:24], choice_3, i_3r1[24:24]);
  AND2 I377 (gtint_3[25:25], choice_3, i_3r1[25:25]);
  AND2 I378 (gtint_3[26:26], choice_3, i_3r1[26:26]);
  AND2 I379 (gtint_3[27:27], choice_3, i_3r1[27:27]);
  AND2 I380 (gtint_3[28:28], choice_3, i_3r1[28:28]);
  AND2 I381 (gtint_3[29:29], choice_3, i_3r1[29:29]);
  AND2 I382 (gtint_3[30:30], choice_3, i_3r1[30:30]);
  AND2 I383 (gtint_3[31:31], choice_3, i_3r1[31:31]);
  AND2 I384 (gtint_4[0:0], choice_4, i_4r1[0:0]);
  AND2 I385 (gtint_4[1:1], choice_4, i_4r1[1:1]);
  AND2 I386 (gtint_4[2:2], choice_4, i_4r1[2:2]);
  AND2 I387 (gtint_4[3:3], choice_4, i_4r1[3:3]);
  AND2 I388 (gtint_4[4:4], choice_4, i_4r1[4:4]);
  AND2 I389 (gtint_4[5:5], choice_4, i_4r1[5:5]);
  AND2 I390 (gtint_4[6:6], choice_4, i_4r1[6:6]);
  AND2 I391 (gtint_4[7:7], choice_4, i_4r1[7:7]);
  AND2 I392 (gtint_4[8:8], choice_4, i_4r1[8:8]);
  AND2 I393 (gtint_4[9:9], choice_4, i_4r1[9:9]);
  AND2 I394 (gtint_4[10:10], choice_4, i_4r1[10:10]);
  AND2 I395 (gtint_4[11:11], choice_4, i_4r1[11:11]);
  AND2 I396 (gtint_4[12:12], choice_4, i_4r1[12:12]);
  AND2 I397 (gtint_4[13:13], choice_4, i_4r1[13:13]);
  AND2 I398 (gtint_4[14:14], choice_4, i_4r1[14:14]);
  AND2 I399 (gtint_4[15:15], choice_4, i_4r1[15:15]);
  AND2 I400 (gtint_4[16:16], choice_4, i_4r1[16:16]);
  AND2 I401 (gtint_4[17:17], choice_4, i_4r1[17:17]);
  AND2 I402 (gtint_4[18:18], choice_4, i_4r1[18:18]);
  AND2 I403 (gtint_4[19:19], choice_4, i_4r1[19:19]);
  AND2 I404 (gtint_4[20:20], choice_4, i_4r1[20:20]);
  AND2 I405 (gtint_4[21:21], choice_4, i_4r1[21:21]);
  AND2 I406 (gtint_4[22:22], choice_4, i_4r1[22:22]);
  AND2 I407 (gtint_4[23:23], choice_4, i_4r1[23:23]);
  AND2 I408 (gtint_4[24:24], choice_4, i_4r1[24:24]);
  AND2 I409 (gtint_4[25:25], choice_4, i_4r1[25:25]);
  AND2 I410 (gtint_4[26:26], choice_4, i_4r1[26:26]);
  AND2 I411 (gtint_4[27:27], choice_4, i_4r1[27:27]);
  AND2 I412 (gtint_4[28:28], choice_4, i_4r1[28:28]);
  AND2 I413 (gtint_4[29:29], choice_4, i_4r1[29:29]);
  AND2 I414 (gtint_4[30:30], choice_4, i_4r1[30:30]);
  AND2 I415 (gtint_4[31:31], choice_4, i_4r1[31:31]);
  AND2 I416 (gtint_5[0:0], choice_5, i_5r1[0:0]);
  AND2 I417 (gtint_5[1:1], choice_5, i_5r1[1:1]);
  AND2 I418 (gtint_5[2:2], choice_5, i_5r1[2:2]);
  AND2 I419 (gtint_5[3:3], choice_5, i_5r1[3:3]);
  AND2 I420 (gtint_5[4:4], choice_5, i_5r1[4:4]);
  AND2 I421 (gtint_5[5:5], choice_5, i_5r1[5:5]);
  AND2 I422 (gtint_5[6:6], choice_5, i_5r1[6:6]);
  AND2 I423 (gtint_5[7:7], choice_5, i_5r1[7:7]);
  AND2 I424 (gtint_5[8:8], choice_5, i_5r1[8:8]);
  AND2 I425 (gtint_5[9:9], choice_5, i_5r1[9:9]);
  AND2 I426 (gtint_5[10:10], choice_5, i_5r1[10:10]);
  AND2 I427 (gtint_5[11:11], choice_5, i_5r1[11:11]);
  AND2 I428 (gtint_5[12:12], choice_5, i_5r1[12:12]);
  AND2 I429 (gtint_5[13:13], choice_5, i_5r1[13:13]);
  AND2 I430 (gtint_5[14:14], choice_5, i_5r1[14:14]);
  AND2 I431 (gtint_5[15:15], choice_5, i_5r1[15:15]);
  AND2 I432 (gtint_5[16:16], choice_5, i_5r1[16:16]);
  AND2 I433 (gtint_5[17:17], choice_5, i_5r1[17:17]);
  AND2 I434 (gtint_5[18:18], choice_5, i_5r1[18:18]);
  AND2 I435 (gtint_5[19:19], choice_5, i_5r1[19:19]);
  AND2 I436 (gtint_5[20:20], choice_5, i_5r1[20:20]);
  AND2 I437 (gtint_5[21:21], choice_5, i_5r1[21:21]);
  AND2 I438 (gtint_5[22:22], choice_5, i_5r1[22:22]);
  AND2 I439 (gtint_5[23:23], choice_5, i_5r1[23:23]);
  AND2 I440 (gtint_5[24:24], choice_5, i_5r1[24:24]);
  AND2 I441 (gtint_5[25:25], choice_5, i_5r1[25:25]);
  AND2 I442 (gtint_5[26:26], choice_5, i_5r1[26:26]);
  AND2 I443 (gtint_5[27:27], choice_5, i_5r1[27:27]);
  AND2 I444 (gtint_5[28:28], choice_5, i_5r1[28:28]);
  AND2 I445 (gtint_5[29:29], choice_5, i_5r1[29:29]);
  AND2 I446 (gtint_5[30:30], choice_5, i_5r1[30:30]);
  AND2 I447 (gtint_5[31:31], choice_5, i_5r1[31:31]);
  AND2 I448 (gtint_6[0:0], choice_6, i_6r1[0:0]);
  AND2 I449 (gtint_6[1:1], choice_6, i_6r1[1:1]);
  AND2 I450 (gtint_6[2:2], choice_6, i_6r1[2:2]);
  AND2 I451 (gtint_6[3:3], choice_6, i_6r1[3:3]);
  AND2 I452 (gtint_6[4:4], choice_6, i_6r1[4:4]);
  AND2 I453 (gtint_6[5:5], choice_6, i_6r1[5:5]);
  AND2 I454 (gtint_6[6:6], choice_6, i_6r1[6:6]);
  AND2 I455 (gtint_6[7:7], choice_6, i_6r1[7:7]);
  AND2 I456 (gtint_6[8:8], choice_6, i_6r1[8:8]);
  AND2 I457 (gtint_6[9:9], choice_6, i_6r1[9:9]);
  AND2 I458 (gtint_6[10:10], choice_6, i_6r1[10:10]);
  AND2 I459 (gtint_6[11:11], choice_6, i_6r1[11:11]);
  AND2 I460 (gtint_6[12:12], choice_6, i_6r1[12:12]);
  AND2 I461 (gtint_6[13:13], choice_6, i_6r1[13:13]);
  AND2 I462 (gtint_6[14:14], choice_6, i_6r1[14:14]);
  AND2 I463 (gtint_6[15:15], choice_6, i_6r1[15:15]);
  AND2 I464 (gtint_6[16:16], choice_6, i_6r1[16:16]);
  AND2 I465 (gtint_6[17:17], choice_6, i_6r1[17:17]);
  AND2 I466 (gtint_6[18:18], choice_6, i_6r1[18:18]);
  AND2 I467 (gtint_6[19:19], choice_6, i_6r1[19:19]);
  AND2 I468 (gtint_6[20:20], choice_6, i_6r1[20:20]);
  AND2 I469 (gtint_6[21:21], choice_6, i_6r1[21:21]);
  AND2 I470 (gtint_6[22:22], choice_6, i_6r1[22:22]);
  AND2 I471 (gtint_6[23:23], choice_6, i_6r1[23:23]);
  AND2 I472 (gtint_6[24:24], choice_6, i_6r1[24:24]);
  AND2 I473 (gtint_6[25:25], choice_6, i_6r1[25:25]);
  AND2 I474 (gtint_6[26:26], choice_6, i_6r1[26:26]);
  AND2 I475 (gtint_6[27:27], choice_6, i_6r1[27:27]);
  AND2 I476 (gtint_6[28:28], choice_6, i_6r1[28:28]);
  AND2 I477 (gtint_6[29:29], choice_6, i_6r1[29:29]);
  AND2 I478 (gtint_6[30:30], choice_6, i_6r1[30:30]);
  AND2 I479 (gtint_6[31:31], choice_6, i_6r1[31:31]);
  AND2 I480 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I481 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I482 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I483 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I484 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I485 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I486 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I487 (gfint_0[7:7], choice_0, i_0r0[7:7]);
  AND2 I488 (gfint_0[8:8], choice_0, i_0r0[8:8]);
  AND2 I489 (gfint_0[9:9], choice_0, i_0r0[9:9]);
  AND2 I490 (gfint_0[10:10], choice_0, i_0r0[10:10]);
  AND2 I491 (gfint_0[11:11], choice_0, i_0r0[11:11]);
  AND2 I492 (gfint_0[12:12], choice_0, i_0r0[12:12]);
  AND2 I493 (gfint_0[13:13], choice_0, i_0r0[13:13]);
  AND2 I494 (gfint_0[14:14], choice_0, i_0r0[14:14]);
  AND2 I495 (gfint_0[15:15], choice_0, i_0r0[15:15]);
  AND2 I496 (gfint_0[16:16], choice_0, i_0r0[16:16]);
  AND2 I497 (gfint_0[17:17], choice_0, i_0r0[17:17]);
  AND2 I498 (gfint_0[18:18], choice_0, i_0r0[18:18]);
  AND2 I499 (gfint_0[19:19], choice_0, i_0r0[19:19]);
  AND2 I500 (gfint_0[20:20], choice_0, i_0r0[20:20]);
  AND2 I501 (gfint_0[21:21], choice_0, i_0r0[21:21]);
  AND2 I502 (gfint_0[22:22], choice_0, i_0r0[22:22]);
  AND2 I503 (gfint_0[23:23], choice_0, i_0r0[23:23]);
  AND2 I504 (gfint_0[24:24], choice_0, i_0r0[24:24]);
  AND2 I505 (gfint_0[25:25], choice_0, i_0r0[25:25]);
  AND2 I506 (gfint_0[26:26], choice_0, i_0r0[26:26]);
  AND2 I507 (gfint_0[27:27], choice_0, i_0r0[27:27]);
  AND2 I508 (gfint_0[28:28], choice_0, i_0r0[28:28]);
  AND2 I509 (gfint_0[29:29], choice_0, i_0r0[29:29]);
  AND2 I510 (gfint_0[30:30], choice_0, i_0r0[30:30]);
  AND2 I511 (gfint_0[31:31], choice_0, i_0r0[31:31]);
  AND2 I512 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I513 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I514 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I515 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I516 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I517 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I518 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I519 (gfint_1[7:7], choice_1, i_1r0[7:7]);
  AND2 I520 (gfint_1[8:8], choice_1, i_1r0[8:8]);
  AND2 I521 (gfint_1[9:9], choice_1, i_1r0[9:9]);
  AND2 I522 (gfint_1[10:10], choice_1, i_1r0[10:10]);
  AND2 I523 (gfint_1[11:11], choice_1, i_1r0[11:11]);
  AND2 I524 (gfint_1[12:12], choice_1, i_1r0[12:12]);
  AND2 I525 (gfint_1[13:13], choice_1, i_1r0[13:13]);
  AND2 I526 (gfint_1[14:14], choice_1, i_1r0[14:14]);
  AND2 I527 (gfint_1[15:15], choice_1, i_1r0[15:15]);
  AND2 I528 (gfint_1[16:16], choice_1, i_1r0[16:16]);
  AND2 I529 (gfint_1[17:17], choice_1, i_1r0[17:17]);
  AND2 I530 (gfint_1[18:18], choice_1, i_1r0[18:18]);
  AND2 I531 (gfint_1[19:19], choice_1, i_1r0[19:19]);
  AND2 I532 (gfint_1[20:20], choice_1, i_1r0[20:20]);
  AND2 I533 (gfint_1[21:21], choice_1, i_1r0[21:21]);
  AND2 I534 (gfint_1[22:22], choice_1, i_1r0[22:22]);
  AND2 I535 (gfint_1[23:23], choice_1, i_1r0[23:23]);
  AND2 I536 (gfint_1[24:24], choice_1, i_1r0[24:24]);
  AND2 I537 (gfint_1[25:25], choice_1, i_1r0[25:25]);
  AND2 I538 (gfint_1[26:26], choice_1, i_1r0[26:26]);
  AND2 I539 (gfint_1[27:27], choice_1, i_1r0[27:27]);
  AND2 I540 (gfint_1[28:28], choice_1, i_1r0[28:28]);
  AND2 I541 (gfint_1[29:29], choice_1, i_1r0[29:29]);
  AND2 I542 (gfint_1[30:30], choice_1, i_1r0[30:30]);
  AND2 I543 (gfint_1[31:31], choice_1, i_1r0[31:31]);
  AND2 I544 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I545 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I546 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I547 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AND2 I548 (gfint_2[4:4], choice_2, i_2r0[4:4]);
  AND2 I549 (gfint_2[5:5], choice_2, i_2r0[5:5]);
  AND2 I550 (gfint_2[6:6], choice_2, i_2r0[6:6]);
  AND2 I551 (gfint_2[7:7], choice_2, i_2r0[7:7]);
  AND2 I552 (gfint_2[8:8], choice_2, i_2r0[8:8]);
  AND2 I553 (gfint_2[9:9], choice_2, i_2r0[9:9]);
  AND2 I554 (gfint_2[10:10], choice_2, i_2r0[10:10]);
  AND2 I555 (gfint_2[11:11], choice_2, i_2r0[11:11]);
  AND2 I556 (gfint_2[12:12], choice_2, i_2r0[12:12]);
  AND2 I557 (gfint_2[13:13], choice_2, i_2r0[13:13]);
  AND2 I558 (gfint_2[14:14], choice_2, i_2r0[14:14]);
  AND2 I559 (gfint_2[15:15], choice_2, i_2r0[15:15]);
  AND2 I560 (gfint_2[16:16], choice_2, i_2r0[16:16]);
  AND2 I561 (gfint_2[17:17], choice_2, i_2r0[17:17]);
  AND2 I562 (gfint_2[18:18], choice_2, i_2r0[18:18]);
  AND2 I563 (gfint_2[19:19], choice_2, i_2r0[19:19]);
  AND2 I564 (gfint_2[20:20], choice_2, i_2r0[20:20]);
  AND2 I565 (gfint_2[21:21], choice_2, i_2r0[21:21]);
  AND2 I566 (gfint_2[22:22], choice_2, i_2r0[22:22]);
  AND2 I567 (gfint_2[23:23], choice_2, i_2r0[23:23]);
  AND2 I568 (gfint_2[24:24], choice_2, i_2r0[24:24]);
  AND2 I569 (gfint_2[25:25], choice_2, i_2r0[25:25]);
  AND2 I570 (gfint_2[26:26], choice_2, i_2r0[26:26]);
  AND2 I571 (gfint_2[27:27], choice_2, i_2r0[27:27]);
  AND2 I572 (gfint_2[28:28], choice_2, i_2r0[28:28]);
  AND2 I573 (gfint_2[29:29], choice_2, i_2r0[29:29]);
  AND2 I574 (gfint_2[30:30], choice_2, i_2r0[30:30]);
  AND2 I575 (gfint_2[31:31], choice_2, i_2r0[31:31]);
  AND2 I576 (gfint_3[0:0], choice_3, i_3r0[0:0]);
  AND2 I577 (gfint_3[1:1], choice_3, i_3r0[1:1]);
  AND2 I578 (gfint_3[2:2], choice_3, i_3r0[2:2]);
  AND2 I579 (gfint_3[3:3], choice_3, i_3r0[3:3]);
  AND2 I580 (gfint_3[4:4], choice_3, i_3r0[4:4]);
  AND2 I581 (gfint_3[5:5], choice_3, i_3r0[5:5]);
  AND2 I582 (gfint_3[6:6], choice_3, i_3r0[6:6]);
  AND2 I583 (gfint_3[7:7], choice_3, i_3r0[7:7]);
  AND2 I584 (gfint_3[8:8], choice_3, i_3r0[8:8]);
  AND2 I585 (gfint_3[9:9], choice_3, i_3r0[9:9]);
  AND2 I586 (gfint_3[10:10], choice_3, i_3r0[10:10]);
  AND2 I587 (gfint_3[11:11], choice_3, i_3r0[11:11]);
  AND2 I588 (gfint_3[12:12], choice_3, i_3r0[12:12]);
  AND2 I589 (gfint_3[13:13], choice_3, i_3r0[13:13]);
  AND2 I590 (gfint_3[14:14], choice_3, i_3r0[14:14]);
  AND2 I591 (gfint_3[15:15], choice_3, i_3r0[15:15]);
  AND2 I592 (gfint_3[16:16], choice_3, i_3r0[16:16]);
  AND2 I593 (gfint_3[17:17], choice_3, i_3r0[17:17]);
  AND2 I594 (gfint_3[18:18], choice_3, i_3r0[18:18]);
  AND2 I595 (gfint_3[19:19], choice_3, i_3r0[19:19]);
  AND2 I596 (gfint_3[20:20], choice_3, i_3r0[20:20]);
  AND2 I597 (gfint_3[21:21], choice_3, i_3r0[21:21]);
  AND2 I598 (gfint_3[22:22], choice_3, i_3r0[22:22]);
  AND2 I599 (gfint_3[23:23], choice_3, i_3r0[23:23]);
  AND2 I600 (gfint_3[24:24], choice_3, i_3r0[24:24]);
  AND2 I601 (gfint_3[25:25], choice_3, i_3r0[25:25]);
  AND2 I602 (gfint_3[26:26], choice_3, i_3r0[26:26]);
  AND2 I603 (gfint_3[27:27], choice_3, i_3r0[27:27]);
  AND2 I604 (gfint_3[28:28], choice_3, i_3r0[28:28]);
  AND2 I605 (gfint_3[29:29], choice_3, i_3r0[29:29]);
  AND2 I606 (gfint_3[30:30], choice_3, i_3r0[30:30]);
  AND2 I607 (gfint_3[31:31], choice_3, i_3r0[31:31]);
  AND2 I608 (gfint_4[0:0], choice_4, i_4r0[0:0]);
  AND2 I609 (gfint_4[1:1], choice_4, i_4r0[1:1]);
  AND2 I610 (gfint_4[2:2], choice_4, i_4r0[2:2]);
  AND2 I611 (gfint_4[3:3], choice_4, i_4r0[3:3]);
  AND2 I612 (gfint_4[4:4], choice_4, i_4r0[4:4]);
  AND2 I613 (gfint_4[5:5], choice_4, i_4r0[5:5]);
  AND2 I614 (gfint_4[6:6], choice_4, i_4r0[6:6]);
  AND2 I615 (gfint_4[7:7], choice_4, i_4r0[7:7]);
  AND2 I616 (gfint_4[8:8], choice_4, i_4r0[8:8]);
  AND2 I617 (gfint_4[9:9], choice_4, i_4r0[9:9]);
  AND2 I618 (gfint_4[10:10], choice_4, i_4r0[10:10]);
  AND2 I619 (gfint_4[11:11], choice_4, i_4r0[11:11]);
  AND2 I620 (gfint_4[12:12], choice_4, i_4r0[12:12]);
  AND2 I621 (gfint_4[13:13], choice_4, i_4r0[13:13]);
  AND2 I622 (gfint_4[14:14], choice_4, i_4r0[14:14]);
  AND2 I623 (gfint_4[15:15], choice_4, i_4r0[15:15]);
  AND2 I624 (gfint_4[16:16], choice_4, i_4r0[16:16]);
  AND2 I625 (gfint_4[17:17], choice_4, i_4r0[17:17]);
  AND2 I626 (gfint_4[18:18], choice_4, i_4r0[18:18]);
  AND2 I627 (gfint_4[19:19], choice_4, i_4r0[19:19]);
  AND2 I628 (gfint_4[20:20], choice_4, i_4r0[20:20]);
  AND2 I629 (gfint_4[21:21], choice_4, i_4r0[21:21]);
  AND2 I630 (gfint_4[22:22], choice_4, i_4r0[22:22]);
  AND2 I631 (gfint_4[23:23], choice_4, i_4r0[23:23]);
  AND2 I632 (gfint_4[24:24], choice_4, i_4r0[24:24]);
  AND2 I633 (gfint_4[25:25], choice_4, i_4r0[25:25]);
  AND2 I634 (gfint_4[26:26], choice_4, i_4r0[26:26]);
  AND2 I635 (gfint_4[27:27], choice_4, i_4r0[27:27]);
  AND2 I636 (gfint_4[28:28], choice_4, i_4r0[28:28]);
  AND2 I637 (gfint_4[29:29], choice_4, i_4r0[29:29]);
  AND2 I638 (gfint_4[30:30], choice_4, i_4r0[30:30]);
  AND2 I639 (gfint_4[31:31], choice_4, i_4r0[31:31]);
  AND2 I640 (gfint_5[0:0], choice_5, i_5r0[0:0]);
  AND2 I641 (gfint_5[1:1], choice_5, i_5r0[1:1]);
  AND2 I642 (gfint_5[2:2], choice_5, i_5r0[2:2]);
  AND2 I643 (gfint_5[3:3], choice_5, i_5r0[3:3]);
  AND2 I644 (gfint_5[4:4], choice_5, i_5r0[4:4]);
  AND2 I645 (gfint_5[5:5], choice_5, i_5r0[5:5]);
  AND2 I646 (gfint_5[6:6], choice_5, i_5r0[6:6]);
  AND2 I647 (gfint_5[7:7], choice_5, i_5r0[7:7]);
  AND2 I648 (gfint_5[8:8], choice_5, i_5r0[8:8]);
  AND2 I649 (gfint_5[9:9], choice_5, i_5r0[9:9]);
  AND2 I650 (gfint_5[10:10], choice_5, i_5r0[10:10]);
  AND2 I651 (gfint_5[11:11], choice_5, i_5r0[11:11]);
  AND2 I652 (gfint_5[12:12], choice_5, i_5r0[12:12]);
  AND2 I653 (gfint_5[13:13], choice_5, i_5r0[13:13]);
  AND2 I654 (gfint_5[14:14], choice_5, i_5r0[14:14]);
  AND2 I655 (gfint_5[15:15], choice_5, i_5r0[15:15]);
  AND2 I656 (gfint_5[16:16], choice_5, i_5r0[16:16]);
  AND2 I657 (gfint_5[17:17], choice_5, i_5r0[17:17]);
  AND2 I658 (gfint_5[18:18], choice_5, i_5r0[18:18]);
  AND2 I659 (gfint_5[19:19], choice_5, i_5r0[19:19]);
  AND2 I660 (gfint_5[20:20], choice_5, i_5r0[20:20]);
  AND2 I661 (gfint_5[21:21], choice_5, i_5r0[21:21]);
  AND2 I662 (gfint_5[22:22], choice_5, i_5r0[22:22]);
  AND2 I663 (gfint_5[23:23], choice_5, i_5r0[23:23]);
  AND2 I664 (gfint_5[24:24], choice_5, i_5r0[24:24]);
  AND2 I665 (gfint_5[25:25], choice_5, i_5r0[25:25]);
  AND2 I666 (gfint_5[26:26], choice_5, i_5r0[26:26]);
  AND2 I667 (gfint_5[27:27], choice_5, i_5r0[27:27]);
  AND2 I668 (gfint_5[28:28], choice_5, i_5r0[28:28]);
  AND2 I669 (gfint_5[29:29], choice_5, i_5r0[29:29]);
  AND2 I670 (gfint_5[30:30], choice_5, i_5r0[30:30]);
  AND2 I671 (gfint_5[31:31], choice_5, i_5r0[31:31]);
  AND2 I672 (gfint_6[0:0], choice_6, i_6r0[0:0]);
  AND2 I673 (gfint_6[1:1], choice_6, i_6r0[1:1]);
  AND2 I674 (gfint_6[2:2], choice_6, i_6r0[2:2]);
  AND2 I675 (gfint_6[3:3], choice_6, i_6r0[3:3]);
  AND2 I676 (gfint_6[4:4], choice_6, i_6r0[4:4]);
  AND2 I677 (gfint_6[5:5], choice_6, i_6r0[5:5]);
  AND2 I678 (gfint_6[6:6], choice_6, i_6r0[6:6]);
  AND2 I679 (gfint_6[7:7], choice_6, i_6r0[7:7]);
  AND2 I680 (gfint_6[8:8], choice_6, i_6r0[8:8]);
  AND2 I681 (gfint_6[9:9], choice_6, i_6r0[9:9]);
  AND2 I682 (gfint_6[10:10], choice_6, i_6r0[10:10]);
  AND2 I683 (gfint_6[11:11], choice_6, i_6r0[11:11]);
  AND2 I684 (gfint_6[12:12], choice_6, i_6r0[12:12]);
  AND2 I685 (gfint_6[13:13], choice_6, i_6r0[13:13]);
  AND2 I686 (gfint_6[14:14], choice_6, i_6r0[14:14]);
  AND2 I687 (gfint_6[15:15], choice_6, i_6r0[15:15]);
  AND2 I688 (gfint_6[16:16], choice_6, i_6r0[16:16]);
  AND2 I689 (gfint_6[17:17], choice_6, i_6r0[17:17]);
  AND2 I690 (gfint_6[18:18], choice_6, i_6r0[18:18]);
  AND2 I691 (gfint_6[19:19], choice_6, i_6r0[19:19]);
  AND2 I692 (gfint_6[20:20], choice_6, i_6r0[20:20]);
  AND2 I693 (gfint_6[21:21], choice_6, i_6r0[21:21]);
  AND2 I694 (gfint_6[22:22], choice_6, i_6r0[22:22]);
  AND2 I695 (gfint_6[23:23], choice_6, i_6r0[23:23]);
  AND2 I696 (gfint_6[24:24], choice_6, i_6r0[24:24]);
  AND2 I697 (gfint_6[25:25], choice_6, i_6r0[25:25]);
  AND2 I698 (gfint_6[26:26], choice_6, i_6r0[26:26]);
  AND2 I699 (gfint_6[27:27], choice_6, i_6r0[27:27]);
  AND2 I700 (gfint_6[28:28], choice_6, i_6r0[28:28]);
  AND2 I701 (gfint_6[29:29], choice_6, i_6r0[29:29]);
  AND2 I702 (gfint_6[30:30], choice_6, i_6r0[30:30]);
  AND2 I703 (gfint_6[31:31], choice_6, i_6r0[31:31]);
  OR2 I704 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I705 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I706 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I707 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I708 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I709 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I710 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I711 (comp0_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I712 (comp0_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I713 (comp0_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I714 (comp0_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I715 (comp0_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I716 (comp0_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I717 (comp0_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I718 (comp0_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I719 (comp0_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I720 (comp0_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I721 (comp0_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I722 (comp0_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I723 (comp0_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I724 (comp0_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I725 (comp0_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I726 (comp0_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I727 (comp0_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I728 (comp0_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I729 (comp0_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I730 (comp0_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I731 (comp0_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I732 (comp0_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I733 (comp0_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I734 (comp0_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I735 (comp0_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  C3 I736 (simp5751_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I737 (simp5751_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I738 (simp5751_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I739 (simp5751_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I740 (simp5751_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I741 (simp5751_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I742 (simp5751_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I743 (simp5751_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I744 (simp5751_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I745 (simp5751_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I746 (simp5751_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I747 (simp5752_0[0:0], simp5751_0[0:0], simp5751_0[1:1], simp5751_0[2:2]);
  C3 I748 (simp5752_0[1:1], simp5751_0[3:3], simp5751_0[4:4], simp5751_0[5:5]);
  C3 I749 (simp5752_0[2:2], simp5751_0[6:6], simp5751_0[7:7], simp5751_0[8:8]);
  C2 I750 (simp5752_0[3:3], simp5751_0[9:9], simp5751_0[10:10]);
  C3 I751 (simp5753_0[0:0], simp5752_0[0:0], simp5752_0[1:1], simp5752_0[2:2]);
  BUFF I752 (simp5753_0[1:1], simp5752_0[3:3]);
  C2 I753 (icomp_0, simp5753_0[0:0], simp5753_0[1:1]);
  OR2 I754 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I755 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I756 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I757 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I758 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I759 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I760 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  OR2 I761 (comp1_0[7:7], i_1r0[7:7], i_1r1[7:7]);
  OR2 I762 (comp1_0[8:8], i_1r0[8:8], i_1r1[8:8]);
  OR2 I763 (comp1_0[9:9], i_1r0[9:9], i_1r1[9:9]);
  OR2 I764 (comp1_0[10:10], i_1r0[10:10], i_1r1[10:10]);
  OR2 I765 (comp1_0[11:11], i_1r0[11:11], i_1r1[11:11]);
  OR2 I766 (comp1_0[12:12], i_1r0[12:12], i_1r1[12:12]);
  OR2 I767 (comp1_0[13:13], i_1r0[13:13], i_1r1[13:13]);
  OR2 I768 (comp1_0[14:14], i_1r0[14:14], i_1r1[14:14]);
  OR2 I769 (comp1_0[15:15], i_1r0[15:15], i_1r1[15:15]);
  OR2 I770 (comp1_0[16:16], i_1r0[16:16], i_1r1[16:16]);
  OR2 I771 (comp1_0[17:17], i_1r0[17:17], i_1r1[17:17]);
  OR2 I772 (comp1_0[18:18], i_1r0[18:18], i_1r1[18:18]);
  OR2 I773 (comp1_0[19:19], i_1r0[19:19], i_1r1[19:19]);
  OR2 I774 (comp1_0[20:20], i_1r0[20:20], i_1r1[20:20]);
  OR2 I775 (comp1_0[21:21], i_1r0[21:21], i_1r1[21:21]);
  OR2 I776 (comp1_0[22:22], i_1r0[22:22], i_1r1[22:22]);
  OR2 I777 (comp1_0[23:23], i_1r0[23:23], i_1r1[23:23]);
  OR2 I778 (comp1_0[24:24], i_1r0[24:24], i_1r1[24:24]);
  OR2 I779 (comp1_0[25:25], i_1r0[25:25], i_1r1[25:25]);
  OR2 I780 (comp1_0[26:26], i_1r0[26:26], i_1r1[26:26]);
  OR2 I781 (comp1_0[27:27], i_1r0[27:27], i_1r1[27:27]);
  OR2 I782 (comp1_0[28:28], i_1r0[28:28], i_1r1[28:28]);
  OR2 I783 (comp1_0[29:29], i_1r0[29:29], i_1r1[29:29]);
  OR2 I784 (comp1_0[30:30], i_1r0[30:30], i_1r1[30:30]);
  OR2 I785 (comp1_0[31:31], i_1r0[31:31], i_1r1[31:31]);
  C3 I786 (simp6091_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I787 (simp6091_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  C3 I788 (simp6091_0[2:2], comp1_0[6:6], comp1_0[7:7], comp1_0[8:8]);
  C3 I789 (simp6091_0[3:3], comp1_0[9:9], comp1_0[10:10], comp1_0[11:11]);
  C3 I790 (simp6091_0[4:4], comp1_0[12:12], comp1_0[13:13], comp1_0[14:14]);
  C3 I791 (simp6091_0[5:5], comp1_0[15:15], comp1_0[16:16], comp1_0[17:17]);
  C3 I792 (simp6091_0[6:6], comp1_0[18:18], comp1_0[19:19], comp1_0[20:20]);
  C3 I793 (simp6091_0[7:7], comp1_0[21:21], comp1_0[22:22], comp1_0[23:23]);
  C3 I794 (simp6091_0[8:8], comp1_0[24:24], comp1_0[25:25], comp1_0[26:26]);
  C3 I795 (simp6091_0[9:9], comp1_0[27:27], comp1_0[28:28], comp1_0[29:29]);
  C2 I796 (simp6091_0[10:10], comp1_0[30:30], comp1_0[31:31]);
  C3 I797 (simp6092_0[0:0], simp6091_0[0:0], simp6091_0[1:1], simp6091_0[2:2]);
  C3 I798 (simp6092_0[1:1], simp6091_0[3:3], simp6091_0[4:4], simp6091_0[5:5]);
  C3 I799 (simp6092_0[2:2], simp6091_0[6:6], simp6091_0[7:7], simp6091_0[8:8]);
  C2 I800 (simp6092_0[3:3], simp6091_0[9:9], simp6091_0[10:10]);
  C3 I801 (simp6093_0[0:0], simp6092_0[0:0], simp6092_0[1:1], simp6092_0[2:2]);
  BUFF I802 (simp6093_0[1:1], simp6092_0[3:3]);
  C2 I803 (icomp_1, simp6093_0[0:0], simp6093_0[1:1]);
  OR2 I804 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I805 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I806 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2 I807 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  OR2 I808 (comp2_0[4:4], i_2r0[4:4], i_2r1[4:4]);
  OR2 I809 (comp2_0[5:5], i_2r0[5:5], i_2r1[5:5]);
  OR2 I810 (comp2_0[6:6], i_2r0[6:6], i_2r1[6:6]);
  OR2 I811 (comp2_0[7:7], i_2r0[7:7], i_2r1[7:7]);
  OR2 I812 (comp2_0[8:8], i_2r0[8:8], i_2r1[8:8]);
  OR2 I813 (comp2_0[9:9], i_2r0[9:9], i_2r1[9:9]);
  OR2 I814 (comp2_0[10:10], i_2r0[10:10], i_2r1[10:10]);
  OR2 I815 (comp2_0[11:11], i_2r0[11:11], i_2r1[11:11]);
  OR2 I816 (comp2_0[12:12], i_2r0[12:12], i_2r1[12:12]);
  OR2 I817 (comp2_0[13:13], i_2r0[13:13], i_2r1[13:13]);
  OR2 I818 (comp2_0[14:14], i_2r0[14:14], i_2r1[14:14]);
  OR2 I819 (comp2_0[15:15], i_2r0[15:15], i_2r1[15:15]);
  OR2 I820 (comp2_0[16:16], i_2r0[16:16], i_2r1[16:16]);
  OR2 I821 (comp2_0[17:17], i_2r0[17:17], i_2r1[17:17]);
  OR2 I822 (comp2_0[18:18], i_2r0[18:18], i_2r1[18:18]);
  OR2 I823 (comp2_0[19:19], i_2r0[19:19], i_2r1[19:19]);
  OR2 I824 (comp2_0[20:20], i_2r0[20:20], i_2r1[20:20]);
  OR2 I825 (comp2_0[21:21], i_2r0[21:21], i_2r1[21:21]);
  OR2 I826 (comp2_0[22:22], i_2r0[22:22], i_2r1[22:22]);
  OR2 I827 (comp2_0[23:23], i_2r0[23:23], i_2r1[23:23]);
  OR2 I828 (comp2_0[24:24], i_2r0[24:24], i_2r1[24:24]);
  OR2 I829 (comp2_0[25:25], i_2r0[25:25], i_2r1[25:25]);
  OR2 I830 (comp2_0[26:26], i_2r0[26:26], i_2r1[26:26]);
  OR2 I831 (comp2_0[27:27], i_2r0[27:27], i_2r1[27:27]);
  OR2 I832 (comp2_0[28:28], i_2r0[28:28], i_2r1[28:28]);
  OR2 I833 (comp2_0[29:29], i_2r0[29:29], i_2r1[29:29]);
  OR2 I834 (comp2_0[30:30], i_2r0[30:30], i_2r1[30:30]);
  OR2 I835 (comp2_0[31:31], i_2r0[31:31], i_2r1[31:31]);
  C3 I836 (simp6431_0[0:0], comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C3 I837 (simp6431_0[1:1], comp2_0[3:3], comp2_0[4:4], comp2_0[5:5]);
  C3 I838 (simp6431_0[2:2], comp2_0[6:6], comp2_0[7:7], comp2_0[8:8]);
  C3 I839 (simp6431_0[3:3], comp2_0[9:9], comp2_0[10:10], comp2_0[11:11]);
  C3 I840 (simp6431_0[4:4], comp2_0[12:12], comp2_0[13:13], comp2_0[14:14]);
  C3 I841 (simp6431_0[5:5], comp2_0[15:15], comp2_0[16:16], comp2_0[17:17]);
  C3 I842 (simp6431_0[6:6], comp2_0[18:18], comp2_0[19:19], comp2_0[20:20]);
  C3 I843 (simp6431_0[7:7], comp2_0[21:21], comp2_0[22:22], comp2_0[23:23]);
  C3 I844 (simp6431_0[8:8], comp2_0[24:24], comp2_0[25:25], comp2_0[26:26]);
  C3 I845 (simp6431_0[9:9], comp2_0[27:27], comp2_0[28:28], comp2_0[29:29]);
  C2 I846 (simp6431_0[10:10], comp2_0[30:30], comp2_0[31:31]);
  C3 I847 (simp6432_0[0:0], simp6431_0[0:0], simp6431_0[1:1], simp6431_0[2:2]);
  C3 I848 (simp6432_0[1:1], simp6431_0[3:3], simp6431_0[4:4], simp6431_0[5:5]);
  C3 I849 (simp6432_0[2:2], simp6431_0[6:6], simp6431_0[7:7], simp6431_0[8:8]);
  C2 I850 (simp6432_0[3:3], simp6431_0[9:9], simp6431_0[10:10]);
  C3 I851 (simp6433_0[0:0], simp6432_0[0:0], simp6432_0[1:1], simp6432_0[2:2]);
  BUFF I852 (simp6433_0[1:1], simp6432_0[3:3]);
  C2 I853 (icomp_2, simp6433_0[0:0], simp6433_0[1:1]);
  OR2 I854 (comp3_0[0:0], i_3r0[0:0], i_3r1[0:0]);
  OR2 I855 (comp3_0[1:1], i_3r0[1:1], i_3r1[1:1]);
  OR2 I856 (comp3_0[2:2], i_3r0[2:2], i_3r1[2:2]);
  OR2 I857 (comp3_0[3:3], i_3r0[3:3], i_3r1[3:3]);
  OR2 I858 (comp3_0[4:4], i_3r0[4:4], i_3r1[4:4]);
  OR2 I859 (comp3_0[5:5], i_3r0[5:5], i_3r1[5:5]);
  OR2 I860 (comp3_0[6:6], i_3r0[6:6], i_3r1[6:6]);
  OR2 I861 (comp3_0[7:7], i_3r0[7:7], i_3r1[7:7]);
  OR2 I862 (comp3_0[8:8], i_3r0[8:8], i_3r1[8:8]);
  OR2 I863 (comp3_0[9:9], i_3r0[9:9], i_3r1[9:9]);
  OR2 I864 (comp3_0[10:10], i_3r0[10:10], i_3r1[10:10]);
  OR2 I865 (comp3_0[11:11], i_3r0[11:11], i_3r1[11:11]);
  OR2 I866 (comp3_0[12:12], i_3r0[12:12], i_3r1[12:12]);
  OR2 I867 (comp3_0[13:13], i_3r0[13:13], i_3r1[13:13]);
  OR2 I868 (comp3_0[14:14], i_3r0[14:14], i_3r1[14:14]);
  OR2 I869 (comp3_0[15:15], i_3r0[15:15], i_3r1[15:15]);
  OR2 I870 (comp3_0[16:16], i_3r0[16:16], i_3r1[16:16]);
  OR2 I871 (comp3_0[17:17], i_3r0[17:17], i_3r1[17:17]);
  OR2 I872 (comp3_0[18:18], i_3r0[18:18], i_3r1[18:18]);
  OR2 I873 (comp3_0[19:19], i_3r0[19:19], i_3r1[19:19]);
  OR2 I874 (comp3_0[20:20], i_3r0[20:20], i_3r1[20:20]);
  OR2 I875 (comp3_0[21:21], i_3r0[21:21], i_3r1[21:21]);
  OR2 I876 (comp3_0[22:22], i_3r0[22:22], i_3r1[22:22]);
  OR2 I877 (comp3_0[23:23], i_3r0[23:23], i_3r1[23:23]);
  OR2 I878 (comp3_0[24:24], i_3r0[24:24], i_3r1[24:24]);
  OR2 I879 (comp3_0[25:25], i_3r0[25:25], i_3r1[25:25]);
  OR2 I880 (comp3_0[26:26], i_3r0[26:26], i_3r1[26:26]);
  OR2 I881 (comp3_0[27:27], i_3r0[27:27], i_3r1[27:27]);
  OR2 I882 (comp3_0[28:28], i_3r0[28:28], i_3r1[28:28]);
  OR2 I883 (comp3_0[29:29], i_3r0[29:29], i_3r1[29:29]);
  OR2 I884 (comp3_0[30:30], i_3r0[30:30], i_3r1[30:30]);
  OR2 I885 (comp3_0[31:31], i_3r0[31:31], i_3r1[31:31]);
  C3 I886 (simp6771_0[0:0], comp3_0[0:0], comp3_0[1:1], comp3_0[2:2]);
  C3 I887 (simp6771_0[1:1], comp3_0[3:3], comp3_0[4:4], comp3_0[5:5]);
  C3 I888 (simp6771_0[2:2], comp3_0[6:6], comp3_0[7:7], comp3_0[8:8]);
  C3 I889 (simp6771_0[3:3], comp3_0[9:9], comp3_0[10:10], comp3_0[11:11]);
  C3 I890 (simp6771_0[4:4], comp3_0[12:12], comp3_0[13:13], comp3_0[14:14]);
  C3 I891 (simp6771_0[5:5], comp3_0[15:15], comp3_0[16:16], comp3_0[17:17]);
  C3 I892 (simp6771_0[6:6], comp3_0[18:18], comp3_0[19:19], comp3_0[20:20]);
  C3 I893 (simp6771_0[7:7], comp3_0[21:21], comp3_0[22:22], comp3_0[23:23]);
  C3 I894 (simp6771_0[8:8], comp3_0[24:24], comp3_0[25:25], comp3_0[26:26]);
  C3 I895 (simp6771_0[9:9], comp3_0[27:27], comp3_0[28:28], comp3_0[29:29]);
  C2 I896 (simp6771_0[10:10], comp3_0[30:30], comp3_0[31:31]);
  C3 I897 (simp6772_0[0:0], simp6771_0[0:0], simp6771_0[1:1], simp6771_0[2:2]);
  C3 I898 (simp6772_0[1:1], simp6771_0[3:3], simp6771_0[4:4], simp6771_0[5:5]);
  C3 I899 (simp6772_0[2:2], simp6771_0[6:6], simp6771_0[7:7], simp6771_0[8:8]);
  C2 I900 (simp6772_0[3:3], simp6771_0[9:9], simp6771_0[10:10]);
  C3 I901 (simp6773_0[0:0], simp6772_0[0:0], simp6772_0[1:1], simp6772_0[2:2]);
  BUFF I902 (simp6773_0[1:1], simp6772_0[3:3]);
  C2 I903 (icomp_3, simp6773_0[0:0], simp6773_0[1:1]);
  OR2 I904 (comp4_0[0:0], i_4r0[0:0], i_4r1[0:0]);
  OR2 I905 (comp4_0[1:1], i_4r0[1:1], i_4r1[1:1]);
  OR2 I906 (comp4_0[2:2], i_4r0[2:2], i_4r1[2:2]);
  OR2 I907 (comp4_0[3:3], i_4r0[3:3], i_4r1[3:3]);
  OR2 I908 (comp4_0[4:4], i_4r0[4:4], i_4r1[4:4]);
  OR2 I909 (comp4_0[5:5], i_4r0[5:5], i_4r1[5:5]);
  OR2 I910 (comp4_0[6:6], i_4r0[6:6], i_4r1[6:6]);
  OR2 I911 (comp4_0[7:7], i_4r0[7:7], i_4r1[7:7]);
  OR2 I912 (comp4_0[8:8], i_4r0[8:8], i_4r1[8:8]);
  OR2 I913 (comp4_0[9:9], i_4r0[9:9], i_4r1[9:9]);
  OR2 I914 (comp4_0[10:10], i_4r0[10:10], i_4r1[10:10]);
  OR2 I915 (comp4_0[11:11], i_4r0[11:11], i_4r1[11:11]);
  OR2 I916 (comp4_0[12:12], i_4r0[12:12], i_4r1[12:12]);
  OR2 I917 (comp4_0[13:13], i_4r0[13:13], i_4r1[13:13]);
  OR2 I918 (comp4_0[14:14], i_4r0[14:14], i_4r1[14:14]);
  OR2 I919 (comp4_0[15:15], i_4r0[15:15], i_4r1[15:15]);
  OR2 I920 (comp4_0[16:16], i_4r0[16:16], i_4r1[16:16]);
  OR2 I921 (comp4_0[17:17], i_4r0[17:17], i_4r1[17:17]);
  OR2 I922 (comp4_0[18:18], i_4r0[18:18], i_4r1[18:18]);
  OR2 I923 (comp4_0[19:19], i_4r0[19:19], i_4r1[19:19]);
  OR2 I924 (comp4_0[20:20], i_4r0[20:20], i_4r1[20:20]);
  OR2 I925 (comp4_0[21:21], i_4r0[21:21], i_4r1[21:21]);
  OR2 I926 (comp4_0[22:22], i_4r0[22:22], i_4r1[22:22]);
  OR2 I927 (comp4_0[23:23], i_4r0[23:23], i_4r1[23:23]);
  OR2 I928 (comp4_0[24:24], i_4r0[24:24], i_4r1[24:24]);
  OR2 I929 (comp4_0[25:25], i_4r0[25:25], i_4r1[25:25]);
  OR2 I930 (comp4_0[26:26], i_4r0[26:26], i_4r1[26:26]);
  OR2 I931 (comp4_0[27:27], i_4r0[27:27], i_4r1[27:27]);
  OR2 I932 (comp4_0[28:28], i_4r0[28:28], i_4r1[28:28]);
  OR2 I933 (comp4_0[29:29], i_4r0[29:29], i_4r1[29:29]);
  OR2 I934 (comp4_0[30:30], i_4r0[30:30], i_4r1[30:30]);
  OR2 I935 (comp4_0[31:31], i_4r0[31:31], i_4r1[31:31]);
  C3 I936 (simp7111_0[0:0], comp4_0[0:0], comp4_0[1:1], comp4_0[2:2]);
  C3 I937 (simp7111_0[1:1], comp4_0[3:3], comp4_0[4:4], comp4_0[5:5]);
  C3 I938 (simp7111_0[2:2], comp4_0[6:6], comp4_0[7:7], comp4_0[8:8]);
  C3 I939 (simp7111_0[3:3], comp4_0[9:9], comp4_0[10:10], comp4_0[11:11]);
  C3 I940 (simp7111_0[4:4], comp4_0[12:12], comp4_0[13:13], comp4_0[14:14]);
  C3 I941 (simp7111_0[5:5], comp4_0[15:15], comp4_0[16:16], comp4_0[17:17]);
  C3 I942 (simp7111_0[6:6], comp4_0[18:18], comp4_0[19:19], comp4_0[20:20]);
  C3 I943 (simp7111_0[7:7], comp4_0[21:21], comp4_0[22:22], comp4_0[23:23]);
  C3 I944 (simp7111_0[8:8], comp4_0[24:24], comp4_0[25:25], comp4_0[26:26]);
  C3 I945 (simp7111_0[9:9], comp4_0[27:27], comp4_0[28:28], comp4_0[29:29]);
  C2 I946 (simp7111_0[10:10], comp4_0[30:30], comp4_0[31:31]);
  C3 I947 (simp7112_0[0:0], simp7111_0[0:0], simp7111_0[1:1], simp7111_0[2:2]);
  C3 I948 (simp7112_0[1:1], simp7111_0[3:3], simp7111_0[4:4], simp7111_0[5:5]);
  C3 I949 (simp7112_0[2:2], simp7111_0[6:6], simp7111_0[7:7], simp7111_0[8:8]);
  C2 I950 (simp7112_0[3:3], simp7111_0[9:9], simp7111_0[10:10]);
  C3 I951 (simp7113_0[0:0], simp7112_0[0:0], simp7112_0[1:1], simp7112_0[2:2]);
  BUFF I952 (simp7113_0[1:1], simp7112_0[3:3]);
  C2 I953 (icomp_4, simp7113_0[0:0], simp7113_0[1:1]);
  OR2 I954 (comp5_0[0:0], i_5r0[0:0], i_5r1[0:0]);
  OR2 I955 (comp5_0[1:1], i_5r0[1:1], i_5r1[1:1]);
  OR2 I956 (comp5_0[2:2], i_5r0[2:2], i_5r1[2:2]);
  OR2 I957 (comp5_0[3:3], i_5r0[3:3], i_5r1[3:3]);
  OR2 I958 (comp5_0[4:4], i_5r0[4:4], i_5r1[4:4]);
  OR2 I959 (comp5_0[5:5], i_5r0[5:5], i_5r1[5:5]);
  OR2 I960 (comp5_0[6:6], i_5r0[6:6], i_5r1[6:6]);
  OR2 I961 (comp5_0[7:7], i_5r0[7:7], i_5r1[7:7]);
  OR2 I962 (comp5_0[8:8], i_5r0[8:8], i_5r1[8:8]);
  OR2 I963 (comp5_0[9:9], i_5r0[9:9], i_5r1[9:9]);
  OR2 I964 (comp5_0[10:10], i_5r0[10:10], i_5r1[10:10]);
  OR2 I965 (comp5_0[11:11], i_5r0[11:11], i_5r1[11:11]);
  OR2 I966 (comp5_0[12:12], i_5r0[12:12], i_5r1[12:12]);
  OR2 I967 (comp5_0[13:13], i_5r0[13:13], i_5r1[13:13]);
  OR2 I968 (comp5_0[14:14], i_5r0[14:14], i_5r1[14:14]);
  OR2 I969 (comp5_0[15:15], i_5r0[15:15], i_5r1[15:15]);
  OR2 I970 (comp5_0[16:16], i_5r0[16:16], i_5r1[16:16]);
  OR2 I971 (comp5_0[17:17], i_5r0[17:17], i_5r1[17:17]);
  OR2 I972 (comp5_0[18:18], i_5r0[18:18], i_5r1[18:18]);
  OR2 I973 (comp5_0[19:19], i_5r0[19:19], i_5r1[19:19]);
  OR2 I974 (comp5_0[20:20], i_5r0[20:20], i_5r1[20:20]);
  OR2 I975 (comp5_0[21:21], i_5r0[21:21], i_5r1[21:21]);
  OR2 I976 (comp5_0[22:22], i_5r0[22:22], i_5r1[22:22]);
  OR2 I977 (comp5_0[23:23], i_5r0[23:23], i_5r1[23:23]);
  OR2 I978 (comp5_0[24:24], i_5r0[24:24], i_5r1[24:24]);
  OR2 I979 (comp5_0[25:25], i_5r0[25:25], i_5r1[25:25]);
  OR2 I980 (comp5_0[26:26], i_5r0[26:26], i_5r1[26:26]);
  OR2 I981 (comp5_0[27:27], i_5r0[27:27], i_5r1[27:27]);
  OR2 I982 (comp5_0[28:28], i_5r0[28:28], i_5r1[28:28]);
  OR2 I983 (comp5_0[29:29], i_5r0[29:29], i_5r1[29:29]);
  OR2 I984 (comp5_0[30:30], i_5r0[30:30], i_5r1[30:30]);
  OR2 I985 (comp5_0[31:31], i_5r0[31:31], i_5r1[31:31]);
  C3 I986 (simp7451_0[0:0], comp5_0[0:0], comp5_0[1:1], comp5_0[2:2]);
  C3 I987 (simp7451_0[1:1], comp5_0[3:3], comp5_0[4:4], comp5_0[5:5]);
  C3 I988 (simp7451_0[2:2], comp5_0[6:6], comp5_0[7:7], comp5_0[8:8]);
  C3 I989 (simp7451_0[3:3], comp5_0[9:9], comp5_0[10:10], comp5_0[11:11]);
  C3 I990 (simp7451_0[4:4], comp5_0[12:12], comp5_0[13:13], comp5_0[14:14]);
  C3 I991 (simp7451_0[5:5], comp5_0[15:15], comp5_0[16:16], comp5_0[17:17]);
  C3 I992 (simp7451_0[6:6], comp5_0[18:18], comp5_0[19:19], comp5_0[20:20]);
  C3 I993 (simp7451_0[7:7], comp5_0[21:21], comp5_0[22:22], comp5_0[23:23]);
  C3 I994 (simp7451_0[8:8], comp5_0[24:24], comp5_0[25:25], comp5_0[26:26]);
  C3 I995 (simp7451_0[9:9], comp5_0[27:27], comp5_0[28:28], comp5_0[29:29]);
  C2 I996 (simp7451_0[10:10], comp5_0[30:30], comp5_0[31:31]);
  C3 I997 (simp7452_0[0:0], simp7451_0[0:0], simp7451_0[1:1], simp7451_0[2:2]);
  C3 I998 (simp7452_0[1:1], simp7451_0[3:3], simp7451_0[4:4], simp7451_0[5:5]);
  C3 I999 (simp7452_0[2:2], simp7451_0[6:6], simp7451_0[7:7], simp7451_0[8:8]);
  C2 I1000 (simp7452_0[3:3], simp7451_0[9:9], simp7451_0[10:10]);
  C3 I1001 (simp7453_0[0:0], simp7452_0[0:0], simp7452_0[1:1], simp7452_0[2:2]);
  BUFF I1002 (simp7453_0[1:1], simp7452_0[3:3]);
  C2 I1003 (icomp_5, simp7453_0[0:0], simp7453_0[1:1]);
  OR2 I1004 (comp6_0[0:0], i_6r0[0:0], i_6r1[0:0]);
  OR2 I1005 (comp6_0[1:1], i_6r0[1:1], i_6r1[1:1]);
  OR2 I1006 (comp6_0[2:2], i_6r0[2:2], i_6r1[2:2]);
  OR2 I1007 (comp6_0[3:3], i_6r0[3:3], i_6r1[3:3]);
  OR2 I1008 (comp6_0[4:4], i_6r0[4:4], i_6r1[4:4]);
  OR2 I1009 (comp6_0[5:5], i_6r0[5:5], i_6r1[5:5]);
  OR2 I1010 (comp6_0[6:6], i_6r0[6:6], i_6r1[6:6]);
  OR2 I1011 (comp6_0[7:7], i_6r0[7:7], i_6r1[7:7]);
  OR2 I1012 (comp6_0[8:8], i_6r0[8:8], i_6r1[8:8]);
  OR2 I1013 (comp6_0[9:9], i_6r0[9:9], i_6r1[9:9]);
  OR2 I1014 (comp6_0[10:10], i_6r0[10:10], i_6r1[10:10]);
  OR2 I1015 (comp6_0[11:11], i_6r0[11:11], i_6r1[11:11]);
  OR2 I1016 (comp6_0[12:12], i_6r0[12:12], i_6r1[12:12]);
  OR2 I1017 (comp6_0[13:13], i_6r0[13:13], i_6r1[13:13]);
  OR2 I1018 (comp6_0[14:14], i_6r0[14:14], i_6r1[14:14]);
  OR2 I1019 (comp6_0[15:15], i_6r0[15:15], i_6r1[15:15]);
  OR2 I1020 (comp6_0[16:16], i_6r0[16:16], i_6r1[16:16]);
  OR2 I1021 (comp6_0[17:17], i_6r0[17:17], i_6r1[17:17]);
  OR2 I1022 (comp6_0[18:18], i_6r0[18:18], i_6r1[18:18]);
  OR2 I1023 (comp6_0[19:19], i_6r0[19:19], i_6r1[19:19]);
  OR2 I1024 (comp6_0[20:20], i_6r0[20:20], i_6r1[20:20]);
  OR2 I1025 (comp6_0[21:21], i_6r0[21:21], i_6r1[21:21]);
  OR2 I1026 (comp6_0[22:22], i_6r0[22:22], i_6r1[22:22]);
  OR2 I1027 (comp6_0[23:23], i_6r0[23:23], i_6r1[23:23]);
  OR2 I1028 (comp6_0[24:24], i_6r0[24:24], i_6r1[24:24]);
  OR2 I1029 (comp6_0[25:25], i_6r0[25:25], i_6r1[25:25]);
  OR2 I1030 (comp6_0[26:26], i_6r0[26:26], i_6r1[26:26]);
  OR2 I1031 (comp6_0[27:27], i_6r0[27:27], i_6r1[27:27]);
  OR2 I1032 (comp6_0[28:28], i_6r0[28:28], i_6r1[28:28]);
  OR2 I1033 (comp6_0[29:29], i_6r0[29:29], i_6r1[29:29]);
  OR2 I1034 (comp6_0[30:30], i_6r0[30:30], i_6r1[30:30]);
  OR2 I1035 (comp6_0[31:31], i_6r0[31:31], i_6r1[31:31]);
  C3 I1036 (simp7791_0[0:0], comp6_0[0:0], comp6_0[1:1], comp6_0[2:2]);
  C3 I1037 (simp7791_0[1:1], comp6_0[3:3], comp6_0[4:4], comp6_0[5:5]);
  C3 I1038 (simp7791_0[2:2], comp6_0[6:6], comp6_0[7:7], comp6_0[8:8]);
  C3 I1039 (simp7791_0[3:3], comp6_0[9:9], comp6_0[10:10], comp6_0[11:11]);
  C3 I1040 (simp7791_0[4:4], comp6_0[12:12], comp6_0[13:13], comp6_0[14:14]);
  C3 I1041 (simp7791_0[5:5], comp6_0[15:15], comp6_0[16:16], comp6_0[17:17]);
  C3 I1042 (simp7791_0[6:6], comp6_0[18:18], comp6_0[19:19], comp6_0[20:20]);
  C3 I1043 (simp7791_0[7:7], comp6_0[21:21], comp6_0[22:22], comp6_0[23:23]);
  C3 I1044 (simp7791_0[8:8], comp6_0[24:24], comp6_0[25:25], comp6_0[26:26]);
  C3 I1045 (simp7791_0[9:9], comp6_0[27:27], comp6_0[28:28], comp6_0[29:29]);
  C2 I1046 (simp7791_0[10:10], comp6_0[30:30], comp6_0[31:31]);
  C3 I1047 (simp7792_0[0:0], simp7791_0[0:0], simp7791_0[1:1], simp7791_0[2:2]);
  C3 I1048 (simp7792_0[1:1], simp7791_0[3:3], simp7791_0[4:4], simp7791_0[5:5]);
  C3 I1049 (simp7792_0[2:2], simp7791_0[6:6], simp7791_0[7:7], simp7791_0[8:8]);
  C2 I1050 (simp7792_0[3:3], simp7791_0[9:9], simp7791_0[10:10]);
  C3 I1051 (simp7793_0[0:0], simp7792_0[0:0], simp7792_0[1:1], simp7792_0[2:2]);
  BUFF I1052 (simp7793_0[1:1], simp7792_0[3:3]);
  C2 I1053 (icomp_6, simp7793_0[0:0], simp7793_0[1:1]);
  C2R I1054 (choice_0, icomp_0, nchosen_0, reset);
  C2R I1055 (choice_1, icomp_1, nchosen_0, reset);
  C2R I1056 (choice_2, icomp_2, nchosen_0, reset);
  C2R I1057 (choice_3, icomp_3, nchosen_0, reset);
  C2R I1058 (choice_4, icomp_4, nchosen_0, reset);
  C2R I1059 (choice_5, icomp_5, nchosen_0, reset);
  C2R I1060 (choice_6, icomp_6, nchosen_0, reset);
  NOR3 I1061 (simp7871_0[0:0], choice_0, choice_1, choice_2);
  NOR3 I1062 (simp7871_0[1:1], choice_3, choice_4, choice_5);
  INV I1063 (simp7871_0[2:2], choice_6);
  NAND3 I1064 (anychoice_0, simp7871_0[0:0], simp7871_0[1:1], simp7871_0[2:2]);
  NOR2 I1065 (nchosen_0, anychoice_0, o_0a);
  C2R I1066 (i_0a, choice_0, o_0a, reset);
  C2R I1067 (i_1a, choice_1, o_0a, reset);
  C2R I1068 (i_2a, choice_2, o_0a, reset);
  C2R I1069 (i_3a, choice_3, o_0a, reset);
  C2R I1070 (i_4a, choice_4, o_0a, reset);
  C2R I1071 (i_5a, choice_5, o_0a, reset);
  C2R I1072 (i_6a, choice_6, o_0a, reset);
endmodule

// tkj4m3_1 TeakJ [Many [3,1],One 4]
module tkj4m3_1 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  input i_1r0;
  input i_1r1;
  output i_1a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [3:0] joinf_0;
  wire [3:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_1r0);
  BUFF I4 (joint_0[0:0], i_0r1[0:0]);
  BUFF I5 (joint_0[1:1], i_0r1[1:1]);
  BUFF I6 (joint_0[2:2], i_0r1[2:2]);
  BUFF I7 (joint_0[3:3], i_1r1);
  OR2 I8 (dcomplete_0, i_1r0, i_1r1);
  BUFF I9 (icomplete_0, dcomplete_0);
  C2 I10 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I11 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I12 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I13 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I14 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I15 (o_0r1[1:1], joint_0[1:1]);
  BUFF I16 (o_0r1[2:2], joint_0[2:2]);
  BUFF I17 (o_0r1[3:3], joint_0[3:3]);
  BUFF I18 (i_0a, o_0a);
  BUFF I19 (i_1a, o_0a);
endmodule

// tkf4mo0w3 TeakF [0] [One 4,Many [3]]
module tkf4mo0w3 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  wire ucomplete_0;
  wire comp_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (comp_0, i_0r0[3:3], i_0r1[3:3]);
  BUFF I2 (ucomplete_0, comp_0);
  C2 I3 (acomplete_0, ucomplete_0, icomplete_0);
  C2 I4 (o_0r0[0:0], i_0r0[0:0], icomplete_0);
  BUFF I5 (o_0r0[1:1], i_0r0[1:1]);
  BUFF I6 (o_0r0[2:2], i_0r0[2:2]);
  C2 I7 (o_0r1[0:0], i_0r1[0:0], icomplete_0);
  BUFF I8 (o_0r1[1:1], i_0r1[1:1]);
  BUFF I9 (o_0r1[2:2], i_0r1[2:2]);
  C2 I10 (i_0a, acomplete_0, o_0a);
endmodule

// tks3_o0w3_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0 TeakS (0+:3) [([Imp 0 0],0),([Imp 1 0],0),
//   ([Imp 2 0],0),([Imp 3 0],0),([Imp 4 0],0),([Imp 5 0],0),([Imp 6 0],0),([Imp 7 0],0)] [One 3,Many [0,
//   0,0,0,0,0,0,0]]
module tks3_o0w3_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, o_5r, o_5a, o_6r, o_6a, o_7r, o_7a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  output o_7r;
  input o_7a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire sel_4;
  wire sel_5;
  wire sel_6;
  wire sel_7;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire gsel_4;
  wire gsel_5;
  wire gsel_6;
  wire gsel_7;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire match2_0;
  wire match3_0;
  wire match4_0;
  wire match5_0;
  wire match6_0;
  wire match7_0;
  wire [2:0] comp_0;
  wire [2:0] simp631_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (match0_0, i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I2 (sel_1, match1_0);
  C3 I3 (match1_0, i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I4 (sel_2, match2_0);
  C3 I5 (match2_0, i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I6 (sel_3, match3_0);
  C3 I7 (match3_0, i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I8 (sel_4, match4_0);
  C3 I9 (match4_0, i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I10 (sel_5, match5_0);
  C3 I11 (match5_0, i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I12 (sel_6, match6_0);
  C3 I13 (match6_0, i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I14 (sel_7, match7_0);
  C3 I15 (match7_0, i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  C2 I16 (gsel_0, sel_0, icomplete_0);
  C2 I17 (gsel_1, sel_1, icomplete_0);
  C2 I18 (gsel_2, sel_2, icomplete_0);
  C2 I19 (gsel_3, sel_3, icomplete_0);
  C2 I20 (gsel_4, sel_4, icomplete_0);
  C2 I21 (gsel_5, sel_5, icomplete_0);
  C2 I22 (gsel_6, sel_6, icomplete_0);
  C2 I23 (gsel_7, sel_7, icomplete_0);
  OR2 I24 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I25 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I26 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I27 (icomplete_0, comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  BUFF I28 (o_0r, gsel_0);
  BUFF I29 (o_1r, gsel_1);
  BUFF I30 (o_2r, gsel_2);
  BUFF I31 (o_3r, gsel_3);
  BUFF I32 (o_4r, gsel_4);
  BUFF I33 (o_5r, gsel_5);
  BUFF I34 (o_6r, gsel_6);
  BUFF I35 (o_7r, gsel_7);
  NOR3 I36 (simp631_0[0:0], o_0a, o_1a, o_2a);
  NOR3 I37 (simp631_0[1:1], o_3a, o_4a, o_5a);
  NOR2 I38 (simp631_0[2:2], o_6a, o_7a);
  NAND3 I39 (oack_0, simp631_0[0:0], simp631_0[1:1], simp631_0[2:2]);
  C2 I40 (i_0a, oack_0, icomplete_0);
endmodule

// tkm8x32b TeakM [Many [32,32,32,32,32,32,32,32],One 32]
module tkm8x32b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, i_4r0, i_4r1, i_4a, i_5r0, i_5r1, i_5a, i_6r0, i_6r1, i_6a, i_7r0, i_7r1, i_7a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  input [31:0] i_2r0;
  input [31:0] i_2r1;
  output i_2a;
  input [31:0] i_3r0;
  input [31:0] i_3r1;
  output i_3a;
  input [31:0] i_4r0;
  input [31:0] i_4r1;
  output i_4a;
  input [31:0] i_5r0;
  input [31:0] i_5r1;
  output i_5a;
  input [31:0] i_6r0;
  input [31:0] i_6r1;
  output i_6a;
  input [31:0] i_7r0;
  input [31:0] i_7r1;
  output i_7a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire [31:0] gfint_0;
  wire [31:0] gfint_1;
  wire [31:0] gfint_2;
  wire [31:0] gfint_3;
  wire [31:0] gfint_4;
  wire [31:0] gfint_5;
  wire [31:0] gfint_6;
  wire [31:0] gfint_7;
  wire [31:0] gtint_0;
  wire [31:0] gtint_1;
  wire [31:0] gtint_2;
  wire [31:0] gtint_3;
  wire [31:0] gtint_4;
  wire [31:0] gtint_5;
  wire [31:0] gtint_6;
  wire [31:0] gtint_7;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire choice_4;
  wire choice_5;
  wire choice_6;
  wire choice_7;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire icomp_3;
  wire icomp_4;
  wire icomp_5;
  wire icomp_6;
  wire icomp_7;
  wire nchosen_0;
  wire [2:0] simp341_0;
  wire [2:0] simp351_0;
  wire [2:0] simp361_0;
  wire [2:0] simp371_0;
  wire [2:0] simp381_0;
  wire [2:0] simp391_0;
  wire [2:0] simp401_0;
  wire [2:0] simp411_0;
  wire [2:0] simp421_0;
  wire [2:0] simp431_0;
  wire [2:0] simp441_0;
  wire [2:0] simp451_0;
  wire [2:0] simp461_0;
  wire [2:0] simp471_0;
  wire [2:0] simp481_0;
  wire [2:0] simp491_0;
  wire [2:0] simp501_0;
  wire [2:0] simp511_0;
  wire [2:0] simp521_0;
  wire [2:0] simp531_0;
  wire [2:0] simp541_0;
  wire [2:0] simp551_0;
  wire [2:0] simp561_0;
  wire [2:0] simp571_0;
  wire [2:0] simp581_0;
  wire [2:0] simp591_0;
  wire [2:0] simp601_0;
  wire [2:0] simp611_0;
  wire [2:0] simp621_0;
  wire [2:0] simp631_0;
  wire [2:0] simp641_0;
  wire [2:0] simp651_0;
  wire [2:0] simp661_0;
  wire [2:0] simp671_0;
  wire [2:0] simp681_0;
  wire [2:0] simp691_0;
  wire [2:0] simp701_0;
  wire [2:0] simp711_0;
  wire [2:0] simp721_0;
  wire [2:0] simp731_0;
  wire [2:0] simp741_0;
  wire [2:0] simp751_0;
  wire [2:0] simp761_0;
  wire [2:0] simp771_0;
  wire [2:0] simp781_0;
  wire [2:0] simp791_0;
  wire [2:0] simp801_0;
  wire [2:0] simp811_0;
  wire [2:0] simp821_0;
  wire [2:0] simp831_0;
  wire [2:0] simp841_0;
  wire [2:0] simp851_0;
  wire [2:0] simp861_0;
  wire [2:0] simp871_0;
  wire [2:0] simp881_0;
  wire [2:0] simp891_0;
  wire [2:0] simp901_0;
  wire [2:0] simp911_0;
  wire [2:0] simp921_0;
  wire [2:0] simp931_0;
  wire [2:0] simp941_0;
  wire [2:0] simp951_0;
  wire [2:0] simp961_0;
  wire [2:0] simp971_0;
  wire [31:0] comp0_0;
  wire [10:0] simp6431_0;
  wire [3:0] simp6432_0;
  wire [1:0] simp6433_0;
  wire [31:0] comp1_0;
  wire [10:0] simp6771_0;
  wire [3:0] simp6772_0;
  wire [1:0] simp6773_0;
  wire [31:0] comp2_0;
  wire [10:0] simp7111_0;
  wire [3:0] simp7112_0;
  wire [1:0] simp7113_0;
  wire [31:0] comp3_0;
  wire [10:0] simp7451_0;
  wire [3:0] simp7452_0;
  wire [1:0] simp7453_0;
  wire [31:0] comp4_0;
  wire [10:0] simp7791_0;
  wire [3:0] simp7792_0;
  wire [1:0] simp7793_0;
  wire [31:0] comp5_0;
  wire [10:0] simp8131_0;
  wire [3:0] simp8132_0;
  wire [1:0] simp8133_0;
  wire [31:0] comp6_0;
  wire [10:0] simp8471_0;
  wire [3:0] simp8472_0;
  wire [1:0] simp8473_0;
  wire [31:0] comp7_0;
  wire [10:0] simp8811_0;
  wire [3:0] simp8812_0;
  wire [1:0] simp8813_0;
  wire [2:0] simp8901_0;
  NOR3 I0 (simp341_0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  NOR3 I1 (simp341_0[1:1], gfint_3[0:0], gfint_4[0:0], gfint_5[0:0]);
  NOR2 I2 (simp341_0[2:2], gfint_6[0:0], gfint_7[0:0]);
  NAND3 I3 (o_0r0[0:0], simp341_0[0:0], simp341_0[1:1], simp341_0[2:2]);
  NOR3 I4 (simp351_0[0:0], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  NOR3 I5 (simp351_0[1:1], gfint_3[1:1], gfint_4[1:1], gfint_5[1:1]);
  NOR2 I6 (simp351_0[2:2], gfint_6[1:1], gfint_7[1:1]);
  NAND3 I7 (o_0r0[1:1], simp351_0[0:0], simp351_0[1:1], simp351_0[2:2]);
  NOR3 I8 (simp361_0[0:0], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  NOR3 I9 (simp361_0[1:1], gfint_3[2:2], gfint_4[2:2], gfint_5[2:2]);
  NOR2 I10 (simp361_0[2:2], gfint_6[2:2], gfint_7[2:2]);
  NAND3 I11 (o_0r0[2:2], simp361_0[0:0], simp361_0[1:1], simp361_0[2:2]);
  NOR3 I12 (simp371_0[0:0], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  NOR3 I13 (simp371_0[1:1], gfint_3[3:3], gfint_4[3:3], gfint_5[3:3]);
  NOR2 I14 (simp371_0[2:2], gfint_6[3:3], gfint_7[3:3]);
  NAND3 I15 (o_0r0[3:3], simp371_0[0:0], simp371_0[1:1], simp371_0[2:2]);
  NOR3 I16 (simp381_0[0:0], gfint_0[4:4], gfint_1[4:4], gfint_2[4:4]);
  NOR3 I17 (simp381_0[1:1], gfint_3[4:4], gfint_4[4:4], gfint_5[4:4]);
  NOR2 I18 (simp381_0[2:2], gfint_6[4:4], gfint_7[4:4]);
  NAND3 I19 (o_0r0[4:4], simp381_0[0:0], simp381_0[1:1], simp381_0[2:2]);
  NOR3 I20 (simp391_0[0:0], gfint_0[5:5], gfint_1[5:5], gfint_2[5:5]);
  NOR3 I21 (simp391_0[1:1], gfint_3[5:5], gfint_4[5:5], gfint_5[5:5]);
  NOR2 I22 (simp391_0[2:2], gfint_6[5:5], gfint_7[5:5]);
  NAND3 I23 (o_0r0[5:5], simp391_0[0:0], simp391_0[1:1], simp391_0[2:2]);
  NOR3 I24 (simp401_0[0:0], gfint_0[6:6], gfint_1[6:6], gfint_2[6:6]);
  NOR3 I25 (simp401_0[1:1], gfint_3[6:6], gfint_4[6:6], gfint_5[6:6]);
  NOR2 I26 (simp401_0[2:2], gfint_6[6:6], gfint_7[6:6]);
  NAND3 I27 (o_0r0[6:6], simp401_0[0:0], simp401_0[1:1], simp401_0[2:2]);
  NOR3 I28 (simp411_0[0:0], gfint_0[7:7], gfint_1[7:7], gfint_2[7:7]);
  NOR3 I29 (simp411_0[1:1], gfint_3[7:7], gfint_4[7:7], gfint_5[7:7]);
  NOR2 I30 (simp411_0[2:2], gfint_6[7:7], gfint_7[7:7]);
  NAND3 I31 (o_0r0[7:7], simp411_0[0:0], simp411_0[1:1], simp411_0[2:2]);
  NOR3 I32 (simp421_0[0:0], gfint_0[8:8], gfint_1[8:8], gfint_2[8:8]);
  NOR3 I33 (simp421_0[1:1], gfint_3[8:8], gfint_4[8:8], gfint_5[8:8]);
  NOR2 I34 (simp421_0[2:2], gfint_6[8:8], gfint_7[8:8]);
  NAND3 I35 (o_0r0[8:8], simp421_0[0:0], simp421_0[1:1], simp421_0[2:2]);
  NOR3 I36 (simp431_0[0:0], gfint_0[9:9], gfint_1[9:9], gfint_2[9:9]);
  NOR3 I37 (simp431_0[1:1], gfint_3[9:9], gfint_4[9:9], gfint_5[9:9]);
  NOR2 I38 (simp431_0[2:2], gfint_6[9:9], gfint_7[9:9]);
  NAND3 I39 (o_0r0[9:9], simp431_0[0:0], simp431_0[1:1], simp431_0[2:2]);
  NOR3 I40 (simp441_0[0:0], gfint_0[10:10], gfint_1[10:10], gfint_2[10:10]);
  NOR3 I41 (simp441_0[1:1], gfint_3[10:10], gfint_4[10:10], gfint_5[10:10]);
  NOR2 I42 (simp441_0[2:2], gfint_6[10:10], gfint_7[10:10]);
  NAND3 I43 (o_0r0[10:10], simp441_0[0:0], simp441_0[1:1], simp441_0[2:2]);
  NOR3 I44 (simp451_0[0:0], gfint_0[11:11], gfint_1[11:11], gfint_2[11:11]);
  NOR3 I45 (simp451_0[1:1], gfint_3[11:11], gfint_4[11:11], gfint_5[11:11]);
  NOR2 I46 (simp451_0[2:2], gfint_6[11:11], gfint_7[11:11]);
  NAND3 I47 (o_0r0[11:11], simp451_0[0:0], simp451_0[1:1], simp451_0[2:2]);
  NOR3 I48 (simp461_0[0:0], gfint_0[12:12], gfint_1[12:12], gfint_2[12:12]);
  NOR3 I49 (simp461_0[1:1], gfint_3[12:12], gfint_4[12:12], gfint_5[12:12]);
  NOR2 I50 (simp461_0[2:2], gfint_6[12:12], gfint_7[12:12]);
  NAND3 I51 (o_0r0[12:12], simp461_0[0:0], simp461_0[1:1], simp461_0[2:2]);
  NOR3 I52 (simp471_0[0:0], gfint_0[13:13], gfint_1[13:13], gfint_2[13:13]);
  NOR3 I53 (simp471_0[1:1], gfint_3[13:13], gfint_4[13:13], gfint_5[13:13]);
  NOR2 I54 (simp471_0[2:2], gfint_6[13:13], gfint_7[13:13]);
  NAND3 I55 (o_0r0[13:13], simp471_0[0:0], simp471_0[1:1], simp471_0[2:2]);
  NOR3 I56 (simp481_0[0:0], gfint_0[14:14], gfint_1[14:14], gfint_2[14:14]);
  NOR3 I57 (simp481_0[1:1], gfint_3[14:14], gfint_4[14:14], gfint_5[14:14]);
  NOR2 I58 (simp481_0[2:2], gfint_6[14:14], gfint_7[14:14]);
  NAND3 I59 (o_0r0[14:14], simp481_0[0:0], simp481_0[1:1], simp481_0[2:2]);
  NOR3 I60 (simp491_0[0:0], gfint_0[15:15], gfint_1[15:15], gfint_2[15:15]);
  NOR3 I61 (simp491_0[1:1], gfint_3[15:15], gfint_4[15:15], gfint_5[15:15]);
  NOR2 I62 (simp491_0[2:2], gfint_6[15:15], gfint_7[15:15]);
  NAND3 I63 (o_0r0[15:15], simp491_0[0:0], simp491_0[1:1], simp491_0[2:2]);
  NOR3 I64 (simp501_0[0:0], gfint_0[16:16], gfint_1[16:16], gfint_2[16:16]);
  NOR3 I65 (simp501_0[1:1], gfint_3[16:16], gfint_4[16:16], gfint_5[16:16]);
  NOR2 I66 (simp501_0[2:2], gfint_6[16:16], gfint_7[16:16]);
  NAND3 I67 (o_0r0[16:16], simp501_0[0:0], simp501_0[1:1], simp501_0[2:2]);
  NOR3 I68 (simp511_0[0:0], gfint_0[17:17], gfint_1[17:17], gfint_2[17:17]);
  NOR3 I69 (simp511_0[1:1], gfint_3[17:17], gfint_4[17:17], gfint_5[17:17]);
  NOR2 I70 (simp511_0[2:2], gfint_6[17:17], gfint_7[17:17]);
  NAND3 I71 (o_0r0[17:17], simp511_0[0:0], simp511_0[1:1], simp511_0[2:2]);
  NOR3 I72 (simp521_0[0:0], gfint_0[18:18], gfint_1[18:18], gfint_2[18:18]);
  NOR3 I73 (simp521_0[1:1], gfint_3[18:18], gfint_4[18:18], gfint_5[18:18]);
  NOR2 I74 (simp521_0[2:2], gfint_6[18:18], gfint_7[18:18]);
  NAND3 I75 (o_0r0[18:18], simp521_0[0:0], simp521_0[1:1], simp521_0[2:2]);
  NOR3 I76 (simp531_0[0:0], gfint_0[19:19], gfint_1[19:19], gfint_2[19:19]);
  NOR3 I77 (simp531_0[1:1], gfint_3[19:19], gfint_4[19:19], gfint_5[19:19]);
  NOR2 I78 (simp531_0[2:2], gfint_6[19:19], gfint_7[19:19]);
  NAND3 I79 (o_0r0[19:19], simp531_0[0:0], simp531_0[1:1], simp531_0[2:2]);
  NOR3 I80 (simp541_0[0:0], gfint_0[20:20], gfint_1[20:20], gfint_2[20:20]);
  NOR3 I81 (simp541_0[1:1], gfint_3[20:20], gfint_4[20:20], gfint_5[20:20]);
  NOR2 I82 (simp541_0[2:2], gfint_6[20:20], gfint_7[20:20]);
  NAND3 I83 (o_0r0[20:20], simp541_0[0:0], simp541_0[1:1], simp541_0[2:2]);
  NOR3 I84 (simp551_0[0:0], gfint_0[21:21], gfint_1[21:21], gfint_2[21:21]);
  NOR3 I85 (simp551_0[1:1], gfint_3[21:21], gfint_4[21:21], gfint_5[21:21]);
  NOR2 I86 (simp551_0[2:2], gfint_6[21:21], gfint_7[21:21]);
  NAND3 I87 (o_0r0[21:21], simp551_0[0:0], simp551_0[1:1], simp551_0[2:2]);
  NOR3 I88 (simp561_0[0:0], gfint_0[22:22], gfint_1[22:22], gfint_2[22:22]);
  NOR3 I89 (simp561_0[1:1], gfint_3[22:22], gfint_4[22:22], gfint_5[22:22]);
  NOR2 I90 (simp561_0[2:2], gfint_6[22:22], gfint_7[22:22]);
  NAND3 I91 (o_0r0[22:22], simp561_0[0:0], simp561_0[1:1], simp561_0[2:2]);
  NOR3 I92 (simp571_0[0:0], gfint_0[23:23], gfint_1[23:23], gfint_2[23:23]);
  NOR3 I93 (simp571_0[1:1], gfint_3[23:23], gfint_4[23:23], gfint_5[23:23]);
  NOR2 I94 (simp571_0[2:2], gfint_6[23:23], gfint_7[23:23]);
  NAND3 I95 (o_0r0[23:23], simp571_0[0:0], simp571_0[1:1], simp571_0[2:2]);
  NOR3 I96 (simp581_0[0:0], gfint_0[24:24], gfint_1[24:24], gfint_2[24:24]);
  NOR3 I97 (simp581_0[1:1], gfint_3[24:24], gfint_4[24:24], gfint_5[24:24]);
  NOR2 I98 (simp581_0[2:2], gfint_6[24:24], gfint_7[24:24]);
  NAND3 I99 (o_0r0[24:24], simp581_0[0:0], simp581_0[1:1], simp581_0[2:2]);
  NOR3 I100 (simp591_0[0:0], gfint_0[25:25], gfint_1[25:25], gfint_2[25:25]);
  NOR3 I101 (simp591_0[1:1], gfint_3[25:25], gfint_4[25:25], gfint_5[25:25]);
  NOR2 I102 (simp591_0[2:2], gfint_6[25:25], gfint_7[25:25]);
  NAND3 I103 (o_0r0[25:25], simp591_0[0:0], simp591_0[1:1], simp591_0[2:2]);
  NOR3 I104 (simp601_0[0:0], gfint_0[26:26], gfint_1[26:26], gfint_2[26:26]);
  NOR3 I105 (simp601_0[1:1], gfint_3[26:26], gfint_4[26:26], gfint_5[26:26]);
  NOR2 I106 (simp601_0[2:2], gfint_6[26:26], gfint_7[26:26]);
  NAND3 I107 (o_0r0[26:26], simp601_0[0:0], simp601_0[1:1], simp601_0[2:2]);
  NOR3 I108 (simp611_0[0:0], gfint_0[27:27], gfint_1[27:27], gfint_2[27:27]);
  NOR3 I109 (simp611_0[1:1], gfint_3[27:27], gfint_4[27:27], gfint_5[27:27]);
  NOR2 I110 (simp611_0[2:2], gfint_6[27:27], gfint_7[27:27]);
  NAND3 I111 (o_0r0[27:27], simp611_0[0:0], simp611_0[1:1], simp611_0[2:2]);
  NOR3 I112 (simp621_0[0:0], gfint_0[28:28], gfint_1[28:28], gfint_2[28:28]);
  NOR3 I113 (simp621_0[1:1], gfint_3[28:28], gfint_4[28:28], gfint_5[28:28]);
  NOR2 I114 (simp621_0[2:2], gfint_6[28:28], gfint_7[28:28]);
  NAND3 I115 (o_0r0[28:28], simp621_0[0:0], simp621_0[1:1], simp621_0[2:2]);
  NOR3 I116 (simp631_0[0:0], gfint_0[29:29], gfint_1[29:29], gfint_2[29:29]);
  NOR3 I117 (simp631_0[1:1], gfint_3[29:29], gfint_4[29:29], gfint_5[29:29]);
  NOR2 I118 (simp631_0[2:2], gfint_6[29:29], gfint_7[29:29]);
  NAND3 I119 (o_0r0[29:29], simp631_0[0:0], simp631_0[1:1], simp631_0[2:2]);
  NOR3 I120 (simp641_0[0:0], gfint_0[30:30], gfint_1[30:30], gfint_2[30:30]);
  NOR3 I121 (simp641_0[1:1], gfint_3[30:30], gfint_4[30:30], gfint_5[30:30]);
  NOR2 I122 (simp641_0[2:2], gfint_6[30:30], gfint_7[30:30]);
  NAND3 I123 (o_0r0[30:30], simp641_0[0:0], simp641_0[1:1], simp641_0[2:2]);
  NOR3 I124 (simp651_0[0:0], gfint_0[31:31], gfint_1[31:31], gfint_2[31:31]);
  NOR3 I125 (simp651_0[1:1], gfint_3[31:31], gfint_4[31:31], gfint_5[31:31]);
  NOR2 I126 (simp651_0[2:2], gfint_6[31:31], gfint_7[31:31]);
  NAND3 I127 (o_0r0[31:31], simp651_0[0:0], simp651_0[1:1], simp651_0[2:2]);
  NOR3 I128 (simp661_0[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  NOR3 I129 (simp661_0[1:1], gtint_3[0:0], gtint_4[0:0], gtint_5[0:0]);
  NOR2 I130 (simp661_0[2:2], gtint_6[0:0], gtint_7[0:0]);
  NAND3 I131 (o_0r1[0:0], simp661_0[0:0], simp661_0[1:1], simp661_0[2:2]);
  NOR3 I132 (simp671_0[0:0], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  NOR3 I133 (simp671_0[1:1], gtint_3[1:1], gtint_4[1:1], gtint_5[1:1]);
  NOR2 I134 (simp671_0[2:2], gtint_6[1:1], gtint_7[1:1]);
  NAND3 I135 (o_0r1[1:1], simp671_0[0:0], simp671_0[1:1], simp671_0[2:2]);
  NOR3 I136 (simp681_0[0:0], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  NOR3 I137 (simp681_0[1:1], gtint_3[2:2], gtint_4[2:2], gtint_5[2:2]);
  NOR2 I138 (simp681_0[2:2], gtint_6[2:2], gtint_7[2:2]);
  NAND3 I139 (o_0r1[2:2], simp681_0[0:0], simp681_0[1:1], simp681_0[2:2]);
  NOR3 I140 (simp691_0[0:0], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  NOR3 I141 (simp691_0[1:1], gtint_3[3:3], gtint_4[3:3], gtint_5[3:3]);
  NOR2 I142 (simp691_0[2:2], gtint_6[3:3], gtint_7[3:3]);
  NAND3 I143 (o_0r1[3:3], simp691_0[0:0], simp691_0[1:1], simp691_0[2:2]);
  NOR3 I144 (simp701_0[0:0], gtint_0[4:4], gtint_1[4:4], gtint_2[4:4]);
  NOR3 I145 (simp701_0[1:1], gtint_3[4:4], gtint_4[4:4], gtint_5[4:4]);
  NOR2 I146 (simp701_0[2:2], gtint_6[4:4], gtint_7[4:4]);
  NAND3 I147 (o_0r1[4:4], simp701_0[0:0], simp701_0[1:1], simp701_0[2:2]);
  NOR3 I148 (simp711_0[0:0], gtint_0[5:5], gtint_1[5:5], gtint_2[5:5]);
  NOR3 I149 (simp711_0[1:1], gtint_3[5:5], gtint_4[5:5], gtint_5[5:5]);
  NOR2 I150 (simp711_0[2:2], gtint_6[5:5], gtint_7[5:5]);
  NAND3 I151 (o_0r1[5:5], simp711_0[0:0], simp711_0[1:1], simp711_0[2:2]);
  NOR3 I152 (simp721_0[0:0], gtint_0[6:6], gtint_1[6:6], gtint_2[6:6]);
  NOR3 I153 (simp721_0[1:1], gtint_3[6:6], gtint_4[6:6], gtint_5[6:6]);
  NOR2 I154 (simp721_0[2:2], gtint_6[6:6], gtint_7[6:6]);
  NAND3 I155 (o_0r1[6:6], simp721_0[0:0], simp721_0[1:1], simp721_0[2:2]);
  NOR3 I156 (simp731_0[0:0], gtint_0[7:7], gtint_1[7:7], gtint_2[7:7]);
  NOR3 I157 (simp731_0[1:1], gtint_3[7:7], gtint_4[7:7], gtint_5[7:7]);
  NOR2 I158 (simp731_0[2:2], gtint_6[7:7], gtint_7[7:7]);
  NAND3 I159 (o_0r1[7:7], simp731_0[0:0], simp731_0[1:1], simp731_0[2:2]);
  NOR3 I160 (simp741_0[0:0], gtint_0[8:8], gtint_1[8:8], gtint_2[8:8]);
  NOR3 I161 (simp741_0[1:1], gtint_3[8:8], gtint_4[8:8], gtint_5[8:8]);
  NOR2 I162 (simp741_0[2:2], gtint_6[8:8], gtint_7[8:8]);
  NAND3 I163 (o_0r1[8:8], simp741_0[0:0], simp741_0[1:1], simp741_0[2:2]);
  NOR3 I164 (simp751_0[0:0], gtint_0[9:9], gtint_1[9:9], gtint_2[9:9]);
  NOR3 I165 (simp751_0[1:1], gtint_3[9:9], gtint_4[9:9], gtint_5[9:9]);
  NOR2 I166 (simp751_0[2:2], gtint_6[9:9], gtint_7[9:9]);
  NAND3 I167 (o_0r1[9:9], simp751_0[0:0], simp751_0[1:1], simp751_0[2:2]);
  NOR3 I168 (simp761_0[0:0], gtint_0[10:10], gtint_1[10:10], gtint_2[10:10]);
  NOR3 I169 (simp761_0[1:1], gtint_3[10:10], gtint_4[10:10], gtint_5[10:10]);
  NOR2 I170 (simp761_0[2:2], gtint_6[10:10], gtint_7[10:10]);
  NAND3 I171 (o_0r1[10:10], simp761_0[0:0], simp761_0[1:1], simp761_0[2:2]);
  NOR3 I172 (simp771_0[0:0], gtint_0[11:11], gtint_1[11:11], gtint_2[11:11]);
  NOR3 I173 (simp771_0[1:1], gtint_3[11:11], gtint_4[11:11], gtint_5[11:11]);
  NOR2 I174 (simp771_0[2:2], gtint_6[11:11], gtint_7[11:11]);
  NAND3 I175 (o_0r1[11:11], simp771_0[0:0], simp771_0[1:1], simp771_0[2:2]);
  NOR3 I176 (simp781_0[0:0], gtint_0[12:12], gtint_1[12:12], gtint_2[12:12]);
  NOR3 I177 (simp781_0[1:1], gtint_3[12:12], gtint_4[12:12], gtint_5[12:12]);
  NOR2 I178 (simp781_0[2:2], gtint_6[12:12], gtint_7[12:12]);
  NAND3 I179 (o_0r1[12:12], simp781_0[0:0], simp781_0[1:1], simp781_0[2:2]);
  NOR3 I180 (simp791_0[0:0], gtint_0[13:13], gtint_1[13:13], gtint_2[13:13]);
  NOR3 I181 (simp791_0[1:1], gtint_3[13:13], gtint_4[13:13], gtint_5[13:13]);
  NOR2 I182 (simp791_0[2:2], gtint_6[13:13], gtint_7[13:13]);
  NAND3 I183 (o_0r1[13:13], simp791_0[0:0], simp791_0[1:1], simp791_0[2:2]);
  NOR3 I184 (simp801_0[0:0], gtint_0[14:14], gtint_1[14:14], gtint_2[14:14]);
  NOR3 I185 (simp801_0[1:1], gtint_3[14:14], gtint_4[14:14], gtint_5[14:14]);
  NOR2 I186 (simp801_0[2:2], gtint_6[14:14], gtint_7[14:14]);
  NAND3 I187 (o_0r1[14:14], simp801_0[0:0], simp801_0[1:1], simp801_0[2:2]);
  NOR3 I188 (simp811_0[0:0], gtint_0[15:15], gtint_1[15:15], gtint_2[15:15]);
  NOR3 I189 (simp811_0[1:1], gtint_3[15:15], gtint_4[15:15], gtint_5[15:15]);
  NOR2 I190 (simp811_0[2:2], gtint_6[15:15], gtint_7[15:15]);
  NAND3 I191 (o_0r1[15:15], simp811_0[0:0], simp811_0[1:1], simp811_0[2:2]);
  NOR3 I192 (simp821_0[0:0], gtint_0[16:16], gtint_1[16:16], gtint_2[16:16]);
  NOR3 I193 (simp821_0[1:1], gtint_3[16:16], gtint_4[16:16], gtint_5[16:16]);
  NOR2 I194 (simp821_0[2:2], gtint_6[16:16], gtint_7[16:16]);
  NAND3 I195 (o_0r1[16:16], simp821_0[0:0], simp821_0[1:1], simp821_0[2:2]);
  NOR3 I196 (simp831_0[0:0], gtint_0[17:17], gtint_1[17:17], gtint_2[17:17]);
  NOR3 I197 (simp831_0[1:1], gtint_3[17:17], gtint_4[17:17], gtint_5[17:17]);
  NOR2 I198 (simp831_0[2:2], gtint_6[17:17], gtint_7[17:17]);
  NAND3 I199 (o_0r1[17:17], simp831_0[0:0], simp831_0[1:1], simp831_0[2:2]);
  NOR3 I200 (simp841_0[0:0], gtint_0[18:18], gtint_1[18:18], gtint_2[18:18]);
  NOR3 I201 (simp841_0[1:1], gtint_3[18:18], gtint_4[18:18], gtint_5[18:18]);
  NOR2 I202 (simp841_0[2:2], gtint_6[18:18], gtint_7[18:18]);
  NAND3 I203 (o_0r1[18:18], simp841_0[0:0], simp841_0[1:1], simp841_0[2:2]);
  NOR3 I204 (simp851_0[0:0], gtint_0[19:19], gtint_1[19:19], gtint_2[19:19]);
  NOR3 I205 (simp851_0[1:1], gtint_3[19:19], gtint_4[19:19], gtint_5[19:19]);
  NOR2 I206 (simp851_0[2:2], gtint_6[19:19], gtint_7[19:19]);
  NAND3 I207 (o_0r1[19:19], simp851_0[0:0], simp851_0[1:1], simp851_0[2:2]);
  NOR3 I208 (simp861_0[0:0], gtint_0[20:20], gtint_1[20:20], gtint_2[20:20]);
  NOR3 I209 (simp861_0[1:1], gtint_3[20:20], gtint_4[20:20], gtint_5[20:20]);
  NOR2 I210 (simp861_0[2:2], gtint_6[20:20], gtint_7[20:20]);
  NAND3 I211 (o_0r1[20:20], simp861_0[0:0], simp861_0[1:1], simp861_0[2:2]);
  NOR3 I212 (simp871_0[0:0], gtint_0[21:21], gtint_1[21:21], gtint_2[21:21]);
  NOR3 I213 (simp871_0[1:1], gtint_3[21:21], gtint_4[21:21], gtint_5[21:21]);
  NOR2 I214 (simp871_0[2:2], gtint_6[21:21], gtint_7[21:21]);
  NAND3 I215 (o_0r1[21:21], simp871_0[0:0], simp871_0[1:1], simp871_0[2:2]);
  NOR3 I216 (simp881_0[0:0], gtint_0[22:22], gtint_1[22:22], gtint_2[22:22]);
  NOR3 I217 (simp881_0[1:1], gtint_3[22:22], gtint_4[22:22], gtint_5[22:22]);
  NOR2 I218 (simp881_0[2:2], gtint_6[22:22], gtint_7[22:22]);
  NAND3 I219 (o_0r1[22:22], simp881_0[0:0], simp881_0[1:1], simp881_0[2:2]);
  NOR3 I220 (simp891_0[0:0], gtint_0[23:23], gtint_1[23:23], gtint_2[23:23]);
  NOR3 I221 (simp891_0[1:1], gtint_3[23:23], gtint_4[23:23], gtint_5[23:23]);
  NOR2 I222 (simp891_0[2:2], gtint_6[23:23], gtint_7[23:23]);
  NAND3 I223 (o_0r1[23:23], simp891_0[0:0], simp891_0[1:1], simp891_0[2:2]);
  NOR3 I224 (simp901_0[0:0], gtint_0[24:24], gtint_1[24:24], gtint_2[24:24]);
  NOR3 I225 (simp901_0[1:1], gtint_3[24:24], gtint_4[24:24], gtint_5[24:24]);
  NOR2 I226 (simp901_0[2:2], gtint_6[24:24], gtint_7[24:24]);
  NAND3 I227 (o_0r1[24:24], simp901_0[0:0], simp901_0[1:1], simp901_0[2:2]);
  NOR3 I228 (simp911_0[0:0], gtint_0[25:25], gtint_1[25:25], gtint_2[25:25]);
  NOR3 I229 (simp911_0[1:1], gtint_3[25:25], gtint_4[25:25], gtint_5[25:25]);
  NOR2 I230 (simp911_0[2:2], gtint_6[25:25], gtint_7[25:25]);
  NAND3 I231 (o_0r1[25:25], simp911_0[0:0], simp911_0[1:1], simp911_0[2:2]);
  NOR3 I232 (simp921_0[0:0], gtint_0[26:26], gtint_1[26:26], gtint_2[26:26]);
  NOR3 I233 (simp921_0[1:1], gtint_3[26:26], gtint_4[26:26], gtint_5[26:26]);
  NOR2 I234 (simp921_0[2:2], gtint_6[26:26], gtint_7[26:26]);
  NAND3 I235 (o_0r1[26:26], simp921_0[0:0], simp921_0[1:1], simp921_0[2:2]);
  NOR3 I236 (simp931_0[0:0], gtint_0[27:27], gtint_1[27:27], gtint_2[27:27]);
  NOR3 I237 (simp931_0[1:1], gtint_3[27:27], gtint_4[27:27], gtint_5[27:27]);
  NOR2 I238 (simp931_0[2:2], gtint_6[27:27], gtint_7[27:27]);
  NAND3 I239 (o_0r1[27:27], simp931_0[0:0], simp931_0[1:1], simp931_0[2:2]);
  NOR3 I240 (simp941_0[0:0], gtint_0[28:28], gtint_1[28:28], gtint_2[28:28]);
  NOR3 I241 (simp941_0[1:1], gtint_3[28:28], gtint_4[28:28], gtint_5[28:28]);
  NOR2 I242 (simp941_0[2:2], gtint_6[28:28], gtint_7[28:28]);
  NAND3 I243 (o_0r1[28:28], simp941_0[0:0], simp941_0[1:1], simp941_0[2:2]);
  NOR3 I244 (simp951_0[0:0], gtint_0[29:29], gtint_1[29:29], gtint_2[29:29]);
  NOR3 I245 (simp951_0[1:1], gtint_3[29:29], gtint_4[29:29], gtint_5[29:29]);
  NOR2 I246 (simp951_0[2:2], gtint_6[29:29], gtint_7[29:29]);
  NAND3 I247 (o_0r1[29:29], simp951_0[0:0], simp951_0[1:1], simp951_0[2:2]);
  NOR3 I248 (simp961_0[0:0], gtint_0[30:30], gtint_1[30:30], gtint_2[30:30]);
  NOR3 I249 (simp961_0[1:1], gtint_3[30:30], gtint_4[30:30], gtint_5[30:30]);
  NOR2 I250 (simp961_0[2:2], gtint_6[30:30], gtint_7[30:30]);
  NAND3 I251 (o_0r1[30:30], simp961_0[0:0], simp961_0[1:1], simp961_0[2:2]);
  NOR3 I252 (simp971_0[0:0], gtint_0[31:31], gtint_1[31:31], gtint_2[31:31]);
  NOR3 I253 (simp971_0[1:1], gtint_3[31:31], gtint_4[31:31], gtint_5[31:31]);
  NOR2 I254 (simp971_0[2:2], gtint_6[31:31], gtint_7[31:31]);
  NAND3 I255 (o_0r1[31:31], simp971_0[0:0], simp971_0[1:1], simp971_0[2:2]);
  AND2 I256 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I257 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I258 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I259 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I260 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I261 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I262 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I263 (gtint_0[7:7], choice_0, i_0r1[7:7]);
  AND2 I264 (gtint_0[8:8], choice_0, i_0r1[8:8]);
  AND2 I265 (gtint_0[9:9], choice_0, i_0r1[9:9]);
  AND2 I266 (gtint_0[10:10], choice_0, i_0r1[10:10]);
  AND2 I267 (gtint_0[11:11], choice_0, i_0r1[11:11]);
  AND2 I268 (gtint_0[12:12], choice_0, i_0r1[12:12]);
  AND2 I269 (gtint_0[13:13], choice_0, i_0r1[13:13]);
  AND2 I270 (gtint_0[14:14], choice_0, i_0r1[14:14]);
  AND2 I271 (gtint_0[15:15], choice_0, i_0r1[15:15]);
  AND2 I272 (gtint_0[16:16], choice_0, i_0r1[16:16]);
  AND2 I273 (gtint_0[17:17], choice_0, i_0r1[17:17]);
  AND2 I274 (gtint_0[18:18], choice_0, i_0r1[18:18]);
  AND2 I275 (gtint_0[19:19], choice_0, i_0r1[19:19]);
  AND2 I276 (gtint_0[20:20], choice_0, i_0r1[20:20]);
  AND2 I277 (gtint_0[21:21], choice_0, i_0r1[21:21]);
  AND2 I278 (gtint_0[22:22], choice_0, i_0r1[22:22]);
  AND2 I279 (gtint_0[23:23], choice_0, i_0r1[23:23]);
  AND2 I280 (gtint_0[24:24], choice_0, i_0r1[24:24]);
  AND2 I281 (gtint_0[25:25], choice_0, i_0r1[25:25]);
  AND2 I282 (gtint_0[26:26], choice_0, i_0r1[26:26]);
  AND2 I283 (gtint_0[27:27], choice_0, i_0r1[27:27]);
  AND2 I284 (gtint_0[28:28], choice_0, i_0r1[28:28]);
  AND2 I285 (gtint_0[29:29], choice_0, i_0r1[29:29]);
  AND2 I286 (gtint_0[30:30], choice_0, i_0r1[30:30]);
  AND2 I287 (gtint_0[31:31], choice_0, i_0r1[31:31]);
  AND2 I288 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I289 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I290 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I291 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I292 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I293 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I294 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I295 (gtint_1[7:7], choice_1, i_1r1[7:7]);
  AND2 I296 (gtint_1[8:8], choice_1, i_1r1[8:8]);
  AND2 I297 (gtint_1[9:9], choice_1, i_1r1[9:9]);
  AND2 I298 (gtint_1[10:10], choice_1, i_1r1[10:10]);
  AND2 I299 (gtint_1[11:11], choice_1, i_1r1[11:11]);
  AND2 I300 (gtint_1[12:12], choice_1, i_1r1[12:12]);
  AND2 I301 (gtint_1[13:13], choice_1, i_1r1[13:13]);
  AND2 I302 (gtint_1[14:14], choice_1, i_1r1[14:14]);
  AND2 I303 (gtint_1[15:15], choice_1, i_1r1[15:15]);
  AND2 I304 (gtint_1[16:16], choice_1, i_1r1[16:16]);
  AND2 I305 (gtint_1[17:17], choice_1, i_1r1[17:17]);
  AND2 I306 (gtint_1[18:18], choice_1, i_1r1[18:18]);
  AND2 I307 (gtint_1[19:19], choice_1, i_1r1[19:19]);
  AND2 I308 (gtint_1[20:20], choice_1, i_1r1[20:20]);
  AND2 I309 (gtint_1[21:21], choice_1, i_1r1[21:21]);
  AND2 I310 (gtint_1[22:22], choice_1, i_1r1[22:22]);
  AND2 I311 (gtint_1[23:23], choice_1, i_1r1[23:23]);
  AND2 I312 (gtint_1[24:24], choice_1, i_1r1[24:24]);
  AND2 I313 (gtint_1[25:25], choice_1, i_1r1[25:25]);
  AND2 I314 (gtint_1[26:26], choice_1, i_1r1[26:26]);
  AND2 I315 (gtint_1[27:27], choice_1, i_1r1[27:27]);
  AND2 I316 (gtint_1[28:28], choice_1, i_1r1[28:28]);
  AND2 I317 (gtint_1[29:29], choice_1, i_1r1[29:29]);
  AND2 I318 (gtint_1[30:30], choice_1, i_1r1[30:30]);
  AND2 I319 (gtint_1[31:31], choice_1, i_1r1[31:31]);
  AND2 I320 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I321 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I322 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I323 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AND2 I324 (gtint_2[4:4], choice_2, i_2r1[4:4]);
  AND2 I325 (gtint_2[5:5], choice_2, i_2r1[5:5]);
  AND2 I326 (gtint_2[6:6], choice_2, i_2r1[6:6]);
  AND2 I327 (gtint_2[7:7], choice_2, i_2r1[7:7]);
  AND2 I328 (gtint_2[8:8], choice_2, i_2r1[8:8]);
  AND2 I329 (gtint_2[9:9], choice_2, i_2r1[9:9]);
  AND2 I330 (gtint_2[10:10], choice_2, i_2r1[10:10]);
  AND2 I331 (gtint_2[11:11], choice_2, i_2r1[11:11]);
  AND2 I332 (gtint_2[12:12], choice_2, i_2r1[12:12]);
  AND2 I333 (gtint_2[13:13], choice_2, i_2r1[13:13]);
  AND2 I334 (gtint_2[14:14], choice_2, i_2r1[14:14]);
  AND2 I335 (gtint_2[15:15], choice_2, i_2r1[15:15]);
  AND2 I336 (gtint_2[16:16], choice_2, i_2r1[16:16]);
  AND2 I337 (gtint_2[17:17], choice_2, i_2r1[17:17]);
  AND2 I338 (gtint_2[18:18], choice_2, i_2r1[18:18]);
  AND2 I339 (gtint_2[19:19], choice_2, i_2r1[19:19]);
  AND2 I340 (gtint_2[20:20], choice_2, i_2r1[20:20]);
  AND2 I341 (gtint_2[21:21], choice_2, i_2r1[21:21]);
  AND2 I342 (gtint_2[22:22], choice_2, i_2r1[22:22]);
  AND2 I343 (gtint_2[23:23], choice_2, i_2r1[23:23]);
  AND2 I344 (gtint_2[24:24], choice_2, i_2r1[24:24]);
  AND2 I345 (gtint_2[25:25], choice_2, i_2r1[25:25]);
  AND2 I346 (gtint_2[26:26], choice_2, i_2r1[26:26]);
  AND2 I347 (gtint_2[27:27], choice_2, i_2r1[27:27]);
  AND2 I348 (gtint_2[28:28], choice_2, i_2r1[28:28]);
  AND2 I349 (gtint_2[29:29], choice_2, i_2r1[29:29]);
  AND2 I350 (gtint_2[30:30], choice_2, i_2r1[30:30]);
  AND2 I351 (gtint_2[31:31], choice_2, i_2r1[31:31]);
  AND2 I352 (gtint_3[0:0], choice_3, i_3r1[0:0]);
  AND2 I353 (gtint_3[1:1], choice_3, i_3r1[1:1]);
  AND2 I354 (gtint_3[2:2], choice_3, i_3r1[2:2]);
  AND2 I355 (gtint_3[3:3], choice_3, i_3r1[3:3]);
  AND2 I356 (gtint_3[4:4], choice_3, i_3r1[4:4]);
  AND2 I357 (gtint_3[5:5], choice_3, i_3r1[5:5]);
  AND2 I358 (gtint_3[6:6], choice_3, i_3r1[6:6]);
  AND2 I359 (gtint_3[7:7], choice_3, i_3r1[7:7]);
  AND2 I360 (gtint_3[8:8], choice_3, i_3r1[8:8]);
  AND2 I361 (gtint_3[9:9], choice_3, i_3r1[9:9]);
  AND2 I362 (gtint_3[10:10], choice_3, i_3r1[10:10]);
  AND2 I363 (gtint_3[11:11], choice_3, i_3r1[11:11]);
  AND2 I364 (gtint_3[12:12], choice_3, i_3r1[12:12]);
  AND2 I365 (gtint_3[13:13], choice_3, i_3r1[13:13]);
  AND2 I366 (gtint_3[14:14], choice_3, i_3r1[14:14]);
  AND2 I367 (gtint_3[15:15], choice_3, i_3r1[15:15]);
  AND2 I368 (gtint_3[16:16], choice_3, i_3r1[16:16]);
  AND2 I369 (gtint_3[17:17], choice_3, i_3r1[17:17]);
  AND2 I370 (gtint_3[18:18], choice_3, i_3r1[18:18]);
  AND2 I371 (gtint_3[19:19], choice_3, i_3r1[19:19]);
  AND2 I372 (gtint_3[20:20], choice_3, i_3r1[20:20]);
  AND2 I373 (gtint_3[21:21], choice_3, i_3r1[21:21]);
  AND2 I374 (gtint_3[22:22], choice_3, i_3r1[22:22]);
  AND2 I375 (gtint_3[23:23], choice_3, i_3r1[23:23]);
  AND2 I376 (gtint_3[24:24], choice_3, i_3r1[24:24]);
  AND2 I377 (gtint_3[25:25], choice_3, i_3r1[25:25]);
  AND2 I378 (gtint_3[26:26], choice_3, i_3r1[26:26]);
  AND2 I379 (gtint_3[27:27], choice_3, i_3r1[27:27]);
  AND2 I380 (gtint_3[28:28], choice_3, i_3r1[28:28]);
  AND2 I381 (gtint_3[29:29], choice_3, i_3r1[29:29]);
  AND2 I382 (gtint_3[30:30], choice_3, i_3r1[30:30]);
  AND2 I383 (gtint_3[31:31], choice_3, i_3r1[31:31]);
  AND2 I384 (gtint_4[0:0], choice_4, i_4r1[0:0]);
  AND2 I385 (gtint_4[1:1], choice_4, i_4r1[1:1]);
  AND2 I386 (gtint_4[2:2], choice_4, i_4r1[2:2]);
  AND2 I387 (gtint_4[3:3], choice_4, i_4r1[3:3]);
  AND2 I388 (gtint_4[4:4], choice_4, i_4r1[4:4]);
  AND2 I389 (gtint_4[5:5], choice_4, i_4r1[5:5]);
  AND2 I390 (gtint_4[6:6], choice_4, i_4r1[6:6]);
  AND2 I391 (gtint_4[7:7], choice_4, i_4r1[7:7]);
  AND2 I392 (gtint_4[8:8], choice_4, i_4r1[8:8]);
  AND2 I393 (gtint_4[9:9], choice_4, i_4r1[9:9]);
  AND2 I394 (gtint_4[10:10], choice_4, i_4r1[10:10]);
  AND2 I395 (gtint_4[11:11], choice_4, i_4r1[11:11]);
  AND2 I396 (gtint_4[12:12], choice_4, i_4r1[12:12]);
  AND2 I397 (gtint_4[13:13], choice_4, i_4r1[13:13]);
  AND2 I398 (gtint_4[14:14], choice_4, i_4r1[14:14]);
  AND2 I399 (gtint_4[15:15], choice_4, i_4r1[15:15]);
  AND2 I400 (gtint_4[16:16], choice_4, i_4r1[16:16]);
  AND2 I401 (gtint_4[17:17], choice_4, i_4r1[17:17]);
  AND2 I402 (gtint_4[18:18], choice_4, i_4r1[18:18]);
  AND2 I403 (gtint_4[19:19], choice_4, i_4r1[19:19]);
  AND2 I404 (gtint_4[20:20], choice_4, i_4r1[20:20]);
  AND2 I405 (gtint_4[21:21], choice_4, i_4r1[21:21]);
  AND2 I406 (gtint_4[22:22], choice_4, i_4r1[22:22]);
  AND2 I407 (gtint_4[23:23], choice_4, i_4r1[23:23]);
  AND2 I408 (gtint_4[24:24], choice_4, i_4r1[24:24]);
  AND2 I409 (gtint_4[25:25], choice_4, i_4r1[25:25]);
  AND2 I410 (gtint_4[26:26], choice_4, i_4r1[26:26]);
  AND2 I411 (gtint_4[27:27], choice_4, i_4r1[27:27]);
  AND2 I412 (gtint_4[28:28], choice_4, i_4r1[28:28]);
  AND2 I413 (gtint_4[29:29], choice_4, i_4r1[29:29]);
  AND2 I414 (gtint_4[30:30], choice_4, i_4r1[30:30]);
  AND2 I415 (gtint_4[31:31], choice_4, i_4r1[31:31]);
  AND2 I416 (gtint_5[0:0], choice_5, i_5r1[0:0]);
  AND2 I417 (gtint_5[1:1], choice_5, i_5r1[1:1]);
  AND2 I418 (gtint_5[2:2], choice_5, i_5r1[2:2]);
  AND2 I419 (gtint_5[3:3], choice_5, i_5r1[3:3]);
  AND2 I420 (gtint_5[4:4], choice_5, i_5r1[4:4]);
  AND2 I421 (gtint_5[5:5], choice_5, i_5r1[5:5]);
  AND2 I422 (gtint_5[6:6], choice_5, i_5r1[6:6]);
  AND2 I423 (gtint_5[7:7], choice_5, i_5r1[7:7]);
  AND2 I424 (gtint_5[8:8], choice_5, i_5r1[8:8]);
  AND2 I425 (gtint_5[9:9], choice_5, i_5r1[9:9]);
  AND2 I426 (gtint_5[10:10], choice_5, i_5r1[10:10]);
  AND2 I427 (gtint_5[11:11], choice_5, i_5r1[11:11]);
  AND2 I428 (gtint_5[12:12], choice_5, i_5r1[12:12]);
  AND2 I429 (gtint_5[13:13], choice_5, i_5r1[13:13]);
  AND2 I430 (gtint_5[14:14], choice_5, i_5r1[14:14]);
  AND2 I431 (gtint_5[15:15], choice_5, i_5r1[15:15]);
  AND2 I432 (gtint_5[16:16], choice_5, i_5r1[16:16]);
  AND2 I433 (gtint_5[17:17], choice_5, i_5r1[17:17]);
  AND2 I434 (gtint_5[18:18], choice_5, i_5r1[18:18]);
  AND2 I435 (gtint_5[19:19], choice_5, i_5r1[19:19]);
  AND2 I436 (gtint_5[20:20], choice_5, i_5r1[20:20]);
  AND2 I437 (gtint_5[21:21], choice_5, i_5r1[21:21]);
  AND2 I438 (gtint_5[22:22], choice_5, i_5r1[22:22]);
  AND2 I439 (gtint_5[23:23], choice_5, i_5r1[23:23]);
  AND2 I440 (gtint_5[24:24], choice_5, i_5r1[24:24]);
  AND2 I441 (gtint_5[25:25], choice_5, i_5r1[25:25]);
  AND2 I442 (gtint_5[26:26], choice_5, i_5r1[26:26]);
  AND2 I443 (gtint_5[27:27], choice_5, i_5r1[27:27]);
  AND2 I444 (gtint_5[28:28], choice_5, i_5r1[28:28]);
  AND2 I445 (gtint_5[29:29], choice_5, i_5r1[29:29]);
  AND2 I446 (gtint_5[30:30], choice_5, i_5r1[30:30]);
  AND2 I447 (gtint_5[31:31], choice_5, i_5r1[31:31]);
  AND2 I448 (gtint_6[0:0], choice_6, i_6r1[0:0]);
  AND2 I449 (gtint_6[1:1], choice_6, i_6r1[1:1]);
  AND2 I450 (gtint_6[2:2], choice_6, i_6r1[2:2]);
  AND2 I451 (gtint_6[3:3], choice_6, i_6r1[3:3]);
  AND2 I452 (gtint_6[4:4], choice_6, i_6r1[4:4]);
  AND2 I453 (gtint_6[5:5], choice_6, i_6r1[5:5]);
  AND2 I454 (gtint_6[6:6], choice_6, i_6r1[6:6]);
  AND2 I455 (gtint_6[7:7], choice_6, i_6r1[7:7]);
  AND2 I456 (gtint_6[8:8], choice_6, i_6r1[8:8]);
  AND2 I457 (gtint_6[9:9], choice_6, i_6r1[9:9]);
  AND2 I458 (gtint_6[10:10], choice_6, i_6r1[10:10]);
  AND2 I459 (gtint_6[11:11], choice_6, i_6r1[11:11]);
  AND2 I460 (gtint_6[12:12], choice_6, i_6r1[12:12]);
  AND2 I461 (gtint_6[13:13], choice_6, i_6r1[13:13]);
  AND2 I462 (gtint_6[14:14], choice_6, i_6r1[14:14]);
  AND2 I463 (gtint_6[15:15], choice_6, i_6r1[15:15]);
  AND2 I464 (gtint_6[16:16], choice_6, i_6r1[16:16]);
  AND2 I465 (gtint_6[17:17], choice_6, i_6r1[17:17]);
  AND2 I466 (gtint_6[18:18], choice_6, i_6r1[18:18]);
  AND2 I467 (gtint_6[19:19], choice_6, i_6r1[19:19]);
  AND2 I468 (gtint_6[20:20], choice_6, i_6r1[20:20]);
  AND2 I469 (gtint_6[21:21], choice_6, i_6r1[21:21]);
  AND2 I470 (gtint_6[22:22], choice_6, i_6r1[22:22]);
  AND2 I471 (gtint_6[23:23], choice_6, i_6r1[23:23]);
  AND2 I472 (gtint_6[24:24], choice_6, i_6r1[24:24]);
  AND2 I473 (gtint_6[25:25], choice_6, i_6r1[25:25]);
  AND2 I474 (gtint_6[26:26], choice_6, i_6r1[26:26]);
  AND2 I475 (gtint_6[27:27], choice_6, i_6r1[27:27]);
  AND2 I476 (gtint_6[28:28], choice_6, i_6r1[28:28]);
  AND2 I477 (gtint_6[29:29], choice_6, i_6r1[29:29]);
  AND2 I478 (gtint_6[30:30], choice_6, i_6r1[30:30]);
  AND2 I479 (gtint_6[31:31], choice_6, i_6r1[31:31]);
  AND2 I480 (gtint_7[0:0], choice_7, i_7r1[0:0]);
  AND2 I481 (gtint_7[1:1], choice_7, i_7r1[1:1]);
  AND2 I482 (gtint_7[2:2], choice_7, i_7r1[2:2]);
  AND2 I483 (gtint_7[3:3], choice_7, i_7r1[3:3]);
  AND2 I484 (gtint_7[4:4], choice_7, i_7r1[4:4]);
  AND2 I485 (gtint_7[5:5], choice_7, i_7r1[5:5]);
  AND2 I486 (gtint_7[6:6], choice_7, i_7r1[6:6]);
  AND2 I487 (gtint_7[7:7], choice_7, i_7r1[7:7]);
  AND2 I488 (gtint_7[8:8], choice_7, i_7r1[8:8]);
  AND2 I489 (gtint_7[9:9], choice_7, i_7r1[9:9]);
  AND2 I490 (gtint_7[10:10], choice_7, i_7r1[10:10]);
  AND2 I491 (gtint_7[11:11], choice_7, i_7r1[11:11]);
  AND2 I492 (gtint_7[12:12], choice_7, i_7r1[12:12]);
  AND2 I493 (gtint_7[13:13], choice_7, i_7r1[13:13]);
  AND2 I494 (gtint_7[14:14], choice_7, i_7r1[14:14]);
  AND2 I495 (gtint_7[15:15], choice_7, i_7r1[15:15]);
  AND2 I496 (gtint_7[16:16], choice_7, i_7r1[16:16]);
  AND2 I497 (gtint_7[17:17], choice_7, i_7r1[17:17]);
  AND2 I498 (gtint_7[18:18], choice_7, i_7r1[18:18]);
  AND2 I499 (gtint_7[19:19], choice_7, i_7r1[19:19]);
  AND2 I500 (gtint_7[20:20], choice_7, i_7r1[20:20]);
  AND2 I501 (gtint_7[21:21], choice_7, i_7r1[21:21]);
  AND2 I502 (gtint_7[22:22], choice_7, i_7r1[22:22]);
  AND2 I503 (gtint_7[23:23], choice_7, i_7r1[23:23]);
  AND2 I504 (gtint_7[24:24], choice_7, i_7r1[24:24]);
  AND2 I505 (gtint_7[25:25], choice_7, i_7r1[25:25]);
  AND2 I506 (gtint_7[26:26], choice_7, i_7r1[26:26]);
  AND2 I507 (gtint_7[27:27], choice_7, i_7r1[27:27]);
  AND2 I508 (gtint_7[28:28], choice_7, i_7r1[28:28]);
  AND2 I509 (gtint_7[29:29], choice_7, i_7r1[29:29]);
  AND2 I510 (gtint_7[30:30], choice_7, i_7r1[30:30]);
  AND2 I511 (gtint_7[31:31], choice_7, i_7r1[31:31]);
  AND2 I512 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I513 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I514 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I515 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I516 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I517 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I518 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I519 (gfint_0[7:7], choice_0, i_0r0[7:7]);
  AND2 I520 (gfint_0[8:8], choice_0, i_0r0[8:8]);
  AND2 I521 (gfint_0[9:9], choice_0, i_0r0[9:9]);
  AND2 I522 (gfint_0[10:10], choice_0, i_0r0[10:10]);
  AND2 I523 (gfint_0[11:11], choice_0, i_0r0[11:11]);
  AND2 I524 (gfint_0[12:12], choice_0, i_0r0[12:12]);
  AND2 I525 (gfint_0[13:13], choice_0, i_0r0[13:13]);
  AND2 I526 (gfint_0[14:14], choice_0, i_0r0[14:14]);
  AND2 I527 (gfint_0[15:15], choice_0, i_0r0[15:15]);
  AND2 I528 (gfint_0[16:16], choice_0, i_0r0[16:16]);
  AND2 I529 (gfint_0[17:17], choice_0, i_0r0[17:17]);
  AND2 I530 (gfint_0[18:18], choice_0, i_0r0[18:18]);
  AND2 I531 (gfint_0[19:19], choice_0, i_0r0[19:19]);
  AND2 I532 (gfint_0[20:20], choice_0, i_0r0[20:20]);
  AND2 I533 (gfint_0[21:21], choice_0, i_0r0[21:21]);
  AND2 I534 (gfint_0[22:22], choice_0, i_0r0[22:22]);
  AND2 I535 (gfint_0[23:23], choice_0, i_0r0[23:23]);
  AND2 I536 (gfint_0[24:24], choice_0, i_0r0[24:24]);
  AND2 I537 (gfint_0[25:25], choice_0, i_0r0[25:25]);
  AND2 I538 (gfint_0[26:26], choice_0, i_0r0[26:26]);
  AND2 I539 (gfint_0[27:27], choice_0, i_0r0[27:27]);
  AND2 I540 (gfint_0[28:28], choice_0, i_0r0[28:28]);
  AND2 I541 (gfint_0[29:29], choice_0, i_0r0[29:29]);
  AND2 I542 (gfint_0[30:30], choice_0, i_0r0[30:30]);
  AND2 I543 (gfint_0[31:31], choice_0, i_0r0[31:31]);
  AND2 I544 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I545 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I546 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I547 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I548 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I549 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I550 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I551 (gfint_1[7:7], choice_1, i_1r0[7:7]);
  AND2 I552 (gfint_1[8:8], choice_1, i_1r0[8:8]);
  AND2 I553 (gfint_1[9:9], choice_1, i_1r0[9:9]);
  AND2 I554 (gfint_1[10:10], choice_1, i_1r0[10:10]);
  AND2 I555 (gfint_1[11:11], choice_1, i_1r0[11:11]);
  AND2 I556 (gfint_1[12:12], choice_1, i_1r0[12:12]);
  AND2 I557 (gfint_1[13:13], choice_1, i_1r0[13:13]);
  AND2 I558 (gfint_1[14:14], choice_1, i_1r0[14:14]);
  AND2 I559 (gfint_1[15:15], choice_1, i_1r0[15:15]);
  AND2 I560 (gfint_1[16:16], choice_1, i_1r0[16:16]);
  AND2 I561 (gfint_1[17:17], choice_1, i_1r0[17:17]);
  AND2 I562 (gfint_1[18:18], choice_1, i_1r0[18:18]);
  AND2 I563 (gfint_1[19:19], choice_1, i_1r0[19:19]);
  AND2 I564 (gfint_1[20:20], choice_1, i_1r0[20:20]);
  AND2 I565 (gfint_1[21:21], choice_1, i_1r0[21:21]);
  AND2 I566 (gfint_1[22:22], choice_1, i_1r0[22:22]);
  AND2 I567 (gfint_1[23:23], choice_1, i_1r0[23:23]);
  AND2 I568 (gfint_1[24:24], choice_1, i_1r0[24:24]);
  AND2 I569 (gfint_1[25:25], choice_1, i_1r0[25:25]);
  AND2 I570 (gfint_1[26:26], choice_1, i_1r0[26:26]);
  AND2 I571 (gfint_1[27:27], choice_1, i_1r0[27:27]);
  AND2 I572 (gfint_1[28:28], choice_1, i_1r0[28:28]);
  AND2 I573 (gfint_1[29:29], choice_1, i_1r0[29:29]);
  AND2 I574 (gfint_1[30:30], choice_1, i_1r0[30:30]);
  AND2 I575 (gfint_1[31:31], choice_1, i_1r0[31:31]);
  AND2 I576 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I577 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I578 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I579 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AND2 I580 (gfint_2[4:4], choice_2, i_2r0[4:4]);
  AND2 I581 (gfint_2[5:5], choice_2, i_2r0[5:5]);
  AND2 I582 (gfint_2[6:6], choice_2, i_2r0[6:6]);
  AND2 I583 (gfint_2[7:7], choice_2, i_2r0[7:7]);
  AND2 I584 (gfint_2[8:8], choice_2, i_2r0[8:8]);
  AND2 I585 (gfint_2[9:9], choice_2, i_2r0[9:9]);
  AND2 I586 (gfint_2[10:10], choice_2, i_2r0[10:10]);
  AND2 I587 (gfint_2[11:11], choice_2, i_2r0[11:11]);
  AND2 I588 (gfint_2[12:12], choice_2, i_2r0[12:12]);
  AND2 I589 (gfint_2[13:13], choice_2, i_2r0[13:13]);
  AND2 I590 (gfint_2[14:14], choice_2, i_2r0[14:14]);
  AND2 I591 (gfint_2[15:15], choice_2, i_2r0[15:15]);
  AND2 I592 (gfint_2[16:16], choice_2, i_2r0[16:16]);
  AND2 I593 (gfint_2[17:17], choice_2, i_2r0[17:17]);
  AND2 I594 (gfint_2[18:18], choice_2, i_2r0[18:18]);
  AND2 I595 (gfint_2[19:19], choice_2, i_2r0[19:19]);
  AND2 I596 (gfint_2[20:20], choice_2, i_2r0[20:20]);
  AND2 I597 (gfint_2[21:21], choice_2, i_2r0[21:21]);
  AND2 I598 (gfint_2[22:22], choice_2, i_2r0[22:22]);
  AND2 I599 (gfint_2[23:23], choice_2, i_2r0[23:23]);
  AND2 I600 (gfint_2[24:24], choice_2, i_2r0[24:24]);
  AND2 I601 (gfint_2[25:25], choice_2, i_2r0[25:25]);
  AND2 I602 (gfint_2[26:26], choice_2, i_2r0[26:26]);
  AND2 I603 (gfint_2[27:27], choice_2, i_2r0[27:27]);
  AND2 I604 (gfint_2[28:28], choice_2, i_2r0[28:28]);
  AND2 I605 (gfint_2[29:29], choice_2, i_2r0[29:29]);
  AND2 I606 (gfint_2[30:30], choice_2, i_2r0[30:30]);
  AND2 I607 (gfint_2[31:31], choice_2, i_2r0[31:31]);
  AND2 I608 (gfint_3[0:0], choice_3, i_3r0[0:0]);
  AND2 I609 (gfint_3[1:1], choice_3, i_3r0[1:1]);
  AND2 I610 (gfint_3[2:2], choice_3, i_3r0[2:2]);
  AND2 I611 (gfint_3[3:3], choice_3, i_3r0[3:3]);
  AND2 I612 (gfint_3[4:4], choice_3, i_3r0[4:4]);
  AND2 I613 (gfint_3[5:5], choice_3, i_3r0[5:5]);
  AND2 I614 (gfint_3[6:6], choice_3, i_3r0[6:6]);
  AND2 I615 (gfint_3[7:7], choice_3, i_3r0[7:7]);
  AND2 I616 (gfint_3[8:8], choice_3, i_3r0[8:8]);
  AND2 I617 (gfint_3[9:9], choice_3, i_3r0[9:9]);
  AND2 I618 (gfint_3[10:10], choice_3, i_3r0[10:10]);
  AND2 I619 (gfint_3[11:11], choice_3, i_3r0[11:11]);
  AND2 I620 (gfint_3[12:12], choice_3, i_3r0[12:12]);
  AND2 I621 (gfint_3[13:13], choice_3, i_3r0[13:13]);
  AND2 I622 (gfint_3[14:14], choice_3, i_3r0[14:14]);
  AND2 I623 (gfint_3[15:15], choice_3, i_3r0[15:15]);
  AND2 I624 (gfint_3[16:16], choice_3, i_3r0[16:16]);
  AND2 I625 (gfint_3[17:17], choice_3, i_3r0[17:17]);
  AND2 I626 (gfint_3[18:18], choice_3, i_3r0[18:18]);
  AND2 I627 (gfint_3[19:19], choice_3, i_3r0[19:19]);
  AND2 I628 (gfint_3[20:20], choice_3, i_3r0[20:20]);
  AND2 I629 (gfint_3[21:21], choice_3, i_3r0[21:21]);
  AND2 I630 (gfint_3[22:22], choice_3, i_3r0[22:22]);
  AND2 I631 (gfint_3[23:23], choice_3, i_3r0[23:23]);
  AND2 I632 (gfint_3[24:24], choice_3, i_3r0[24:24]);
  AND2 I633 (gfint_3[25:25], choice_3, i_3r0[25:25]);
  AND2 I634 (gfint_3[26:26], choice_3, i_3r0[26:26]);
  AND2 I635 (gfint_3[27:27], choice_3, i_3r0[27:27]);
  AND2 I636 (gfint_3[28:28], choice_3, i_3r0[28:28]);
  AND2 I637 (gfint_3[29:29], choice_3, i_3r0[29:29]);
  AND2 I638 (gfint_3[30:30], choice_3, i_3r0[30:30]);
  AND2 I639 (gfint_3[31:31], choice_3, i_3r0[31:31]);
  AND2 I640 (gfint_4[0:0], choice_4, i_4r0[0:0]);
  AND2 I641 (gfint_4[1:1], choice_4, i_4r0[1:1]);
  AND2 I642 (gfint_4[2:2], choice_4, i_4r0[2:2]);
  AND2 I643 (gfint_4[3:3], choice_4, i_4r0[3:3]);
  AND2 I644 (gfint_4[4:4], choice_4, i_4r0[4:4]);
  AND2 I645 (gfint_4[5:5], choice_4, i_4r0[5:5]);
  AND2 I646 (gfint_4[6:6], choice_4, i_4r0[6:6]);
  AND2 I647 (gfint_4[7:7], choice_4, i_4r0[7:7]);
  AND2 I648 (gfint_4[8:8], choice_4, i_4r0[8:8]);
  AND2 I649 (gfint_4[9:9], choice_4, i_4r0[9:9]);
  AND2 I650 (gfint_4[10:10], choice_4, i_4r0[10:10]);
  AND2 I651 (gfint_4[11:11], choice_4, i_4r0[11:11]);
  AND2 I652 (gfint_4[12:12], choice_4, i_4r0[12:12]);
  AND2 I653 (gfint_4[13:13], choice_4, i_4r0[13:13]);
  AND2 I654 (gfint_4[14:14], choice_4, i_4r0[14:14]);
  AND2 I655 (gfint_4[15:15], choice_4, i_4r0[15:15]);
  AND2 I656 (gfint_4[16:16], choice_4, i_4r0[16:16]);
  AND2 I657 (gfint_4[17:17], choice_4, i_4r0[17:17]);
  AND2 I658 (gfint_4[18:18], choice_4, i_4r0[18:18]);
  AND2 I659 (gfint_4[19:19], choice_4, i_4r0[19:19]);
  AND2 I660 (gfint_4[20:20], choice_4, i_4r0[20:20]);
  AND2 I661 (gfint_4[21:21], choice_4, i_4r0[21:21]);
  AND2 I662 (gfint_4[22:22], choice_4, i_4r0[22:22]);
  AND2 I663 (gfint_4[23:23], choice_4, i_4r0[23:23]);
  AND2 I664 (gfint_4[24:24], choice_4, i_4r0[24:24]);
  AND2 I665 (gfint_4[25:25], choice_4, i_4r0[25:25]);
  AND2 I666 (gfint_4[26:26], choice_4, i_4r0[26:26]);
  AND2 I667 (gfint_4[27:27], choice_4, i_4r0[27:27]);
  AND2 I668 (gfint_4[28:28], choice_4, i_4r0[28:28]);
  AND2 I669 (gfint_4[29:29], choice_4, i_4r0[29:29]);
  AND2 I670 (gfint_4[30:30], choice_4, i_4r0[30:30]);
  AND2 I671 (gfint_4[31:31], choice_4, i_4r0[31:31]);
  AND2 I672 (gfint_5[0:0], choice_5, i_5r0[0:0]);
  AND2 I673 (gfint_5[1:1], choice_5, i_5r0[1:1]);
  AND2 I674 (gfint_5[2:2], choice_5, i_5r0[2:2]);
  AND2 I675 (gfint_5[3:3], choice_5, i_5r0[3:3]);
  AND2 I676 (gfint_5[4:4], choice_5, i_5r0[4:4]);
  AND2 I677 (gfint_5[5:5], choice_5, i_5r0[5:5]);
  AND2 I678 (gfint_5[6:6], choice_5, i_5r0[6:6]);
  AND2 I679 (gfint_5[7:7], choice_5, i_5r0[7:7]);
  AND2 I680 (gfint_5[8:8], choice_5, i_5r0[8:8]);
  AND2 I681 (gfint_5[9:9], choice_5, i_5r0[9:9]);
  AND2 I682 (gfint_5[10:10], choice_5, i_5r0[10:10]);
  AND2 I683 (gfint_5[11:11], choice_5, i_5r0[11:11]);
  AND2 I684 (gfint_5[12:12], choice_5, i_5r0[12:12]);
  AND2 I685 (gfint_5[13:13], choice_5, i_5r0[13:13]);
  AND2 I686 (gfint_5[14:14], choice_5, i_5r0[14:14]);
  AND2 I687 (gfint_5[15:15], choice_5, i_5r0[15:15]);
  AND2 I688 (gfint_5[16:16], choice_5, i_5r0[16:16]);
  AND2 I689 (gfint_5[17:17], choice_5, i_5r0[17:17]);
  AND2 I690 (gfint_5[18:18], choice_5, i_5r0[18:18]);
  AND2 I691 (gfint_5[19:19], choice_5, i_5r0[19:19]);
  AND2 I692 (gfint_5[20:20], choice_5, i_5r0[20:20]);
  AND2 I693 (gfint_5[21:21], choice_5, i_5r0[21:21]);
  AND2 I694 (gfint_5[22:22], choice_5, i_5r0[22:22]);
  AND2 I695 (gfint_5[23:23], choice_5, i_5r0[23:23]);
  AND2 I696 (gfint_5[24:24], choice_5, i_5r0[24:24]);
  AND2 I697 (gfint_5[25:25], choice_5, i_5r0[25:25]);
  AND2 I698 (gfint_5[26:26], choice_5, i_5r0[26:26]);
  AND2 I699 (gfint_5[27:27], choice_5, i_5r0[27:27]);
  AND2 I700 (gfint_5[28:28], choice_5, i_5r0[28:28]);
  AND2 I701 (gfint_5[29:29], choice_5, i_5r0[29:29]);
  AND2 I702 (gfint_5[30:30], choice_5, i_5r0[30:30]);
  AND2 I703 (gfint_5[31:31], choice_5, i_5r0[31:31]);
  AND2 I704 (gfint_6[0:0], choice_6, i_6r0[0:0]);
  AND2 I705 (gfint_6[1:1], choice_6, i_6r0[1:1]);
  AND2 I706 (gfint_6[2:2], choice_6, i_6r0[2:2]);
  AND2 I707 (gfint_6[3:3], choice_6, i_6r0[3:3]);
  AND2 I708 (gfint_6[4:4], choice_6, i_6r0[4:4]);
  AND2 I709 (gfint_6[5:5], choice_6, i_6r0[5:5]);
  AND2 I710 (gfint_6[6:6], choice_6, i_6r0[6:6]);
  AND2 I711 (gfint_6[7:7], choice_6, i_6r0[7:7]);
  AND2 I712 (gfint_6[8:8], choice_6, i_6r0[8:8]);
  AND2 I713 (gfint_6[9:9], choice_6, i_6r0[9:9]);
  AND2 I714 (gfint_6[10:10], choice_6, i_6r0[10:10]);
  AND2 I715 (gfint_6[11:11], choice_6, i_6r0[11:11]);
  AND2 I716 (gfint_6[12:12], choice_6, i_6r0[12:12]);
  AND2 I717 (gfint_6[13:13], choice_6, i_6r0[13:13]);
  AND2 I718 (gfint_6[14:14], choice_6, i_6r0[14:14]);
  AND2 I719 (gfint_6[15:15], choice_6, i_6r0[15:15]);
  AND2 I720 (gfint_6[16:16], choice_6, i_6r0[16:16]);
  AND2 I721 (gfint_6[17:17], choice_6, i_6r0[17:17]);
  AND2 I722 (gfint_6[18:18], choice_6, i_6r0[18:18]);
  AND2 I723 (gfint_6[19:19], choice_6, i_6r0[19:19]);
  AND2 I724 (gfint_6[20:20], choice_6, i_6r0[20:20]);
  AND2 I725 (gfint_6[21:21], choice_6, i_6r0[21:21]);
  AND2 I726 (gfint_6[22:22], choice_6, i_6r0[22:22]);
  AND2 I727 (gfint_6[23:23], choice_6, i_6r0[23:23]);
  AND2 I728 (gfint_6[24:24], choice_6, i_6r0[24:24]);
  AND2 I729 (gfint_6[25:25], choice_6, i_6r0[25:25]);
  AND2 I730 (gfint_6[26:26], choice_6, i_6r0[26:26]);
  AND2 I731 (gfint_6[27:27], choice_6, i_6r0[27:27]);
  AND2 I732 (gfint_6[28:28], choice_6, i_6r0[28:28]);
  AND2 I733 (gfint_6[29:29], choice_6, i_6r0[29:29]);
  AND2 I734 (gfint_6[30:30], choice_6, i_6r0[30:30]);
  AND2 I735 (gfint_6[31:31], choice_6, i_6r0[31:31]);
  AND2 I736 (gfint_7[0:0], choice_7, i_7r0[0:0]);
  AND2 I737 (gfint_7[1:1], choice_7, i_7r0[1:1]);
  AND2 I738 (gfint_7[2:2], choice_7, i_7r0[2:2]);
  AND2 I739 (gfint_7[3:3], choice_7, i_7r0[3:3]);
  AND2 I740 (gfint_7[4:4], choice_7, i_7r0[4:4]);
  AND2 I741 (gfint_7[5:5], choice_7, i_7r0[5:5]);
  AND2 I742 (gfint_7[6:6], choice_7, i_7r0[6:6]);
  AND2 I743 (gfint_7[7:7], choice_7, i_7r0[7:7]);
  AND2 I744 (gfint_7[8:8], choice_7, i_7r0[8:8]);
  AND2 I745 (gfint_7[9:9], choice_7, i_7r0[9:9]);
  AND2 I746 (gfint_7[10:10], choice_7, i_7r0[10:10]);
  AND2 I747 (gfint_7[11:11], choice_7, i_7r0[11:11]);
  AND2 I748 (gfint_7[12:12], choice_7, i_7r0[12:12]);
  AND2 I749 (gfint_7[13:13], choice_7, i_7r0[13:13]);
  AND2 I750 (gfint_7[14:14], choice_7, i_7r0[14:14]);
  AND2 I751 (gfint_7[15:15], choice_7, i_7r0[15:15]);
  AND2 I752 (gfint_7[16:16], choice_7, i_7r0[16:16]);
  AND2 I753 (gfint_7[17:17], choice_7, i_7r0[17:17]);
  AND2 I754 (gfint_7[18:18], choice_7, i_7r0[18:18]);
  AND2 I755 (gfint_7[19:19], choice_7, i_7r0[19:19]);
  AND2 I756 (gfint_7[20:20], choice_7, i_7r0[20:20]);
  AND2 I757 (gfint_7[21:21], choice_7, i_7r0[21:21]);
  AND2 I758 (gfint_7[22:22], choice_7, i_7r0[22:22]);
  AND2 I759 (gfint_7[23:23], choice_7, i_7r0[23:23]);
  AND2 I760 (gfint_7[24:24], choice_7, i_7r0[24:24]);
  AND2 I761 (gfint_7[25:25], choice_7, i_7r0[25:25]);
  AND2 I762 (gfint_7[26:26], choice_7, i_7r0[26:26]);
  AND2 I763 (gfint_7[27:27], choice_7, i_7r0[27:27]);
  AND2 I764 (gfint_7[28:28], choice_7, i_7r0[28:28]);
  AND2 I765 (gfint_7[29:29], choice_7, i_7r0[29:29]);
  AND2 I766 (gfint_7[30:30], choice_7, i_7r0[30:30]);
  AND2 I767 (gfint_7[31:31], choice_7, i_7r0[31:31]);
  OR2 I768 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I769 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I770 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I771 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I772 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I773 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I774 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I775 (comp0_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I776 (comp0_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I777 (comp0_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I778 (comp0_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I779 (comp0_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I780 (comp0_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I781 (comp0_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I782 (comp0_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I783 (comp0_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I784 (comp0_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I785 (comp0_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I786 (comp0_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I787 (comp0_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I788 (comp0_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I789 (comp0_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I790 (comp0_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I791 (comp0_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I792 (comp0_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I793 (comp0_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I794 (comp0_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I795 (comp0_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I796 (comp0_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I797 (comp0_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I798 (comp0_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I799 (comp0_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  C3 I800 (simp6431_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I801 (simp6431_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I802 (simp6431_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I803 (simp6431_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I804 (simp6431_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I805 (simp6431_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I806 (simp6431_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I807 (simp6431_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I808 (simp6431_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I809 (simp6431_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I810 (simp6431_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I811 (simp6432_0[0:0], simp6431_0[0:0], simp6431_0[1:1], simp6431_0[2:2]);
  C3 I812 (simp6432_0[1:1], simp6431_0[3:3], simp6431_0[4:4], simp6431_0[5:5]);
  C3 I813 (simp6432_0[2:2], simp6431_0[6:6], simp6431_0[7:7], simp6431_0[8:8]);
  C2 I814 (simp6432_0[3:3], simp6431_0[9:9], simp6431_0[10:10]);
  C3 I815 (simp6433_0[0:0], simp6432_0[0:0], simp6432_0[1:1], simp6432_0[2:2]);
  BUFF I816 (simp6433_0[1:1], simp6432_0[3:3]);
  C2 I817 (icomp_0, simp6433_0[0:0], simp6433_0[1:1]);
  OR2 I818 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I819 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I820 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I821 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I822 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I823 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I824 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  OR2 I825 (comp1_0[7:7], i_1r0[7:7], i_1r1[7:7]);
  OR2 I826 (comp1_0[8:8], i_1r0[8:8], i_1r1[8:8]);
  OR2 I827 (comp1_0[9:9], i_1r0[9:9], i_1r1[9:9]);
  OR2 I828 (comp1_0[10:10], i_1r0[10:10], i_1r1[10:10]);
  OR2 I829 (comp1_0[11:11], i_1r0[11:11], i_1r1[11:11]);
  OR2 I830 (comp1_0[12:12], i_1r0[12:12], i_1r1[12:12]);
  OR2 I831 (comp1_0[13:13], i_1r0[13:13], i_1r1[13:13]);
  OR2 I832 (comp1_0[14:14], i_1r0[14:14], i_1r1[14:14]);
  OR2 I833 (comp1_0[15:15], i_1r0[15:15], i_1r1[15:15]);
  OR2 I834 (comp1_0[16:16], i_1r0[16:16], i_1r1[16:16]);
  OR2 I835 (comp1_0[17:17], i_1r0[17:17], i_1r1[17:17]);
  OR2 I836 (comp1_0[18:18], i_1r0[18:18], i_1r1[18:18]);
  OR2 I837 (comp1_0[19:19], i_1r0[19:19], i_1r1[19:19]);
  OR2 I838 (comp1_0[20:20], i_1r0[20:20], i_1r1[20:20]);
  OR2 I839 (comp1_0[21:21], i_1r0[21:21], i_1r1[21:21]);
  OR2 I840 (comp1_0[22:22], i_1r0[22:22], i_1r1[22:22]);
  OR2 I841 (comp1_0[23:23], i_1r0[23:23], i_1r1[23:23]);
  OR2 I842 (comp1_0[24:24], i_1r0[24:24], i_1r1[24:24]);
  OR2 I843 (comp1_0[25:25], i_1r0[25:25], i_1r1[25:25]);
  OR2 I844 (comp1_0[26:26], i_1r0[26:26], i_1r1[26:26]);
  OR2 I845 (comp1_0[27:27], i_1r0[27:27], i_1r1[27:27]);
  OR2 I846 (comp1_0[28:28], i_1r0[28:28], i_1r1[28:28]);
  OR2 I847 (comp1_0[29:29], i_1r0[29:29], i_1r1[29:29]);
  OR2 I848 (comp1_0[30:30], i_1r0[30:30], i_1r1[30:30]);
  OR2 I849 (comp1_0[31:31], i_1r0[31:31], i_1r1[31:31]);
  C3 I850 (simp6771_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I851 (simp6771_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  C3 I852 (simp6771_0[2:2], comp1_0[6:6], comp1_0[7:7], comp1_0[8:8]);
  C3 I853 (simp6771_0[3:3], comp1_0[9:9], comp1_0[10:10], comp1_0[11:11]);
  C3 I854 (simp6771_0[4:4], comp1_0[12:12], comp1_0[13:13], comp1_0[14:14]);
  C3 I855 (simp6771_0[5:5], comp1_0[15:15], comp1_0[16:16], comp1_0[17:17]);
  C3 I856 (simp6771_0[6:6], comp1_0[18:18], comp1_0[19:19], comp1_0[20:20]);
  C3 I857 (simp6771_0[7:7], comp1_0[21:21], comp1_0[22:22], comp1_0[23:23]);
  C3 I858 (simp6771_0[8:8], comp1_0[24:24], comp1_0[25:25], comp1_0[26:26]);
  C3 I859 (simp6771_0[9:9], comp1_0[27:27], comp1_0[28:28], comp1_0[29:29]);
  C2 I860 (simp6771_0[10:10], comp1_0[30:30], comp1_0[31:31]);
  C3 I861 (simp6772_0[0:0], simp6771_0[0:0], simp6771_0[1:1], simp6771_0[2:2]);
  C3 I862 (simp6772_0[1:1], simp6771_0[3:3], simp6771_0[4:4], simp6771_0[5:5]);
  C3 I863 (simp6772_0[2:2], simp6771_0[6:6], simp6771_0[7:7], simp6771_0[8:8]);
  C2 I864 (simp6772_0[3:3], simp6771_0[9:9], simp6771_0[10:10]);
  C3 I865 (simp6773_0[0:0], simp6772_0[0:0], simp6772_0[1:1], simp6772_0[2:2]);
  BUFF I866 (simp6773_0[1:1], simp6772_0[3:3]);
  C2 I867 (icomp_1, simp6773_0[0:0], simp6773_0[1:1]);
  OR2 I868 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I869 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I870 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2 I871 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  OR2 I872 (comp2_0[4:4], i_2r0[4:4], i_2r1[4:4]);
  OR2 I873 (comp2_0[5:5], i_2r0[5:5], i_2r1[5:5]);
  OR2 I874 (comp2_0[6:6], i_2r0[6:6], i_2r1[6:6]);
  OR2 I875 (comp2_0[7:7], i_2r0[7:7], i_2r1[7:7]);
  OR2 I876 (comp2_0[8:8], i_2r0[8:8], i_2r1[8:8]);
  OR2 I877 (comp2_0[9:9], i_2r0[9:9], i_2r1[9:9]);
  OR2 I878 (comp2_0[10:10], i_2r0[10:10], i_2r1[10:10]);
  OR2 I879 (comp2_0[11:11], i_2r0[11:11], i_2r1[11:11]);
  OR2 I880 (comp2_0[12:12], i_2r0[12:12], i_2r1[12:12]);
  OR2 I881 (comp2_0[13:13], i_2r0[13:13], i_2r1[13:13]);
  OR2 I882 (comp2_0[14:14], i_2r0[14:14], i_2r1[14:14]);
  OR2 I883 (comp2_0[15:15], i_2r0[15:15], i_2r1[15:15]);
  OR2 I884 (comp2_0[16:16], i_2r0[16:16], i_2r1[16:16]);
  OR2 I885 (comp2_0[17:17], i_2r0[17:17], i_2r1[17:17]);
  OR2 I886 (comp2_0[18:18], i_2r0[18:18], i_2r1[18:18]);
  OR2 I887 (comp2_0[19:19], i_2r0[19:19], i_2r1[19:19]);
  OR2 I888 (comp2_0[20:20], i_2r0[20:20], i_2r1[20:20]);
  OR2 I889 (comp2_0[21:21], i_2r0[21:21], i_2r1[21:21]);
  OR2 I890 (comp2_0[22:22], i_2r0[22:22], i_2r1[22:22]);
  OR2 I891 (comp2_0[23:23], i_2r0[23:23], i_2r1[23:23]);
  OR2 I892 (comp2_0[24:24], i_2r0[24:24], i_2r1[24:24]);
  OR2 I893 (comp2_0[25:25], i_2r0[25:25], i_2r1[25:25]);
  OR2 I894 (comp2_0[26:26], i_2r0[26:26], i_2r1[26:26]);
  OR2 I895 (comp2_0[27:27], i_2r0[27:27], i_2r1[27:27]);
  OR2 I896 (comp2_0[28:28], i_2r0[28:28], i_2r1[28:28]);
  OR2 I897 (comp2_0[29:29], i_2r0[29:29], i_2r1[29:29]);
  OR2 I898 (comp2_0[30:30], i_2r0[30:30], i_2r1[30:30]);
  OR2 I899 (comp2_0[31:31], i_2r0[31:31], i_2r1[31:31]);
  C3 I900 (simp7111_0[0:0], comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C3 I901 (simp7111_0[1:1], comp2_0[3:3], comp2_0[4:4], comp2_0[5:5]);
  C3 I902 (simp7111_0[2:2], comp2_0[6:6], comp2_0[7:7], comp2_0[8:8]);
  C3 I903 (simp7111_0[3:3], comp2_0[9:9], comp2_0[10:10], comp2_0[11:11]);
  C3 I904 (simp7111_0[4:4], comp2_0[12:12], comp2_0[13:13], comp2_0[14:14]);
  C3 I905 (simp7111_0[5:5], comp2_0[15:15], comp2_0[16:16], comp2_0[17:17]);
  C3 I906 (simp7111_0[6:6], comp2_0[18:18], comp2_0[19:19], comp2_0[20:20]);
  C3 I907 (simp7111_0[7:7], comp2_0[21:21], comp2_0[22:22], comp2_0[23:23]);
  C3 I908 (simp7111_0[8:8], comp2_0[24:24], comp2_0[25:25], comp2_0[26:26]);
  C3 I909 (simp7111_0[9:9], comp2_0[27:27], comp2_0[28:28], comp2_0[29:29]);
  C2 I910 (simp7111_0[10:10], comp2_0[30:30], comp2_0[31:31]);
  C3 I911 (simp7112_0[0:0], simp7111_0[0:0], simp7111_0[1:1], simp7111_0[2:2]);
  C3 I912 (simp7112_0[1:1], simp7111_0[3:3], simp7111_0[4:4], simp7111_0[5:5]);
  C3 I913 (simp7112_0[2:2], simp7111_0[6:6], simp7111_0[7:7], simp7111_0[8:8]);
  C2 I914 (simp7112_0[3:3], simp7111_0[9:9], simp7111_0[10:10]);
  C3 I915 (simp7113_0[0:0], simp7112_0[0:0], simp7112_0[1:1], simp7112_0[2:2]);
  BUFF I916 (simp7113_0[1:1], simp7112_0[3:3]);
  C2 I917 (icomp_2, simp7113_0[0:0], simp7113_0[1:1]);
  OR2 I918 (comp3_0[0:0], i_3r0[0:0], i_3r1[0:0]);
  OR2 I919 (comp3_0[1:1], i_3r0[1:1], i_3r1[1:1]);
  OR2 I920 (comp3_0[2:2], i_3r0[2:2], i_3r1[2:2]);
  OR2 I921 (comp3_0[3:3], i_3r0[3:3], i_3r1[3:3]);
  OR2 I922 (comp3_0[4:4], i_3r0[4:4], i_3r1[4:4]);
  OR2 I923 (comp3_0[5:5], i_3r0[5:5], i_3r1[5:5]);
  OR2 I924 (comp3_0[6:6], i_3r0[6:6], i_3r1[6:6]);
  OR2 I925 (comp3_0[7:7], i_3r0[7:7], i_3r1[7:7]);
  OR2 I926 (comp3_0[8:8], i_3r0[8:8], i_3r1[8:8]);
  OR2 I927 (comp3_0[9:9], i_3r0[9:9], i_3r1[9:9]);
  OR2 I928 (comp3_0[10:10], i_3r0[10:10], i_3r1[10:10]);
  OR2 I929 (comp3_0[11:11], i_3r0[11:11], i_3r1[11:11]);
  OR2 I930 (comp3_0[12:12], i_3r0[12:12], i_3r1[12:12]);
  OR2 I931 (comp3_0[13:13], i_3r0[13:13], i_3r1[13:13]);
  OR2 I932 (comp3_0[14:14], i_3r0[14:14], i_3r1[14:14]);
  OR2 I933 (comp3_0[15:15], i_3r0[15:15], i_3r1[15:15]);
  OR2 I934 (comp3_0[16:16], i_3r0[16:16], i_3r1[16:16]);
  OR2 I935 (comp3_0[17:17], i_3r0[17:17], i_3r1[17:17]);
  OR2 I936 (comp3_0[18:18], i_3r0[18:18], i_3r1[18:18]);
  OR2 I937 (comp3_0[19:19], i_3r0[19:19], i_3r1[19:19]);
  OR2 I938 (comp3_0[20:20], i_3r0[20:20], i_3r1[20:20]);
  OR2 I939 (comp3_0[21:21], i_3r0[21:21], i_3r1[21:21]);
  OR2 I940 (comp3_0[22:22], i_3r0[22:22], i_3r1[22:22]);
  OR2 I941 (comp3_0[23:23], i_3r0[23:23], i_3r1[23:23]);
  OR2 I942 (comp3_0[24:24], i_3r0[24:24], i_3r1[24:24]);
  OR2 I943 (comp3_0[25:25], i_3r0[25:25], i_3r1[25:25]);
  OR2 I944 (comp3_0[26:26], i_3r0[26:26], i_3r1[26:26]);
  OR2 I945 (comp3_0[27:27], i_3r0[27:27], i_3r1[27:27]);
  OR2 I946 (comp3_0[28:28], i_3r0[28:28], i_3r1[28:28]);
  OR2 I947 (comp3_0[29:29], i_3r0[29:29], i_3r1[29:29]);
  OR2 I948 (comp3_0[30:30], i_3r0[30:30], i_3r1[30:30]);
  OR2 I949 (comp3_0[31:31], i_3r0[31:31], i_3r1[31:31]);
  C3 I950 (simp7451_0[0:0], comp3_0[0:0], comp3_0[1:1], comp3_0[2:2]);
  C3 I951 (simp7451_0[1:1], comp3_0[3:3], comp3_0[4:4], comp3_0[5:5]);
  C3 I952 (simp7451_0[2:2], comp3_0[6:6], comp3_0[7:7], comp3_0[8:8]);
  C3 I953 (simp7451_0[3:3], comp3_0[9:9], comp3_0[10:10], comp3_0[11:11]);
  C3 I954 (simp7451_0[4:4], comp3_0[12:12], comp3_0[13:13], comp3_0[14:14]);
  C3 I955 (simp7451_0[5:5], comp3_0[15:15], comp3_0[16:16], comp3_0[17:17]);
  C3 I956 (simp7451_0[6:6], comp3_0[18:18], comp3_0[19:19], comp3_0[20:20]);
  C3 I957 (simp7451_0[7:7], comp3_0[21:21], comp3_0[22:22], comp3_0[23:23]);
  C3 I958 (simp7451_0[8:8], comp3_0[24:24], comp3_0[25:25], comp3_0[26:26]);
  C3 I959 (simp7451_0[9:9], comp3_0[27:27], comp3_0[28:28], comp3_0[29:29]);
  C2 I960 (simp7451_0[10:10], comp3_0[30:30], comp3_0[31:31]);
  C3 I961 (simp7452_0[0:0], simp7451_0[0:0], simp7451_0[1:1], simp7451_0[2:2]);
  C3 I962 (simp7452_0[1:1], simp7451_0[3:3], simp7451_0[4:4], simp7451_0[5:5]);
  C3 I963 (simp7452_0[2:2], simp7451_0[6:6], simp7451_0[7:7], simp7451_0[8:8]);
  C2 I964 (simp7452_0[3:3], simp7451_0[9:9], simp7451_0[10:10]);
  C3 I965 (simp7453_0[0:0], simp7452_0[0:0], simp7452_0[1:1], simp7452_0[2:2]);
  BUFF I966 (simp7453_0[1:1], simp7452_0[3:3]);
  C2 I967 (icomp_3, simp7453_0[0:0], simp7453_0[1:1]);
  OR2 I968 (comp4_0[0:0], i_4r0[0:0], i_4r1[0:0]);
  OR2 I969 (comp4_0[1:1], i_4r0[1:1], i_4r1[1:1]);
  OR2 I970 (comp4_0[2:2], i_4r0[2:2], i_4r1[2:2]);
  OR2 I971 (comp4_0[3:3], i_4r0[3:3], i_4r1[3:3]);
  OR2 I972 (comp4_0[4:4], i_4r0[4:4], i_4r1[4:4]);
  OR2 I973 (comp4_0[5:5], i_4r0[5:5], i_4r1[5:5]);
  OR2 I974 (comp4_0[6:6], i_4r0[6:6], i_4r1[6:6]);
  OR2 I975 (comp4_0[7:7], i_4r0[7:7], i_4r1[7:7]);
  OR2 I976 (comp4_0[8:8], i_4r0[8:8], i_4r1[8:8]);
  OR2 I977 (comp4_0[9:9], i_4r0[9:9], i_4r1[9:9]);
  OR2 I978 (comp4_0[10:10], i_4r0[10:10], i_4r1[10:10]);
  OR2 I979 (comp4_0[11:11], i_4r0[11:11], i_4r1[11:11]);
  OR2 I980 (comp4_0[12:12], i_4r0[12:12], i_4r1[12:12]);
  OR2 I981 (comp4_0[13:13], i_4r0[13:13], i_4r1[13:13]);
  OR2 I982 (comp4_0[14:14], i_4r0[14:14], i_4r1[14:14]);
  OR2 I983 (comp4_0[15:15], i_4r0[15:15], i_4r1[15:15]);
  OR2 I984 (comp4_0[16:16], i_4r0[16:16], i_4r1[16:16]);
  OR2 I985 (comp4_0[17:17], i_4r0[17:17], i_4r1[17:17]);
  OR2 I986 (comp4_0[18:18], i_4r0[18:18], i_4r1[18:18]);
  OR2 I987 (comp4_0[19:19], i_4r0[19:19], i_4r1[19:19]);
  OR2 I988 (comp4_0[20:20], i_4r0[20:20], i_4r1[20:20]);
  OR2 I989 (comp4_0[21:21], i_4r0[21:21], i_4r1[21:21]);
  OR2 I990 (comp4_0[22:22], i_4r0[22:22], i_4r1[22:22]);
  OR2 I991 (comp4_0[23:23], i_4r0[23:23], i_4r1[23:23]);
  OR2 I992 (comp4_0[24:24], i_4r0[24:24], i_4r1[24:24]);
  OR2 I993 (comp4_0[25:25], i_4r0[25:25], i_4r1[25:25]);
  OR2 I994 (comp4_0[26:26], i_4r0[26:26], i_4r1[26:26]);
  OR2 I995 (comp4_0[27:27], i_4r0[27:27], i_4r1[27:27]);
  OR2 I996 (comp4_0[28:28], i_4r0[28:28], i_4r1[28:28]);
  OR2 I997 (comp4_0[29:29], i_4r0[29:29], i_4r1[29:29]);
  OR2 I998 (comp4_0[30:30], i_4r0[30:30], i_4r1[30:30]);
  OR2 I999 (comp4_0[31:31], i_4r0[31:31], i_4r1[31:31]);
  C3 I1000 (simp7791_0[0:0], comp4_0[0:0], comp4_0[1:1], comp4_0[2:2]);
  C3 I1001 (simp7791_0[1:1], comp4_0[3:3], comp4_0[4:4], comp4_0[5:5]);
  C3 I1002 (simp7791_0[2:2], comp4_0[6:6], comp4_0[7:7], comp4_0[8:8]);
  C3 I1003 (simp7791_0[3:3], comp4_0[9:9], comp4_0[10:10], comp4_0[11:11]);
  C3 I1004 (simp7791_0[4:4], comp4_0[12:12], comp4_0[13:13], comp4_0[14:14]);
  C3 I1005 (simp7791_0[5:5], comp4_0[15:15], comp4_0[16:16], comp4_0[17:17]);
  C3 I1006 (simp7791_0[6:6], comp4_0[18:18], comp4_0[19:19], comp4_0[20:20]);
  C3 I1007 (simp7791_0[7:7], comp4_0[21:21], comp4_0[22:22], comp4_0[23:23]);
  C3 I1008 (simp7791_0[8:8], comp4_0[24:24], comp4_0[25:25], comp4_0[26:26]);
  C3 I1009 (simp7791_0[9:9], comp4_0[27:27], comp4_0[28:28], comp4_0[29:29]);
  C2 I1010 (simp7791_0[10:10], comp4_0[30:30], comp4_0[31:31]);
  C3 I1011 (simp7792_0[0:0], simp7791_0[0:0], simp7791_0[1:1], simp7791_0[2:2]);
  C3 I1012 (simp7792_0[1:1], simp7791_0[3:3], simp7791_0[4:4], simp7791_0[5:5]);
  C3 I1013 (simp7792_0[2:2], simp7791_0[6:6], simp7791_0[7:7], simp7791_0[8:8]);
  C2 I1014 (simp7792_0[3:3], simp7791_0[9:9], simp7791_0[10:10]);
  C3 I1015 (simp7793_0[0:0], simp7792_0[0:0], simp7792_0[1:1], simp7792_0[2:2]);
  BUFF I1016 (simp7793_0[1:1], simp7792_0[3:3]);
  C2 I1017 (icomp_4, simp7793_0[0:0], simp7793_0[1:1]);
  OR2 I1018 (comp5_0[0:0], i_5r0[0:0], i_5r1[0:0]);
  OR2 I1019 (comp5_0[1:1], i_5r0[1:1], i_5r1[1:1]);
  OR2 I1020 (comp5_0[2:2], i_5r0[2:2], i_5r1[2:2]);
  OR2 I1021 (comp5_0[3:3], i_5r0[3:3], i_5r1[3:3]);
  OR2 I1022 (comp5_0[4:4], i_5r0[4:4], i_5r1[4:4]);
  OR2 I1023 (comp5_0[5:5], i_5r0[5:5], i_5r1[5:5]);
  OR2 I1024 (comp5_0[6:6], i_5r0[6:6], i_5r1[6:6]);
  OR2 I1025 (comp5_0[7:7], i_5r0[7:7], i_5r1[7:7]);
  OR2 I1026 (comp5_0[8:8], i_5r0[8:8], i_5r1[8:8]);
  OR2 I1027 (comp5_0[9:9], i_5r0[9:9], i_5r1[9:9]);
  OR2 I1028 (comp5_0[10:10], i_5r0[10:10], i_5r1[10:10]);
  OR2 I1029 (comp5_0[11:11], i_5r0[11:11], i_5r1[11:11]);
  OR2 I1030 (comp5_0[12:12], i_5r0[12:12], i_5r1[12:12]);
  OR2 I1031 (comp5_0[13:13], i_5r0[13:13], i_5r1[13:13]);
  OR2 I1032 (comp5_0[14:14], i_5r0[14:14], i_5r1[14:14]);
  OR2 I1033 (comp5_0[15:15], i_5r0[15:15], i_5r1[15:15]);
  OR2 I1034 (comp5_0[16:16], i_5r0[16:16], i_5r1[16:16]);
  OR2 I1035 (comp5_0[17:17], i_5r0[17:17], i_5r1[17:17]);
  OR2 I1036 (comp5_0[18:18], i_5r0[18:18], i_5r1[18:18]);
  OR2 I1037 (comp5_0[19:19], i_5r0[19:19], i_5r1[19:19]);
  OR2 I1038 (comp5_0[20:20], i_5r0[20:20], i_5r1[20:20]);
  OR2 I1039 (comp5_0[21:21], i_5r0[21:21], i_5r1[21:21]);
  OR2 I1040 (comp5_0[22:22], i_5r0[22:22], i_5r1[22:22]);
  OR2 I1041 (comp5_0[23:23], i_5r0[23:23], i_5r1[23:23]);
  OR2 I1042 (comp5_0[24:24], i_5r0[24:24], i_5r1[24:24]);
  OR2 I1043 (comp5_0[25:25], i_5r0[25:25], i_5r1[25:25]);
  OR2 I1044 (comp5_0[26:26], i_5r0[26:26], i_5r1[26:26]);
  OR2 I1045 (comp5_0[27:27], i_5r0[27:27], i_5r1[27:27]);
  OR2 I1046 (comp5_0[28:28], i_5r0[28:28], i_5r1[28:28]);
  OR2 I1047 (comp5_0[29:29], i_5r0[29:29], i_5r1[29:29]);
  OR2 I1048 (comp5_0[30:30], i_5r0[30:30], i_5r1[30:30]);
  OR2 I1049 (comp5_0[31:31], i_5r0[31:31], i_5r1[31:31]);
  C3 I1050 (simp8131_0[0:0], comp5_0[0:0], comp5_0[1:1], comp5_0[2:2]);
  C3 I1051 (simp8131_0[1:1], comp5_0[3:3], comp5_0[4:4], comp5_0[5:5]);
  C3 I1052 (simp8131_0[2:2], comp5_0[6:6], comp5_0[7:7], comp5_0[8:8]);
  C3 I1053 (simp8131_0[3:3], comp5_0[9:9], comp5_0[10:10], comp5_0[11:11]);
  C3 I1054 (simp8131_0[4:4], comp5_0[12:12], comp5_0[13:13], comp5_0[14:14]);
  C3 I1055 (simp8131_0[5:5], comp5_0[15:15], comp5_0[16:16], comp5_0[17:17]);
  C3 I1056 (simp8131_0[6:6], comp5_0[18:18], comp5_0[19:19], comp5_0[20:20]);
  C3 I1057 (simp8131_0[7:7], comp5_0[21:21], comp5_0[22:22], comp5_0[23:23]);
  C3 I1058 (simp8131_0[8:8], comp5_0[24:24], comp5_0[25:25], comp5_0[26:26]);
  C3 I1059 (simp8131_0[9:9], comp5_0[27:27], comp5_0[28:28], comp5_0[29:29]);
  C2 I1060 (simp8131_0[10:10], comp5_0[30:30], comp5_0[31:31]);
  C3 I1061 (simp8132_0[0:0], simp8131_0[0:0], simp8131_0[1:1], simp8131_0[2:2]);
  C3 I1062 (simp8132_0[1:1], simp8131_0[3:3], simp8131_0[4:4], simp8131_0[5:5]);
  C3 I1063 (simp8132_0[2:2], simp8131_0[6:6], simp8131_0[7:7], simp8131_0[8:8]);
  C2 I1064 (simp8132_0[3:3], simp8131_0[9:9], simp8131_0[10:10]);
  C3 I1065 (simp8133_0[0:0], simp8132_0[0:0], simp8132_0[1:1], simp8132_0[2:2]);
  BUFF I1066 (simp8133_0[1:1], simp8132_0[3:3]);
  C2 I1067 (icomp_5, simp8133_0[0:0], simp8133_0[1:1]);
  OR2 I1068 (comp6_0[0:0], i_6r0[0:0], i_6r1[0:0]);
  OR2 I1069 (comp6_0[1:1], i_6r0[1:1], i_6r1[1:1]);
  OR2 I1070 (comp6_0[2:2], i_6r0[2:2], i_6r1[2:2]);
  OR2 I1071 (comp6_0[3:3], i_6r0[3:3], i_6r1[3:3]);
  OR2 I1072 (comp6_0[4:4], i_6r0[4:4], i_6r1[4:4]);
  OR2 I1073 (comp6_0[5:5], i_6r0[5:5], i_6r1[5:5]);
  OR2 I1074 (comp6_0[6:6], i_6r0[6:6], i_6r1[6:6]);
  OR2 I1075 (comp6_0[7:7], i_6r0[7:7], i_6r1[7:7]);
  OR2 I1076 (comp6_0[8:8], i_6r0[8:8], i_6r1[8:8]);
  OR2 I1077 (comp6_0[9:9], i_6r0[9:9], i_6r1[9:9]);
  OR2 I1078 (comp6_0[10:10], i_6r0[10:10], i_6r1[10:10]);
  OR2 I1079 (comp6_0[11:11], i_6r0[11:11], i_6r1[11:11]);
  OR2 I1080 (comp6_0[12:12], i_6r0[12:12], i_6r1[12:12]);
  OR2 I1081 (comp6_0[13:13], i_6r0[13:13], i_6r1[13:13]);
  OR2 I1082 (comp6_0[14:14], i_6r0[14:14], i_6r1[14:14]);
  OR2 I1083 (comp6_0[15:15], i_6r0[15:15], i_6r1[15:15]);
  OR2 I1084 (comp6_0[16:16], i_6r0[16:16], i_6r1[16:16]);
  OR2 I1085 (comp6_0[17:17], i_6r0[17:17], i_6r1[17:17]);
  OR2 I1086 (comp6_0[18:18], i_6r0[18:18], i_6r1[18:18]);
  OR2 I1087 (comp6_0[19:19], i_6r0[19:19], i_6r1[19:19]);
  OR2 I1088 (comp6_0[20:20], i_6r0[20:20], i_6r1[20:20]);
  OR2 I1089 (comp6_0[21:21], i_6r0[21:21], i_6r1[21:21]);
  OR2 I1090 (comp6_0[22:22], i_6r0[22:22], i_6r1[22:22]);
  OR2 I1091 (comp6_0[23:23], i_6r0[23:23], i_6r1[23:23]);
  OR2 I1092 (comp6_0[24:24], i_6r0[24:24], i_6r1[24:24]);
  OR2 I1093 (comp6_0[25:25], i_6r0[25:25], i_6r1[25:25]);
  OR2 I1094 (comp6_0[26:26], i_6r0[26:26], i_6r1[26:26]);
  OR2 I1095 (comp6_0[27:27], i_6r0[27:27], i_6r1[27:27]);
  OR2 I1096 (comp6_0[28:28], i_6r0[28:28], i_6r1[28:28]);
  OR2 I1097 (comp6_0[29:29], i_6r0[29:29], i_6r1[29:29]);
  OR2 I1098 (comp6_0[30:30], i_6r0[30:30], i_6r1[30:30]);
  OR2 I1099 (comp6_0[31:31], i_6r0[31:31], i_6r1[31:31]);
  C3 I1100 (simp8471_0[0:0], comp6_0[0:0], comp6_0[1:1], comp6_0[2:2]);
  C3 I1101 (simp8471_0[1:1], comp6_0[3:3], comp6_0[4:4], comp6_0[5:5]);
  C3 I1102 (simp8471_0[2:2], comp6_0[6:6], comp6_0[7:7], comp6_0[8:8]);
  C3 I1103 (simp8471_0[3:3], comp6_0[9:9], comp6_0[10:10], comp6_0[11:11]);
  C3 I1104 (simp8471_0[4:4], comp6_0[12:12], comp6_0[13:13], comp6_0[14:14]);
  C3 I1105 (simp8471_0[5:5], comp6_0[15:15], comp6_0[16:16], comp6_0[17:17]);
  C3 I1106 (simp8471_0[6:6], comp6_0[18:18], comp6_0[19:19], comp6_0[20:20]);
  C3 I1107 (simp8471_0[7:7], comp6_0[21:21], comp6_0[22:22], comp6_0[23:23]);
  C3 I1108 (simp8471_0[8:8], comp6_0[24:24], comp6_0[25:25], comp6_0[26:26]);
  C3 I1109 (simp8471_0[9:9], comp6_0[27:27], comp6_0[28:28], comp6_0[29:29]);
  C2 I1110 (simp8471_0[10:10], comp6_0[30:30], comp6_0[31:31]);
  C3 I1111 (simp8472_0[0:0], simp8471_0[0:0], simp8471_0[1:1], simp8471_0[2:2]);
  C3 I1112 (simp8472_0[1:1], simp8471_0[3:3], simp8471_0[4:4], simp8471_0[5:5]);
  C3 I1113 (simp8472_0[2:2], simp8471_0[6:6], simp8471_0[7:7], simp8471_0[8:8]);
  C2 I1114 (simp8472_0[3:3], simp8471_0[9:9], simp8471_0[10:10]);
  C3 I1115 (simp8473_0[0:0], simp8472_0[0:0], simp8472_0[1:1], simp8472_0[2:2]);
  BUFF I1116 (simp8473_0[1:1], simp8472_0[3:3]);
  C2 I1117 (icomp_6, simp8473_0[0:0], simp8473_0[1:1]);
  OR2 I1118 (comp7_0[0:0], i_7r0[0:0], i_7r1[0:0]);
  OR2 I1119 (comp7_0[1:1], i_7r0[1:1], i_7r1[1:1]);
  OR2 I1120 (comp7_0[2:2], i_7r0[2:2], i_7r1[2:2]);
  OR2 I1121 (comp7_0[3:3], i_7r0[3:3], i_7r1[3:3]);
  OR2 I1122 (comp7_0[4:4], i_7r0[4:4], i_7r1[4:4]);
  OR2 I1123 (comp7_0[5:5], i_7r0[5:5], i_7r1[5:5]);
  OR2 I1124 (comp7_0[6:6], i_7r0[6:6], i_7r1[6:6]);
  OR2 I1125 (comp7_0[7:7], i_7r0[7:7], i_7r1[7:7]);
  OR2 I1126 (comp7_0[8:8], i_7r0[8:8], i_7r1[8:8]);
  OR2 I1127 (comp7_0[9:9], i_7r0[9:9], i_7r1[9:9]);
  OR2 I1128 (comp7_0[10:10], i_7r0[10:10], i_7r1[10:10]);
  OR2 I1129 (comp7_0[11:11], i_7r0[11:11], i_7r1[11:11]);
  OR2 I1130 (comp7_0[12:12], i_7r0[12:12], i_7r1[12:12]);
  OR2 I1131 (comp7_0[13:13], i_7r0[13:13], i_7r1[13:13]);
  OR2 I1132 (comp7_0[14:14], i_7r0[14:14], i_7r1[14:14]);
  OR2 I1133 (comp7_0[15:15], i_7r0[15:15], i_7r1[15:15]);
  OR2 I1134 (comp7_0[16:16], i_7r0[16:16], i_7r1[16:16]);
  OR2 I1135 (comp7_0[17:17], i_7r0[17:17], i_7r1[17:17]);
  OR2 I1136 (comp7_0[18:18], i_7r0[18:18], i_7r1[18:18]);
  OR2 I1137 (comp7_0[19:19], i_7r0[19:19], i_7r1[19:19]);
  OR2 I1138 (comp7_0[20:20], i_7r0[20:20], i_7r1[20:20]);
  OR2 I1139 (comp7_0[21:21], i_7r0[21:21], i_7r1[21:21]);
  OR2 I1140 (comp7_0[22:22], i_7r0[22:22], i_7r1[22:22]);
  OR2 I1141 (comp7_0[23:23], i_7r0[23:23], i_7r1[23:23]);
  OR2 I1142 (comp7_0[24:24], i_7r0[24:24], i_7r1[24:24]);
  OR2 I1143 (comp7_0[25:25], i_7r0[25:25], i_7r1[25:25]);
  OR2 I1144 (comp7_0[26:26], i_7r0[26:26], i_7r1[26:26]);
  OR2 I1145 (comp7_0[27:27], i_7r0[27:27], i_7r1[27:27]);
  OR2 I1146 (comp7_0[28:28], i_7r0[28:28], i_7r1[28:28]);
  OR2 I1147 (comp7_0[29:29], i_7r0[29:29], i_7r1[29:29]);
  OR2 I1148 (comp7_0[30:30], i_7r0[30:30], i_7r1[30:30]);
  OR2 I1149 (comp7_0[31:31], i_7r0[31:31], i_7r1[31:31]);
  C3 I1150 (simp8811_0[0:0], comp7_0[0:0], comp7_0[1:1], comp7_0[2:2]);
  C3 I1151 (simp8811_0[1:1], comp7_0[3:3], comp7_0[4:4], comp7_0[5:5]);
  C3 I1152 (simp8811_0[2:2], comp7_0[6:6], comp7_0[7:7], comp7_0[8:8]);
  C3 I1153 (simp8811_0[3:3], comp7_0[9:9], comp7_0[10:10], comp7_0[11:11]);
  C3 I1154 (simp8811_0[4:4], comp7_0[12:12], comp7_0[13:13], comp7_0[14:14]);
  C3 I1155 (simp8811_0[5:5], comp7_0[15:15], comp7_0[16:16], comp7_0[17:17]);
  C3 I1156 (simp8811_0[6:6], comp7_0[18:18], comp7_0[19:19], comp7_0[20:20]);
  C3 I1157 (simp8811_0[7:7], comp7_0[21:21], comp7_0[22:22], comp7_0[23:23]);
  C3 I1158 (simp8811_0[8:8], comp7_0[24:24], comp7_0[25:25], comp7_0[26:26]);
  C3 I1159 (simp8811_0[9:9], comp7_0[27:27], comp7_0[28:28], comp7_0[29:29]);
  C2 I1160 (simp8811_0[10:10], comp7_0[30:30], comp7_0[31:31]);
  C3 I1161 (simp8812_0[0:0], simp8811_0[0:0], simp8811_0[1:1], simp8811_0[2:2]);
  C3 I1162 (simp8812_0[1:1], simp8811_0[3:3], simp8811_0[4:4], simp8811_0[5:5]);
  C3 I1163 (simp8812_0[2:2], simp8811_0[6:6], simp8811_0[7:7], simp8811_0[8:8]);
  C2 I1164 (simp8812_0[3:3], simp8811_0[9:9], simp8811_0[10:10]);
  C3 I1165 (simp8813_0[0:0], simp8812_0[0:0], simp8812_0[1:1], simp8812_0[2:2]);
  BUFF I1166 (simp8813_0[1:1], simp8812_0[3:3]);
  C2 I1167 (icomp_7, simp8813_0[0:0], simp8813_0[1:1]);
  C2R I1168 (choice_0, icomp_0, nchosen_0, reset);
  C2R I1169 (choice_1, icomp_1, nchosen_0, reset);
  C2R I1170 (choice_2, icomp_2, nchosen_0, reset);
  C2R I1171 (choice_3, icomp_3, nchosen_0, reset);
  C2R I1172 (choice_4, icomp_4, nchosen_0, reset);
  C2R I1173 (choice_5, icomp_5, nchosen_0, reset);
  C2R I1174 (choice_6, icomp_6, nchosen_0, reset);
  C2R I1175 (choice_7, icomp_7, nchosen_0, reset);
  NOR3 I1176 (simp8901_0[0:0], choice_0, choice_1, choice_2);
  NOR3 I1177 (simp8901_0[1:1], choice_3, choice_4, choice_5);
  NOR2 I1178 (simp8901_0[2:2], choice_6, choice_7);
  NAND3 I1179 (anychoice_0, simp8901_0[0:0], simp8901_0[1:1], simp8901_0[2:2]);
  NOR2 I1180 (nchosen_0, anychoice_0, o_0a);
  C2R I1181 (i_0a, choice_0, o_0a, reset);
  C2R I1182 (i_1a, choice_1, o_0a, reset);
  C2R I1183 (i_2a, choice_2, o_0a, reset);
  C2R I1184 (i_3a, choice_3, o_0a, reset);
  C2R I1185 (i_4a, choice_4, o_0a, reset);
  C2R I1186 (i_5a, choice_5, o_0a, reset);
  C2R I1187 (i_6a, choice_6, o_0a, reset);
  C2R I1188 (i_7a, choice_7, o_0a, reset);
endmodule

// tko2m2_1api0w1b_2api1w1b_3nm1b0_4apt1o0w1bt3o0w1b_5nm1b0_6apt2o0w1bt5o0w1b_7addt4o0w2bt6o0w2b TeakO 
//   [
//     (1,TeakOAppend 1 [(0,0+:1)]),
//     (2,TeakOAppend 1 [(0,1+:1)]),
//     (3,TeakOConstant 1 0),
//     (4,TeakOAppend 1 [(1,0+:1),(3,0+:1)]),
//     (5,TeakOConstant 1 0),
//     (6,TeakOAppend 1 [(2,0+:1),(5,0+:1)]),
//     (7,TeakOp TeakOpAdd [(4,0+:2),(6,0+:2)])] [One 2,One 2]
module tko2m2_1api0w1b_2api1w1b_3nm1b0_4apt1o0w1bt3o0w1b_5nm1b0_6apt2o0w1bt5o0w1b_7addt4o0w2bt6o0w2b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [1:0] gocomp_0;
  wire termf_1;
  wire termf_2;
  wire termf_3;
  wire [1:0] termf_4;
  wire termf_5;
  wire [1:0] termf_6;
  wire termt_1;
  wire termt_2;
  wire termt_3;
  wire [1:0] termt_4;
  wire termt_5;
  wire [1:0] termt_6;
  wire [1:0] cf7__0;
  wire [1:0] ct7__0;
  wire [3:0] ha7__0;
  wire [7:0] fa7_1min_0;
  wire [1:0] simp551_0;
  wire [1:0] simp561_0;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  C2 I2 (go_0, gocomp_0[0:0], gocomp_0[1:1]);
  BUFF I3 (termf_1, i_0r0[0:0]);
  BUFF I4 (termt_1, i_0r1[0:0]);
  BUFF I5 (termf_2, i_0r0[1:1]);
  BUFF I6 (termt_2, i_0r1[1:1]);
  BUFF I7 (termf_3, go_0);
  GND I8 (termt_3);
  BUFF I9 (termf_4[0:0], termf_1);
  BUFF I10 (termf_4[1:1], termf_3);
  BUFF I11 (termt_4[0:0], termt_1);
  BUFF I12 (termt_4[1:1], termt_3);
  BUFF I13 (termf_5, go_0);
  GND I14 (termt_5);
  BUFF I15 (termf_6[0:0], termf_2);
  BUFF I16 (termf_6[1:1], termf_5);
  BUFF I17 (termt_6[0:0], termt_2);
  BUFF I18 (termt_6[1:1], termt_5);
  C2 I19 (ha7__0[0:0], termf_6[0:0], termf_4[0:0]);
  C2 I20 (ha7__0[1:1], termf_6[0:0], termt_4[0:0]);
  C2 I21 (ha7__0[2:2], termt_6[0:0], termf_4[0:0]);
  C2 I22 (ha7__0[3:3], termt_6[0:0], termt_4[0:0]);
  OR3 I23 (cf7__0[0:0], ha7__0[0:0], ha7__0[1:1], ha7__0[2:2]);
  BUFF I24 (ct7__0[0:0], ha7__0[3:3]);
  OR2 I25 (o_0r0[0:0], ha7__0[0:0], ha7__0[3:3]);
  OR2 I26 (o_0r1[0:0], ha7__0[1:1], ha7__0[2:2]);
  C3 I27 (fa7_1min_0[0:0], cf7__0[0:0], termf_6[1:1], termf_4[1:1]);
  C3 I28 (fa7_1min_0[1:1], cf7__0[0:0], termf_6[1:1], termt_4[1:1]);
  C3 I29 (fa7_1min_0[2:2], cf7__0[0:0], termt_6[1:1], termf_4[1:1]);
  C3 I30 (fa7_1min_0[3:3], cf7__0[0:0], termt_6[1:1], termt_4[1:1]);
  C3 I31 (fa7_1min_0[4:4], ct7__0[0:0], termf_6[1:1], termf_4[1:1]);
  C3 I32 (fa7_1min_0[5:5], ct7__0[0:0], termf_6[1:1], termt_4[1:1]);
  C3 I33 (fa7_1min_0[6:6], ct7__0[0:0], termt_6[1:1], termf_4[1:1]);
  C3 I34 (fa7_1min_0[7:7], ct7__0[0:0], termt_6[1:1], termt_4[1:1]);
  NOR3 I35 (simp551_0[0:0], fa7_1min_0[0:0], fa7_1min_0[3:3], fa7_1min_0[5:5]);
  INV I36 (simp551_0[1:1], fa7_1min_0[6:6]);
  NAND2 I37 (o_0r0[1:1], simp551_0[0:0], simp551_0[1:1]);
  NOR3 I38 (simp561_0[0:0], fa7_1min_0[1:1], fa7_1min_0[2:2], fa7_1min_0[4:4]);
  INV I39 (simp561_0[1:1], fa7_1min_0[7:7]);
  NAND2 I40 (o_0r1[1:1], simp561_0[0:0], simp561_0[1:1]);
  AO222 I41 (ct7__0[1:1], termt_4[1:1], termt_6[1:1], termt_4[1:1], ct7__0[0:0], termt_6[1:1], ct7__0[0:0]);
  AO222 I42 (cf7__0[1:1], termf_4[1:1], termf_6[1:1], termf_4[1:1], cf7__0[0:0], termf_6[1:1], cf7__0[0:0]);
  BUFF I43 (i_0a, o_0a);
endmodule

// tkf2mo0w1 TeakF [0] [One 2,Many [1]]
module tkf2mo0w1 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  wire ucomplete_0;
  wire comp_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (comp_0, i_0r0[1:1], i_0r1[1:1]);
  BUFF I2 (ucomplete_0, comp_0);
  C2 I3 (acomplete_0, ucomplete_0, icomplete_0);
  C2 I4 (o_0r0, i_0r0[0:0], icomplete_0);
  C2 I5 (o_0r1, i_0r1[0:0], icomplete_0);
  C2 I6 (i_0a, acomplete_0, o_0a);
endmodule

// tks5_o0w5_0o0w0_1m2c1m4c3o0w0_8c7o0w0_10c7o0w0_18c7o0w0 TeakS (0+:5) [([Imp 0 0],0),([Imp 1 0,Imp 2 
//   1,Imp 4 3],0),([Imp 8 7],0),([Imp 16 7],0),([Imp 24 7],0)] [One 5,Many [0,0,0,0,0]]
module tks5_o0w5_0o0w0_1m2c1m4c3o0w0_8c7o0w0_10c7o0w0_18c7o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, reset);
  input [4:0] i_0r0;
  input [4:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire sel_4;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire gsel_4;
  wire oack_0;
  wire match0_0;
  wire [1:0] simp141_0;
  wire [2:0] match1_0;
  wire [1:0] simp171_0;
  wire [1:0] simp181_0;
  wire match2_0;
  wire match3_0;
  wire match4_0;
  wire [4:0] comp_0;
  wire [1:0] simp401_0;
  wire [1:0] simp461_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (simp141_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C2 I2 (simp141_0[1:1], i_0r0[3:3], i_0r0[4:4]);
  C2 I3 (match0_0, simp141_0[0:0], simp141_0[1:1]);
  OR3 I4 (sel_1, match1_0[0:0], match1_0[1:1], match1_0[2:2]);
  C3 I5 (simp171_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C2 I6 (simp171_0[1:1], i_0r0[3:3], i_0r0[4:4]);
  C2 I7 (match1_0[0:0], simp171_0[0:0], simp171_0[1:1]);
  C3 I8 (simp181_0[0:0], i_0r1[1:1], i_0r0[2:2], i_0r0[3:3]);
  BUFF I9 (simp181_0[1:1], i_0r0[4:4]);
  C2 I10 (match1_0[1:1], simp181_0[0:0], simp181_0[1:1]);
  C3 I11 (match1_0[2:2], i_0r1[2:2], i_0r0[3:3], i_0r0[4:4]);
  BUFF I12 (sel_2, match2_0);
  C2 I13 (match2_0, i_0r1[3:3], i_0r0[4:4]);
  BUFF I14 (sel_3, match3_0);
  C2 I15 (match3_0, i_0r0[3:3], i_0r1[4:4]);
  BUFF I16 (sel_4, match4_0);
  C2 I17 (match4_0, i_0r1[3:3], i_0r1[4:4]);
  C2 I18 (gsel_0, sel_0, icomplete_0);
  C2 I19 (gsel_1, sel_1, icomplete_0);
  C2 I20 (gsel_2, sel_2, icomplete_0);
  C2 I21 (gsel_3, sel_3, icomplete_0);
  C2 I22 (gsel_4, sel_4, icomplete_0);
  OR2 I23 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I24 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I25 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I26 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I27 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  C3 I28 (simp401_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C2 I29 (simp401_0[1:1], comp_0[3:3], comp_0[4:4]);
  C2 I30 (icomplete_0, simp401_0[0:0], simp401_0[1:1]);
  BUFF I31 (o_0r, gsel_0);
  BUFF I32 (o_1r, gsel_1);
  BUFF I33 (o_2r, gsel_2);
  BUFF I34 (o_3r, gsel_3);
  BUFF I35 (o_4r, gsel_4);
  NOR3 I36 (simp461_0[0:0], o_0a, o_1a, o_2a);
  NOR2 I37 (simp461_0[1:1], o_3a, o_4a);
  NAND2 I38 (oack_0, simp461_0[0:0], simp461_0[1:1]);
  C2 I39 (i_0a, oack_0, icomplete_0);
endmodule

// tkm5x0b TeakM [Many [0,0,0,0,0],One 0]
module tkm5x0b (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, i_3r, i_3a, i_4r, i_4a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  input i_4r;
  output i_4a;
  output o_0r;
  input o_0a;
  input reset;
  wire nchosen_0;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire choice_4;
  wire [1:0] simp121_0;
  C2R I0 (choice_0, i_0r, nchosen_0, reset);
  C2R I1 (choice_1, i_1r, nchosen_0, reset);
  C2R I2 (choice_2, i_2r, nchosen_0, reset);
  C2R I3 (choice_3, i_3r, nchosen_0, reset);
  C2R I4 (choice_4, i_4r, nchosen_0, reset);
  NOR2 I5 (nchosen_0, o_0r, o_0a);
  NOR3 I6 (simp121_0[0:0], choice_0, choice_1, choice_2);
  NOR2 I7 (simp121_0[1:1], choice_3, choice_4);
  NAND2 I8 (o_0r, simp121_0[0:0], simp121_0[1:1]);
  C2R I9 (i_0a, choice_0, o_0a, reset);
  C2R I10 (i_1a, choice_1, o_0a, reset);
  C2R I11 (i_2a, choice_2, o_0a, reset);
  C2R I12 (i_3a, choice_3, o_0a, reset);
  C2R I13 (i_4a, choice_4, o_0a, reset);
endmodule

// tkvsel5_wo0w5_ro0w5o0w3o0w3o0w3o0w3 TeakV "sel" 5 [] [0] [0,0,0,0,0] [Many [5],Many [0],Many [0,0,0,
//   0,0],Many [5,3,3,3,3]]
module tkvsel5_wo0w5_ro0w5o0w3o0w3o0w3o0w3 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, reset);
  input [4:0] wg_0r0;
  input [4:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  output [4:0] rd_0r0;
  output [4:0] rd_0r1;
  input rd_0a;
  output [2:0] rd_1r0;
  output [2:0] rd_1r1;
  input rd_1a;
  output [2:0] rd_2r0;
  output [2:0] rd_2r1;
  input rd_2a;
  output [2:0] rd_3r0;
  output [2:0] rd_3r1;
  input rd_3a;
  output [2:0] rd_4r0;
  output [2:0] rd_4r1;
  input rd_4a;
  input reset;
  wire [4:0] wf_0;
  wire [4:0] wt_0;
  wire [4:0] df_0;
  wire [4:0] dt_0;
  wire wc_0;
  wire [4:0] wacks_0;
  wire [4:0] wenr_0;
  wire [4:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [4:0] drlgf_0;
  wire [4:0] drlgt_0;
  wire [4:0] comp0_0;
  wire [1:0] simp491_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [4:0] conwgit_0;
  wire [4:0] conwgif_0;
  wire conwig_0;
  wire [1:0] simp831_0;
  wire [3:0] simp1181_0;
  wire [1:0] simp1182_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I7 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I8 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I9 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I10 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I11 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I12 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I13 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I14 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I15 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  NOR2 I16 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I17 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I18 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I19 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I20 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR3 I21 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I22 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I23 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I24 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I25 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  AO22 I26 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I27 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I28 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I29 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I30 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  OR2 I31 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I32 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I33 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I34 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I35 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  C3 I36 (simp491_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C2 I37 (simp491_0[1:1], comp0_0[3:3], comp0_0[4:4]);
  C2 I38 (wc_0, simp491_0[0:0], simp491_0[1:1]);
  AND2 I39 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I40 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I41 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I42 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I43 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I44 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I45 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I46 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I47 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I48 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  BUFF I49 (conwigc_0, wc_0);
  AO22 I50 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I51 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I52 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I53 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I54 (wenr_0[0:0], wc_0);
  BUFF I55 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I56 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I57 (wenr_0[1:1], wc_0);
  BUFF I58 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I59 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I60 (wenr_0[2:2], wc_0);
  BUFF I61 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I62 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I63 (wenr_0[3:3], wc_0);
  BUFF I64 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I65 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I66 (wenr_0[4:4], wc_0);
  C3 I67 (simp831_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I68 (simp831_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C2 I69 (wd_0r, simp831_0[0:0], simp831_0[1:1]);
  AND2 I70 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I71 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I72 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I73 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I74 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I75 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I76 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I77 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I78 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I79 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I80 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I81 (rd_3r0[0:0], df_0[0:0], rg_3r);
  AND2 I82 (rd_3r0[1:1], df_0[1:1], rg_3r);
  AND2 I83 (rd_3r0[2:2], df_0[2:2], rg_3r);
  AND2 I84 (rd_4r0[0:0], df_0[0:0], rg_4r);
  AND2 I85 (rd_4r0[1:1], df_0[1:1], rg_4r);
  AND2 I86 (rd_4r0[2:2], df_0[2:2], rg_4r);
  AND2 I87 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I88 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I89 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I90 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I91 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I92 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I93 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I94 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I95 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I96 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I97 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I98 (rd_3r1[0:0], dt_0[0:0], rg_3r);
  AND2 I99 (rd_3r1[1:1], dt_0[1:1], rg_3r);
  AND2 I100 (rd_3r1[2:2], dt_0[2:2], rg_3r);
  AND2 I101 (rd_4r1[0:0], dt_0[0:0], rg_4r);
  AND2 I102 (rd_4r1[1:1], dt_0[1:1], rg_4r);
  AND2 I103 (rd_4r1[2:2], dt_0[2:2], rg_4r);
  NOR3 I104 (simp1181_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I105 (simp1181_0[1:1], rg_3r, rg_4r, rg_0a);
  NOR3 I106 (simp1181_0[2:2], rg_1a, rg_2a, rg_3a);
  INV I107 (simp1181_0[3:3], rg_4a);
  NAND3 I108 (simp1182_0[0:0], simp1181_0[0:0], simp1181_0[1:1], simp1181_0[2:2]);
  INV I109 (simp1182_0[1:1], simp1181_0[3:3]);
  OR2 I110 (anyread_0, simp1182_0[0:0], simp1182_0[1:1]);
  BUFF I111 (wg_0a, wd_0a);
  BUFF I112 (rg_0a, rd_0a);
  BUFF I113 (rg_1a, rd_1a);
  BUFF I114 (rg_2a, rd_2a);
  BUFF I115 (rg_3a, rd_3a);
  BUFF I116 (rg_4a, rd_4a);
endmodule

// tks35_o32w3_1o0w32_2o0w32_3o0w32_4o0w32_5o0w32_6o0w32_7o0w32 TeakS (32+:3) [([Imp 1 0],0),([Imp 2 0]
//   ,0),([Imp 3 0],0),([Imp 4 0],0),([Imp 5 0],0),([Imp 6 0],0),([Imp 7 0],0)] [One 35,Many [32,32,32,32
//   ,32,32,32]]
module tks35_o32w3_1o0w32_2o0w32_3o0w32_4o0w32_5o0w32_6o0w32_7o0w32 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r0, o_1r1, o_1a, o_2r0, o_2r1, o_2a, o_3r0, o_3r1, o_3a, o_4r0, o_4r1, o_4a, o_5r0, o_5r1, o_5a, o_6r0, o_6r1, o_6a, reset);
  input [34:0] i_0r0;
  input [34:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  output [31:0] o_1r0;
  output [31:0] o_1r1;
  input o_1a;
  output [31:0] o_2r0;
  output [31:0] o_2r1;
  input o_2a;
  output [31:0] o_3r0;
  output [31:0] o_3r1;
  input o_3a;
  output [31:0] o_4r0;
  output [31:0] o_4r1;
  input o_4a;
  output [31:0] o_5r0;
  output [31:0] o_5r1;
  input o_5a;
  output [31:0] o_6r0;
  output [31:0] o_6r1;
  input o_6a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire sel_4;
  wire sel_5;
  wire sel_6;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire gsel_4;
  wire gsel_5;
  wire gsel_6;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire match2_0;
  wire match3_0;
  wire match4_0;
  wire match5_0;
  wire match6_0;
  wire [34:0] comp_0;
  wire [11:0] simp801_0;
  wire [3:0] simp802_0;
  wire [1:0] simp803_0;
  wire [2:0] simp5291_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (match0_0, i_0r1[32:32], i_0r0[33:33], i_0r0[34:34]);
  BUFF I2 (sel_1, match1_0);
  C3 I3 (match1_0, i_0r0[32:32], i_0r1[33:33], i_0r0[34:34]);
  BUFF I4 (sel_2, match2_0);
  C3 I5 (match2_0, i_0r1[32:32], i_0r1[33:33], i_0r0[34:34]);
  BUFF I6 (sel_3, match3_0);
  C3 I7 (match3_0, i_0r0[32:32], i_0r0[33:33], i_0r1[34:34]);
  BUFF I8 (sel_4, match4_0);
  C3 I9 (match4_0, i_0r1[32:32], i_0r0[33:33], i_0r1[34:34]);
  BUFF I10 (sel_5, match5_0);
  C3 I11 (match5_0, i_0r0[32:32], i_0r1[33:33], i_0r1[34:34]);
  BUFF I12 (sel_6, match6_0);
  C3 I13 (match6_0, i_0r1[32:32], i_0r1[33:33], i_0r1[34:34]);
  C2 I14 (gsel_0, sel_0, icomplete_0);
  C2 I15 (gsel_1, sel_1, icomplete_0);
  C2 I16 (gsel_2, sel_2, icomplete_0);
  C2 I17 (gsel_3, sel_3, icomplete_0);
  C2 I18 (gsel_4, sel_4, icomplete_0);
  C2 I19 (gsel_5, sel_5, icomplete_0);
  C2 I20 (gsel_6, sel_6, icomplete_0);
  OR2 I21 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I22 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I23 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I24 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I25 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I26 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I27 (comp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I28 (comp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I29 (comp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I30 (comp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I31 (comp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I32 (comp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I33 (comp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I34 (comp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I35 (comp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I36 (comp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I37 (comp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I38 (comp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I39 (comp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I40 (comp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I41 (comp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I42 (comp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I43 (comp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I44 (comp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I45 (comp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I46 (comp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I47 (comp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I48 (comp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I49 (comp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I50 (comp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I51 (comp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I52 (comp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I53 (comp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  OR2 I54 (comp_0[33:33], i_0r0[33:33], i_0r1[33:33]);
  OR2 I55 (comp_0[34:34], i_0r0[34:34], i_0r1[34:34]);
  C3 I56 (simp801_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I57 (simp801_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C3 I58 (simp801_0[2:2], comp_0[6:6], comp_0[7:7], comp_0[8:8]);
  C3 I59 (simp801_0[3:3], comp_0[9:9], comp_0[10:10], comp_0[11:11]);
  C3 I60 (simp801_0[4:4], comp_0[12:12], comp_0[13:13], comp_0[14:14]);
  C3 I61 (simp801_0[5:5], comp_0[15:15], comp_0[16:16], comp_0[17:17]);
  C3 I62 (simp801_0[6:6], comp_0[18:18], comp_0[19:19], comp_0[20:20]);
  C3 I63 (simp801_0[7:7], comp_0[21:21], comp_0[22:22], comp_0[23:23]);
  C3 I64 (simp801_0[8:8], comp_0[24:24], comp_0[25:25], comp_0[26:26]);
  C3 I65 (simp801_0[9:9], comp_0[27:27], comp_0[28:28], comp_0[29:29]);
  C3 I66 (simp801_0[10:10], comp_0[30:30], comp_0[31:31], comp_0[32:32]);
  C2 I67 (simp801_0[11:11], comp_0[33:33], comp_0[34:34]);
  C3 I68 (simp802_0[0:0], simp801_0[0:0], simp801_0[1:1], simp801_0[2:2]);
  C3 I69 (simp802_0[1:1], simp801_0[3:3], simp801_0[4:4], simp801_0[5:5]);
  C3 I70 (simp802_0[2:2], simp801_0[6:6], simp801_0[7:7], simp801_0[8:8]);
  C3 I71 (simp802_0[3:3], simp801_0[9:9], simp801_0[10:10], simp801_0[11:11]);
  C3 I72 (simp803_0[0:0], simp802_0[0:0], simp802_0[1:1], simp802_0[2:2]);
  BUFF I73 (simp803_0[1:1], simp802_0[3:3]);
  C2 I74 (icomplete_0, simp803_0[0:0], simp803_0[1:1]);
  C2 I75 (o_0r0[0:0], i_0r0[0:0], gsel_0);
  C2 I76 (o_0r0[1:1], i_0r0[1:1], gsel_0);
  C2 I77 (o_0r0[2:2], i_0r0[2:2], gsel_0);
  C2 I78 (o_0r0[3:3], i_0r0[3:3], gsel_0);
  C2 I79 (o_0r0[4:4], i_0r0[4:4], gsel_0);
  C2 I80 (o_0r0[5:5], i_0r0[5:5], gsel_0);
  C2 I81 (o_0r0[6:6], i_0r0[6:6], gsel_0);
  C2 I82 (o_0r0[7:7], i_0r0[7:7], gsel_0);
  C2 I83 (o_0r0[8:8], i_0r0[8:8], gsel_0);
  C2 I84 (o_0r0[9:9], i_0r0[9:9], gsel_0);
  C2 I85 (o_0r0[10:10], i_0r0[10:10], gsel_0);
  C2 I86 (o_0r0[11:11], i_0r0[11:11], gsel_0);
  C2 I87 (o_0r0[12:12], i_0r0[12:12], gsel_0);
  C2 I88 (o_0r0[13:13], i_0r0[13:13], gsel_0);
  C2 I89 (o_0r0[14:14], i_0r0[14:14], gsel_0);
  C2 I90 (o_0r0[15:15], i_0r0[15:15], gsel_0);
  C2 I91 (o_0r0[16:16], i_0r0[16:16], gsel_0);
  C2 I92 (o_0r0[17:17], i_0r0[17:17], gsel_0);
  C2 I93 (o_0r0[18:18], i_0r0[18:18], gsel_0);
  C2 I94 (o_0r0[19:19], i_0r0[19:19], gsel_0);
  C2 I95 (o_0r0[20:20], i_0r0[20:20], gsel_0);
  C2 I96 (o_0r0[21:21], i_0r0[21:21], gsel_0);
  C2 I97 (o_0r0[22:22], i_0r0[22:22], gsel_0);
  C2 I98 (o_0r0[23:23], i_0r0[23:23], gsel_0);
  C2 I99 (o_0r0[24:24], i_0r0[24:24], gsel_0);
  C2 I100 (o_0r0[25:25], i_0r0[25:25], gsel_0);
  C2 I101 (o_0r0[26:26], i_0r0[26:26], gsel_0);
  C2 I102 (o_0r0[27:27], i_0r0[27:27], gsel_0);
  C2 I103 (o_0r0[28:28], i_0r0[28:28], gsel_0);
  C2 I104 (o_0r0[29:29], i_0r0[29:29], gsel_0);
  C2 I105 (o_0r0[30:30], i_0r0[30:30], gsel_0);
  C2 I106 (o_0r0[31:31], i_0r0[31:31], gsel_0);
  C2 I107 (o_1r0[0:0], i_0r0[0:0], gsel_1);
  C2 I108 (o_1r0[1:1], i_0r0[1:1], gsel_1);
  C2 I109 (o_1r0[2:2], i_0r0[2:2], gsel_1);
  C2 I110 (o_1r0[3:3], i_0r0[3:3], gsel_1);
  C2 I111 (o_1r0[4:4], i_0r0[4:4], gsel_1);
  C2 I112 (o_1r0[5:5], i_0r0[5:5], gsel_1);
  C2 I113 (o_1r0[6:6], i_0r0[6:6], gsel_1);
  C2 I114 (o_1r0[7:7], i_0r0[7:7], gsel_1);
  C2 I115 (o_1r0[8:8], i_0r0[8:8], gsel_1);
  C2 I116 (o_1r0[9:9], i_0r0[9:9], gsel_1);
  C2 I117 (o_1r0[10:10], i_0r0[10:10], gsel_1);
  C2 I118 (o_1r0[11:11], i_0r0[11:11], gsel_1);
  C2 I119 (o_1r0[12:12], i_0r0[12:12], gsel_1);
  C2 I120 (o_1r0[13:13], i_0r0[13:13], gsel_1);
  C2 I121 (o_1r0[14:14], i_0r0[14:14], gsel_1);
  C2 I122 (o_1r0[15:15], i_0r0[15:15], gsel_1);
  C2 I123 (o_1r0[16:16], i_0r0[16:16], gsel_1);
  C2 I124 (o_1r0[17:17], i_0r0[17:17], gsel_1);
  C2 I125 (o_1r0[18:18], i_0r0[18:18], gsel_1);
  C2 I126 (o_1r0[19:19], i_0r0[19:19], gsel_1);
  C2 I127 (o_1r0[20:20], i_0r0[20:20], gsel_1);
  C2 I128 (o_1r0[21:21], i_0r0[21:21], gsel_1);
  C2 I129 (o_1r0[22:22], i_0r0[22:22], gsel_1);
  C2 I130 (o_1r0[23:23], i_0r0[23:23], gsel_1);
  C2 I131 (o_1r0[24:24], i_0r0[24:24], gsel_1);
  C2 I132 (o_1r0[25:25], i_0r0[25:25], gsel_1);
  C2 I133 (o_1r0[26:26], i_0r0[26:26], gsel_1);
  C2 I134 (o_1r0[27:27], i_0r0[27:27], gsel_1);
  C2 I135 (o_1r0[28:28], i_0r0[28:28], gsel_1);
  C2 I136 (o_1r0[29:29], i_0r0[29:29], gsel_1);
  C2 I137 (o_1r0[30:30], i_0r0[30:30], gsel_1);
  C2 I138 (o_1r0[31:31], i_0r0[31:31], gsel_1);
  C2 I139 (o_2r0[0:0], i_0r0[0:0], gsel_2);
  C2 I140 (o_2r0[1:1], i_0r0[1:1], gsel_2);
  C2 I141 (o_2r0[2:2], i_0r0[2:2], gsel_2);
  C2 I142 (o_2r0[3:3], i_0r0[3:3], gsel_2);
  C2 I143 (o_2r0[4:4], i_0r0[4:4], gsel_2);
  C2 I144 (o_2r0[5:5], i_0r0[5:5], gsel_2);
  C2 I145 (o_2r0[6:6], i_0r0[6:6], gsel_2);
  C2 I146 (o_2r0[7:7], i_0r0[7:7], gsel_2);
  C2 I147 (o_2r0[8:8], i_0r0[8:8], gsel_2);
  C2 I148 (o_2r0[9:9], i_0r0[9:9], gsel_2);
  C2 I149 (o_2r0[10:10], i_0r0[10:10], gsel_2);
  C2 I150 (o_2r0[11:11], i_0r0[11:11], gsel_2);
  C2 I151 (o_2r0[12:12], i_0r0[12:12], gsel_2);
  C2 I152 (o_2r0[13:13], i_0r0[13:13], gsel_2);
  C2 I153 (o_2r0[14:14], i_0r0[14:14], gsel_2);
  C2 I154 (o_2r0[15:15], i_0r0[15:15], gsel_2);
  C2 I155 (o_2r0[16:16], i_0r0[16:16], gsel_2);
  C2 I156 (o_2r0[17:17], i_0r0[17:17], gsel_2);
  C2 I157 (o_2r0[18:18], i_0r0[18:18], gsel_2);
  C2 I158 (o_2r0[19:19], i_0r0[19:19], gsel_2);
  C2 I159 (o_2r0[20:20], i_0r0[20:20], gsel_2);
  C2 I160 (o_2r0[21:21], i_0r0[21:21], gsel_2);
  C2 I161 (o_2r0[22:22], i_0r0[22:22], gsel_2);
  C2 I162 (o_2r0[23:23], i_0r0[23:23], gsel_2);
  C2 I163 (o_2r0[24:24], i_0r0[24:24], gsel_2);
  C2 I164 (o_2r0[25:25], i_0r0[25:25], gsel_2);
  C2 I165 (o_2r0[26:26], i_0r0[26:26], gsel_2);
  C2 I166 (o_2r0[27:27], i_0r0[27:27], gsel_2);
  C2 I167 (o_2r0[28:28], i_0r0[28:28], gsel_2);
  C2 I168 (o_2r0[29:29], i_0r0[29:29], gsel_2);
  C2 I169 (o_2r0[30:30], i_0r0[30:30], gsel_2);
  C2 I170 (o_2r0[31:31], i_0r0[31:31], gsel_2);
  C2 I171 (o_3r0[0:0], i_0r0[0:0], gsel_3);
  C2 I172 (o_3r0[1:1], i_0r0[1:1], gsel_3);
  C2 I173 (o_3r0[2:2], i_0r0[2:2], gsel_3);
  C2 I174 (o_3r0[3:3], i_0r0[3:3], gsel_3);
  C2 I175 (o_3r0[4:4], i_0r0[4:4], gsel_3);
  C2 I176 (o_3r0[5:5], i_0r0[5:5], gsel_3);
  C2 I177 (o_3r0[6:6], i_0r0[6:6], gsel_3);
  C2 I178 (o_3r0[7:7], i_0r0[7:7], gsel_3);
  C2 I179 (o_3r0[8:8], i_0r0[8:8], gsel_3);
  C2 I180 (o_3r0[9:9], i_0r0[9:9], gsel_3);
  C2 I181 (o_3r0[10:10], i_0r0[10:10], gsel_3);
  C2 I182 (o_3r0[11:11], i_0r0[11:11], gsel_3);
  C2 I183 (o_3r0[12:12], i_0r0[12:12], gsel_3);
  C2 I184 (o_3r0[13:13], i_0r0[13:13], gsel_3);
  C2 I185 (o_3r0[14:14], i_0r0[14:14], gsel_3);
  C2 I186 (o_3r0[15:15], i_0r0[15:15], gsel_3);
  C2 I187 (o_3r0[16:16], i_0r0[16:16], gsel_3);
  C2 I188 (o_3r0[17:17], i_0r0[17:17], gsel_3);
  C2 I189 (o_3r0[18:18], i_0r0[18:18], gsel_3);
  C2 I190 (o_3r0[19:19], i_0r0[19:19], gsel_3);
  C2 I191 (o_3r0[20:20], i_0r0[20:20], gsel_3);
  C2 I192 (o_3r0[21:21], i_0r0[21:21], gsel_3);
  C2 I193 (o_3r0[22:22], i_0r0[22:22], gsel_3);
  C2 I194 (o_3r0[23:23], i_0r0[23:23], gsel_3);
  C2 I195 (o_3r0[24:24], i_0r0[24:24], gsel_3);
  C2 I196 (o_3r0[25:25], i_0r0[25:25], gsel_3);
  C2 I197 (o_3r0[26:26], i_0r0[26:26], gsel_3);
  C2 I198 (o_3r0[27:27], i_0r0[27:27], gsel_3);
  C2 I199 (o_3r0[28:28], i_0r0[28:28], gsel_3);
  C2 I200 (o_3r0[29:29], i_0r0[29:29], gsel_3);
  C2 I201 (o_3r0[30:30], i_0r0[30:30], gsel_3);
  C2 I202 (o_3r0[31:31], i_0r0[31:31], gsel_3);
  C2 I203 (o_4r0[0:0], i_0r0[0:0], gsel_4);
  C2 I204 (o_4r0[1:1], i_0r0[1:1], gsel_4);
  C2 I205 (o_4r0[2:2], i_0r0[2:2], gsel_4);
  C2 I206 (o_4r0[3:3], i_0r0[3:3], gsel_4);
  C2 I207 (o_4r0[4:4], i_0r0[4:4], gsel_4);
  C2 I208 (o_4r0[5:5], i_0r0[5:5], gsel_4);
  C2 I209 (o_4r0[6:6], i_0r0[6:6], gsel_4);
  C2 I210 (o_4r0[7:7], i_0r0[7:7], gsel_4);
  C2 I211 (o_4r0[8:8], i_0r0[8:8], gsel_4);
  C2 I212 (o_4r0[9:9], i_0r0[9:9], gsel_4);
  C2 I213 (o_4r0[10:10], i_0r0[10:10], gsel_4);
  C2 I214 (o_4r0[11:11], i_0r0[11:11], gsel_4);
  C2 I215 (o_4r0[12:12], i_0r0[12:12], gsel_4);
  C2 I216 (o_4r0[13:13], i_0r0[13:13], gsel_4);
  C2 I217 (o_4r0[14:14], i_0r0[14:14], gsel_4);
  C2 I218 (o_4r0[15:15], i_0r0[15:15], gsel_4);
  C2 I219 (o_4r0[16:16], i_0r0[16:16], gsel_4);
  C2 I220 (o_4r0[17:17], i_0r0[17:17], gsel_4);
  C2 I221 (o_4r0[18:18], i_0r0[18:18], gsel_4);
  C2 I222 (o_4r0[19:19], i_0r0[19:19], gsel_4);
  C2 I223 (o_4r0[20:20], i_0r0[20:20], gsel_4);
  C2 I224 (o_4r0[21:21], i_0r0[21:21], gsel_4);
  C2 I225 (o_4r0[22:22], i_0r0[22:22], gsel_4);
  C2 I226 (o_4r0[23:23], i_0r0[23:23], gsel_4);
  C2 I227 (o_4r0[24:24], i_0r0[24:24], gsel_4);
  C2 I228 (o_4r0[25:25], i_0r0[25:25], gsel_4);
  C2 I229 (o_4r0[26:26], i_0r0[26:26], gsel_4);
  C2 I230 (o_4r0[27:27], i_0r0[27:27], gsel_4);
  C2 I231 (o_4r0[28:28], i_0r0[28:28], gsel_4);
  C2 I232 (o_4r0[29:29], i_0r0[29:29], gsel_4);
  C2 I233 (o_4r0[30:30], i_0r0[30:30], gsel_4);
  C2 I234 (o_4r0[31:31], i_0r0[31:31], gsel_4);
  C2 I235 (o_5r0[0:0], i_0r0[0:0], gsel_5);
  C2 I236 (o_5r0[1:1], i_0r0[1:1], gsel_5);
  C2 I237 (o_5r0[2:2], i_0r0[2:2], gsel_5);
  C2 I238 (o_5r0[3:3], i_0r0[3:3], gsel_5);
  C2 I239 (o_5r0[4:4], i_0r0[4:4], gsel_5);
  C2 I240 (o_5r0[5:5], i_0r0[5:5], gsel_5);
  C2 I241 (o_5r0[6:6], i_0r0[6:6], gsel_5);
  C2 I242 (o_5r0[7:7], i_0r0[7:7], gsel_5);
  C2 I243 (o_5r0[8:8], i_0r0[8:8], gsel_5);
  C2 I244 (o_5r0[9:9], i_0r0[9:9], gsel_5);
  C2 I245 (o_5r0[10:10], i_0r0[10:10], gsel_5);
  C2 I246 (o_5r0[11:11], i_0r0[11:11], gsel_5);
  C2 I247 (o_5r0[12:12], i_0r0[12:12], gsel_5);
  C2 I248 (o_5r0[13:13], i_0r0[13:13], gsel_5);
  C2 I249 (o_5r0[14:14], i_0r0[14:14], gsel_5);
  C2 I250 (o_5r0[15:15], i_0r0[15:15], gsel_5);
  C2 I251 (o_5r0[16:16], i_0r0[16:16], gsel_5);
  C2 I252 (o_5r0[17:17], i_0r0[17:17], gsel_5);
  C2 I253 (o_5r0[18:18], i_0r0[18:18], gsel_5);
  C2 I254 (o_5r0[19:19], i_0r0[19:19], gsel_5);
  C2 I255 (o_5r0[20:20], i_0r0[20:20], gsel_5);
  C2 I256 (o_5r0[21:21], i_0r0[21:21], gsel_5);
  C2 I257 (o_5r0[22:22], i_0r0[22:22], gsel_5);
  C2 I258 (o_5r0[23:23], i_0r0[23:23], gsel_5);
  C2 I259 (o_5r0[24:24], i_0r0[24:24], gsel_5);
  C2 I260 (o_5r0[25:25], i_0r0[25:25], gsel_5);
  C2 I261 (o_5r0[26:26], i_0r0[26:26], gsel_5);
  C2 I262 (o_5r0[27:27], i_0r0[27:27], gsel_5);
  C2 I263 (o_5r0[28:28], i_0r0[28:28], gsel_5);
  C2 I264 (o_5r0[29:29], i_0r0[29:29], gsel_5);
  C2 I265 (o_5r0[30:30], i_0r0[30:30], gsel_5);
  C2 I266 (o_5r0[31:31], i_0r0[31:31], gsel_5);
  C2 I267 (o_6r0[0:0], i_0r0[0:0], gsel_6);
  C2 I268 (o_6r0[1:1], i_0r0[1:1], gsel_6);
  C2 I269 (o_6r0[2:2], i_0r0[2:2], gsel_6);
  C2 I270 (o_6r0[3:3], i_0r0[3:3], gsel_6);
  C2 I271 (o_6r0[4:4], i_0r0[4:4], gsel_6);
  C2 I272 (o_6r0[5:5], i_0r0[5:5], gsel_6);
  C2 I273 (o_6r0[6:6], i_0r0[6:6], gsel_6);
  C2 I274 (o_6r0[7:7], i_0r0[7:7], gsel_6);
  C2 I275 (o_6r0[8:8], i_0r0[8:8], gsel_6);
  C2 I276 (o_6r0[9:9], i_0r0[9:9], gsel_6);
  C2 I277 (o_6r0[10:10], i_0r0[10:10], gsel_6);
  C2 I278 (o_6r0[11:11], i_0r0[11:11], gsel_6);
  C2 I279 (o_6r0[12:12], i_0r0[12:12], gsel_6);
  C2 I280 (o_6r0[13:13], i_0r0[13:13], gsel_6);
  C2 I281 (o_6r0[14:14], i_0r0[14:14], gsel_6);
  C2 I282 (o_6r0[15:15], i_0r0[15:15], gsel_6);
  C2 I283 (o_6r0[16:16], i_0r0[16:16], gsel_6);
  C2 I284 (o_6r0[17:17], i_0r0[17:17], gsel_6);
  C2 I285 (o_6r0[18:18], i_0r0[18:18], gsel_6);
  C2 I286 (o_6r0[19:19], i_0r0[19:19], gsel_6);
  C2 I287 (o_6r0[20:20], i_0r0[20:20], gsel_6);
  C2 I288 (o_6r0[21:21], i_0r0[21:21], gsel_6);
  C2 I289 (o_6r0[22:22], i_0r0[22:22], gsel_6);
  C2 I290 (o_6r0[23:23], i_0r0[23:23], gsel_6);
  C2 I291 (o_6r0[24:24], i_0r0[24:24], gsel_6);
  C2 I292 (o_6r0[25:25], i_0r0[25:25], gsel_6);
  C2 I293 (o_6r0[26:26], i_0r0[26:26], gsel_6);
  C2 I294 (o_6r0[27:27], i_0r0[27:27], gsel_6);
  C2 I295 (o_6r0[28:28], i_0r0[28:28], gsel_6);
  C2 I296 (o_6r0[29:29], i_0r0[29:29], gsel_6);
  C2 I297 (o_6r0[30:30], i_0r0[30:30], gsel_6);
  C2 I298 (o_6r0[31:31], i_0r0[31:31], gsel_6);
  C2 I299 (o_0r1[0:0], i_0r1[0:0], gsel_0);
  C2 I300 (o_0r1[1:1], i_0r1[1:1], gsel_0);
  C2 I301 (o_0r1[2:2], i_0r1[2:2], gsel_0);
  C2 I302 (o_0r1[3:3], i_0r1[3:3], gsel_0);
  C2 I303 (o_0r1[4:4], i_0r1[4:4], gsel_0);
  C2 I304 (o_0r1[5:5], i_0r1[5:5], gsel_0);
  C2 I305 (o_0r1[6:6], i_0r1[6:6], gsel_0);
  C2 I306 (o_0r1[7:7], i_0r1[7:7], gsel_0);
  C2 I307 (o_0r1[8:8], i_0r1[8:8], gsel_0);
  C2 I308 (o_0r1[9:9], i_0r1[9:9], gsel_0);
  C2 I309 (o_0r1[10:10], i_0r1[10:10], gsel_0);
  C2 I310 (o_0r1[11:11], i_0r1[11:11], gsel_0);
  C2 I311 (o_0r1[12:12], i_0r1[12:12], gsel_0);
  C2 I312 (o_0r1[13:13], i_0r1[13:13], gsel_0);
  C2 I313 (o_0r1[14:14], i_0r1[14:14], gsel_0);
  C2 I314 (o_0r1[15:15], i_0r1[15:15], gsel_0);
  C2 I315 (o_0r1[16:16], i_0r1[16:16], gsel_0);
  C2 I316 (o_0r1[17:17], i_0r1[17:17], gsel_0);
  C2 I317 (o_0r1[18:18], i_0r1[18:18], gsel_0);
  C2 I318 (o_0r1[19:19], i_0r1[19:19], gsel_0);
  C2 I319 (o_0r1[20:20], i_0r1[20:20], gsel_0);
  C2 I320 (o_0r1[21:21], i_0r1[21:21], gsel_0);
  C2 I321 (o_0r1[22:22], i_0r1[22:22], gsel_0);
  C2 I322 (o_0r1[23:23], i_0r1[23:23], gsel_0);
  C2 I323 (o_0r1[24:24], i_0r1[24:24], gsel_0);
  C2 I324 (o_0r1[25:25], i_0r1[25:25], gsel_0);
  C2 I325 (o_0r1[26:26], i_0r1[26:26], gsel_0);
  C2 I326 (o_0r1[27:27], i_0r1[27:27], gsel_0);
  C2 I327 (o_0r1[28:28], i_0r1[28:28], gsel_0);
  C2 I328 (o_0r1[29:29], i_0r1[29:29], gsel_0);
  C2 I329 (o_0r1[30:30], i_0r1[30:30], gsel_0);
  C2 I330 (o_0r1[31:31], i_0r1[31:31], gsel_0);
  C2 I331 (o_1r1[0:0], i_0r1[0:0], gsel_1);
  C2 I332 (o_1r1[1:1], i_0r1[1:1], gsel_1);
  C2 I333 (o_1r1[2:2], i_0r1[2:2], gsel_1);
  C2 I334 (o_1r1[3:3], i_0r1[3:3], gsel_1);
  C2 I335 (o_1r1[4:4], i_0r1[4:4], gsel_1);
  C2 I336 (o_1r1[5:5], i_0r1[5:5], gsel_1);
  C2 I337 (o_1r1[6:6], i_0r1[6:6], gsel_1);
  C2 I338 (o_1r1[7:7], i_0r1[7:7], gsel_1);
  C2 I339 (o_1r1[8:8], i_0r1[8:8], gsel_1);
  C2 I340 (o_1r1[9:9], i_0r1[9:9], gsel_1);
  C2 I341 (o_1r1[10:10], i_0r1[10:10], gsel_1);
  C2 I342 (o_1r1[11:11], i_0r1[11:11], gsel_1);
  C2 I343 (o_1r1[12:12], i_0r1[12:12], gsel_1);
  C2 I344 (o_1r1[13:13], i_0r1[13:13], gsel_1);
  C2 I345 (o_1r1[14:14], i_0r1[14:14], gsel_1);
  C2 I346 (o_1r1[15:15], i_0r1[15:15], gsel_1);
  C2 I347 (o_1r1[16:16], i_0r1[16:16], gsel_1);
  C2 I348 (o_1r1[17:17], i_0r1[17:17], gsel_1);
  C2 I349 (o_1r1[18:18], i_0r1[18:18], gsel_1);
  C2 I350 (o_1r1[19:19], i_0r1[19:19], gsel_1);
  C2 I351 (o_1r1[20:20], i_0r1[20:20], gsel_1);
  C2 I352 (o_1r1[21:21], i_0r1[21:21], gsel_1);
  C2 I353 (o_1r1[22:22], i_0r1[22:22], gsel_1);
  C2 I354 (o_1r1[23:23], i_0r1[23:23], gsel_1);
  C2 I355 (o_1r1[24:24], i_0r1[24:24], gsel_1);
  C2 I356 (o_1r1[25:25], i_0r1[25:25], gsel_1);
  C2 I357 (o_1r1[26:26], i_0r1[26:26], gsel_1);
  C2 I358 (o_1r1[27:27], i_0r1[27:27], gsel_1);
  C2 I359 (o_1r1[28:28], i_0r1[28:28], gsel_1);
  C2 I360 (o_1r1[29:29], i_0r1[29:29], gsel_1);
  C2 I361 (o_1r1[30:30], i_0r1[30:30], gsel_1);
  C2 I362 (o_1r1[31:31], i_0r1[31:31], gsel_1);
  C2 I363 (o_2r1[0:0], i_0r1[0:0], gsel_2);
  C2 I364 (o_2r1[1:1], i_0r1[1:1], gsel_2);
  C2 I365 (o_2r1[2:2], i_0r1[2:2], gsel_2);
  C2 I366 (o_2r1[3:3], i_0r1[3:3], gsel_2);
  C2 I367 (o_2r1[4:4], i_0r1[4:4], gsel_2);
  C2 I368 (o_2r1[5:5], i_0r1[5:5], gsel_2);
  C2 I369 (o_2r1[6:6], i_0r1[6:6], gsel_2);
  C2 I370 (o_2r1[7:7], i_0r1[7:7], gsel_2);
  C2 I371 (o_2r1[8:8], i_0r1[8:8], gsel_2);
  C2 I372 (o_2r1[9:9], i_0r1[9:9], gsel_2);
  C2 I373 (o_2r1[10:10], i_0r1[10:10], gsel_2);
  C2 I374 (o_2r1[11:11], i_0r1[11:11], gsel_2);
  C2 I375 (o_2r1[12:12], i_0r1[12:12], gsel_2);
  C2 I376 (o_2r1[13:13], i_0r1[13:13], gsel_2);
  C2 I377 (o_2r1[14:14], i_0r1[14:14], gsel_2);
  C2 I378 (o_2r1[15:15], i_0r1[15:15], gsel_2);
  C2 I379 (o_2r1[16:16], i_0r1[16:16], gsel_2);
  C2 I380 (o_2r1[17:17], i_0r1[17:17], gsel_2);
  C2 I381 (o_2r1[18:18], i_0r1[18:18], gsel_2);
  C2 I382 (o_2r1[19:19], i_0r1[19:19], gsel_2);
  C2 I383 (o_2r1[20:20], i_0r1[20:20], gsel_2);
  C2 I384 (o_2r1[21:21], i_0r1[21:21], gsel_2);
  C2 I385 (o_2r1[22:22], i_0r1[22:22], gsel_2);
  C2 I386 (o_2r1[23:23], i_0r1[23:23], gsel_2);
  C2 I387 (o_2r1[24:24], i_0r1[24:24], gsel_2);
  C2 I388 (o_2r1[25:25], i_0r1[25:25], gsel_2);
  C2 I389 (o_2r1[26:26], i_0r1[26:26], gsel_2);
  C2 I390 (o_2r1[27:27], i_0r1[27:27], gsel_2);
  C2 I391 (o_2r1[28:28], i_0r1[28:28], gsel_2);
  C2 I392 (o_2r1[29:29], i_0r1[29:29], gsel_2);
  C2 I393 (o_2r1[30:30], i_0r1[30:30], gsel_2);
  C2 I394 (o_2r1[31:31], i_0r1[31:31], gsel_2);
  C2 I395 (o_3r1[0:0], i_0r1[0:0], gsel_3);
  C2 I396 (o_3r1[1:1], i_0r1[1:1], gsel_3);
  C2 I397 (o_3r1[2:2], i_0r1[2:2], gsel_3);
  C2 I398 (o_3r1[3:3], i_0r1[3:3], gsel_3);
  C2 I399 (o_3r1[4:4], i_0r1[4:4], gsel_3);
  C2 I400 (o_3r1[5:5], i_0r1[5:5], gsel_3);
  C2 I401 (o_3r1[6:6], i_0r1[6:6], gsel_3);
  C2 I402 (o_3r1[7:7], i_0r1[7:7], gsel_3);
  C2 I403 (o_3r1[8:8], i_0r1[8:8], gsel_3);
  C2 I404 (o_3r1[9:9], i_0r1[9:9], gsel_3);
  C2 I405 (o_3r1[10:10], i_0r1[10:10], gsel_3);
  C2 I406 (o_3r1[11:11], i_0r1[11:11], gsel_3);
  C2 I407 (o_3r1[12:12], i_0r1[12:12], gsel_3);
  C2 I408 (o_3r1[13:13], i_0r1[13:13], gsel_3);
  C2 I409 (o_3r1[14:14], i_0r1[14:14], gsel_3);
  C2 I410 (o_3r1[15:15], i_0r1[15:15], gsel_3);
  C2 I411 (o_3r1[16:16], i_0r1[16:16], gsel_3);
  C2 I412 (o_3r1[17:17], i_0r1[17:17], gsel_3);
  C2 I413 (o_3r1[18:18], i_0r1[18:18], gsel_3);
  C2 I414 (o_3r1[19:19], i_0r1[19:19], gsel_3);
  C2 I415 (o_3r1[20:20], i_0r1[20:20], gsel_3);
  C2 I416 (o_3r1[21:21], i_0r1[21:21], gsel_3);
  C2 I417 (o_3r1[22:22], i_0r1[22:22], gsel_3);
  C2 I418 (o_3r1[23:23], i_0r1[23:23], gsel_3);
  C2 I419 (o_3r1[24:24], i_0r1[24:24], gsel_3);
  C2 I420 (o_3r1[25:25], i_0r1[25:25], gsel_3);
  C2 I421 (o_3r1[26:26], i_0r1[26:26], gsel_3);
  C2 I422 (o_3r1[27:27], i_0r1[27:27], gsel_3);
  C2 I423 (o_3r1[28:28], i_0r1[28:28], gsel_3);
  C2 I424 (o_3r1[29:29], i_0r1[29:29], gsel_3);
  C2 I425 (o_3r1[30:30], i_0r1[30:30], gsel_3);
  C2 I426 (o_3r1[31:31], i_0r1[31:31], gsel_3);
  C2 I427 (o_4r1[0:0], i_0r1[0:0], gsel_4);
  C2 I428 (o_4r1[1:1], i_0r1[1:1], gsel_4);
  C2 I429 (o_4r1[2:2], i_0r1[2:2], gsel_4);
  C2 I430 (o_4r1[3:3], i_0r1[3:3], gsel_4);
  C2 I431 (o_4r1[4:4], i_0r1[4:4], gsel_4);
  C2 I432 (o_4r1[5:5], i_0r1[5:5], gsel_4);
  C2 I433 (o_4r1[6:6], i_0r1[6:6], gsel_4);
  C2 I434 (o_4r1[7:7], i_0r1[7:7], gsel_4);
  C2 I435 (o_4r1[8:8], i_0r1[8:8], gsel_4);
  C2 I436 (o_4r1[9:9], i_0r1[9:9], gsel_4);
  C2 I437 (o_4r1[10:10], i_0r1[10:10], gsel_4);
  C2 I438 (o_4r1[11:11], i_0r1[11:11], gsel_4);
  C2 I439 (o_4r1[12:12], i_0r1[12:12], gsel_4);
  C2 I440 (o_4r1[13:13], i_0r1[13:13], gsel_4);
  C2 I441 (o_4r1[14:14], i_0r1[14:14], gsel_4);
  C2 I442 (o_4r1[15:15], i_0r1[15:15], gsel_4);
  C2 I443 (o_4r1[16:16], i_0r1[16:16], gsel_4);
  C2 I444 (o_4r1[17:17], i_0r1[17:17], gsel_4);
  C2 I445 (o_4r1[18:18], i_0r1[18:18], gsel_4);
  C2 I446 (o_4r1[19:19], i_0r1[19:19], gsel_4);
  C2 I447 (o_4r1[20:20], i_0r1[20:20], gsel_4);
  C2 I448 (o_4r1[21:21], i_0r1[21:21], gsel_4);
  C2 I449 (o_4r1[22:22], i_0r1[22:22], gsel_4);
  C2 I450 (o_4r1[23:23], i_0r1[23:23], gsel_4);
  C2 I451 (o_4r1[24:24], i_0r1[24:24], gsel_4);
  C2 I452 (o_4r1[25:25], i_0r1[25:25], gsel_4);
  C2 I453 (o_4r1[26:26], i_0r1[26:26], gsel_4);
  C2 I454 (o_4r1[27:27], i_0r1[27:27], gsel_4);
  C2 I455 (o_4r1[28:28], i_0r1[28:28], gsel_4);
  C2 I456 (o_4r1[29:29], i_0r1[29:29], gsel_4);
  C2 I457 (o_4r1[30:30], i_0r1[30:30], gsel_4);
  C2 I458 (o_4r1[31:31], i_0r1[31:31], gsel_4);
  C2 I459 (o_5r1[0:0], i_0r1[0:0], gsel_5);
  C2 I460 (o_5r1[1:1], i_0r1[1:1], gsel_5);
  C2 I461 (o_5r1[2:2], i_0r1[2:2], gsel_5);
  C2 I462 (o_5r1[3:3], i_0r1[3:3], gsel_5);
  C2 I463 (o_5r1[4:4], i_0r1[4:4], gsel_5);
  C2 I464 (o_5r1[5:5], i_0r1[5:5], gsel_5);
  C2 I465 (o_5r1[6:6], i_0r1[6:6], gsel_5);
  C2 I466 (o_5r1[7:7], i_0r1[7:7], gsel_5);
  C2 I467 (o_5r1[8:8], i_0r1[8:8], gsel_5);
  C2 I468 (o_5r1[9:9], i_0r1[9:9], gsel_5);
  C2 I469 (o_5r1[10:10], i_0r1[10:10], gsel_5);
  C2 I470 (o_5r1[11:11], i_0r1[11:11], gsel_5);
  C2 I471 (o_5r1[12:12], i_0r1[12:12], gsel_5);
  C2 I472 (o_5r1[13:13], i_0r1[13:13], gsel_5);
  C2 I473 (o_5r1[14:14], i_0r1[14:14], gsel_5);
  C2 I474 (o_5r1[15:15], i_0r1[15:15], gsel_5);
  C2 I475 (o_5r1[16:16], i_0r1[16:16], gsel_5);
  C2 I476 (o_5r1[17:17], i_0r1[17:17], gsel_5);
  C2 I477 (o_5r1[18:18], i_0r1[18:18], gsel_5);
  C2 I478 (o_5r1[19:19], i_0r1[19:19], gsel_5);
  C2 I479 (o_5r1[20:20], i_0r1[20:20], gsel_5);
  C2 I480 (o_5r1[21:21], i_0r1[21:21], gsel_5);
  C2 I481 (o_5r1[22:22], i_0r1[22:22], gsel_5);
  C2 I482 (o_5r1[23:23], i_0r1[23:23], gsel_5);
  C2 I483 (o_5r1[24:24], i_0r1[24:24], gsel_5);
  C2 I484 (o_5r1[25:25], i_0r1[25:25], gsel_5);
  C2 I485 (o_5r1[26:26], i_0r1[26:26], gsel_5);
  C2 I486 (o_5r1[27:27], i_0r1[27:27], gsel_5);
  C2 I487 (o_5r1[28:28], i_0r1[28:28], gsel_5);
  C2 I488 (o_5r1[29:29], i_0r1[29:29], gsel_5);
  C2 I489 (o_5r1[30:30], i_0r1[30:30], gsel_5);
  C2 I490 (o_5r1[31:31], i_0r1[31:31], gsel_5);
  C2 I491 (o_6r1[0:0], i_0r1[0:0], gsel_6);
  C2 I492 (o_6r1[1:1], i_0r1[1:1], gsel_6);
  C2 I493 (o_6r1[2:2], i_0r1[2:2], gsel_6);
  C2 I494 (o_6r1[3:3], i_0r1[3:3], gsel_6);
  C2 I495 (o_6r1[4:4], i_0r1[4:4], gsel_6);
  C2 I496 (o_6r1[5:5], i_0r1[5:5], gsel_6);
  C2 I497 (o_6r1[6:6], i_0r1[6:6], gsel_6);
  C2 I498 (o_6r1[7:7], i_0r1[7:7], gsel_6);
  C2 I499 (o_6r1[8:8], i_0r1[8:8], gsel_6);
  C2 I500 (o_6r1[9:9], i_0r1[9:9], gsel_6);
  C2 I501 (o_6r1[10:10], i_0r1[10:10], gsel_6);
  C2 I502 (o_6r1[11:11], i_0r1[11:11], gsel_6);
  C2 I503 (o_6r1[12:12], i_0r1[12:12], gsel_6);
  C2 I504 (o_6r1[13:13], i_0r1[13:13], gsel_6);
  C2 I505 (o_6r1[14:14], i_0r1[14:14], gsel_6);
  C2 I506 (o_6r1[15:15], i_0r1[15:15], gsel_6);
  C2 I507 (o_6r1[16:16], i_0r1[16:16], gsel_6);
  C2 I508 (o_6r1[17:17], i_0r1[17:17], gsel_6);
  C2 I509 (o_6r1[18:18], i_0r1[18:18], gsel_6);
  C2 I510 (o_6r1[19:19], i_0r1[19:19], gsel_6);
  C2 I511 (o_6r1[20:20], i_0r1[20:20], gsel_6);
  C2 I512 (o_6r1[21:21], i_0r1[21:21], gsel_6);
  C2 I513 (o_6r1[22:22], i_0r1[22:22], gsel_6);
  C2 I514 (o_6r1[23:23], i_0r1[23:23], gsel_6);
  C2 I515 (o_6r1[24:24], i_0r1[24:24], gsel_6);
  C2 I516 (o_6r1[25:25], i_0r1[25:25], gsel_6);
  C2 I517 (o_6r1[26:26], i_0r1[26:26], gsel_6);
  C2 I518 (o_6r1[27:27], i_0r1[27:27], gsel_6);
  C2 I519 (o_6r1[28:28], i_0r1[28:28], gsel_6);
  C2 I520 (o_6r1[29:29], i_0r1[29:29], gsel_6);
  C2 I521 (o_6r1[30:30], i_0r1[30:30], gsel_6);
  C2 I522 (o_6r1[31:31], i_0r1[31:31], gsel_6);
  NOR3 I523 (simp5291_0[0:0], o_0a, o_1a, o_2a);
  NOR3 I524 (simp5291_0[1:1], o_3a, o_4a, o_5a);
  INV I525 (simp5291_0[2:2], o_6a);
  NAND3 I526 (oack_0, simp5291_0[0:0], simp5291_0[1:1], simp5291_0[2:2]);
  C2 I527 (i_0a, oack_0, icomplete_0);
endmodule

// tkm7x0b TeakM [Many [0,0,0,0,0,0,0],One 0]
module tkm7x0b (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, i_3r, i_3a, i_4r, i_4a, i_5r, i_5a, i_6r, i_6a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  input i_4r;
  output i_4a;
  input i_5r;
  output i_5a;
  input i_6r;
  output i_6a;
  output o_0r;
  input o_0a;
  input reset;
  wire nchosen_0;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire choice_4;
  wire choice_5;
  wire choice_6;
  wire [2:0] simp161_0;
  C2R I0 (choice_0, i_0r, nchosen_0, reset);
  C2R I1 (choice_1, i_1r, nchosen_0, reset);
  C2R I2 (choice_2, i_2r, nchosen_0, reset);
  C2R I3 (choice_3, i_3r, nchosen_0, reset);
  C2R I4 (choice_4, i_4r, nchosen_0, reset);
  C2R I5 (choice_5, i_5r, nchosen_0, reset);
  C2R I6 (choice_6, i_6r, nchosen_0, reset);
  NOR2 I7 (nchosen_0, o_0r, o_0a);
  NOR3 I8 (simp161_0[0:0], choice_0, choice_1, choice_2);
  NOR3 I9 (simp161_0[1:1], choice_3, choice_4, choice_5);
  INV I10 (simp161_0[2:2], choice_6);
  NAND3 I11 (o_0r, simp161_0[0:0], simp161_0[1:1], simp161_0[2:2]);
  C2R I12 (i_0a, choice_0, o_0a, reset);
  C2R I13 (i_1a, choice_1, o_0a, reset);
  C2R I14 (i_2a, choice_2, o_0a, reset);
  C2R I15 (i_3a, choice_3, o_0a, reset);
  C2R I16 (i_4a, choice_4, o_0a, reset);
  C2R I17 (i_5a, choice_5, o_0a, reset);
  C2R I18 (i_6a, choice_6, o_0a, reset);
endmodule

// tks35_o32w3_0o0w32_1o0w32_2o0w32_3o0w32_4o0w32_5o0w32_6o0w32_7o0w32 TeakS (32+:3) [([Imp 0 0],0),([I
//   mp 1 0],0),([Imp 2 0],0),([Imp 3 0],0),([Imp 4 0],0),([Imp 5 0],0),([Imp 6 0],0),([Imp 7 0],0)] [One
//    35,Many [32,32,32,32,32,32,32,32]]
module tks35_o32w3_0o0w32_1o0w32_2o0w32_3o0w32_4o0w32_5o0w32_6o0w32_7o0w32 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r0, o_1r1, o_1a, o_2r0, o_2r1, o_2a, o_3r0, o_3r1, o_3a, o_4r0, o_4r1, o_4a, o_5r0, o_5r1, o_5a, o_6r0, o_6r1, o_6a, o_7r0, o_7r1, o_7a, reset);
  input [34:0] i_0r0;
  input [34:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  output [31:0] o_1r0;
  output [31:0] o_1r1;
  input o_1a;
  output [31:0] o_2r0;
  output [31:0] o_2r1;
  input o_2a;
  output [31:0] o_3r0;
  output [31:0] o_3r1;
  input o_3a;
  output [31:0] o_4r0;
  output [31:0] o_4r1;
  input o_4a;
  output [31:0] o_5r0;
  output [31:0] o_5r1;
  input o_5a;
  output [31:0] o_6r0;
  output [31:0] o_6r1;
  input o_6a;
  output [31:0] o_7r0;
  output [31:0] o_7r1;
  input o_7a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire sel_4;
  wire sel_5;
  wire sel_6;
  wire sel_7;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire gsel_4;
  wire gsel_5;
  wire gsel_6;
  wire gsel_7;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire match2_0;
  wire match3_0;
  wire match4_0;
  wire match5_0;
  wire match6_0;
  wire match7_0;
  wire [34:0] comp_0;
  wire [11:0] simp861_0;
  wire [3:0] simp862_0;
  wire [1:0] simp863_0;
  wire [2:0] simp5991_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (match0_0, i_0r0[32:32], i_0r0[33:33], i_0r0[34:34]);
  BUFF I2 (sel_1, match1_0);
  C3 I3 (match1_0, i_0r1[32:32], i_0r0[33:33], i_0r0[34:34]);
  BUFF I4 (sel_2, match2_0);
  C3 I5 (match2_0, i_0r0[32:32], i_0r1[33:33], i_0r0[34:34]);
  BUFF I6 (sel_3, match3_0);
  C3 I7 (match3_0, i_0r1[32:32], i_0r1[33:33], i_0r0[34:34]);
  BUFF I8 (sel_4, match4_0);
  C3 I9 (match4_0, i_0r0[32:32], i_0r0[33:33], i_0r1[34:34]);
  BUFF I10 (sel_5, match5_0);
  C3 I11 (match5_0, i_0r1[32:32], i_0r0[33:33], i_0r1[34:34]);
  BUFF I12 (sel_6, match6_0);
  C3 I13 (match6_0, i_0r0[32:32], i_0r1[33:33], i_0r1[34:34]);
  BUFF I14 (sel_7, match7_0);
  C3 I15 (match7_0, i_0r1[32:32], i_0r1[33:33], i_0r1[34:34]);
  C2 I16 (gsel_0, sel_0, icomplete_0);
  C2 I17 (gsel_1, sel_1, icomplete_0);
  C2 I18 (gsel_2, sel_2, icomplete_0);
  C2 I19 (gsel_3, sel_3, icomplete_0);
  C2 I20 (gsel_4, sel_4, icomplete_0);
  C2 I21 (gsel_5, sel_5, icomplete_0);
  C2 I22 (gsel_6, sel_6, icomplete_0);
  C2 I23 (gsel_7, sel_7, icomplete_0);
  OR2 I24 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I25 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I26 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I27 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I28 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I29 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I30 (comp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I31 (comp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I32 (comp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I33 (comp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I34 (comp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I35 (comp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I36 (comp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I37 (comp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I38 (comp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I39 (comp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I40 (comp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I41 (comp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I42 (comp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I43 (comp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I44 (comp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I45 (comp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I46 (comp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I47 (comp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I48 (comp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I49 (comp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I50 (comp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I51 (comp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I52 (comp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I53 (comp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I54 (comp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I55 (comp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I56 (comp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  OR2 I57 (comp_0[33:33], i_0r0[33:33], i_0r1[33:33]);
  OR2 I58 (comp_0[34:34], i_0r0[34:34], i_0r1[34:34]);
  C3 I59 (simp861_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I60 (simp861_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C3 I61 (simp861_0[2:2], comp_0[6:6], comp_0[7:7], comp_0[8:8]);
  C3 I62 (simp861_0[3:3], comp_0[9:9], comp_0[10:10], comp_0[11:11]);
  C3 I63 (simp861_0[4:4], comp_0[12:12], comp_0[13:13], comp_0[14:14]);
  C3 I64 (simp861_0[5:5], comp_0[15:15], comp_0[16:16], comp_0[17:17]);
  C3 I65 (simp861_0[6:6], comp_0[18:18], comp_0[19:19], comp_0[20:20]);
  C3 I66 (simp861_0[7:7], comp_0[21:21], comp_0[22:22], comp_0[23:23]);
  C3 I67 (simp861_0[8:8], comp_0[24:24], comp_0[25:25], comp_0[26:26]);
  C3 I68 (simp861_0[9:9], comp_0[27:27], comp_0[28:28], comp_0[29:29]);
  C3 I69 (simp861_0[10:10], comp_0[30:30], comp_0[31:31], comp_0[32:32]);
  C2 I70 (simp861_0[11:11], comp_0[33:33], comp_0[34:34]);
  C3 I71 (simp862_0[0:0], simp861_0[0:0], simp861_0[1:1], simp861_0[2:2]);
  C3 I72 (simp862_0[1:1], simp861_0[3:3], simp861_0[4:4], simp861_0[5:5]);
  C3 I73 (simp862_0[2:2], simp861_0[6:6], simp861_0[7:7], simp861_0[8:8]);
  C3 I74 (simp862_0[3:3], simp861_0[9:9], simp861_0[10:10], simp861_0[11:11]);
  C3 I75 (simp863_0[0:0], simp862_0[0:0], simp862_0[1:1], simp862_0[2:2]);
  BUFF I76 (simp863_0[1:1], simp862_0[3:3]);
  C2 I77 (icomplete_0, simp863_0[0:0], simp863_0[1:1]);
  C2 I78 (o_0r0[0:0], i_0r0[0:0], gsel_0);
  C2 I79 (o_0r0[1:1], i_0r0[1:1], gsel_0);
  C2 I80 (o_0r0[2:2], i_0r0[2:2], gsel_0);
  C2 I81 (o_0r0[3:3], i_0r0[3:3], gsel_0);
  C2 I82 (o_0r0[4:4], i_0r0[4:4], gsel_0);
  C2 I83 (o_0r0[5:5], i_0r0[5:5], gsel_0);
  C2 I84 (o_0r0[6:6], i_0r0[6:6], gsel_0);
  C2 I85 (o_0r0[7:7], i_0r0[7:7], gsel_0);
  C2 I86 (o_0r0[8:8], i_0r0[8:8], gsel_0);
  C2 I87 (o_0r0[9:9], i_0r0[9:9], gsel_0);
  C2 I88 (o_0r0[10:10], i_0r0[10:10], gsel_0);
  C2 I89 (o_0r0[11:11], i_0r0[11:11], gsel_0);
  C2 I90 (o_0r0[12:12], i_0r0[12:12], gsel_0);
  C2 I91 (o_0r0[13:13], i_0r0[13:13], gsel_0);
  C2 I92 (o_0r0[14:14], i_0r0[14:14], gsel_0);
  C2 I93 (o_0r0[15:15], i_0r0[15:15], gsel_0);
  C2 I94 (o_0r0[16:16], i_0r0[16:16], gsel_0);
  C2 I95 (o_0r0[17:17], i_0r0[17:17], gsel_0);
  C2 I96 (o_0r0[18:18], i_0r0[18:18], gsel_0);
  C2 I97 (o_0r0[19:19], i_0r0[19:19], gsel_0);
  C2 I98 (o_0r0[20:20], i_0r0[20:20], gsel_0);
  C2 I99 (o_0r0[21:21], i_0r0[21:21], gsel_0);
  C2 I100 (o_0r0[22:22], i_0r0[22:22], gsel_0);
  C2 I101 (o_0r0[23:23], i_0r0[23:23], gsel_0);
  C2 I102 (o_0r0[24:24], i_0r0[24:24], gsel_0);
  C2 I103 (o_0r0[25:25], i_0r0[25:25], gsel_0);
  C2 I104 (o_0r0[26:26], i_0r0[26:26], gsel_0);
  C2 I105 (o_0r0[27:27], i_0r0[27:27], gsel_0);
  C2 I106 (o_0r0[28:28], i_0r0[28:28], gsel_0);
  C2 I107 (o_0r0[29:29], i_0r0[29:29], gsel_0);
  C2 I108 (o_0r0[30:30], i_0r0[30:30], gsel_0);
  C2 I109 (o_0r0[31:31], i_0r0[31:31], gsel_0);
  C2 I110 (o_1r0[0:0], i_0r0[0:0], gsel_1);
  C2 I111 (o_1r0[1:1], i_0r0[1:1], gsel_1);
  C2 I112 (o_1r0[2:2], i_0r0[2:2], gsel_1);
  C2 I113 (o_1r0[3:3], i_0r0[3:3], gsel_1);
  C2 I114 (o_1r0[4:4], i_0r0[4:4], gsel_1);
  C2 I115 (o_1r0[5:5], i_0r0[5:5], gsel_1);
  C2 I116 (o_1r0[6:6], i_0r0[6:6], gsel_1);
  C2 I117 (o_1r0[7:7], i_0r0[7:7], gsel_1);
  C2 I118 (o_1r0[8:8], i_0r0[8:8], gsel_1);
  C2 I119 (o_1r0[9:9], i_0r0[9:9], gsel_1);
  C2 I120 (o_1r0[10:10], i_0r0[10:10], gsel_1);
  C2 I121 (o_1r0[11:11], i_0r0[11:11], gsel_1);
  C2 I122 (o_1r0[12:12], i_0r0[12:12], gsel_1);
  C2 I123 (o_1r0[13:13], i_0r0[13:13], gsel_1);
  C2 I124 (o_1r0[14:14], i_0r0[14:14], gsel_1);
  C2 I125 (o_1r0[15:15], i_0r0[15:15], gsel_1);
  C2 I126 (o_1r0[16:16], i_0r0[16:16], gsel_1);
  C2 I127 (o_1r0[17:17], i_0r0[17:17], gsel_1);
  C2 I128 (o_1r0[18:18], i_0r0[18:18], gsel_1);
  C2 I129 (o_1r0[19:19], i_0r0[19:19], gsel_1);
  C2 I130 (o_1r0[20:20], i_0r0[20:20], gsel_1);
  C2 I131 (o_1r0[21:21], i_0r0[21:21], gsel_1);
  C2 I132 (o_1r0[22:22], i_0r0[22:22], gsel_1);
  C2 I133 (o_1r0[23:23], i_0r0[23:23], gsel_1);
  C2 I134 (o_1r0[24:24], i_0r0[24:24], gsel_1);
  C2 I135 (o_1r0[25:25], i_0r0[25:25], gsel_1);
  C2 I136 (o_1r0[26:26], i_0r0[26:26], gsel_1);
  C2 I137 (o_1r0[27:27], i_0r0[27:27], gsel_1);
  C2 I138 (o_1r0[28:28], i_0r0[28:28], gsel_1);
  C2 I139 (o_1r0[29:29], i_0r0[29:29], gsel_1);
  C2 I140 (o_1r0[30:30], i_0r0[30:30], gsel_1);
  C2 I141 (o_1r0[31:31], i_0r0[31:31], gsel_1);
  C2 I142 (o_2r0[0:0], i_0r0[0:0], gsel_2);
  C2 I143 (o_2r0[1:1], i_0r0[1:1], gsel_2);
  C2 I144 (o_2r0[2:2], i_0r0[2:2], gsel_2);
  C2 I145 (o_2r0[3:3], i_0r0[3:3], gsel_2);
  C2 I146 (o_2r0[4:4], i_0r0[4:4], gsel_2);
  C2 I147 (o_2r0[5:5], i_0r0[5:5], gsel_2);
  C2 I148 (o_2r0[6:6], i_0r0[6:6], gsel_2);
  C2 I149 (o_2r0[7:7], i_0r0[7:7], gsel_2);
  C2 I150 (o_2r0[8:8], i_0r0[8:8], gsel_2);
  C2 I151 (o_2r0[9:9], i_0r0[9:9], gsel_2);
  C2 I152 (o_2r0[10:10], i_0r0[10:10], gsel_2);
  C2 I153 (o_2r0[11:11], i_0r0[11:11], gsel_2);
  C2 I154 (o_2r0[12:12], i_0r0[12:12], gsel_2);
  C2 I155 (o_2r0[13:13], i_0r0[13:13], gsel_2);
  C2 I156 (o_2r0[14:14], i_0r0[14:14], gsel_2);
  C2 I157 (o_2r0[15:15], i_0r0[15:15], gsel_2);
  C2 I158 (o_2r0[16:16], i_0r0[16:16], gsel_2);
  C2 I159 (o_2r0[17:17], i_0r0[17:17], gsel_2);
  C2 I160 (o_2r0[18:18], i_0r0[18:18], gsel_2);
  C2 I161 (o_2r0[19:19], i_0r0[19:19], gsel_2);
  C2 I162 (o_2r0[20:20], i_0r0[20:20], gsel_2);
  C2 I163 (o_2r0[21:21], i_0r0[21:21], gsel_2);
  C2 I164 (o_2r0[22:22], i_0r0[22:22], gsel_2);
  C2 I165 (o_2r0[23:23], i_0r0[23:23], gsel_2);
  C2 I166 (o_2r0[24:24], i_0r0[24:24], gsel_2);
  C2 I167 (o_2r0[25:25], i_0r0[25:25], gsel_2);
  C2 I168 (o_2r0[26:26], i_0r0[26:26], gsel_2);
  C2 I169 (o_2r0[27:27], i_0r0[27:27], gsel_2);
  C2 I170 (o_2r0[28:28], i_0r0[28:28], gsel_2);
  C2 I171 (o_2r0[29:29], i_0r0[29:29], gsel_2);
  C2 I172 (o_2r0[30:30], i_0r0[30:30], gsel_2);
  C2 I173 (o_2r0[31:31], i_0r0[31:31], gsel_2);
  C2 I174 (o_3r0[0:0], i_0r0[0:0], gsel_3);
  C2 I175 (o_3r0[1:1], i_0r0[1:1], gsel_3);
  C2 I176 (o_3r0[2:2], i_0r0[2:2], gsel_3);
  C2 I177 (o_3r0[3:3], i_0r0[3:3], gsel_3);
  C2 I178 (o_3r0[4:4], i_0r0[4:4], gsel_3);
  C2 I179 (o_3r0[5:5], i_0r0[5:5], gsel_3);
  C2 I180 (o_3r0[6:6], i_0r0[6:6], gsel_3);
  C2 I181 (o_3r0[7:7], i_0r0[7:7], gsel_3);
  C2 I182 (o_3r0[8:8], i_0r0[8:8], gsel_3);
  C2 I183 (o_3r0[9:9], i_0r0[9:9], gsel_3);
  C2 I184 (o_3r0[10:10], i_0r0[10:10], gsel_3);
  C2 I185 (o_3r0[11:11], i_0r0[11:11], gsel_3);
  C2 I186 (o_3r0[12:12], i_0r0[12:12], gsel_3);
  C2 I187 (o_3r0[13:13], i_0r0[13:13], gsel_3);
  C2 I188 (o_3r0[14:14], i_0r0[14:14], gsel_3);
  C2 I189 (o_3r0[15:15], i_0r0[15:15], gsel_3);
  C2 I190 (o_3r0[16:16], i_0r0[16:16], gsel_3);
  C2 I191 (o_3r0[17:17], i_0r0[17:17], gsel_3);
  C2 I192 (o_3r0[18:18], i_0r0[18:18], gsel_3);
  C2 I193 (o_3r0[19:19], i_0r0[19:19], gsel_3);
  C2 I194 (o_3r0[20:20], i_0r0[20:20], gsel_3);
  C2 I195 (o_3r0[21:21], i_0r0[21:21], gsel_3);
  C2 I196 (o_3r0[22:22], i_0r0[22:22], gsel_3);
  C2 I197 (o_3r0[23:23], i_0r0[23:23], gsel_3);
  C2 I198 (o_3r0[24:24], i_0r0[24:24], gsel_3);
  C2 I199 (o_3r0[25:25], i_0r0[25:25], gsel_3);
  C2 I200 (o_3r0[26:26], i_0r0[26:26], gsel_3);
  C2 I201 (o_3r0[27:27], i_0r0[27:27], gsel_3);
  C2 I202 (o_3r0[28:28], i_0r0[28:28], gsel_3);
  C2 I203 (o_3r0[29:29], i_0r0[29:29], gsel_3);
  C2 I204 (o_3r0[30:30], i_0r0[30:30], gsel_3);
  C2 I205 (o_3r0[31:31], i_0r0[31:31], gsel_3);
  C2 I206 (o_4r0[0:0], i_0r0[0:0], gsel_4);
  C2 I207 (o_4r0[1:1], i_0r0[1:1], gsel_4);
  C2 I208 (o_4r0[2:2], i_0r0[2:2], gsel_4);
  C2 I209 (o_4r0[3:3], i_0r0[3:3], gsel_4);
  C2 I210 (o_4r0[4:4], i_0r0[4:4], gsel_4);
  C2 I211 (o_4r0[5:5], i_0r0[5:5], gsel_4);
  C2 I212 (o_4r0[6:6], i_0r0[6:6], gsel_4);
  C2 I213 (o_4r0[7:7], i_0r0[7:7], gsel_4);
  C2 I214 (o_4r0[8:8], i_0r0[8:8], gsel_4);
  C2 I215 (o_4r0[9:9], i_0r0[9:9], gsel_4);
  C2 I216 (o_4r0[10:10], i_0r0[10:10], gsel_4);
  C2 I217 (o_4r0[11:11], i_0r0[11:11], gsel_4);
  C2 I218 (o_4r0[12:12], i_0r0[12:12], gsel_4);
  C2 I219 (o_4r0[13:13], i_0r0[13:13], gsel_4);
  C2 I220 (o_4r0[14:14], i_0r0[14:14], gsel_4);
  C2 I221 (o_4r0[15:15], i_0r0[15:15], gsel_4);
  C2 I222 (o_4r0[16:16], i_0r0[16:16], gsel_4);
  C2 I223 (o_4r0[17:17], i_0r0[17:17], gsel_4);
  C2 I224 (o_4r0[18:18], i_0r0[18:18], gsel_4);
  C2 I225 (o_4r0[19:19], i_0r0[19:19], gsel_4);
  C2 I226 (o_4r0[20:20], i_0r0[20:20], gsel_4);
  C2 I227 (o_4r0[21:21], i_0r0[21:21], gsel_4);
  C2 I228 (o_4r0[22:22], i_0r0[22:22], gsel_4);
  C2 I229 (o_4r0[23:23], i_0r0[23:23], gsel_4);
  C2 I230 (o_4r0[24:24], i_0r0[24:24], gsel_4);
  C2 I231 (o_4r0[25:25], i_0r0[25:25], gsel_4);
  C2 I232 (o_4r0[26:26], i_0r0[26:26], gsel_4);
  C2 I233 (o_4r0[27:27], i_0r0[27:27], gsel_4);
  C2 I234 (o_4r0[28:28], i_0r0[28:28], gsel_4);
  C2 I235 (o_4r0[29:29], i_0r0[29:29], gsel_4);
  C2 I236 (o_4r0[30:30], i_0r0[30:30], gsel_4);
  C2 I237 (o_4r0[31:31], i_0r0[31:31], gsel_4);
  C2 I238 (o_5r0[0:0], i_0r0[0:0], gsel_5);
  C2 I239 (o_5r0[1:1], i_0r0[1:1], gsel_5);
  C2 I240 (o_5r0[2:2], i_0r0[2:2], gsel_5);
  C2 I241 (o_5r0[3:3], i_0r0[3:3], gsel_5);
  C2 I242 (o_5r0[4:4], i_0r0[4:4], gsel_5);
  C2 I243 (o_5r0[5:5], i_0r0[5:5], gsel_5);
  C2 I244 (o_5r0[6:6], i_0r0[6:6], gsel_5);
  C2 I245 (o_5r0[7:7], i_0r0[7:7], gsel_5);
  C2 I246 (o_5r0[8:8], i_0r0[8:8], gsel_5);
  C2 I247 (o_5r0[9:9], i_0r0[9:9], gsel_5);
  C2 I248 (o_5r0[10:10], i_0r0[10:10], gsel_5);
  C2 I249 (o_5r0[11:11], i_0r0[11:11], gsel_5);
  C2 I250 (o_5r0[12:12], i_0r0[12:12], gsel_5);
  C2 I251 (o_5r0[13:13], i_0r0[13:13], gsel_5);
  C2 I252 (o_5r0[14:14], i_0r0[14:14], gsel_5);
  C2 I253 (o_5r0[15:15], i_0r0[15:15], gsel_5);
  C2 I254 (o_5r0[16:16], i_0r0[16:16], gsel_5);
  C2 I255 (o_5r0[17:17], i_0r0[17:17], gsel_5);
  C2 I256 (o_5r0[18:18], i_0r0[18:18], gsel_5);
  C2 I257 (o_5r0[19:19], i_0r0[19:19], gsel_5);
  C2 I258 (o_5r0[20:20], i_0r0[20:20], gsel_5);
  C2 I259 (o_5r0[21:21], i_0r0[21:21], gsel_5);
  C2 I260 (o_5r0[22:22], i_0r0[22:22], gsel_5);
  C2 I261 (o_5r0[23:23], i_0r0[23:23], gsel_5);
  C2 I262 (o_5r0[24:24], i_0r0[24:24], gsel_5);
  C2 I263 (o_5r0[25:25], i_0r0[25:25], gsel_5);
  C2 I264 (o_5r0[26:26], i_0r0[26:26], gsel_5);
  C2 I265 (o_5r0[27:27], i_0r0[27:27], gsel_5);
  C2 I266 (o_5r0[28:28], i_0r0[28:28], gsel_5);
  C2 I267 (o_5r0[29:29], i_0r0[29:29], gsel_5);
  C2 I268 (o_5r0[30:30], i_0r0[30:30], gsel_5);
  C2 I269 (o_5r0[31:31], i_0r0[31:31], gsel_5);
  C2 I270 (o_6r0[0:0], i_0r0[0:0], gsel_6);
  C2 I271 (o_6r0[1:1], i_0r0[1:1], gsel_6);
  C2 I272 (o_6r0[2:2], i_0r0[2:2], gsel_6);
  C2 I273 (o_6r0[3:3], i_0r0[3:3], gsel_6);
  C2 I274 (o_6r0[4:4], i_0r0[4:4], gsel_6);
  C2 I275 (o_6r0[5:5], i_0r0[5:5], gsel_6);
  C2 I276 (o_6r0[6:6], i_0r0[6:6], gsel_6);
  C2 I277 (o_6r0[7:7], i_0r0[7:7], gsel_6);
  C2 I278 (o_6r0[8:8], i_0r0[8:8], gsel_6);
  C2 I279 (o_6r0[9:9], i_0r0[9:9], gsel_6);
  C2 I280 (o_6r0[10:10], i_0r0[10:10], gsel_6);
  C2 I281 (o_6r0[11:11], i_0r0[11:11], gsel_6);
  C2 I282 (o_6r0[12:12], i_0r0[12:12], gsel_6);
  C2 I283 (o_6r0[13:13], i_0r0[13:13], gsel_6);
  C2 I284 (o_6r0[14:14], i_0r0[14:14], gsel_6);
  C2 I285 (o_6r0[15:15], i_0r0[15:15], gsel_6);
  C2 I286 (o_6r0[16:16], i_0r0[16:16], gsel_6);
  C2 I287 (o_6r0[17:17], i_0r0[17:17], gsel_6);
  C2 I288 (o_6r0[18:18], i_0r0[18:18], gsel_6);
  C2 I289 (o_6r0[19:19], i_0r0[19:19], gsel_6);
  C2 I290 (o_6r0[20:20], i_0r0[20:20], gsel_6);
  C2 I291 (o_6r0[21:21], i_0r0[21:21], gsel_6);
  C2 I292 (o_6r0[22:22], i_0r0[22:22], gsel_6);
  C2 I293 (o_6r0[23:23], i_0r0[23:23], gsel_6);
  C2 I294 (o_6r0[24:24], i_0r0[24:24], gsel_6);
  C2 I295 (o_6r0[25:25], i_0r0[25:25], gsel_6);
  C2 I296 (o_6r0[26:26], i_0r0[26:26], gsel_6);
  C2 I297 (o_6r0[27:27], i_0r0[27:27], gsel_6);
  C2 I298 (o_6r0[28:28], i_0r0[28:28], gsel_6);
  C2 I299 (o_6r0[29:29], i_0r0[29:29], gsel_6);
  C2 I300 (o_6r0[30:30], i_0r0[30:30], gsel_6);
  C2 I301 (o_6r0[31:31], i_0r0[31:31], gsel_6);
  C2 I302 (o_7r0[0:0], i_0r0[0:0], gsel_7);
  C2 I303 (o_7r0[1:1], i_0r0[1:1], gsel_7);
  C2 I304 (o_7r0[2:2], i_0r0[2:2], gsel_7);
  C2 I305 (o_7r0[3:3], i_0r0[3:3], gsel_7);
  C2 I306 (o_7r0[4:4], i_0r0[4:4], gsel_7);
  C2 I307 (o_7r0[5:5], i_0r0[5:5], gsel_7);
  C2 I308 (o_7r0[6:6], i_0r0[6:6], gsel_7);
  C2 I309 (o_7r0[7:7], i_0r0[7:7], gsel_7);
  C2 I310 (o_7r0[8:8], i_0r0[8:8], gsel_7);
  C2 I311 (o_7r0[9:9], i_0r0[9:9], gsel_7);
  C2 I312 (o_7r0[10:10], i_0r0[10:10], gsel_7);
  C2 I313 (o_7r0[11:11], i_0r0[11:11], gsel_7);
  C2 I314 (o_7r0[12:12], i_0r0[12:12], gsel_7);
  C2 I315 (o_7r0[13:13], i_0r0[13:13], gsel_7);
  C2 I316 (o_7r0[14:14], i_0r0[14:14], gsel_7);
  C2 I317 (o_7r0[15:15], i_0r0[15:15], gsel_7);
  C2 I318 (o_7r0[16:16], i_0r0[16:16], gsel_7);
  C2 I319 (o_7r0[17:17], i_0r0[17:17], gsel_7);
  C2 I320 (o_7r0[18:18], i_0r0[18:18], gsel_7);
  C2 I321 (o_7r0[19:19], i_0r0[19:19], gsel_7);
  C2 I322 (o_7r0[20:20], i_0r0[20:20], gsel_7);
  C2 I323 (o_7r0[21:21], i_0r0[21:21], gsel_7);
  C2 I324 (o_7r0[22:22], i_0r0[22:22], gsel_7);
  C2 I325 (o_7r0[23:23], i_0r0[23:23], gsel_7);
  C2 I326 (o_7r0[24:24], i_0r0[24:24], gsel_7);
  C2 I327 (o_7r0[25:25], i_0r0[25:25], gsel_7);
  C2 I328 (o_7r0[26:26], i_0r0[26:26], gsel_7);
  C2 I329 (o_7r0[27:27], i_0r0[27:27], gsel_7);
  C2 I330 (o_7r0[28:28], i_0r0[28:28], gsel_7);
  C2 I331 (o_7r0[29:29], i_0r0[29:29], gsel_7);
  C2 I332 (o_7r0[30:30], i_0r0[30:30], gsel_7);
  C2 I333 (o_7r0[31:31], i_0r0[31:31], gsel_7);
  C2 I334 (o_0r1[0:0], i_0r1[0:0], gsel_0);
  C2 I335 (o_0r1[1:1], i_0r1[1:1], gsel_0);
  C2 I336 (o_0r1[2:2], i_0r1[2:2], gsel_0);
  C2 I337 (o_0r1[3:3], i_0r1[3:3], gsel_0);
  C2 I338 (o_0r1[4:4], i_0r1[4:4], gsel_0);
  C2 I339 (o_0r1[5:5], i_0r1[5:5], gsel_0);
  C2 I340 (o_0r1[6:6], i_0r1[6:6], gsel_0);
  C2 I341 (o_0r1[7:7], i_0r1[7:7], gsel_0);
  C2 I342 (o_0r1[8:8], i_0r1[8:8], gsel_0);
  C2 I343 (o_0r1[9:9], i_0r1[9:9], gsel_0);
  C2 I344 (o_0r1[10:10], i_0r1[10:10], gsel_0);
  C2 I345 (o_0r1[11:11], i_0r1[11:11], gsel_0);
  C2 I346 (o_0r1[12:12], i_0r1[12:12], gsel_0);
  C2 I347 (o_0r1[13:13], i_0r1[13:13], gsel_0);
  C2 I348 (o_0r1[14:14], i_0r1[14:14], gsel_0);
  C2 I349 (o_0r1[15:15], i_0r1[15:15], gsel_0);
  C2 I350 (o_0r1[16:16], i_0r1[16:16], gsel_0);
  C2 I351 (o_0r1[17:17], i_0r1[17:17], gsel_0);
  C2 I352 (o_0r1[18:18], i_0r1[18:18], gsel_0);
  C2 I353 (o_0r1[19:19], i_0r1[19:19], gsel_0);
  C2 I354 (o_0r1[20:20], i_0r1[20:20], gsel_0);
  C2 I355 (o_0r1[21:21], i_0r1[21:21], gsel_0);
  C2 I356 (o_0r1[22:22], i_0r1[22:22], gsel_0);
  C2 I357 (o_0r1[23:23], i_0r1[23:23], gsel_0);
  C2 I358 (o_0r1[24:24], i_0r1[24:24], gsel_0);
  C2 I359 (o_0r1[25:25], i_0r1[25:25], gsel_0);
  C2 I360 (o_0r1[26:26], i_0r1[26:26], gsel_0);
  C2 I361 (o_0r1[27:27], i_0r1[27:27], gsel_0);
  C2 I362 (o_0r1[28:28], i_0r1[28:28], gsel_0);
  C2 I363 (o_0r1[29:29], i_0r1[29:29], gsel_0);
  C2 I364 (o_0r1[30:30], i_0r1[30:30], gsel_0);
  C2 I365 (o_0r1[31:31], i_0r1[31:31], gsel_0);
  C2 I366 (o_1r1[0:0], i_0r1[0:0], gsel_1);
  C2 I367 (o_1r1[1:1], i_0r1[1:1], gsel_1);
  C2 I368 (o_1r1[2:2], i_0r1[2:2], gsel_1);
  C2 I369 (o_1r1[3:3], i_0r1[3:3], gsel_1);
  C2 I370 (o_1r1[4:4], i_0r1[4:4], gsel_1);
  C2 I371 (o_1r1[5:5], i_0r1[5:5], gsel_1);
  C2 I372 (o_1r1[6:6], i_0r1[6:6], gsel_1);
  C2 I373 (o_1r1[7:7], i_0r1[7:7], gsel_1);
  C2 I374 (o_1r1[8:8], i_0r1[8:8], gsel_1);
  C2 I375 (o_1r1[9:9], i_0r1[9:9], gsel_1);
  C2 I376 (o_1r1[10:10], i_0r1[10:10], gsel_1);
  C2 I377 (o_1r1[11:11], i_0r1[11:11], gsel_1);
  C2 I378 (o_1r1[12:12], i_0r1[12:12], gsel_1);
  C2 I379 (o_1r1[13:13], i_0r1[13:13], gsel_1);
  C2 I380 (o_1r1[14:14], i_0r1[14:14], gsel_1);
  C2 I381 (o_1r1[15:15], i_0r1[15:15], gsel_1);
  C2 I382 (o_1r1[16:16], i_0r1[16:16], gsel_1);
  C2 I383 (o_1r1[17:17], i_0r1[17:17], gsel_1);
  C2 I384 (o_1r1[18:18], i_0r1[18:18], gsel_1);
  C2 I385 (o_1r1[19:19], i_0r1[19:19], gsel_1);
  C2 I386 (o_1r1[20:20], i_0r1[20:20], gsel_1);
  C2 I387 (o_1r1[21:21], i_0r1[21:21], gsel_1);
  C2 I388 (o_1r1[22:22], i_0r1[22:22], gsel_1);
  C2 I389 (o_1r1[23:23], i_0r1[23:23], gsel_1);
  C2 I390 (o_1r1[24:24], i_0r1[24:24], gsel_1);
  C2 I391 (o_1r1[25:25], i_0r1[25:25], gsel_1);
  C2 I392 (o_1r1[26:26], i_0r1[26:26], gsel_1);
  C2 I393 (o_1r1[27:27], i_0r1[27:27], gsel_1);
  C2 I394 (o_1r1[28:28], i_0r1[28:28], gsel_1);
  C2 I395 (o_1r1[29:29], i_0r1[29:29], gsel_1);
  C2 I396 (o_1r1[30:30], i_0r1[30:30], gsel_1);
  C2 I397 (o_1r1[31:31], i_0r1[31:31], gsel_1);
  C2 I398 (o_2r1[0:0], i_0r1[0:0], gsel_2);
  C2 I399 (o_2r1[1:1], i_0r1[1:1], gsel_2);
  C2 I400 (o_2r1[2:2], i_0r1[2:2], gsel_2);
  C2 I401 (o_2r1[3:3], i_0r1[3:3], gsel_2);
  C2 I402 (o_2r1[4:4], i_0r1[4:4], gsel_2);
  C2 I403 (o_2r1[5:5], i_0r1[5:5], gsel_2);
  C2 I404 (o_2r1[6:6], i_0r1[6:6], gsel_2);
  C2 I405 (o_2r1[7:7], i_0r1[7:7], gsel_2);
  C2 I406 (o_2r1[8:8], i_0r1[8:8], gsel_2);
  C2 I407 (o_2r1[9:9], i_0r1[9:9], gsel_2);
  C2 I408 (o_2r1[10:10], i_0r1[10:10], gsel_2);
  C2 I409 (o_2r1[11:11], i_0r1[11:11], gsel_2);
  C2 I410 (o_2r1[12:12], i_0r1[12:12], gsel_2);
  C2 I411 (o_2r1[13:13], i_0r1[13:13], gsel_2);
  C2 I412 (o_2r1[14:14], i_0r1[14:14], gsel_2);
  C2 I413 (o_2r1[15:15], i_0r1[15:15], gsel_2);
  C2 I414 (o_2r1[16:16], i_0r1[16:16], gsel_2);
  C2 I415 (o_2r1[17:17], i_0r1[17:17], gsel_2);
  C2 I416 (o_2r1[18:18], i_0r1[18:18], gsel_2);
  C2 I417 (o_2r1[19:19], i_0r1[19:19], gsel_2);
  C2 I418 (o_2r1[20:20], i_0r1[20:20], gsel_2);
  C2 I419 (o_2r1[21:21], i_0r1[21:21], gsel_2);
  C2 I420 (o_2r1[22:22], i_0r1[22:22], gsel_2);
  C2 I421 (o_2r1[23:23], i_0r1[23:23], gsel_2);
  C2 I422 (o_2r1[24:24], i_0r1[24:24], gsel_2);
  C2 I423 (o_2r1[25:25], i_0r1[25:25], gsel_2);
  C2 I424 (o_2r1[26:26], i_0r1[26:26], gsel_2);
  C2 I425 (o_2r1[27:27], i_0r1[27:27], gsel_2);
  C2 I426 (o_2r1[28:28], i_0r1[28:28], gsel_2);
  C2 I427 (o_2r1[29:29], i_0r1[29:29], gsel_2);
  C2 I428 (o_2r1[30:30], i_0r1[30:30], gsel_2);
  C2 I429 (o_2r1[31:31], i_0r1[31:31], gsel_2);
  C2 I430 (o_3r1[0:0], i_0r1[0:0], gsel_3);
  C2 I431 (o_3r1[1:1], i_0r1[1:1], gsel_3);
  C2 I432 (o_3r1[2:2], i_0r1[2:2], gsel_3);
  C2 I433 (o_3r1[3:3], i_0r1[3:3], gsel_3);
  C2 I434 (o_3r1[4:4], i_0r1[4:4], gsel_3);
  C2 I435 (o_3r1[5:5], i_0r1[5:5], gsel_3);
  C2 I436 (o_3r1[6:6], i_0r1[6:6], gsel_3);
  C2 I437 (o_3r1[7:7], i_0r1[7:7], gsel_3);
  C2 I438 (o_3r1[8:8], i_0r1[8:8], gsel_3);
  C2 I439 (o_3r1[9:9], i_0r1[9:9], gsel_3);
  C2 I440 (o_3r1[10:10], i_0r1[10:10], gsel_3);
  C2 I441 (o_3r1[11:11], i_0r1[11:11], gsel_3);
  C2 I442 (o_3r1[12:12], i_0r1[12:12], gsel_3);
  C2 I443 (o_3r1[13:13], i_0r1[13:13], gsel_3);
  C2 I444 (o_3r1[14:14], i_0r1[14:14], gsel_3);
  C2 I445 (o_3r1[15:15], i_0r1[15:15], gsel_3);
  C2 I446 (o_3r1[16:16], i_0r1[16:16], gsel_3);
  C2 I447 (o_3r1[17:17], i_0r1[17:17], gsel_3);
  C2 I448 (o_3r1[18:18], i_0r1[18:18], gsel_3);
  C2 I449 (o_3r1[19:19], i_0r1[19:19], gsel_3);
  C2 I450 (o_3r1[20:20], i_0r1[20:20], gsel_3);
  C2 I451 (o_3r1[21:21], i_0r1[21:21], gsel_3);
  C2 I452 (o_3r1[22:22], i_0r1[22:22], gsel_3);
  C2 I453 (o_3r1[23:23], i_0r1[23:23], gsel_3);
  C2 I454 (o_3r1[24:24], i_0r1[24:24], gsel_3);
  C2 I455 (o_3r1[25:25], i_0r1[25:25], gsel_3);
  C2 I456 (o_3r1[26:26], i_0r1[26:26], gsel_3);
  C2 I457 (o_3r1[27:27], i_0r1[27:27], gsel_3);
  C2 I458 (o_3r1[28:28], i_0r1[28:28], gsel_3);
  C2 I459 (o_3r1[29:29], i_0r1[29:29], gsel_3);
  C2 I460 (o_3r1[30:30], i_0r1[30:30], gsel_3);
  C2 I461 (o_3r1[31:31], i_0r1[31:31], gsel_3);
  C2 I462 (o_4r1[0:0], i_0r1[0:0], gsel_4);
  C2 I463 (o_4r1[1:1], i_0r1[1:1], gsel_4);
  C2 I464 (o_4r1[2:2], i_0r1[2:2], gsel_4);
  C2 I465 (o_4r1[3:3], i_0r1[3:3], gsel_4);
  C2 I466 (o_4r1[4:4], i_0r1[4:4], gsel_4);
  C2 I467 (o_4r1[5:5], i_0r1[5:5], gsel_4);
  C2 I468 (o_4r1[6:6], i_0r1[6:6], gsel_4);
  C2 I469 (o_4r1[7:7], i_0r1[7:7], gsel_4);
  C2 I470 (o_4r1[8:8], i_0r1[8:8], gsel_4);
  C2 I471 (o_4r1[9:9], i_0r1[9:9], gsel_4);
  C2 I472 (o_4r1[10:10], i_0r1[10:10], gsel_4);
  C2 I473 (o_4r1[11:11], i_0r1[11:11], gsel_4);
  C2 I474 (o_4r1[12:12], i_0r1[12:12], gsel_4);
  C2 I475 (o_4r1[13:13], i_0r1[13:13], gsel_4);
  C2 I476 (o_4r1[14:14], i_0r1[14:14], gsel_4);
  C2 I477 (o_4r1[15:15], i_0r1[15:15], gsel_4);
  C2 I478 (o_4r1[16:16], i_0r1[16:16], gsel_4);
  C2 I479 (o_4r1[17:17], i_0r1[17:17], gsel_4);
  C2 I480 (o_4r1[18:18], i_0r1[18:18], gsel_4);
  C2 I481 (o_4r1[19:19], i_0r1[19:19], gsel_4);
  C2 I482 (o_4r1[20:20], i_0r1[20:20], gsel_4);
  C2 I483 (o_4r1[21:21], i_0r1[21:21], gsel_4);
  C2 I484 (o_4r1[22:22], i_0r1[22:22], gsel_4);
  C2 I485 (o_4r1[23:23], i_0r1[23:23], gsel_4);
  C2 I486 (o_4r1[24:24], i_0r1[24:24], gsel_4);
  C2 I487 (o_4r1[25:25], i_0r1[25:25], gsel_4);
  C2 I488 (o_4r1[26:26], i_0r1[26:26], gsel_4);
  C2 I489 (o_4r1[27:27], i_0r1[27:27], gsel_4);
  C2 I490 (o_4r1[28:28], i_0r1[28:28], gsel_4);
  C2 I491 (o_4r1[29:29], i_0r1[29:29], gsel_4);
  C2 I492 (o_4r1[30:30], i_0r1[30:30], gsel_4);
  C2 I493 (o_4r1[31:31], i_0r1[31:31], gsel_4);
  C2 I494 (o_5r1[0:0], i_0r1[0:0], gsel_5);
  C2 I495 (o_5r1[1:1], i_0r1[1:1], gsel_5);
  C2 I496 (o_5r1[2:2], i_0r1[2:2], gsel_5);
  C2 I497 (o_5r1[3:3], i_0r1[3:3], gsel_5);
  C2 I498 (o_5r1[4:4], i_0r1[4:4], gsel_5);
  C2 I499 (o_5r1[5:5], i_0r1[5:5], gsel_5);
  C2 I500 (o_5r1[6:6], i_0r1[6:6], gsel_5);
  C2 I501 (o_5r1[7:7], i_0r1[7:7], gsel_5);
  C2 I502 (o_5r1[8:8], i_0r1[8:8], gsel_5);
  C2 I503 (o_5r1[9:9], i_0r1[9:9], gsel_5);
  C2 I504 (o_5r1[10:10], i_0r1[10:10], gsel_5);
  C2 I505 (o_5r1[11:11], i_0r1[11:11], gsel_5);
  C2 I506 (o_5r1[12:12], i_0r1[12:12], gsel_5);
  C2 I507 (o_5r1[13:13], i_0r1[13:13], gsel_5);
  C2 I508 (o_5r1[14:14], i_0r1[14:14], gsel_5);
  C2 I509 (o_5r1[15:15], i_0r1[15:15], gsel_5);
  C2 I510 (o_5r1[16:16], i_0r1[16:16], gsel_5);
  C2 I511 (o_5r1[17:17], i_0r1[17:17], gsel_5);
  C2 I512 (o_5r1[18:18], i_0r1[18:18], gsel_5);
  C2 I513 (o_5r1[19:19], i_0r1[19:19], gsel_5);
  C2 I514 (o_5r1[20:20], i_0r1[20:20], gsel_5);
  C2 I515 (o_5r1[21:21], i_0r1[21:21], gsel_5);
  C2 I516 (o_5r1[22:22], i_0r1[22:22], gsel_5);
  C2 I517 (o_5r1[23:23], i_0r1[23:23], gsel_5);
  C2 I518 (o_5r1[24:24], i_0r1[24:24], gsel_5);
  C2 I519 (o_5r1[25:25], i_0r1[25:25], gsel_5);
  C2 I520 (o_5r1[26:26], i_0r1[26:26], gsel_5);
  C2 I521 (o_5r1[27:27], i_0r1[27:27], gsel_5);
  C2 I522 (o_5r1[28:28], i_0r1[28:28], gsel_5);
  C2 I523 (o_5r1[29:29], i_0r1[29:29], gsel_5);
  C2 I524 (o_5r1[30:30], i_0r1[30:30], gsel_5);
  C2 I525 (o_5r1[31:31], i_0r1[31:31], gsel_5);
  C2 I526 (o_6r1[0:0], i_0r1[0:0], gsel_6);
  C2 I527 (o_6r1[1:1], i_0r1[1:1], gsel_6);
  C2 I528 (o_6r1[2:2], i_0r1[2:2], gsel_6);
  C2 I529 (o_6r1[3:3], i_0r1[3:3], gsel_6);
  C2 I530 (o_6r1[4:4], i_0r1[4:4], gsel_6);
  C2 I531 (o_6r1[5:5], i_0r1[5:5], gsel_6);
  C2 I532 (o_6r1[6:6], i_0r1[6:6], gsel_6);
  C2 I533 (o_6r1[7:7], i_0r1[7:7], gsel_6);
  C2 I534 (o_6r1[8:8], i_0r1[8:8], gsel_6);
  C2 I535 (o_6r1[9:9], i_0r1[9:9], gsel_6);
  C2 I536 (o_6r1[10:10], i_0r1[10:10], gsel_6);
  C2 I537 (o_6r1[11:11], i_0r1[11:11], gsel_6);
  C2 I538 (o_6r1[12:12], i_0r1[12:12], gsel_6);
  C2 I539 (o_6r1[13:13], i_0r1[13:13], gsel_6);
  C2 I540 (o_6r1[14:14], i_0r1[14:14], gsel_6);
  C2 I541 (o_6r1[15:15], i_0r1[15:15], gsel_6);
  C2 I542 (o_6r1[16:16], i_0r1[16:16], gsel_6);
  C2 I543 (o_6r1[17:17], i_0r1[17:17], gsel_6);
  C2 I544 (o_6r1[18:18], i_0r1[18:18], gsel_6);
  C2 I545 (o_6r1[19:19], i_0r1[19:19], gsel_6);
  C2 I546 (o_6r1[20:20], i_0r1[20:20], gsel_6);
  C2 I547 (o_6r1[21:21], i_0r1[21:21], gsel_6);
  C2 I548 (o_6r1[22:22], i_0r1[22:22], gsel_6);
  C2 I549 (o_6r1[23:23], i_0r1[23:23], gsel_6);
  C2 I550 (o_6r1[24:24], i_0r1[24:24], gsel_6);
  C2 I551 (o_6r1[25:25], i_0r1[25:25], gsel_6);
  C2 I552 (o_6r1[26:26], i_0r1[26:26], gsel_6);
  C2 I553 (o_6r1[27:27], i_0r1[27:27], gsel_6);
  C2 I554 (o_6r1[28:28], i_0r1[28:28], gsel_6);
  C2 I555 (o_6r1[29:29], i_0r1[29:29], gsel_6);
  C2 I556 (o_6r1[30:30], i_0r1[30:30], gsel_6);
  C2 I557 (o_6r1[31:31], i_0r1[31:31], gsel_6);
  C2 I558 (o_7r1[0:0], i_0r1[0:0], gsel_7);
  C2 I559 (o_7r1[1:1], i_0r1[1:1], gsel_7);
  C2 I560 (o_7r1[2:2], i_0r1[2:2], gsel_7);
  C2 I561 (o_7r1[3:3], i_0r1[3:3], gsel_7);
  C2 I562 (o_7r1[4:4], i_0r1[4:4], gsel_7);
  C2 I563 (o_7r1[5:5], i_0r1[5:5], gsel_7);
  C2 I564 (o_7r1[6:6], i_0r1[6:6], gsel_7);
  C2 I565 (o_7r1[7:7], i_0r1[7:7], gsel_7);
  C2 I566 (o_7r1[8:8], i_0r1[8:8], gsel_7);
  C2 I567 (o_7r1[9:9], i_0r1[9:9], gsel_7);
  C2 I568 (o_7r1[10:10], i_0r1[10:10], gsel_7);
  C2 I569 (o_7r1[11:11], i_0r1[11:11], gsel_7);
  C2 I570 (o_7r1[12:12], i_0r1[12:12], gsel_7);
  C2 I571 (o_7r1[13:13], i_0r1[13:13], gsel_7);
  C2 I572 (o_7r1[14:14], i_0r1[14:14], gsel_7);
  C2 I573 (o_7r1[15:15], i_0r1[15:15], gsel_7);
  C2 I574 (o_7r1[16:16], i_0r1[16:16], gsel_7);
  C2 I575 (o_7r1[17:17], i_0r1[17:17], gsel_7);
  C2 I576 (o_7r1[18:18], i_0r1[18:18], gsel_7);
  C2 I577 (o_7r1[19:19], i_0r1[19:19], gsel_7);
  C2 I578 (o_7r1[20:20], i_0r1[20:20], gsel_7);
  C2 I579 (o_7r1[21:21], i_0r1[21:21], gsel_7);
  C2 I580 (o_7r1[22:22], i_0r1[22:22], gsel_7);
  C2 I581 (o_7r1[23:23], i_0r1[23:23], gsel_7);
  C2 I582 (o_7r1[24:24], i_0r1[24:24], gsel_7);
  C2 I583 (o_7r1[25:25], i_0r1[25:25], gsel_7);
  C2 I584 (o_7r1[26:26], i_0r1[26:26], gsel_7);
  C2 I585 (o_7r1[27:27], i_0r1[27:27], gsel_7);
  C2 I586 (o_7r1[28:28], i_0r1[28:28], gsel_7);
  C2 I587 (o_7r1[29:29], i_0r1[29:29], gsel_7);
  C2 I588 (o_7r1[30:30], i_0r1[30:30], gsel_7);
  C2 I589 (o_7r1[31:31], i_0r1[31:31], gsel_7);
  NOR3 I590 (simp5991_0[0:0], o_0a, o_1a, o_2a);
  NOR3 I591 (simp5991_0[1:1], o_3a, o_4a, o_5a);
  NOR2 I592 (simp5991_0[2:2], o_6a, o_7a);
  NAND3 I593 (oack_0, simp5991_0[0:0], simp5991_0[1:1], simp5991_0[2:2]);
  C2 I594 (i_0a, oack_0, icomplete_0);
endmodule

// tkvw32_wo0w32_ro0w32o0w32o0w32o0w32 TeakV "w" 32 [] [0] [0,0,0,0] [Many [32],Many [0],Many [0,0,0,0]
//   ,Many [32,32,32,32]]
module tkvw32_wo0w32_ro0w32o0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  output [31:0] rd_3r0;
  output [31:0] rd_3r1;
  input rd_3a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [2:0] simp6641_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_3r0[0:0], df_0[0:0], rg_3r);
  AND2 I521 (rd_3r0[1:1], df_0[1:1], rg_3r);
  AND2 I522 (rd_3r0[2:2], df_0[2:2], rg_3r);
  AND2 I523 (rd_3r0[3:3], df_0[3:3], rg_3r);
  AND2 I524 (rd_3r0[4:4], df_0[4:4], rg_3r);
  AND2 I525 (rd_3r0[5:5], df_0[5:5], rg_3r);
  AND2 I526 (rd_3r0[6:6], df_0[6:6], rg_3r);
  AND2 I527 (rd_3r0[7:7], df_0[7:7], rg_3r);
  AND2 I528 (rd_3r0[8:8], df_0[8:8], rg_3r);
  AND2 I529 (rd_3r0[9:9], df_0[9:9], rg_3r);
  AND2 I530 (rd_3r0[10:10], df_0[10:10], rg_3r);
  AND2 I531 (rd_3r0[11:11], df_0[11:11], rg_3r);
  AND2 I532 (rd_3r0[12:12], df_0[12:12], rg_3r);
  AND2 I533 (rd_3r0[13:13], df_0[13:13], rg_3r);
  AND2 I534 (rd_3r0[14:14], df_0[14:14], rg_3r);
  AND2 I535 (rd_3r0[15:15], df_0[15:15], rg_3r);
  AND2 I536 (rd_3r0[16:16], df_0[16:16], rg_3r);
  AND2 I537 (rd_3r0[17:17], df_0[17:17], rg_3r);
  AND2 I538 (rd_3r0[18:18], df_0[18:18], rg_3r);
  AND2 I539 (rd_3r0[19:19], df_0[19:19], rg_3r);
  AND2 I540 (rd_3r0[20:20], df_0[20:20], rg_3r);
  AND2 I541 (rd_3r0[21:21], df_0[21:21], rg_3r);
  AND2 I542 (rd_3r0[22:22], df_0[22:22], rg_3r);
  AND2 I543 (rd_3r0[23:23], df_0[23:23], rg_3r);
  AND2 I544 (rd_3r0[24:24], df_0[24:24], rg_3r);
  AND2 I545 (rd_3r0[25:25], df_0[25:25], rg_3r);
  AND2 I546 (rd_3r0[26:26], df_0[26:26], rg_3r);
  AND2 I547 (rd_3r0[27:27], df_0[27:27], rg_3r);
  AND2 I548 (rd_3r0[28:28], df_0[28:28], rg_3r);
  AND2 I549 (rd_3r0[29:29], df_0[29:29], rg_3r);
  AND2 I550 (rd_3r0[30:30], df_0[30:30], rg_3r);
  AND2 I551 (rd_3r0[31:31], df_0[31:31], rg_3r);
  AND2 I552 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I553 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I554 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I555 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I556 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I557 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I558 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I559 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I560 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I561 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I562 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I563 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I564 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I565 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I566 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I567 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I568 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I569 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I570 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I571 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I572 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I573 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I574 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I575 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I576 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I577 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I578 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I579 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I580 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I581 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I582 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I583 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I584 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I585 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I586 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I587 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I588 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I589 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I590 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I591 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I592 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I593 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I594 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I595 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I596 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I597 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I598 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I599 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I600 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I601 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I602 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I603 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I604 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I605 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I606 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I607 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I608 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I609 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I610 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I611 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I612 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I613 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I614 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I615 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I616 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I617 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I618 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I619 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I620 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I621 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I622 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I623 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I624 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I625 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I626 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I627 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I628 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I629 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I630 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I631 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I632 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I633 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I634 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I635 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I636 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I637 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I638 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I639 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I640 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I641 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I642 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I643 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I644 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I645 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I646 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I647 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  AND2 I648 (rd_3r1[0:0], dt_0[0:0], rg_3r);
  AND2 I649 (rd_3r1[1:1], dt_0[1:1], rg_3r);
  AND2 I650 (rd_3r1[2:2], dt_0[2:2], rg_3r);
  AND2 I651 (rd_3r1[3:3], dt_0[3:3], rg_3r);
  AND2 I652 (rd_3r1[4:4], dt_0[4:4], rg_3r);
  AND2 I653 (rd_3r1[5:5], dt_0[5:5], rg_3r);
  AND2 I654 (rd_3r1[6:6], dt_0[6:6], rg_3r);
  AND2 I655 (rd_3r1[7:7], dt_0[7:7], rg_3r);
  AND2 I656 (rd_3r1[8:8], dt_0[8:8], rg_3r);
  AND2 I657 (rd_3r1[9:9], dt_0[9:9], rg_3r);
  AND2 I658 (rd_3r1[10:10], dt_0[10:10], rg_3r);
  AND2 I659 (rd_3r1[11:11], dt_0[11:11], rg_3r);
  AND2 I660 (rd_3r1[12:12], dt_0[12:12], rg_3r);
  AND2 I661 (rd_3r1[13:13], dt_0[13:13], rg_3r);
  AND2 I662 (rd_3r1[14:14], dt_0[14:14], rg_3r);
  AND2 I663 (rd_3r1[15:15], dt_0[15:15], rg_3r);
  AND2 I664 (rd_3r1[16:16], dt_0[16:16], rg_3r);
  AND2 I665 (rd_3r1[17:17], dt_0[17:17], rg_3r);
  AND2 I666 (rd_3r1[18:18], dt_0[18:18], rg_3r);
  AND2 I667 (rd_3r1[19:19], dt_0[19:19], rg_3r);
  AND2 I668 (rd_3r1[20:20], dt_0[20:20], rg_3r);
  AND2 I669 (rd_3r1[21:21], dt_0[21:21], rg_3r);
  AND2 I670 (rd_3r1[22:22], dt_0[22:22], rg_3r);
  AND2 I671 (rd_3r1[23:23], dt_0[23:23], rg_3r);
  AND2 I672 (rd_3r1[24:24], dt_0[24:24], rg_3r);
  AND2 I673 (rd_3r1[25:25], dt_0[25:25], rg_3r);
  AND2 I674 (rd_3r1[26:26], dt_0[26:26], rg_3r);
  AND2 I675 (rd_3r1[27:27], dt_0[27:27], rg_3r);
  AND2 I676 (rd_3r1[28:28], dt_0[28:28], rg_3r);
  AND2 I677 (rd_3r1[29:29], dt_0[29:29], rg_3r);
  AND2 I678 (rd_3r1[30:30], dt_0[30:30], rg_3r);
  AND2 I679 (rd_3r1[31:31], dt_0[31:31], rg_3r);
  NOR3 I680 (simp6641_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I681 (simp6641_0[1:1], rg_3r, rg_0a, rg_1a);
  NOR2 I682 (simp6641_0[2:2], rg_2a, rg_3a);
  NAND3 I683 (anyread_0, simp6641_0[0:0], simp6641_0[1:1], simp6641_0[2:2]);
  BUFF I684 (wg_0a, wd_0a);
  BUFF I685 (rg_0a, rd_0a);
  BUFF I686 (rg_1a, rd_1a);
  BUFF I687 (rg_2a, rd_2a);
  BUFF I688 (rg_3a, rd_3a);
endmodule

// tkvwindow1_wo0w1_ro0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1 TeakV "window" 1 [] [0] [0,0,0,0,
//   0,0,0,0,0,0,0,0] [Many [1],Many [0],Many [0,0,0,0,0,0,0,0,0,0,0,0],Many [1,1,1,1,1,1,1,1,1,1,1,1]]
module tkvwindow1_wo0w1_ro0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rg_5r, rg_5a, rg_6r, rg_6a, rg_7r, rg_7a, rg_8r, rg_8a, rg_9r, rg_9a, rg_10r, rg_10a, rg_11r, rg_11a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, rd_5r0, rd_5r1, rd_5a, rd_6r0, rd_6r1, rd_6a, rd_7r0, rd_7r1, rd_7a, rd_8r0, rd_8r1, rd_8a, rd_9r0, rd_9r1, rd_9a, rd_10r0, rd_10r1, rd_10a, rd_11r0, rd_11r1, rd_11a, reset);
  input wg_0r0;
  input wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  input rg_5r;
  output rg_5a;
  input rg_6r;
  output rg_6a;
  input rg_7r;
  output rg_7a;
  input rg_8r;
  output rg_8a;
  input rg_9r;
  output rg_9a;
  input rg_10r;
  output rg_10a;
  input rg_11r;
  output rg_11a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  output rd_1r0;
  output rd_1r1;
  input rd_1a;
  output rd_2r0;
  output rd_2r1;
  input rd_2a;
  output rd_3r0;
  output rd_3r1;
  input rd_3a;
  output rd_4r0;
  output rd_4r1;
  input rd_4a;
  output rd_5r0;
  output rd_5r1;
  input rd_5a;
  output rd_6r0;
  output rd_6r1;
  input rd_6a;
  output rd_7r0;
  output rd_7r1;
  input rd_7a;
  output rd_8r0;
  output rd_8r1;
  input rd_8a;
  output rd_9r0;
  output rd_9r1;
  input rd_9a;
  output rd_10r0;
  output rd_10r1;
  input rd_10a;
  output rd_11r0;
  output rd_11r1;
  input rd_11a;
  input reset;
  wire wf_0;
  wire wt_0;
  wire df_0;
  wire dt_0;
  wire wc_0;
  wire wacks_0;
  wire wenr_0;
  wire wen_0;
  wire anyread_0;
  wire nreset_0;
  wire drlgf_0;
  wire drlgt_0;
  wire comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire conwgit_0;
  wire conwgif_0;
  wire conwig_0;
  wire [7:0] simp601_0;
  wire [2:0] simp602_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0, wenr_0, nreset_0);
  AND2 I2 (drlgf_0, wf_0, wen_0);
  AND2 I3 (drlgt_0, wt_0, wen_0);
  NOR2 I4 (df_0, dt_0, drlgt_0);
  NOR3 I5 (dt_0, df_0, drlgf_0, reset);
  AO22 I6 (wacks_0, drlgf_0, df_0, drlgt_0, dt_0);
  OR2 I7 (comp0_0, wg_0r0, wg_0r1);
  BUFF I8 (wc_0, comp0_0);
  AND2 I9 (conwgif_0, wg_0r0, conwig_0);
  AND2 I10 (conwgit_0, wg_0r1, conwig_0);
  BUFF I11 (conwigc_0, wc_0);
  AO22 I12 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I13 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I14 (wf_0, conwgif_0);
  BUFF I15 (wt_0, conwgit_0);
  BUFF I16 (wenr_0, wc_0);
  C2 I17 (wd_0r, conwig_0, wacks_0);
  AND2 I18 (rd_0r0, df_0, rg_0r);
  AND2 I19 (rd_1r0, df_0, rg_1r);
  AND2 I20 (rd_2r0, df_0, rg_2r);
  AND2 I21 (rd_3r0, df_0, rg_3r);
  AND2 I22 (rd_4r0, df_0, rg_4r);
  AND2 I23 (rd_5r0, df_0, rg_5r);
  AND2 I24 (rd_6r0, df_0, rg_6r);
  AND2 I25 (rd_7r0, df_0, rg_7r);
  AND2 I26 (rd_8r0, df_0, rg_8r);
  AND2 I27 (rd_9r0, df_0, rg_9r);
  AND2 I28 (rd_10r0, df_0, rg_10r);
  AND2 I29 (rd_11r0, df_0, rg_11r);
  AND2 I30 (rd_0r1, dt_0, rg_0r);
  AND2 I31 (rd_1r1, dt_0, rg_1r);
  AND2 I32 (rd_2r1, dt_0, rg_2r);
  AND2 I33 (rd_3r1, dt_0, rg_3r);
  AND2 I34 (rd_4r1, dt_0, rg_4r);
  AND2 I35 (rd_5r1, dt_0, rg_5r);
  AND2 I36 (rd_6r1, dt_0, rg_6r);
  AND2 I37 (rd_7r1, dt_0, rg_7r);
  AND2 I38 (rd_8r1, dt_0, rg_8r);
  AND2 I39 (rd_9r1, dt_0, rg_9r);
  AND2 I40 (rd_10r1, dt_0, rg_10r);
  AND2 I41 (rd_11r1, dt_0, rg_11r);
  NOR3 I42 (simp601_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I43 (simp601_0[1:1], rg_3r, rg_4r, rg_5r);
  NOR3 I44 (simp601_0[2:2], rg_6r, rg_7r, rg_8r);
  NOR3 I45 (simp601_0[3:3], rg_9r, rg_10r, rg_11r);
  NOR3 I46 (simp601_0[4:4], rg_0a, rg_1a, rg_2a);
  NOR3 I47 (simp601_0[5:5], rg_3a, rg_4a, rg_5a);
  NOR3 I48 (simp601_0[6:6], rg_6a, rg_7a, rg_8a);
  NOR3 I49 (simp601_0[7:7], rg_9a, rg_10a, rg_11a);
  NAND3 I50 (simp602_0[0:0], simp601_0[0:0], simp601_0[1:1], simp601_0[2:2]);
  NAND3 I51 (simp602_0[1:1], simp601_0[3:3], simp601_0[4:4], simp601_0[5:5]);
  NAND2 I52 (simp602_0[2:2], simp601_0[6:6], simp601_0[7:7]);
  OR3 I53 (anyread_0, simp602_0[0:0], simp602_0[1:1], simp602_0[2:2]);
  BUFF I54 (wg_0a, wd_0a);
  BUFF I55 (rg_0a, rd_0a);
  BUFF I56 (rg_1a, rd_1a);
  BUFF I57 (rg_2a, rd_2a);
  BUFF I58 (rg_3a, rd_3a);
  BUFF I59 (rg_4a, rd_4a);
  BUFF I60 (rg_5a, rd_5a);
  BUFF I61 (rg_6a, rd_6a);
  BUFF I62 (rg_7a, rd_7a);
  BUFF I63 (rg_8a, rd_8a);
  BUFF I64 (rg_9a, rd_9a);
  BUFF I65 (rg_10a, rd_10a);
  BUFF I66 (rg_11a, rd_11a);
endmodule

// tkvrEn3_wo0w3_ro0w1o1w1o2w1 TeakV "rEn" 3 [] [0] [0,1,2] [Many [3],Many [0],Many [0,0,0],Many [1,1,1
//   ]]
module tkvrEn3_wo0w3_ro0w1o1w1o2w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [2:0] wg_0r0;
  input [2:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  output rd_1r0;
  output rd_1r1;
  input rd_1a;
  output rd_2r0;
  output rd_2r1;
  input rd_2a;
  input reset;
  wire [2:0] wf_0;
  wire [2:0] wt_0;
  wire [2:0] df_0;
  wire [2:0] dt_0;
  wire wc_0;
  wire [2:0] wacks_0;
  wire [2:0] wenr_0;
  wire [2:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [2:0] drlgf_0;
  wire [2:0] drlgt_0;
  wire [2:0] comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [2:0] conwgit_0;
  wire [2:0] conwgif_0;
  wire conwig_0;
  wire [1:0] simp591_0;
  wire [1:0] simp661_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I5 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I6 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I7 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I8 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I9 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  NOR2 I10 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I11 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I12 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR3 I13 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I14 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I15 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  AO22 I16 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I17 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I18 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  OR2 I19 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I20 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I21 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  C3 I22 (wc_0, comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  AND2 I23 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I24 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I25 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I26 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I27 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I28 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  BUFF I29 (conwigc_0, wc_0);
  AO22 I30 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I31 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I32 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I33 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I34 (wenr_0[0:0], wc_0);
  BUFF I35 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I36 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I37 (wenr_0[1:1], wc_0);
  BUFF I38 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I39 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I40 (wenr_0[2:2], wc_0);
  C3 I41 (simp591_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  BUFF I42 (simp591_0[1:1], wacks_0[2:2]);
  C2 I43 (wd_0r, simp591_0[0:0], simp591_0[1:1]);
  AND2 I44 (rd_0r0, df_0[0:0], rg_0r);
  AND2 I45 (rd_1r0, df_0[1:1], rg_1r);
  AND2 I46 (rd_2r0, df_0[2:2], rg_2r);
  AND2 I47 (rd_0r1, dt_0[0:0], rg_0r);
  AND2 I48 (rd_1r1, dt_0[1:1], rg_1r);
  AND2 I49 (rd_2r1, dt_0[2:2], rg_2r);
  NOR3 I50 (simp661_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I51 (simp661_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I52 (anyread_0, simp661_0[0:0], simp661_0[1:1]);
  BUFF I53 (wg_0a, wd_0a);
  BUFF I54 (rg_0a, rd_0a);
  BUFF I55 (rg_1a, rd_1a);
  BUFF I56 (rg_2a, rd_2a);
endmodule

// tkvwEn1_wo0w1_ro0w1 TeakV "wEn" 1 [] [0] [0] [Many [1],Many [0],Many [0],Many [1]]
module tkvwEn1_wo0w1_ro0w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input wg_0r0;
  input wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  input reset;
  wire wf_0;
  wire wt_0;
  wire df_0;
  wire dt_0;
  wire wc_0;
  wire wacks_0;
  wire wenr_0;
  wire wen_0;
  wire anyread_0;
  wire nreset_0;
  wire drlgf_0;
  wire drlgt_0;
  wire comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire conwgit_0;
  wire conwgif_0;
  wire conwig_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0, wenr_0, nreset_0);
  AND2 I2 (drlgf_0, wf_0, wen_0);
  AND2 I3 (drlgt_0, wt_0, wen_0);
  NOR2 I4 (df_0, dt_0, drlgt_0);
  NOR3 I5 (dt_0, df_0, drlgf_0, reset);
  AO22 I6 (wacks_0, drlgf_0, df_0, drlgt_0, dt_0);
  OR2 I7 (comp0_0, wg_0r0, wg_0r1);
  BUFF I8 (wc_0, comp0_0);
  AND2 I9 (conwgif_0, wg_0r0, conwig_0);
  AND2 I10 (conwgit_0, wg_0r1, conwig_0);
  BUFF I11 (conwigc_0, wc_0);
  AO22 I12 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I13 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I14 (wf_0, conwgif_0);
  BUFF I15 (wt_0, conwgit_0);
  BUFF I16 (wenr_0, wc_0);
  C2 I17 (wd_0r, conwig_0, wacks_0);
  AND2 I18 (rd_0r0, df_0, rg_0r);
  AND2 I19 (rd_0r1, dt_0, rg_0r);
  OR2 I20 (anyread_0, rg_0r, rg_0a);
  BUFF I21 (wg_0a, wd_0a);
  BUFF I22 (rg_0a, rd_0a);
endmodule

// tkvinouts_31032_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 TeakV "inouts[31:0]" 32 [] [0] [0,0,0,0,0,0] 
//   [Many [32],Many [0],Many [0,0,0,0,0,0],Many [32,32,32,32,32,32]]
module tkvinouts_31032_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rg_5r, rg_5a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, rd_5r0, rd_5r1, rd_5a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  input rg_5r;
  output rg_5a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  output [31:0] rd_3r0;
  output [31:0] rd_3r1;
  input rd_3a;
  output [31:0] rd_4r0;
  output [31:0] rd_4r1;
  input rd_4a;
  output [31:0] rd_5r0;
  output [31:0] rd_5r1;
  input rd_5a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [3:0] simp7921_0;
  wire [1:0] simp7922_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_3r0[0:0], df_0[0:0], rg_3r);
  AND2 I521 (rd_3r0[1:1], df_0[1:1], rg_3r);
  AND2 I522 (rd_3r0[2:2], df_0[2:2], rg_3r);
  AND2 I523 (rd_3r0[3:3], df_0[3:3], rg_3r);
  AND2 I524 (rd_3r0[4:4], df_0[4:4], rg_3r);
  AND2 I525 (rd_3r0[5:5], df_0[5:5], rg_3r);
  AND2 I526 (rd_3r0[6:6], df_0[6:6], rg_3r);
  AND2 I527 (rd_3r0[7:7], df_0[7:7], rg_3r);
  AND2 I528 (rd_3r0[8:8], df_0[8:8], rg_3r);
  AND2 I529 (rd_3r0[9:9], df_0[9:9], rg_3r);
  AND2 I530 (rd_3r0[10:10], df_0[10:10], rg_3r);
  AND2 I531 (rd_3r0[11:11], df_0[11:11], rg_3r);
  AND2 I532 (rd_3r0[12:12], df_0[12:12], rg_3r);
  AND2 I533 (rd_3r0[13:13], df_0[13:13], rg_3r);
  AND2 I534 (rd_3r0[14:14], df_0[14:14], rg_3r);
  AND2 I535 (rd_3r0[15:15], df_0[15:15], rg_3r);
  AND2 I536 (rd_3r0[16:16], df_0[16:16], rg_3r);
  AND2 I537 (rd_3r0[17:17], df_0[17:17], rg_3r);
  AND2 I538 (rd_3r0[18:18], df_0[18:18], rg_3r);
  AND2 I539 (rd_3r0[19:19], df_0[19:19], rg_3r);
  AND2 I540 (rd_3r0[20:20], df_0[20:20], rg_3r);
  AND2 I541 (rd_3r0[21:21], df_0[21:21], rg_3r);
  AND2 I542 (rd_3r0[22:22], df_0[22:22], rg_3r);
  AND2 I543 (rd_3r0[23:23], df_0[23:23], rg_3r);
  AND2 I544 (rd_3r0[24:24], df_0[24:24], rg_3r);
  AND2 I545 (rd_3r0[25:25], df_0[25:25], rg_3r);
  AND2 I546 (rd_3r0[26:26], df_0[26:26], rg_3r);
  AND2 I547 (rd_3r0[27:27], df_0[27:27], rg_3r);
  AND2 I548 (rd_3r0[28:28], df_0[28:28], rg_3r);
  AND2 I549 (rd_3r0[29:29], df_0[29:29], rg_3r);
  AND2 I550 (rd_3r0[30:30], df_0[30:30], rg_3r);
  AND2 I551 (rd_3r0[31:31], df_0[31:31], rg_3r);
  AND2 I552 (rd_4r0[0:0], df_0[0:0], rg_4r);
  AND2 I553 (rd_4r0[1:1], df_0[1:1], rg_4r);
  AND2 I554 (rd_4r0[2:2], df_0[2:2], rg_4r);
  AND2 I555 (rd_4r0[3:3], df_0[3:3], rg_4r);
  AND2 I556 (rd_4r0[4:4], df_0[4:4], rg_4r);
  AND2 I557 (rd_4r0[5:5], df_0[5:5], rg_4r);
  AND2 I558 (rd_4r0[6:6], df_0[6:6], rg_4r);
  AND2 I559 (rd_4r0[7:7], df_0[7:7], rg_4r);
  AND2 I560 (rd_4r0[8:8], df_0[8:8], rg_4r);
  AND2 I561 (rd_4r0[9:9], df_0[9:9], rg_4r);
  AND2 I562 (rd_4r0[10:10], df_0[10:10], rg_4r);
  AND2 I563 (rd_4r0[11:11], df_0[11:11], rg_4r);
  AND2 I564 (rd_4r0[12:12], df_0[12:12], rg_4r);
  AND2 I565 (rd_4r0[13:13], df_0[13:13], rg_4r);
  AND2 I566 (rd_4r0[14:14], df_0[14:14], rg_4r);
  AND2 I567 (rd_4r0[15:15], df_0[15:15], rg_4r);
  AND2 I568 (rd_4r0[16:16], df_0[16:16], rg_4r);
  AND2 I569 (rd_4r0[17:17], df_0[17:17], rg_4r);
  AND2 I570 (rd_4r0[18:18], df_0[18:18], rg_4r);
  AND2 I571 (rd_4r0[19:19], df_0[19:19], rg_4r);
  AND2 I572 (rd_4r0[20:20], df_0[20:20], rg_4r);
  AND2 I573 (rd_4r0[21:21], df_0[21:21], rg_4r);
  AND2 I574 (rd_4r0[22:22], df_0[22:22], rg_4r);
  AND2 I575 (rd_4r0[23:23], df_0[23:23], rg_4r);
  AND2 I576 (rd_4r0[24:24], df_0[24:24], rg_4r);
  AND2 I577 (rd_4r0[25:25], df_0[25:25], rg_4r);
  AND2 I578 (rd_4r0[26:26], df_0[26:26], rg_4r);
  AND2 I579 (rd_4r0[27:27], df_0[27:27], rg_4r);
  AND2 I580 (rd_4r0[28:28], df_0[28:28], rg_4r);
  AND2 I581 (rd_4r0[29:29], df_0[29:29], rg_4r);
  AND2 I582 (rd_4r0[30:30], df_0[30:30], rg_4r);
  AND2 I583 (rd_4r0[31:31], df_0[31:31], rg_4r);
  AND2 I584 (rd_5r0[0:0], df_0[0:0], rg_5r);
  AND2 I585 (rd_5r0[1:1], df_0[1:1], rg_5r);
  AND2 I586 (rd_5r0[2:2], df_0[2:2], rg_5r);
  AND2 I587 (rd_5r0[3:3], df_0[3:3], rg_5r);
  AND2 I588 (rd_5r0[4:4], df_0[4:4], rg_5r);
  AND2 I589 (rd_5r0[5:5], df_0[5:5], rg_5r);
  AND2 I590 (rd_5r0[6:6], df_0[6:6], rg_5r);
  AND2 I591 (rd_5r0[7:7], df_0[7:7], rg_5r);
  AND2 I592 (rd_5r0[8:8], df_0[8:8], rg_5r);
  AND2 I593 (rd_5r0[9:9], df_0[9:9], rg_5r);
  AND2 I594 (rd_5r0[10:10], df_0[10:10], rg_5r);
  AND2 I595 (rd_5r0[11:11], df_0[11:11], rg_5r);
  AND2 I596 (rd_5r0[12:12], df_0[12:12], rg_5r);
  AND2 I597 (rd_5r0[13:13], df_0[13:13], rg_5r);
  AND2 I598 (rd_5r0[14:14], df_0[14:14], rg_5r);
  AND2 I599 (rd_5r0[15:15], df_0[15:15], rg_5r);
  AND2 I600 (rd_5r0[16:16], df_0[16:16], rg_5r);
  AND2 I601 (rd_5r0[17:17], df_0[17:17], rg_5r);
  AND2 I602 (rd_5r0[18:18], df_0[18:18], rg_5r);
  AND2 I603 (rd_5r0[19:19], df_0[19:19], rg_5r);
  AND2 I604 (rd_5r0[20:20], df_0[20:20], rg_5r);
  AND2 I605 (rd_5r0[21:21], df_0[21:21], rg_5r);
  AND2 I606 (rd_5r0[22:22], df_0[22:22], rg_5r);
  AND2 I607 (rd_5r0[23:23], df_0[23:23], rg_5r);
  AND2 I608 (rd_5r0[24:24], df_0[24:24], rg_5r);
  AND2 I609 (rd_5r0[25:25], df_0[25:25], rg_5r);
  AND2 I610 (rd_5r0[26:26], df_0[26:26], rg_5r);
  AND2 I611 (rd_5r0[27:27], df_0[27:27], rg_5r);
  AND2 I612 (rd_5r0[28:28], df_0[28:28], rg_5r);
  AND2 I613 (rd_5r0[29:29], df_0[29:29], rg_5r);
  AND2 I614 (rd_5r0[30:30], df_0[30:30], rg_5r);
  AND2 I615 (rd_5r0[31:31], df_0[31:31], rg_5r);
  AND2 I616 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I617 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I618 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I619 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I620 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I621 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I622 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I623 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I624 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I625 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I626 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I627 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I628 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I629 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I630 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I631 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I632 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I633 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I634 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I635 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I636 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I637 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I638 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I639 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I640 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I641 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I642 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I643 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I644 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I645 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I646 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I647 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I648 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I649 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I650 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I651 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I652 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I653 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I654 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I655 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I656 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I657 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I658 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I659 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I660 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I661 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I662 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I663 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I664 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I665 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I666 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I667 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I668 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I669 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I670 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I671 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I672 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I673 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I674 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I675 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I676 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I677 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I678 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I679 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I680 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I681 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I682 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I683 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I684 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I685 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I686 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I687 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I688 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I689 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I690 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I691 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I692 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I693 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I694 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I695 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I696 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I697 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I698 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I699 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I700 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I701 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I702 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I703 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I704 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I705 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I706 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I707 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I708 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I709 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I710 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I711 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  AND2 I712 (rd_3r1[0:0], dt_0[0:0], rg_3r);
  AND2 I713 (rd_3r1[1:1], dt_0[1:1], rg_3r);
  AND2 I714 (rd_3r1[2:2], dt_0[2:2], rg_3r);
  AND2 I715 (rd_3r1[3:3], dt_0[3:3], rg_3r);
  AND2 I716 (rd_3r1[4:4], dt_0[4:4], rg_3r);
  AND2 I717 (rd_3r1[5:5], dt_0[5:5], rg_3r);
  AND2 I718 (rd_3r1[6:6], dt_0[6:6], rg_3r);
  AND2 I719 (rd_3r1[7:7], dt_0[7:7], rg_3r);
  AND2 I720 (rd_3r1[8:8], dt_0[8:8], rg_3r);
  AND2 I721 (rd_3r1[9:9], dt_0[9:9], rg_3r);
  AND2 I722 (rd_3r1[10:10], dt_0[10:10], rg_3r);
  AND2 I723 (rd_3r1[11:11], dt_0[11:11], rg_3r);
  AND2 I724 (rd_3r1[12:12], dt_0[12:12], rg_3r);
  AND2 I725 (rd_3r1[13:13], dt_0[13:13], rg_3r);
  AND2 I726 (rd_3r1[14:14], dt_0[14:14], rg_3r);
  AND2 I727 (rd_3r1[15:15], dt_0[15:15], rg_3r);
  AND2 I728 (rd_3r1[16:16], dt_0[16:16], rg_3r);
  AND2 I729 (rd_3r1[17:17], dt_0[17:17], rg_3r);
  AND2 I730 (rd_3r1[18:18], dt_0[18:18], rg_3r);
  AND2 I731 (rd_3r1[19:19], dt_0[19:19], rg_3r);
  AND2 I732 (rd_3r1[20:20], dt_0[20:20], rg_3r);
  AND2 I733 (rd_3r1[21:21], dt_0[21:21], rg_3r);
  AND2 I734 (rd_3r1[22:22], dt_0[22:22], rg_3r);
  AND2 I735 (rd_3r1[23:23], dt_0[23:23], rg_3r);
  AND2 I736 (rd_3r1[24:24], dt_0[24:24], rg_3r);
  AND2 I737 (rd_3r1[25:25], dt_0[25:25], rg_3r);
  AND2 I738 (rd_3r1[26:26], dt_0[26:26], rg_3r);
  AND2 I739 (rd_3r1[27:27], dt_0[27:27], rg_3r);
  AND2 I740 (rd_3r1[28:28], dt_0[28:28], rg_3r);
  AND2 I741 (rd_3r1[29:29], dt_0[29:29], rg_3r);
  AND2 I742 (rd_3r1[30:30], dt_0[30:30], rg_3r);
  AND2 I743 (rd_3r1[31:31], dt_0[31:31], rg_3r);
  AND2 I744 (rd_4r1[0:0], dt_0[0:0], rg_4r);
  AND2 I745 (rd_4r1[1:1], dt_0[1:1], rg_4r);
  AND2 I746 (rd_4r1[2:2], dt_0[2:2], rg_4r);
  AND2 I747 (rd_4r1[3:3], dt_0[3:3], rg_4r);
  AND2 I748 (rd_4r1[4:4], dt_0[4:4], rg_4r);
  AND2 I749 (rd_4r1[5:5], dt_0[5:5], rg_4r);
  AND2 I750 (rd_4r1[6:6], dt_0[6:6], rg_4r);
  AND2 I751 (rd_4r1[7:7], dt_0[7:7], rg_4r);
  AND2 I752 (rd_4r1[8:8], dt_0[8:8], rg_4r);
  AND2 I753 (rd_4r1[9:9], dt_0[9:9], rg_4r);
  AND2 I754 (rd_4r1[10:10], dt_0[10:10], rg_4r);
  AND2 I755 (rd_4r1[11:11], dt_0[11:11], rg_4r);
  AND2 I756 (rd_4r1[12:12], dt_0[12:12], rg_4r);
  AND2 I757 (rd_4r1[13:13], dt_0[13:13], rg_4r);
  AND2 I758 (rd_4r1[14:14], dt_0[14:14], rg_4r);
  AND2 I759 (rd_4r1[15:15], dt_0[15:15], rg_4r);
  AND2 I760 (rd_4r1[16:16], dt_0[16:16], rg_4r);
  AND2 I761 (rd_4r1[17:17], dt_0[17:17], rg_4r);
  AND2 I762 (rd_4r1[18:18], dt_0[18:18], rg_4r);
  AND2 I763 (rd_4r1[19:19], dt_0[19:19], rg_4r);
  AND2 I764 (rd_4r1[20:20], dt_0[20:20], rg_4r);
  AND2 I765 (rd_4r1[21:21], dt_0[21:21], rg_4r);
  AND2 I766 (rd_4r1[22:22], dt_0[22:22], rg_4r);
  AND2 I767 (rd_4r1[23:23], dt_0[23:23], rg_4r);
  AND2 I768 (rd_4r1[24:24], dt_0[24:24], rg_4r);
  AND2 I769 (rd_4r1[25:25], dt_0[25:25], rg_4r);
  AND2 I770 (rd_4r1[26:26], dt_0[26:26], rg_4r);
  AND2 I771 (rd_4r1[27:27], dt_0[27:27], rg_4r);
  AND2 I772 (rd_4r1[28:28], dt_0[28:28], rg_4r);
  AND2 I773 (rd_4r1[29:29], dt_0[29:29], rg_4r);
  AND2 I774 (rd_4r1[30:30], dt_0[30:30], rg_4r);
  AND2 I775 (rd_4r1[31:31], dt_0[31:31], rg_4r);
  AND2 I776 (rd_5r1[0:0], dt_0[0:0], rg_5r);
  AND2 I777 (rd_5r1[1:1], dt_0[1:1], rg_5r);
  AND2 I778 (rd_5r1[2:2], dt_0[2:2], rg_5r);
  AND2 I779 (rd_5r1[3:3], dt_0[3:3], rg_5r);
  AND2 I780 (rd_5r1[4:4], dt_0[4:4], rg_5r);
  AND2 I781 (rd_5r1[5:5], dt_0[5:5], rg_5r);
  AND2 I782 (rd_5r1[6:6], dt_0[6:6], rg_5r);
  AND2 I783 (rd_5r1[7:7], dt_0[7:7], rg_5r);
  AND2 I784 (rd_5r1[8:8], dt_0[8:8], rg_5r);
  AND2 I785 (rd_5r1[9:9], dt_0[9:9], rg_5r);
  AND2 I786 (rd_5r1[10:10], dt_0[10:10], rg_5r);
  AND2 I787 (rd_5r1[11:11], dt_0[11:11], rg_5r);
  AND2 I788 (rd_5r1[12:12], dt_0[12:12], rg_5r);
  AND2 I789 (rd_5r1[13:13], dt_0[13:13], rg_5r);
  AND2 I790 (rd_5r1[14:14], dt_0[14:14], rg_5r);
  AND2 I791 (rd_5r1[15:15], dt_0[15:15], rg_5r);
  AND2 I792 (rd_5r1[16:16], dt_0[16:16], rg_5r);
  AND2 I793 (rd_5r1[17:17], dt_0[17:17], rg_5r);
  AND2 I794 (rd_5r1[18:18], dt_0[18:18], rg_5r);
  AND2 I795 (rd_5r1[19:19], dt_0[19:19], rg_5r);
  AND2 I796 (rd_5r1[20:20], dt_0[20:20], rg_5r);
  AND2 I797 (rd_5r1[21:21], dt_0[21:21], rg_5r);
  AND2 I798 (rd_5r1[22:22], dt_0[22:22], rg_5r);
  AND2 I799 (rd_5r1[23:23], dt_0[23:23], rg_5r);
  AND2 I800 (rd_5r1[24:24], dt_0[24:24], rg_5r);
  AND2 I801 (rd_5r1[25:25], dt_0[25:25], rg_5r);
  AND2 I802 (rd_5r1[26:26], dt_0[26:26], rg_5r);
  AND2 I803 (rd_5r1[27:27], dt_0[27:27], rg_5r);
  AND2 I804 (rd_5r1[28:28], dt_0[28:28], rg_5r);
  AND2 I805 (rd_5r1[29:29], dt_0[29:29], rg_5r);
  AND2 I806 (rd_5r1[30:30], dt_0[30:30], rg_5r);
  AND2 I807 (rd_5r1[31:31], dt_0[31:31], rg_5r);
  NOR3 I808 (simp7921_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I809 (simp7921_0[1:1], rg_3r, rg_4r, rg_5r);
  NOR3 I810 (simp7921_0[2:2], rg_0a, rg_1a, rg_2a);
  NOR3 I811 (simp7921_0[3:3], rg_3a, rg_4a, rg_5a);
  NAND3 I812 (simp7922_0[0:0], simp7921_0[0:0], simp7921_0[1:1], simp7921_0[2:2]);
  INV I813 (simp7922_0[1:1], simp7921_0[3:3]);
  OR2 I814 (anyread_0, simp7922_0[0:0], simp7922_0[1:1]);
  BUFF I815 (wg_0a, wd_0a);
  BUFF I816 (rg_0a, rd_0a);
  BUFF I817 (rg_1a, rd_1a);
  BUFF I818 (rg_2a, rd_2a);
  BUFF I819 (rg_3a, rd_3a);
  BUFF I820 (rg_4a, rd_4a);
  BUFF I821 (rg_5a, rd_5a);
endmodule

// tkvinouts_633232_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 TeakV "inouts[63:32]" 32 [] [0] [0,0,0,0,0,0
//   ] [Many [32],Many [0],Many [0,0,0,0,0,0],Many [32,32,32,32,32,32]]
module tkvinouts_633232_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rg_5r, rg_5a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, rd_5r0, rd_5r1, rd_5a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  input rg_5r;
  output rg_5a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  output [31:0] rd_3r0;
  output [31:0] rd_3r1;
  input rd_3a;
  output [31:0] rd_4r0;
  output [31:0] rd_4r1;
  input rd_4a;
  output [31:0] rd_5r0;
  output [31:0] rd_5r1;
  input rd_5a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [3:0] simp7921_0;
  wire [1:0] simp7922_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_3r0[0:0], df_0[0:0], rg_3r);
  AND2 I521 (rd_3r0[1:1], df_0[1:1], rg_3r);
  AND2 I522 (rd_3r0[2:2], df_0[2:2], rg_3r);
  AND2 I523 (rd_3r0[3:3], df_0[3:3], rg_3r);
  AND2 I524 (rd_3r0[4:4], df_0[4:4], rg_3r);
  AND2 I525 (rd_3r0[5:5], df_0[5:5], rg_3r);
  AND2 I526 (rd_3r0[6:6], df_0[6:6], rg_3r);
  AND2 I527 (rd_3r0[7:7], df_0[7:7], rg_3r);
  AND2 I528 (rd_3r0[8:8], df_0[8:8], rg_3r);
  AND2 I529 (rd_3r0[9:9], df_0[9:9], rg_3r);
  AND2 I530 (rd_3r0[10:10], df_0[10:10], rg_3r);
  AND2 I531 (rd_3r0[11:11], df_0[11:11], rg_3r);
  AND2 I532 (rd_3r0[12:12], df_0[12:12], rg_3r);
  AND2 I533 (rd_3r0[13:13], df_0[13:13], rg_3r);
  AND2 I534 (rd_3r0[14:14], df_0[14:14], rg_3r);
  AND2 I535 (rd_3r0[15:15], df_0[15:15], rg_3r);
  AND2 I536 (rd_3r0[16:16], df_0[16:16], rg_3r);
  AND2 I537 (rd_3r0[17:17], df_0[17:17], rg_3r);
  AND2 I538 (rd_3r0[18:18], df_0[18:18], rg_3r);
  AND2 I539 (rd_3r0[19:19], df_0[19:19], rg_3r);
  AND2 I540 (rd_3r0[20:20], df_0[20:20], rg_3r);
  AND2 I541 (rd_3r0[21:21], df_0[21:21], rg_3r);
  AND2 I542 (rd_3r0[22:22], df_0[22:22], rg_3r);
  AND2 I543 (rd_3r0[23:23], df_0[23:23], rg_3r);
  AND2 I544 (rd_3r0[24:24], df_0[24:24], rg_3r);
  AND2 I545 (rd_3r0[25:25], df_0[25:25], rg_3r);
  AND2 I546 (rd_3r0[26:26], df_0[26:26], rg_3r);
  AND2 I547 (rd_3r0[27:27], df_0[27:27], rg_3r);
  AND2 I548 (rd_3r0[28:28], df_0[28:28], rg_3r);
  AND2 I549 (rd_3r0[29:29], df_0[29:29], rg_3r);
  AND2 I550 (rd_3r0[30:30], df_0[30:30], rg_3r);
  AND2 I551 (rd_3r0[31:31], df_0[31:31], rg_3r);
  AND2 I552 (rd_4r0[0:0], df_0[0:0], rg_4r);
  AND2 I553 (rd_4r0[1:1], df_0[1:1], rg_4r);
  AND2 I554 (rd_4r0[2:2], df_0[2:2], rg_4r);
  AND2 I555 (rd_4r0[3:3], df_0[3:3], rg_4r);
  AND2 I556 (rd_4r0[4:4], df_0[4:4], rg_4r);
  AND2 I557 (rd_4r0[5:5], df_0[5:5], rg_4r);
  AND2 I558 (rd_4r0[6:6], df_0[6:6], rg_4r);
  AND2 I559 (rd_4r0[7:7], df_0[7:7], rg_4r);
  AND2 I560 (rd_4r0[8:8], df_0[8:8], rg_4r);
  AND2 I561 (rd_4r0[9:9], df_0[9:9], rg_4r);
  AND2 I562 (rd_4r0[10:10], df_0[10:10], rg_4r);
  AND2 I563 (rd_4r0[11:11], df_0[11:11], rg_4r);
  AND2 I564 (rd_4r0[12:12], df_0[12:12], rg_4r);
  AND2 I565 (rd_4r0[13:13], df_0[13:13], rg_4r);
  AND2 I566 (rd_4r0[14:14], df_0[14:14], rg_4r);
  AND2 I567 (rd_4r0[15:15], df_0[15:15], rg_4r);
  AND2 I568 (rd_4r0[16:16], df_0[16:16], rg_4r);
  AND2 I569 (rd_4r0[17:17], df_0[17:17], rg_4r);
  AND2 I570 (rd_4r0[18:18], df_0[18:18], rg_4r);
  AND2 I571 (rd_4r0[19:19], df_0[19:19], rg_4r);
  AND2 I572 (rd_4r0[20:20], df_0[20:20], rg_4r);
  AND2 I573 (rd_4r0[21:21], df_0[21:21], rg_4r);
  AND2 I574 (rd_4r0[22:22], df_0[22:22], rg_4r);
  AND2 I575 (rd_4r0[23:23], df_0[23:23], rg_4r);
  AND2 I576 (rd_4r0[24:24], df_0[24:24], rg_4r);
  AND2 I577 (rd_4r0[25:25], df_0[25:25], rg_4r);
  AND2 I578 (rd_4r0[26:26], df_0[26:26], rg_4r);
  AND2 I579 (rd_4r0[27:27], df_0[27:27], rg_4r);
  AND2 I580 (rd_4r0[28:28], df_0[28:28], rg_4r);
  AND2 I581 (rd_4r0[29:29], df_0[29:29], rg_4r);
  AND2 I582 (rd_4r0[30:30], df_0[30:30], rg_4r);
  AND2 I583 (rd_4r0[31:31], df_0[31:31], rg_4r);
  AND2 I584 (rd_5r0[0:0], df_0[0:0], rg_5r);
  AND2 I585 (rd_5r0[1:1], df_0[1:1], rg_5r);
  AND2 I586 (rd_5r0[2:2], df_0[2:2], rg_5r);
  AND2 I587 (rd_5r0[3:3], df_0[3:3], rg_5r);
  AND2 I588 (rd_5r0[4:4], df_0[4:4], rg_5r);
  AND2 I589 (rd_5r0[5:5], df_0[5:5], rg_5r);
  AND2 I590 (rd_5r0[6:6], df_0[6:6], rg_5r);
  AND2 I591 (rd_5r0[7:7], df_0[7:7], rg_5r);
  AND2 I592 (rd_5r0[8:8], df_0[8:8], rg_5r);
  AND2 I593 (rd_5r0[9:9], df_0[9:9], rg_5r);
  AND2 I594 (rd_5r0[10:10], df_0[10:10], rg_5r);
  AND2 I595 (rd_5r0[11:11], df_0[11:11], rg_5r);
  AND2 I596 (rd_5r0[12:12], df_0[12:12], rg_5r);
  AND2 I597 (rd_5r0[13:13], df_0[13:13], rg_5r);
  AND2 I598 (rd_5r0[14:14], df_0[14:14], rg_5r);
  AND2 I599 (rd_5r0[15:15], df_0[15:15], rg_5r);
  AND2 I600 (rd_5r0[16:16], df_0[16:16], rg_5r);
  AND2 I601 (rd_5r0[17:17], df_0[17:17], rg_5r);
  AND2 I602 (rd_5r0[18:18], df_0[18:18], rg_5r);
  AND2 I603 (rd_5r0[19:19], df_0[19:19], rg_5r);
  AND2 I604 (rd_5r0[20:20], df_0[20:20], rg_5r);
  AND2 I605 (rd_5r0[21:21], df_0[21:21], rg_5r);
  AND2 I606 (rd_5r0[22:22], df_0[22:22], rg_5r);
  AND2 I607 (rd_5r0[23:23], df_0[23:23], rg_5r);
  AND2 I608 (rd_5r0[24:24], df_0[24:24], rg_5r);
  AND2 I609 (rd_5r0[25:25], df_0[25:25], rg_5r);
  AND2 I610 (rd_5r0[26:26], df_0[26:26], rg_5r);
  AND2 I611 (rd_5r0[27:27], df_0[27:27], rg_5r);
  AND2 I612 (rd_5r0[28:28], df_0[28:28], rg_5r);
  AND2 I613 (rd_5r0[29:29], df_0[29:29], rg_5r);
  AND2 I614 (rd_5r0[30:30], df_0[30:30], rg_5r);
  AND2 I615 (rd_5r0[31:31], df_0[31:31], rg_5r);
  AND2 I616 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I617 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I618 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I619 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I620 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I621 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I622 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I623 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I624 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I625 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I626 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I627 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I628 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I629 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I630 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I631 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I632 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I633 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I634 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I635 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I636 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I637 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I638 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I639 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I640 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I641 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I642 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I643 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I644 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I645 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I646 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I647 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I648 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I649 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I650 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I651 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I652 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I653 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I654 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I655 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I656 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I657 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I658 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I659 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I660 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I661 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I662 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I663 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I664 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I665 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I666 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I667 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I668 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I669 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I670 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I671 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I672 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I673 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I674 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I675 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I676 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I677 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I678 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I679 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I680 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I681 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I682 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I683 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I684 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I685 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I686 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I687 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I688 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I689 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I690 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I691 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I692 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I693 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I694 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I695 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I696 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I697 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I698 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I699 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I700 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I701 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I702 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I703 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I704 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I705 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I706 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I707 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I708 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I709 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I710 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I711 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  AND2 I712 (rd_3r1[0:0], dt_0[0:0], rg_3r);
  AND2 I713 (rd_3r1[1:1], dt_0[1:1], rg_3r);
  AND2 I714 (rd_3r1[2:2], dt_0[2:2], rg_3r);
  AND2 I715 (rd_3r1[3:3], dt_0[3:3], rg_3r);
  AND2 I716 (rd_3r1[4:4], dt_0[4:4], rg_3r);
  AND2 I717 (rd_3r1[5:5], dt_0[5:5], rg_3r);
  AND2 I718 (rd_3r1[6:6], dt_0[6:6], rg_3r);
  AND2 I719 (rd_3r1[7:7], dt_0[7:7], rg_3r);
  AND2 I720 (rd_3r1[8:8], dt_0[8:8], rg_3r);
  AND2 I721 (rd_3r1[9:9], dt_0[9:9], rg_3r);
  AND2 I722 (rd_3r1[10:10], dt_0[10:10], rg_3r);
  AND2 I723 (rd_3r1[11:11], dt_0[11:11], rg_3r);
  AND2 I724 (rd_3r1[12:12], dt_0[12:12], rg_3r);
  AND2 I725 (rd_3r1[13:13], dt_0[13:13], rg_3r);
  AND2 I726 (rd_3r1[14:14], dt_0[14:14], rg_3r);
  AND2 I727 (rd_3r1[15:15], dt_0[15:15], rg_3r);
  AND2 I728 (rd_3r1[16:16], dt_0[16:16], rg_3r);
  AND2 I729 (rd_3r1[17:17], dt_0[17:17], rg_3r);
  AND2 I730 (rd_3r1[18:18], dt_0[18:18], rg_3r);
  AND2 I731 (rd_3r1[19:19], dt_0[19:19], rg_3r);
  AND2 I732 (rd_3r1[20:20], dt_0[20:20], rg_3r);
  AND2 I733 (rd_3r1[21:21], dt_0[21:21], rg_3r);
  AND2 I734 (rd_3r1[22:22], dt_0[22:22], rg_3r);
  AND2 I735 (rd_3r1[23:23], dt_0[23:23], rg_3r);
  AND2 I736 (rd_3r1[24:24], dt_0[24:24], rg_3r);
  AND2 I737 (rd_3r1[25:25], dt_0[25:25], rg_3r);
  AND2 I738 (rd_3r1[26:26], dt_0[26:26], rg_3r);
  AND2 I739 (rd_3r1[27:27], dt_0[27:27], rg_3r);
  AND2 I740 (rd_3r1[28:28], dt_0[28:28], rg_3r);
  AND2 I741 (rd_3r1[29:29], dt_0[29:29], rg_3r);
  AND2 I742 (rd_3r1[30:30], dt_0[30:30], rg_3r);
  AND2 I743 (rd_3r1[31:31], dt_0[31:31], rg_3r);
  AND2 I744 (rd_4r1[0:0], dt_0[0:0], rg_4r);
  AND2 I745 (rd_4r1[1:1], dt_0[1:1], rg_4r);
  AND2 I746 (rd_4r1[2:2], dt_0[2:2], rg_4r);
  AND2 I747 (rd_4r1[3:3], dt_0[3:3], rg_4r);
  AND2 I748 (rd_4r1[4:4], dt_0[4:4], rg_4r);
  AND2 I749 (rd_4r1[5:5], dt_0[5:5], rg_4r);
  AND2 I750 (rd_4r1[6:6], dt_0[6:6], rg_4r);
  AND2 I751 (rd_4r1[7:7], dt_0[7:7], rg_4r);
  AND2 I752 (rd_4r1[8:8], dt_0[8:8], rg_4r);
  AND2 I753 (rd_4r1[9:9], dt_0[9:9], rg_4r);
  AND2 I754 (rd_4r1[10:10], dt_0[10:10], rg_4r);
  AND2 I755 (rd_4r1[11:11], dt_0[11:11], rg_4r);
  AND2 I756 (rd_4r1[12:12], dt_0[12:12], rg_4r);
  AND2 I757 (rd_4r1[13:13], dt_0[13:13], rg_4r);
  AND2 I758 (rd_4r1[14:14], dt_0[14:14], rg_4r);
  AND2 I759 (rd_4r1[15:15], dt_0[15:15], rg_4r);
  AND2 I760 (rd_4r1[16:16], dt_0[16:16], rg_4r);
  AND2 I761 (rd_4r1[17:17], dt_0[17:17], rg_4r);
  AND2 I762 (rd_4r1[18:18], dt_0[18:18], rg_4r);
  AND2 I763 (rd_4r1[19:19], dt_0[19:19], rg_4r);
  AND2 I764 (rd_4r1[20:20], dt_0[20:20], rg_4r);
  AND2 I765 (rd_4r1[21:21], dt_0[21:21], rg_4r);
  AND2 I766 (rd_4r1[22:22], dt_0[22:22], rg_4r);
  AND2 I767 (rd_4r1[23:23], dt_0[23:23], rg_4r);
  AND2 I768 (rd_4r1[24:24], dt_0[24:24], rg_4r);
  AND2 I769 (rd_4r1[25:25], dt_0[25:25], rg_4r);
  AND2 I770 (rd_4r1[26:26], dt_0[26:26], rg_4r);
  AND2 I771 (rd_4r1[27:27], dt_0[27:27], rg_4r);
  AND2 I772 (rd_4r1[28:28], dt_0[28:28], rg_4r);
  AND2 I773 (rd_4r1[29:29], dt_0[29:29], rg_4r);
  AND2 I774 (rd_4r1[30:30], dt_0[30:30], rg_4r);
  AND2 I775 (rd_4r1[31:31], dt_0[31:31], rg_4r);
  AND2 I776 (rd_5r1[0:0], dt_0[0:0], rg_5r);
  AND2 I777 (rd_5r1[1:1], dt_0[1:1], rg_5r);
  AND2 I778 (rd_5r1[2:2], dt_0[2:2], rg_5r);
  AND2 I779 (rd_5r1[3:3], dt_0[3:3], rg_5r);
  AND2 I780 (rd_5r1[4:4], dt_0[4:4], rg_5r);
  AND2 I781 (rd_5r1[5:5], dt_0[5:5], rg_5r);
  AND2 I782 (rd_5r1[6:6], dt_0[6:6], rg_5r);
  AND2 I783 (rd_5r1[7:7], dt_0[7:7], rg_5r);
  AND2 I784 (rd_5r1[8:8], dt_0[8:8], rg_5r);
  AND2 I785 (rd_5r1[9:9], dt_0[9:9], rg_5r);
  AND2 I786 (rd_5r1[10:10], dt_0[10:10], rg_5r);
  AND2 I787 (rd_5r1[11:11], dt_0[11:11], rg_5r);
  AND2 I788 (rd_5r1[12:12], dt_0[12:12], rg_5r);
  AND2 I789 (rd_5r1[13:13], dt_0[13:13], rg_5r);
  AND2 I790 (rd_5r1[14:14], dt_0[14:14], rg_5r);
  AND2 I791 (rd_5r1[15:15], dt_0[15:15], rg_5r);
  AND2 I792 (rd_5r1[16:16], dt_0[16:16], rg_5r);
  AND2 I793 (rd_5r1[17:17], dt_0[17:17], rg_5r);
  AND2 I794 (rd_5r1[18:18], dt_0[18:18], rg_5r);
  AND2 I795 (rd_5r1[19:19], dt_0[19:19], rg_5r);
  AND2 I796 (rd_5r1[20:20], dt_0[20:20], rg_5r);
  AND2 I797 (rd_5r1[21:21], dt_0[21:21], rg_5r);
  AND2 I798 (rd_5r1[22:22], dt_0[22:22], rg_5r);
  AND2 I799 (rd_5r1[23:23], dt_0[23:23], rg_5r);
  AND2 I800 (rd_5r1[24:24], dt_0[24:24], rg_5r);
  AND2 I801 (rd_5r1[25:25], dt_0[25:25], rg_5r);
  AND2 I802 (rd_5r1[26:26], dt_0[26:26], rg_5r);
  AND2 I803 (rd_5r1[27:27], dt_0[27:27], rg_5r);
  AND2 I804 (rd_5r1[28:28], dt_0[28:28], rg_5r);
  AND2 I805 (rd_5r1[29:29], dt_0[29:29], rg_5r);
  AND2 I806 (rd_5r1[30:30], dt_0[30:30], rg_5r);
  AND2 I807 (rd_5r1[31:31], dt_0[31:31], rg_5r);
  NOR3 I808 (simp7921_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I809 (simp7921_0[1:1], rg_3r, rg_4r, rg_5r);
  NOR3 I810 (simp7921_0[2:2], rg_0a, rg_1a, rg_2a);
  NOR3 I811 (simp7921_0[3:3], rg_3a, rg_4a, rg_5a);
  NAND3 I812 (simp7922_0[0:0], simp7921_0[0:0], simp7921_0[1:1], simp7921_0[2:2]);
  INV I813 (simp7922_0[1:1], simp7921_0[3:3]);
  OR2 I814 (anyread_0, simp7922_0[0:0], simp7922_0[1:1]);
  BUFF I815 (wg_0a, wd_0a);
  BUFF I816 (rg_0a, rd_0a);
  BUFF I817 (rg_1a, rd_1a);
  BUFF I818 (rg_2a, rd_2a);
  BUFF I819 (rg_3a, rd_3a);
  BUFF I820 (rg_4a, rd_4a);
  BUFF I821 (rg_5a, rd_5a);
endmodule

// tkvinouts_956432_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 TeakV "inouts[95:64]" 32 [] [0] [0,0,0,0,0,0
//   ] [Many [32],Many [0],Many [0,0,0,0,0,0],Many [32,32,32,32,32,32]]
module tkvinouts_956432_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rg_5r, rg_5a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, rd_5r0, rd_5r1, rd_5a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  input rg_5r;
  output rg_5a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  output [31:0] rd_3r0;
  output [31:0] rd_3r1;
  input rd_3a;
  output [31:0] rd_4r0;
  output [31:0] rd_4r1;
  input rd_4a;
  output [31:0] rd_5r0;
  output [31:0] rd_5r1;
  input rd_5a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [3:0] simp7921_0;
  wire [1:0] simp7922_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_3r0[0:0], df_0[0:0], rg_3r);
  AND2 I521 (rd_3r0[1:1], df_0[1:1], rg_3r);
  AND2 I522 (rd_3r0[2:2], df_0[2:2], rg_3r);
  AND2 I523 (rd_3r0[3:3], df_0[3:3], rg_3r);
  AND2 I524 (rd_3r0[4:4], df_0[4:4], rg_3r);
  AND2 I525 (rd_3r0[5:5], df_0[5:5], rg_3r);
  AND2 I526 (rd_3r0[6:6], df_0[6:6], rg_3r);
  AND2 I527 (rd_3r0[7:7], df_0[7:7], rg_3r);
  AND2 I528 (rd_3r0[8:8], df_0[8:8], rg_3r);
  AND2 I529 (rd_3r0[9:9], df_0[9:9], rg_3r);
  AND2 I530 (rd_3r0[10:10], df_0[10:10], rg_3r);
  AND2 I531 (rd_3r0[11:11], df_0[11:11], rg_3r);
  AND2 I532 (rd_3r0[12:12], df_0[12:12], rg_3r);
  AND2 I533 (rd_3r0[13:13], df_0[13:13], rg_3r);
  AND2 I534 (rd_3r0[14:14], df_0[14:14], rg_3r);
  AND2 I535 (rd_3r0[15:15], df_0[15:15], rg_3r);
  AND2 I536 (rd_3r0[16:16], df_0[16:16], rg_3r);
  AND2 I537 (rd_3r0[17:17], df_0[17:17], rg_3r);
  AND2 I538 (rd_3r0[18:18], df_0[18:18], rg_3r);
  AND2 I539 (rd_3r0[19:19], df_0[19:19], rg_3r);
  AND2 I540 (rd_3r0[20:20], df_0[20:20], rg_3r);
  AND2 I541 (rd_3r0[21:21], df_0[21:21], rg_3r);
  AND2 I542 (rd_3r0[22:22], df_0[22:22], rg_3r);
  AND2 I543 (rd_3r0[23:23], df_0[23:23], rg_3r);
  AND2 I544 (rd_3r0[24:24], df_0[24:24], rg_3r);
  AND2 I545 (rd_3r0[25:25], df_0[25:25], rg_3r);
  AND2 I546 (rd_3r0[26:26], df_0[26:26], rg_3r);
  AND2 I547 (rd_3r0[27:27], df_0[27:27], rg_3r);
  AND2 I548 (rd_3r0[28:28], df_0[28:28], rg_3r);
  AND2 I549 (rd_3r0[29:29], df_0[29:29], rg_3r);
  AND2 I550 (rd_3r0[30:30], df_0[30:30], rg_3r);
  AND2 I551 (rd_3r0[31:31], df_0[31:31], rg_3r);
  AND2 I552 (rd_4r0[0:0], df_0[0:0], rg_4r);
  AND2 I553 (rd_4r0[1:1], df_0[1:1], rg_4r);
  AND2 I554 (rd_4r0[2:2], df_0[2:2], rg_4r);
  AND2 I555 (rd_4r0[3:3], df_0[3:3], rg_4r);
  AND2 I556 (rd_4r0[4:4], df_0[4:4], rg_4r);
  AND2 I557 (rd_4r0[5:5], df_0[5:5], rg_4r);
  AND2 I558 (rd_4r0[6:6], df_0[6:6], rg_4r);
  AND2 I559 (rd_4r0[7:7], df_0[7:7], rg_4r);
  AND2 I560 (rd_4r0[8:8], df_0[8:8], rg_4r);
  AND2 I561 (rd_4r0[9:9], df_0[9:9], rg_4r);
  AND2 I562 (rd_4r0[10:10], df_0[10:10], rg_4r);
  AND2 I563 (rd_4r0[11:11], df_0[11:11], rg_4r);
  AND2 I564 (rd_4r0[12:12], df_0[12:12], rg_4r);
  AND2 I565 (rd_4r0[13:13], df_0[13:13], rg_4r);
  AND2 I566 (rd_4r0[14:14], df_0[14:14], rg_4r);
  AND2 I567 (rd_4r0[15:15], df_0[15:15], rg_4r);
  AND2 I568 (rd_4r0[16:16], df_0[16:16], rg_4r);
  AND2 I569 (rd_4r0[17:17], df_0[17:17], rg_4r);
  AND2 I570 (rd_4r0[18:18], df_0[18:18], rg_4r);
  AND2 I571 (rd_4r0[19:19], df_0[19:19], rg_4r);
  AND2 I572 (rd_4r0[20:20], df_0[20:20], rg_4r);
  AND2 I573 (rd_4r0[21:21], df_0[21:21], rg_4r);
  AND2 I574 (rd_4r0[22:22], df_0[22:22], rg_4r);
  AND2 I575 (rd_4r0[23:23], df_0[23:23], rg_4r);
  AND2 I576 (rd_4r0[24:24], df_0[24:24], rg_4r);
  AND2 I577 (rd_4r0[25:25], df_0[25:25], rg_4r);
  AND2 I578 (rd_4r0[26:26], df_0[26:26], rg_4r);
  AND2 I579 (rd_4r0[27:27], df_0[27:27], rg_4r);
  AND2 I580 (rd_4r0[28:28], df_0[28:28], rg_4r);
  AND2 I581 (rd_4r0[29:29], df_0[29:29], rg_4r);
  AND2 I582 (rd_4r0[30:30], df_0[30:30], rg_4r);
  AND2 I583 (rd_4r0[31:31], df_0[31:31], rg_4r);
  AND2 I584 (rd_5r0[0:0], df_0[0:0], rg_5r);
  AND2 I585 (rd_5r0[1:1], df_0[1:1], rg_5r);
  AND2 I586 (rd_5r0[2:2], df_0[2:2], rg_5r);
  AND2 I587 (rd_5r0[3:3], df_0[3:3], rg_5r);
  AND2 I588 (rd_5r0[4:4], df_0[4:4], rg_5r);
  AND2 I589 (rd_5r0[5:5], df_0[5:5], rg_5r);
  AND2 I590 (rd_5r0[6:6], df_0[6:6], rg_5r);
  AND2 I591 (rd_5r0[7:7], df_0[7:7], rg_5r);
  AND2 I592 (rd_5r0[8:8], df_0[8:8], rg_5r);
  AND2 I593 (rd_5r0[9:9], df_0[9:9], rg_5r);
  AND2 I594 (rd_5r0[10:10], df_0[10:10], rg_5r);
  AND2 I595 (rd_5r0[11:11], df_0[11:11], rg_5r);
  AND2 I596 (rd_5r0[12:12], df_0[12:12], rg_5r);
  AND2 I597 (rd_5r0[13:13], df_0[13:13], rg_5r);
  AND2 I598 (rd_5r0[14:14], df_0[14:14], rg_5r);
  AND2 I599 (rd_5r0[15:15], df_0[15:15], rg_5r);
  AND2 I600 (rd_5r0[16:16], df_0[16:16], rg_5r);
  AND2 I601 (rd_5r0[17:17], df_0[17:17], rg_5r);
  AND2 I602 (rd_5r0[18:18], df_0[18:18], rg_5r);
  AND2 I603 (rd_5r0[19:19], df_0[19:19], rg_5r);
  AND2 I604 (rd_5r0[20:20], df_0[20:20], rg_5r);
  AND2 I605 (rd_5r0[21:21], df_0[21:21], rg_5r);
  AND2 I606 (rd_5r0[22:22], df_0[22:22], rg_5r);
  AND2 I607 (rd_5r0[23:23], df_0[23:23], rg_5r);
  AND2 I608 (rd_5r0[24:24], df_0[24:24], rg_5r);
  AND2 I609 (rd_5r0[25:25], df_0[25:25], rg_5r);
  AND2 I610 (rd_5r0[26:26], df_0[26:26], rg_5r);
  AND2 I611 (rd_5r0[27:27], df_0[27:27], rg_5r);
  AND2 I612 (rd_5r0[28:28], df_0[28:28], rg_5r);
  AND2 I613 (rd_5r0[29:29], df_0[29:29], rg_5r);
  AND2 I614 (rd_5r0[30:30], df_0[30:30], rg_5r);
  AND2 I615 (rd_5r0[31:31], df_0[31:31], rg_5r);
  AND2 I616 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I617 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I618 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I619 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I620 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I621 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I622 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I623 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I624 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I625 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I626 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I627 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I628 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I629 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I630 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I631 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I632 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I633 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I634 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I635 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I636 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I637 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I638 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I639 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I640 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I641 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I642 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I643 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I644 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I645 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I646 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I647 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I648 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I649 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I650 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I651 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I652 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I653 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I654 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I655 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I656 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I657 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I658 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I659 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I660 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I661 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I662 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I663 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I664 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I665 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I666 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I667 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I668 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I669 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I670 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I671 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I672 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I673 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I674 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I675 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I676 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I677 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I678 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I679 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I680 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I681 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I682 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I683 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I684 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I685 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I686 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I687 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I688 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I689 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I690 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I691 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I692 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I693 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I694 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I695 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I696 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I697 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I698 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I699 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I700 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I701 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I702 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I703 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I704 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I705 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I706 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I707 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I708 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I709 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I710 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I711 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  AND2 I712 (rd_3r1[0:0], dt_0[0:0], rg_3r);
  AND2 I713 (rd_3r1[1:1], dt_0[1:1], rg_3r);
  AND2 I714 (rd_3r1[2:2], dt_0[2:2], rg_3r);
  AND2 I715 (rd_3r1[3:3], dt_0[3:3], rg_3r);
  AND2 I716 (rd_3r1[4:4], dt_0[4:4], rg_3r);
  AND2 I717 (rd_3r1[5:5], dt_0[5:5], rg_3r);
  AND2 I718 (rd_3r1[6:6], dt_0[6:6], rg_3r);
  AND2 I719 (rd_3r1[7:7], dt_0[7:7], rg_3r);
  AND2 I720 (rd_3r1[8:8], dt_0[8:8], rg_3r);
  AND2 I721 (rd_3r1[9:9], dt_0[9:9], rg_3r);
  AND2 I722 (rd_3r1[10:10], dt_0[10:10], rg_3r);
  AND2 I723 (rd_3r1[11:11], dt_0[11:11], rg_3r);
  AND2 I724 (rd_3r1[12:12], dt_0[12:12], rg_3r);
  AND2 I725 (rd_3r1[13:13], dt_0[13:13], rg_3r);
  AND2 I726 (rd_3r1[14:14], dt_0[14:14], rg_3r);
  AND2 I727 (rd_3r1[15:15], dt_0[15:15], rg_3r);
  AND2 I728 (rd_3r1[16:16], dt_0[16:16], rg_3r);
  AND2 I729 (rd_3r1[17:17], dt_0[17:17], rg_3r);
  AND2 I730 (rd_3r1[18:18], dt_0[18:18], rg_3r);
  AND2 I731 (rd_3r1[19:19], dt_0[19:19], rg_3r);
  AND2 I732 (rd_3r1[20:20], dt_0[20:20], rg_3r);
  AND2 I733 (rd_3r1[21:21], dt_0[21:21], rg_3r);
  AND2 I734 (rd_3r1[22:22], dt_0[22:22], rg_3r);
  AND2 I735 (rd_3r1[23:23], dt_0[23:23], rg_3r);
  AND2 I736 (rd_3r1[24:24], dt_0[24:24], rg_3r);
  AND2 I737 (rd_3r1[25:25], dt_0[25:25], rg_3r);
  AND2 I738 (rd_3r1[26:26], dt_0[26:26], rg_3r);
  AND2 I739 (rd_3r1[27:27], dt_0[27:27], rg_3r);
  AND2 I740 (rd_3r1[28:28], dt_0[28:28], rg_3r);
  AND2 I741 (rd_3r1[29:29], dt_0[29:29], rg_3r);
  AND2 I742 (rd_3r1[30:30], dt_0[30:30], rg_3r);
  AND2 I743 (rd_3r1[31:31], dt_0[31:31], rg_3r);
  AND2 I744 (rd_4r1[0:0], dt_0[0:0], rg_4r);
  AND2 I745 (rd_4r1[1:1], dt_0[1:1], rg_4r);
  AND2 I746 (rd_4r1[2:2], dt_0[2:2], rg_4r);
  AND2 I747 (rd_4r1[3:3], dt_0[3:3], rg_4r);
  AND2 I748 (rd_4r1[4:4], dt_0[4:4], rg_4r);
  AND2 I749 (rd_4r1[5:5], dt_0[5:5], rg_4r);
  AND2 I750 (rd_4r1[6:6], dt_0[6:6], rg_4r);
  AND2 I751 (rd_4r1[7:7], dt_0[7:7], rg_4r);
  AND2 I752 (rd_4r1[8:8], dt_0[8:8], rg_4r);
  AND2 I753 (rd_4r1[9:9], dt_0[9:9], rg_4r);
  AND2 I754 (rd_4r1[10:10], dt_0[10:10], rg_4r);
  AND2 I755 (rd_4r1[11:11], dt_0[11:11], rg_4r);
  AND2 I756 (rd_4r1[12:12], dt_0[12:12], rg_4r);
  AND2 I757 (rd_4r1[13:13], dt_0[13:13], rg_4r);
  AND2 I758 (rd_4r1[14:14], dt_0[14:14], rg_4r);
  AND2 I759 (rd_4r1[15:15], dt_0[15:15], rg_4r);
  AND2 I760 (rd_4r1[16:16], dt_0[16:16], rg_4r);
  AND2 I761 (rd_4r1[17:17], dt_0[17:17], rg_4r);
  AND2 I762 (rd_4r1[18:18], dt_0[18:18], rg_4r);
  AND2 I763 (rd_4r1[19:19], dt_0[19:19], rg_4r);
  AND2 I764 (rd_4r1[20:20], dt_0[20:20], rg_4r);
  AND2 I765 (rd_4r1[21:21], dt_0[21:21], rg_4r);
  AND2 I766 (rd_4r1[22:22], dt_0[22:22], rg_4r);
  AND2 I767 (rd_4r1[23:23], dt_0[23:23], rg_4r);
  AND2 I768 (rd_4r1[24:24], dt_0[24:24], rg_4r);
  AND2 I769 (rd_4r1[25:25], dt_0[25:25], rg_4r);
  AND2 I770 (rd_4r1[26:26], dt_0[26:26], rg_4r);
  AND2 I771 (rd_4r1[27:27], dt_0[27:27], rg_4r);
  AND2 I772 (rd_4r1[28:28], dt_0[28:28], rg_4r);
  AND2 I773 (rd_4r1[29:29], dt_0[29:29], rg_4r);
  AND2 I774 (rd_4r1[30:30], dt_0[30:30], rg_4r);
  AND2 I775 (rd_4r1[31:31], dt_0[31:31], rg_4r);
  AND2 I776 (rd_5r1[0:0], dt_0[0:0], rg_5r);
  AND2 I777 (rd_5r1[1:1], dt_0[1:1], rg_5r);
  AND2 I778 (rd_5r1[2:2], dt_0[2:2], rg_5r);
  AND2 I779 (rd_5r1[3:3], dt_0[3:3], rg_5r);
  AND2 I780 (rd_5r1[4:4], dt_0[4:4], rg_5r);
  AND2 I781 (rd_5r1[5:5], dt_0[5:5], rg_5r);
  AND2 I782 (rd_5r1[6:6], dt_0[6:6], rg_5r);
  AND2 I783 (rd_5r1[7:7], dt_0[7:7], rg_5r);
  AND2 I784 (rd_5r1[8:8], dt_0[8:8], rg_5r);
  AND2 I785 (rd_5r1[9:9], dt_0[9:9], rg_5r);
  AND2 I786 (rd_5r1[10:10], dt_0[10:10], rg_5r);
  AND2 I787 (rd_5r1[11:11], dt_0[11:11], rg_5r);
  AND2 I788 (rd_5r1[12:12], dt_0[12:12], rg_5r);
  AND2 I789 (rd_5r1[13:13], dt_0[13:13], rg_5r);
  AND2 I790 (rd_5r1[14:14], dt_0[14:14], rg_5r);
  AND2 I791 (rd_5r1[15:15], dt_0[15:15], rg_5r);
  AND2 I792 (rd_5r1[16:16], dt_0[16:16], rg_5r);
  AND2 I793 (rd_5r1[17:17], dt_0[17:17], rg_5r);
  AND2 I794 (rd_5r1[18:18], dt_0[18:18], rg_5r);
  AND2 I795 (rd_5r1[19:19], dt_0[19:19], rg_5r);
  AND2 I796 (rd_5r1[20:20], dt_0[20:20], rg_5r);
  AND2 I797 (rd_5r1[21:21], dt_0[21:21], rg_5r);
  AND2 I798 (rd_5r1[22:22], dt_0[22:22], rg_5r);
  AND2 I799 (rd_5r1[23:23], dt_0[23:23], rg_5r);
  AND2 I800 (rd_5r1[24:24], dt_0[24:24], rg_5r);
  AND2 I801 (rd_5r1[25:25], dt_0[25:25], rg_5r);
  AND2 I802 (rd_5r1[26:26], dt_0[26:26], rg_5r);
  AND2 I803 (rd_5r1[27:27], dt_0[27:27], rg_5r);
  AND2 I804 (rd_5r1[28:28], dt_0[28:28], rg_5r);
  AND2 I805 (rd_5r1[29:29], dt_0[29:29], rg_5r);
  AND2 I806 (rd_5r1[30:30], dt_0[30:30], rg_5r);
  AND2 I807 (rd_5r1[31:31], dt_0[31:31], rg_5r);
  NOR3 I808 (simp7921_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I809 (simp7921_0[1:1], rg_3r, rg_4r, rg_5r);
  NOR3 I810 (simp7921_0[2:2], rg_0a, rg_1a, rg_2a);
  NOR3 I811 (simp7921_0[3:3], rg_3a, rg_4a, rg_5a);
  NAND3 I812 (simp7922_0[0:0], simp7921_0[0:0], simp7921_0[1:1], simp7921_0[2:2]);
  INV I813 (simp7922_0[1:1], simp7921_0[3:3]);
  OR2 I814 (anyread_0, simp7922_0[0:0], simp7922_0[1:1]);
  BUFF I815 (wg_0a, wd_0a);
  BUFF I816 (rg_0a, rd_0a);
  BUFF I817 (rg_1a, rd_1a);
  BUFF I818 (rg_2a, rd_2a);
  BUFF I819 (rg_3a, rd_3a);
  BUFF I820 (rg_4a, rd_4a);
  BUFF I821 (rg_5a, rd_5a);
endmodule

// tkvinouts_1279632_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 TeakV "inouts[127:96]" 32 [] [0] [0,0,0,0,0
//   ,0] [Many [32],Many [0],Many [0,0,0,0,0,0],Many [32,32,32,32,32,32]]
module tkvinouts_1279632_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rg_5r, rg_5a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, rd_5r0, rd_5r1, rd_5a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  input rg_5r;
  output rg_5a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  output [31:0] rd_3r0;
  output [31:0] rd_3r1;
  input rd_3a;
  output [31:0] rd_4r0;
  output [31:0] rd_4r1;
  input rd_4a;
  output [31:0] rd_5r0;
  output [31:0] rd_5r1;
  input rd_5a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [3:0] simp7921_0;
  wire [1:0] simp7922_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_3r0[0:0], df_0[0:0], rg_3r);
  AND2 I521 (rd_3r0[1:1], df_0[1:1], rg_3r);
  AND2 I522 (rd_3r0[2:2], df_0[2:2], rg_3r);
  AND2 I523 (rd_3r0[3:3], df_0[3:3], rg_3r);
  AND2 I524 (rd_3r0[4:4], df_0[4:4], rg_3r);
  AND2 I525 (rd_3r0[5:5], df_0[5:5], rg_3r);
  AND2 I526 (rd_3r0[6:6], df_0[6:6], rg_3r);
  AND2 I527 (rd_3r0[7:7], df_0[7:7], rg_3r);
  AND2 I528 (rd_3r0[8:8], df_0[8:8], rg_3r);
  AND2 I529 (rd_3r0[9:9], df_0[9:9], rg_3r);
  AND2 I530 (rd_3r0[10:10], df_0[10:10], rg_3r);
  AND2 I531 (rd_3r0[11:11], df_0[11:11], rg_3r);
  AND2 I532 (rd_3r0[12:12], df_0[12:12], rg_3r);
  AND2 I533 (rd_3r0[13:13], df_0[13:13], rg_3r);
  AND2 I534 (rd_3r0[14:14], df_0[14:14], rg_3r);
  AND2 I535 (rd_3r0[15:15], df_0[15:15], rg_3r);
  AND2 I536 (rd_3r0[16:16], df_0[16:16], rg_3r);
  AND2 I537 (rd_3r0[17:17], df_0[17:17], rg_3r);
  AND2 I538 (rd_3r0[18:18], df_0[18:18], rg_3r);
  AND2 I539 (rd_3r0[19:19], df_0[19:19], rg_3r);
  AND2 I540 (rd_3r0[20:20], df_0[20:20], rg_3r);
  AND2 I541 (rd_3r0[21:21], df_0[21:21], rg_3r);
  AND2 I542 (rd_3r0[22:22], df_0[22:22], rg_3r);
  AND2 I543 (rd_3r0[23:23], df_0[23:23], rg_3r);
  AND2 I544 (rd_3r0[24:24], df_0[24:24], rg_3r);
  AND2 I545 (rd_3r0[25:25], df_0[25:25], rg_3r);
  AND2 I546 (rd_3r0[26:26], df_0[26:26], rg_3r);
  AND2 I547 (rd_3r0[27:27], df_0[27:27], rg_3r);
  AND2 I548 (rd_3r0[28:28], df_0[28:28], rg_3r);
  AND2 I549 (rd_3r0[29:29], df_0[29:29], rg_3r);
  AND2 I550 (rd_3r0[30:30], df_0[30:30], rg_3r);
  AND2 I551 (rd_3r0[31:31], df_0[31:31], rg_3r);
  AND2 I552 (rd_4r0[0:0], df_0[0:0], rg_4r);
  AND2 I553 (rd_4r0[1:1], df_0[1:1], rg_4r);
  AND2 I554 (rd_4r0[2:2], df_0[2:2], rg_4r);
  AND2 I555 (rd_4r0[3:3], df_0[3:3], rg_4r);
  AND2 I556 (rd_4r0[4:4], df_0[4:4], rg_4r);
  AND2 I557 (rd_4r0[5:5], df_0[5:5], rg_4r);
  AND2 I558 (rd_4r0[6:6], df_0[6:6], rg_4r);
  AND2 I559 (rd_4r0[7:7], df_0[7:7], rg_4r);
  AND2 I560 (rd_4r0[8:8], df_0[8:8], rg_4r);
  AND2 I561 (rd_4r0[9:9], df_0[9:9], rg_4r);
  AND2 I562 (rd_4r0[10:10], df_0[10:10], rg_4r);
  AND2 I563 (rd_4r0[11:11], df_0[11:11], rg_4r);
  AND2 I564 (rd_4r0[12:12], df_0[12:12], rg_4r);
  AND2 I565 (rd_4r0[13:13], df_0[13:13], rg_4r);
  AND2 I566 (rd_4r0[14:14], df_0[14:14], rg_4r);
  AND2 I567 (rd_4r0[15:15], df_0[15:15], rg_4r);
  AND2 I568 (rd_4r0[16:16], df_0[16:16], rg_4r);
  AND2 I569 (rd_4r0[17:17], df_0[17:17], rg_4r);
  AND2 I570 (rd_4r0[18:18], df_0[18:18], rg_4r);
  AND2 I571 (rd_4r0[19:19], df_0[19:19], rg_4r);
  AND2 I572 (rd_4r0[20:20], df_0[20:20], rg_4r);
  AND2 I573 (rd_4r0[21:21], df_0[21:21], rg_4r);
  AND2 I574 (rd_4r0[22:22], df_0[22:22], rg_4r);
  AND2 I575 (rd_4r0[23:23], df_0[23:23], rg_4r);
  AND2 I576 (rd_4r0[24:24], df_0[24:24], rg_4r);
  AND2 I577 (rd_4r0[25:25], df_0[25:25], rg_4r);
  AND2 I578 (rd_4r0[26:26], df_0[26:26], rg_4r);
  AND2 I579 (rd_4r0[27:27], df_0[27:27], rg_4r);
  AND2 I580 (rd_4r0[28:28], df_0[28:28], rg_4r);
  AND2 I581 (rd_4r0[29:29], df_0[29:29], rg_4r);
  AND2 I582 (rd_4r0[30:30], df_0[30:30], rg_4r);
  AND2 I583 (rd_4r0[31:31], df_0[31:31], rg_4r);
  AND2 I584 (rd_5r0[0:0], df_0[0:0], rg_5r);
  AND2 I585 (rd_5r0[1:1], df_0[1:1], rg_5r);
  AND2 I586 (rd_5r0[2:2], df_0[2:2], rg_5r);
  AND2 I587 (rd_5r0[3:3], df_0[3:3], rg_5r);
  AND2 I588 (rd_5r0[4:4], df_0[4:4], rg_5r);
  AND2 I589 (rd_5r0[5:5], df_0[5:5], rg_5r);
  AND2 I590 (rd_5r0[6:6], df_0[6:6], rg_5r);
  AND2 I591 (rd_5r0[7:7], df_0[7:7], rg_5r);
  AND2 I592 (rd_5r0[8:8], df_0[8:8], rg_5r);
  AND2 I593 (rd_5r0[9:9], df_0[9:9], rg_5r);
  AND2 I594 (rd_5r0[10:10], df_0[10:10], rg_5r);
  AND2 I595 (rd_5r0[11:11], df_0[11:11], rg_5r);
  AND2 I596 (rd_5r0[12:12], df_0[12:12], rg_5r);
  AND2 I597 (rd_5r0[13:13], df_0[13:13], rg_5r);
  AND2 I598 (rd_5r0[14:14], df_0[14:14], rg_5r);
  AND2 I599 (rd_5r0[15:15], df_0[15:15], rg_5r);
  AND2 I600 (rd_5r0[16:16], df_0[16:16], rg_5r);
  AND2 I601 (rd_5r0[17:17], df_0[17:17], rg_5r);
  AND2 I602 (rd_5r0[18:18], df_0[18:18], rg_5r);
  AND2 I603 (rd_5r0[19:19], df_0[19:19], rg_5r);
  AND2 I604 (rd_5r0[20:20], df_0[20:20], rg_5r);
  AND2 I605 (rd_5r0[21:21], df_0[21:21], rg_5r);
  AND2 I606 (rd_5r0[22:22], df_0[22:22], rg_5r);
  AND2 I607 (rd_5r0[23:23], df_0[23:23], rg_5r);
  AND2 I608 (rd_5r0[24:24], df_0[24:24], rg_5r);
  AND2 I609 (rd_5r0[25:25], df_0[25:25], rg_5r);
  AND2 I610 (rd_5r0[26:26], df_0[26:26], rg_5r);
  AND2 I611 (rd_5r0[27:27], df_0[27:27], rg_5r);
  AND2 I612 (rd_5r0[28:28], df_0[28:28], rg_5r);
  AND2 I613 (rd_5r0[29:29], df_0[29:29], rg_5r);
  AND2 I614 (rd_5r0[30:30], df_0[30:30], rg_5r);
  AND2 I615 (rd_5r0[31:31], df_0[31:31], rg_5r);
  AND2 I616 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I617 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I618 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I619 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I620 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I621 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I622 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I623 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I624 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I625 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I626 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I627 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I628 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I629 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I630 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I631 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I632 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I633 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I634 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I635 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I636 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I637 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I638 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I639 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I640 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I641 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I642 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I643 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I644 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I645 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I646 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I647 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I648 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I649 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I650 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I651 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I652 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I653 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I654 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I655 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I656 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I657 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I658 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I659 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I660 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I661 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I662 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I663 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I664 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I665 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I666 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I667 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I668 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I669 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I670 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I671 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I672 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I673 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I674 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I675 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I676 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I677 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I678 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I679 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I680 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I681 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I682 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I683 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I684 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I685 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I686 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I687 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I688 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I689 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I690 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I691 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I692 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I693 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I694 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I695 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I696 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I697 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I698 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I699 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I700 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I701 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I702 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I703 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I704 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I705 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I706 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I707 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I708 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I709 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I710 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I711 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  AND2 I712 (rd_3r1[0:0], dt_0[0:0], rg_3r);
  AND2 I713 (rd_3r1[1:1], dt_0[1:1], rg_3r);
  AND2 I714 (rd_3r1[2:2], dt_0[2:2], rg_3r);
  AND2 I715 (rd_3r1[3:3], dt_0[3:3], rg_3r);
  AND2 I716 (rd_3r1[4:4], dt_0[4:4], rg_3r);
  AND2 I717 (rd_3r1[5:5], dt_0[5:5], rg_3r);
  AND2 I718 (rd_3r1[6:6], dt_0[6:6], rg_3r);
  AND2 I719 (rd_3r1[7:7], dt_0[7:7], rg_3r);
  AND2 I720 (rd_3r1[8:8], dt_0[8:8], rg_3r);
  AND2 I721 (rd_3r1[9:9], dt_0[9:9], rg_3r);
  AND2 I722 (rd_3r1[10:10], dt_0[10:10], rg_3r);
  AND2 I723 (rd_3r1[11:11], dt_0[11:11], rg_3r);
  AND2 I724 (rd_3r1[12:12], dt_0[12:12], rg_3r);
  AND2 I725 (rd_3r1[13:13], dt_0[13:13], rg_3r);
  AND2 I726 (rd_3r1[14:14], dt_0[14:14], rg_3r);
  AND2 I727 (rd_3r1[15:15], dt_0[15:15], rg_3r);
  AND2 I728 (rd_3r1[16:16], dt_0[16:16], rg_3r);
  AND2 I729 (rd_3r1[17:17], dt_0[17:17], rg_3r);
  AND2 I730 (rd_3r1[18:18], dt_0[18:18], rg_3r);
  AND2 I731 (rd_3r1[19:19], dt_0[19:19], rg_3r);
  AND2 I732 (rd_3r1[20:20], dt_0[20:20], rg_3r);
  AND2 I733 (rd_3r1[21:21], dt_0[21:21], rg_3r);
  AND2 I734 (rd_3r1[22:22], dt_0[22:22], rg_3r);
  AND2 I735 (rd_3r1[23:23], dt_0[23:23], rg_3r);
  AND2 I736 (rd_3r1[24:24], dt_0[24:24], rg_3r);
  AND2 I737 (rd_3r1[25:25], dt_0[25:25], rg_3r);
  AND2 I738 (rd_3r1[26:26], dt_0[26:26], rg_3r);
  AND2 I739 (rd_3r1[27:27], dt_0[27:27], rg_3r);
  AND2 I740 (rd_3r1[28:28], dt_0[28:28], rg_3r);
  AND2 I741 (rd_3r1[29:29], dt_0[29:29], rg_3r);
  AND2 I742 (rd_3r1[30:30], dt_0[30:30], rg_3r);
  AND2 I743 (rd_3r1[31:31], dt_0[31:31], rg_3r);
  AND2 I744 (rd_4r1[0:0], dt_0[0:0], rg_4r);
  AND2 I745 (rd_4r1[1:1], dt_0[1:1], rg_4r);
  AND2 I746 (rd_4r1[2:2], dt_0[2:2], rg_4r);
  AND2 I747 (rd_4r1[3:3], dt_0[3:3], rg_4r);
  AND2 I748 (rd_4r1[4:4], dt_0[4:4], rg_4r);
  AND2 I749 (rd_4r1[5:5], dt_0[5:5], rg_4r);
  AND2 I750 (rd_4r1[6:6], dt_0[6:6], rg_4r);
  AND2 I751 (rd_4r1[7:7], dt_0[7:7], rg_4r);
  AND2 I752 (rd_4r1[8:8], dt_0[8:8], rg_4r);
  AND2 I753 (rd_4r1[9:9], dt_0[9:9], rg_4r);
  AND2 I754 (rd_4r1[10:10], dt_0[10:10], rg_4r);
  AND2 I755 (rd_4r1[11:11], dt_0[11:11], rg_4r);
  AND2 I756 (rd_4r1[12:12], dt_0[12:12], rg_4r);
  AND2 I757 (rd_4r1[13:13], dt_0[13:13], rg_4r);
  AND2 I758 (rd_4r1[14:14], dt_0[14:14], rg_4r);
  AND2 I759 (rd_4r1[15:15], dt_0[15:15], rg_4r);
  AND2 I760 (rd_4r1[16:16], dt_0[16:16], rg_4r);
  AND2 I761 (rd_4r1[17:17], dt_0[17:17], rg_4r);
  AND2 I762 (rd_4r1[18:18], dt_0[18:18], rg_4r);
  AND2 I763 (rd_4r1[19:19], dt_0[19:19], rg_4r);
  AND2 I764 (rd_4r1[20:20], dt_0[20:20], rg_4r);
  AND2 I765 (rd_4r1[21:21], dt_0[21:21], rg_4r);
  AND2 I766 (rd_4r1[22:22], dt_0[22:22], rg_4r);
  AND2 I767 (rd_4r1[23:23], dt_0[23:23], rg_4r);
  AND2 I768 (rd_4r1[24:24], dt_0[24:24], rg_4r);
  AND2 I769 (rd_4r1[25:25], dt_0[25:25], rg_4r);
  AND2 I770 (rd_4r1[26:26], dt_0[26:26], rg_4r);
  AND2 I771 (rd_4r1[27:27], dt_0[27:27], rg_4r);
  AND2 I772 (rd_4r1[28:28], dt_0[28:28], rg_4r);
  AND2 I773 (rd_4r1[29:29], dt_0[29:29], rg_4r);
  AND2 I774 (rd_4r1[30:30], dt_0[30:30], rg_4r);
  AND2 I775 (rd_4r1[31:31], dt_0[31:31], rg_4r);
  AND2 I776 (rd_5r1[0:0], dt_0[0:0], rg_5r);
  AND2 I777 (rd_5r1[1:1], dt_0[1:1], rg_5r);
  AND2 I778 (rd_5r1[2:2], dt_0[2:2], rg_5r);
  AND2 I779 (rd_5r1[3:3], dt_0[3:3], rg_5r);
  AND2 I780 (rd_5r1[4:4], dt_0[4:4], rg_5r);
  AND2 I781 (rd_5r1[5:5], dt_0[5:5], rg_5r);
  AND2 I782 (rd_5r1[6:6], dt_0[6:6], rg_5r);
  AND2 I783 (rd_5r1[7:7], dt_0[7:7], rg_5r);
  AND2 I784 (rd_5r1[8:8], dt_0[8:8], rg_5r);
  AND2 I785 (rd_5r1[9:9], dt_0[9:9], rg_5r);
  AND2 I786 (rd_5r1[10:10], dt_0[10:10], rg_5r);
  AND2 I787 (rd_5r1[11:11], dt_0[11:11], rg_5r);
  AND2 I788 (rd_5r1[12:12], dt_0[12:12], rg_5r);
  AND2 I789 (rd_5r1[13:13], dt_0[13:13], rg_5r);
  AND2 I790 (rd_5r1[14:14], dt_0[14:14], rg_5r);
  AND2 I791 (rd_5r1[15:15], dt_0[15:15], rg_5r);
  AND2 I792 (rd_5r1[16:16], dt_0[16:16], rg_5r);
  AND2 I793 (rd_5r1[17:17], dt_0[17:17], rg_5r);
  AND2 I794 (rd_5r1[18:18], dt_0[18:18], rg_5r);
  AND2 I795 (rd_5r1[19:19], dt_0[19:19], rg_5r);
  AND2 I796 (rd_5r1[20:20], dt_0[20:20], rg_5r);
  AND2 I797 (rd_5r1[21:21], dt_0[21:21], rg_5r);
  AND2 I798 (rd_5r1[22:22], dt_0[22:22], rg_5r);
  AND2 I799 (rd_5r1[23:23], dt_0[23:23], rg_5r);
  AND2 I800 (rd_5r1[24:24], dt_0[24:24], rg_5r);
  AND2 I801 (rd_5r1[25:25], dt_0[25:25], rg_5r);
  AND2 I802 (rd_5r1[26:26], dt_0[26:26], rg_5r);
  AND2 I803 (rd_5r1[27:27], dt_0[27:27], rg_5r);
  AND2 I804 (rd_5r1[28:28], dt_0[28:28], rg_5r);
  AND2 I805 (rd_5r1[29:29], dt_0[29:29], rg_5r);
  AND2 I806 (rd_5r1[30:30], dt_0[30:30], rg_5r);
  AND2 I807 (rd_5r1[31:31], dt_0[31:31], rg_5r);
  NOR3 I808 (simp7921_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I809 (simp7921_0[1:1], rg_3r, rg_4r, rg_5r);
  NOR3 I810 (simp7921_0[2:2], rg_0a, rg_1a, rg_2a);
  NOR3 I811 (simp7921_0[3:3], rg_3a, rg_4a, rg_5a);
  NAND3 I812 (simp7922_0[0:0], simp7921_0[0:0], simp7921_0[1:1], simp7921_0[2:2]);
  INV I813 (simp7922_0[1:1], simp7921_0[3:3]);
  OR2 I814 (anyread_0, simp7922_0[0:0], simp7922_0[1:1]);
  BUFF I815 (wg_0a, wd_0a);
  BUFF I816 (rg_0a, rd_0a);
  BUFF I817 (rg_1a, rd_1a);
  BUFF I818 (rg_2a, rd_2a);
  BUFF I819 (rg_3a, rd_3a);
  BUFF I820 (rg_4a, rd_4a);
  BUFF I821 (rg_5a, rd_5a);
endmodule

// tkvinouts_15912832_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 TeakV "inouts[159:128]" 32 [] [0] [0,0,0,0
//   ,0,0] [Many [32],Many [0],Many [0,0,0,0,0,0],Many [32,32,32,32,32,32]]
module tkvinouts_15912832_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rg_5r, rg_5a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, rd_5r0, rd_5r1, rd_5a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  input rg_5r;
  output rg_5a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  output [31:0] rd_3r0;
  output [31:0] rd_3r1;
  input rd_3a;
  output [31:0] rd_4r0;
  output [31:0] rd_4r1;
  input rd_4a;
  output [31:0] rd_5r0;
  output [31:0] rd_5r1;
  input rd_5a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [3:0] simp7921_0;
  wire [1:0] simp7922_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_3r0[0:0], df_0[0:0], rg_3r);
  AND2 I521 (rd_3r0[1:1], df_0[1:1], rg_3r);
  AND2 I522 (rd_3r0[2:2], df_0[2:2], rg_3r);
  AND2 I523 (rd_3r0[3:3], df_0[3:3], rg_3r);
  AND2 I524 (rd_3r0[4:4], df_0[4:4], rg_3r);
  AND2 I525 (rd_3r0[5:5], df_0[5:5], rg_3r);
  AND2 I526 (rd_3r0[6:6], df_0[6:6], rg_3r);
  AND2 I527 (rd_3r0[7:7], df_0[7:7], rg_3r);
  AND2 I528 (rd_3r0[8:8], df_0[8:8], rg_3r);
  AND2 I529 (rd_3r0[9:9], df_0[9:9], rg_3r);
  AND2 I530 (rd_3r0[10:10], df_0[10:10], rg_3r);
  AND2 I531 (rd_3r0[11:11], df_0[11:11], rg_3r);
  AND2 I532 (rd_3r0[12:12], df_0[12:12], rg_3r);
  AND2 I533 (rd_3r0[13:13], df_0[13:13], rg_3r);
  AND2 I534 (rd_3r0[14:14], df_0[14:14], rg_3r);
  AND2 I535 (rd_3r0[15:15], df_0[15:15], rg_3r);
  AND2 I536 (rd_3r0[16:16], df_0[16:16], rg_3r);
  AND2 I537 (rd_3r0[17:17], df_0[17:17], rg_3r);
  AND2 I538 (rd_3r0[18:18], df_0[18:18], rg_3r);
  AND2 I539 (rd_3r0[19:19], df_0[19:19], rg_3r);
  AND2 I540 (rd_3r0[20:20], df_0[20:20], rg_3r);
  AND2 I541 (rd_3r0[21:21], df_0[21:21], rg_3r);
  AND2 I542 (rd_3r0[22:22], df_0[22:22], rg_3r);
  AND2 I543 (rd_3r0[23:23], df_0[23:23], rg_3r);
  AND2 I544 (rd_3r0[24:24], df_0[24:24], rg_3r);
  AND2 I545 (rd_3r0[25:25], df_0[25:25], rg_3r);
  AND2 I546 (rd_3r0[26:26], df_0[26:26], rg_3r);
  AND2 I547 (rd_3r0[27:27], df_0[27:27], rg_3r);
  AND2 I548 (rd_3r0[28:28], df_0[28:28], rg_3r);
  AND2 I549 (rd_3r0[29:29], df_0[29:29], rg_3r);
  AND2 I550 (rd_3r0[30:30], df_0[30:30], rg_3r);
  AND2 I551 (rd_3r0[31:31], df_0[31:31], rg_3r);
  AND2 I552 (rd_4r0[0:0], df_0[0:0], rg_4r);
  AND2 I553 (rd_4r0[1:1], df_0[1:1], rg_4r);
  AND2 I554 (rd_4r0[2:2], df_0[2:2], rg_4r);
  AND2 I555 (rd_4r0[3:3], df_0[3:3], rg_4r);
  AND2 I556 (rd_4r0[4:4], df_0[4:4], rg_4r);
  AND2 I557 (rd_4r0[5:5], df_0[5:5], rg_4r);
  AND2 I558 (rd_4r0[6:6], df_0[6:6], rg_4r);
  AND2 I559 (rd_4r0[7:7], df_0[7:7], rg_4r);
  AND2 I560 (rd_4r0[8:8], df_0[8:8], rg_4r);
  AND2 I561 (rd_4r0[9:9], df_0[9:9], rg_4r);
  AND2 I562 (rd_4r0[10:10], df_0[10:10], rg_4r);
  AND2 I563 (rd_4r0[11:11], df_0[11:11], rg_4r);
  AND2 I564 (rd_4r0[12:12], df_0[12:12], rg_4r);
  AND2 I565 (rd_4r0[13:13], df_0[13:13], rg_4r);
  AND2 I566 (rd_4r0[14:14], df_0[14:14], rg_4r);
  AND2 I567 (rd_4r0[15:15], df_0[15:15], rg_4r);
  AND2 I568 (rd_4r0[16:16], df_0[16:16], rg_4r);
  AND2 I569 (rd_4r0[17:17], df_0[17:17], rg_4r);
  AND2 I570 (rd_4r0[18:18], df_0[18:18], rg_4r);
  AND2 I571 (rd_4r0[19:19], df_0[19:19], rg_4r);
  AND2 I572 (rd_4r0[20:20], df_0[20:20], rg_4r);
  AND2 I573 (rd_4r0[21:21], df_0[21:21], rg_4r);
  AND2 I574 (rd_4r0[22:22], df_0[22:22], rg_4r);
  AND2 I575 (rd_4r0[23:23], df_0[23:23], rg_4r);
  AND2 I576 (rd_4r0[24:24], df_0[24:24], rg_4r);
  AND2 I577 (rd_4r0[25:25], df_0[25:25], rg_4r);
  AND2 I578 (rd_4r0[26:26], df_0[26:26], rg_4r);
  AND2 I579 (rd_4r0[27:27], df_0[27:27], rg_4r);
  AND2 I580 (rd_4r0[28:28], df_0[28:28], rg_4r);
  AND2 I581 (rd_4r0[29:29], df_0[29:29], rg_4r);
  AND2 I582 (rd_4r0[30:30], df_0[30:30], rg_4r);
  AND2 I583 (rd_4r0[31:31], df_0[31:31], rg_4r);
  AND2 I584 (rd_5r0[0:0], df_0[0:0], rg_5r);
  AND2 I585 (rd_5r0[1:1], df_0[1:1], rg_5r);
  AND2 I586 (rd_5r0[2:2], df_0[2:2], rg_5r);
  AND2 I587 (rd_5r0[3:3], df_0[3:3], rg_5r);
  AND2 I588 (rd_5r0[4:4], df_0[4:4], rg_5r);
  AND2 I589 (rd_5r0[5:5], df_0[5:5], rg_5r);
  AND2 I590 (rd_5r0[6:6], df_0[6:6], rg_5r);
  AND2 I591 (rd_5r0[7:7], df_0[7:7], rg_5r);
  AND2 I592 (rd_5r0[8:8], df_0[8:8], rg_5r);
  AND2 I593 (rd_5r0[9:9], df_0[9:9], rg_5r);
  AND2 I594 (rd_5r0[10:10], df_0[10:10], rg_5r);
  AND2 I595 (rd_5r0[11:11], df_0[11:11], rg_5r);
  AND2 I596 (rd_5r0[12:12], df_0[12:12], rg_5r);
  AND2 I597 (rd_5r0[13:13], df_0[13:13], rg_5r);
  AND2 I598 (rd_5r0[14:14], df_0[14:14], rg_5r);
  AND2 I599 (rd_5r0[15:15], df_0[15:15], rg_5r);
  AND2 I600 (rd_5r0[16:16], df_0[16:16], rg_5r);
  AND2 I601 (rd_5r0[17:17], df_0[17:17], rg_5r);
  AND2 I602 (rd_5r0[18:18], df_0[18:18], rg_5r);
  AND2 I603 (rd_5r0[19:19], df_0[19:19], rg_5r);
  AND2 I604 (rd_5r0[20:20], df_0[20:20], rg_5r);
  AND2 I605 (rd_5r0[21:21], df_0[21:21], rg_5r);
  AND2 I606 (rd_5r0[22:22], df_0[22:22], rg_5r);
  AND2 I607 (rd_5r0[23:23], df_0[23:23], rg_5r);
  AND2 I608 (rd_5r0[24:24], df_0[24:24], rg_5r);
  AND2 I609 (rd_5r0[25:25], df_0[25:25], rg_5r);
  AND2 I610 (rd_5r0[26:26], df_0[26:26], rg_5r);
  AND2 I611 (rd_5r0[27:27], df_0[27:27], rg_5r);
  AND2 I612 (rd_5r0[28:28], df_0[28:28], rg_5r);
  AND2 I613 (rd_5r0[29:29], df_0[29:29], rg_5r);
  AND2 I614 (rd_5r0[30:30], df_0[30:30], rg_5r);
  AND2 I615 (rd_5r0[31:31], df_0[31:31], rg_5r);
  AND2 I616 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I617 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I618 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I619 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I620 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I621 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I622 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I623 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I624 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I625 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I626 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I627 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I628 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I629 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I630 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I631 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I632 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I633 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I634 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I635 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I636 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I637 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I638 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I639 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I640 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I641 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I642 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I643 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I644 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I645 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I646 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I647 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I648 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I649 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I650 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I651 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I652 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I653 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I654 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I655 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I656 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I657 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I658 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I659 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I660 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I661 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I662 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I663 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I664 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I665 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I666 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I667 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I668 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I669 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I670 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I671 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I672 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I673 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I674 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I675 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I676 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I677 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I678 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I679 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I680 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I681 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I682 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I683 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I684 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I685 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I686 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I687 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I688 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I689 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I690 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I691 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I692 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I693 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I694 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I695 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I696 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I697 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I698 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I699 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I700 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I701 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I702 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I703 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I704 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I705 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I706 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I707 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I708 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I709 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I710 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I711 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  AND2 I712 (rd_3r1[0:0], dt_0[0:0], rg_3r);
  AND2 I713 (rd_3r1[1:1], dt_0[1:1], rg_3r);
  AND2 I714 (rd_3r1[2:2], dt_0[2:2], rg_3r);
  AND2 I715 (rd_3r1[3:3], dt_0[3:3], rg_3r);
  AND2 I716 (rd_3r1[4:4], dt_0[4:4], rg_3r);
  AND2 I717 (rd_3r1[5:5], dt_0[5:5], rg_3r);
  AND2 I718 (rd_3r1[6:6], dt_0[6:6], rg_3r);
  AND2 I719 (rd_3r1[7:7], dt_0[7:7], rg_3r);
  AND2 I720 (rd_3r1[8:8], dt_0[8:8], rg_3r);
  AND2 I721 (rd_3r1[9:9], dt_0[9:9], rg_3r);
  AND2 I722 (rd_3r1[10:10], dt_0[10:10], rg_3r);
  AND2 I723 (rd_3r1[11:11], dt_0[11:11], rg_3r);
  AND2 I724 (rd_3r1[12:12], dt_0[12:12], rg_3r);
  AND2 I725 (rd_3r1[13:13], dt_0[13:13], rg_3r);
  AND2 I726 (rd_3r1[14:14], dt_0[14:14], rg_3r);
  AND2 I727 (rd_3r1[15:15], dt_0[15:15], rg_3r);
  AND2 I728 (rd_3r1[16:16], dt_0[16:16], rg_3r);
  AND2 I729 (rd_3r1[17:17], dt_0[17:17], rg_3r);
  AND2 I730 (rd_3r1[18:18], dt_0[18:18], rg_3r);
  AND2 I731 (rd_3r1[19:19], dt_0[19:19], rg_3r);
  AND2 I732 (rd_3r1[20:20], dt_0[20:20], rg_3r);
  AND2 I733 (rd_3r1[21:21], dt_0[21:21], rg_3r);
  AND2 I734 (rd_3r1[22:22], dt_0[22:22], rg_3r);
  AND2 I735 (rd_3r1[23:23], dt_0[23:23], rg_3r);
  AND2 I736 (rd_3r1[24:24], dt_0[24:24], rg_3r);
  AND2 I737 (rd_3r1[25:25], dt_0[25:25], rg_3r);
  AND2 I738 (rd_3r1[26:26], dt_0[26:26], rg_3r);
  AND2 I739 (rd_3r1[27:27], dt_0[27:27], rg_3r);
  AND2 I740 (rd_3r1[28:28], dt_0[28:28], rg_3r);
  AND2 I741 (rd_3r1[29:29], dt_0[29:29], rg_3r);
  AND2 I742 (rd_3r1[30:30], dt_0[30:30], rg_3r);
  AND2 I743 (rd_3r1[31:31], dt_0[31:31], rg_3r);
  AND2 I744 (rd_4r1[0:0], dt_0[0:0], rg_4r);
  AND2 I745 (rd_4r1[1:1], dt_0[1:1], rg_4r);
  AND2 I746 (rd_4r1[2:2], dt_0[2:2], rg_4r);
  AND2 I747 (rd_4r1[3:3], dt_0[3:3], rg_4r);
  AND2 I748 (rd_4r1[4:4], dt_0[4:4], rg_4r);
  AND2 I749 (rd_4r1[5:5], dt_0[5:5], rg_4r);
  AND2 I750 (rd_4r1[6:6], dt_0[6:6], rg_4r);
  AND2 I751 (rd_4r1[7:7], dt_0[7:7], rg_4r);
  AND2 I752 (rd_4r1[8:8], dt_0[8:8], rg_4r);
  AND2 I753 (rd_4r1[9:9], dt_0[9:9], rg_4r);
  AND2 I754 (rd_4r1[10:10], dt_0[10:10], rg_4r);
  AND2 I755 (rd_4r1[11:11], dt_0[11:11], rg_4r);
  AND2 I756 (rd_4r1[12:12], dt_0[12:12], rg_4r);
  AND2 I757 (rd_4r1[13:13], dt_0[13:13], rg_4r);
  AND2 I758 (rd_4r1[14:14], dt_0[14:14], rg_4r);
  AND2 I759 (rd_4r1[15:15], dt_0[15:15], rg_4r);
  AND2 I760 (rd_4r1[16:16], dt_0[16:16], rg_4r);
  AND2 I761 (rd_4r1[17:17], dt_0[17:17], rg_4r);
  AND2 I762 (rd_4r1[18:18], dt_0[18:18], rg_4r);
  AND2 I763 (rd_4r1[19:19], dt_0[19:19], rg_4r);
  AND2 I764 (rd_4r1[20:20], dt_0[20:20], rg_4r);
  AND2 I765 (rd_4r1[21:21], dt_0[21:21], rg_4r);
  AND2 I766 (rd_4r1[22:22], dt_0[22:22], rg_4r);
  AND2 I767 (rd_4r1[23:23], dt_0[23:23], rg_4r);
  AND2 I768 (rd_4r1[24:24], dt_0[24:24], rg_4r);
  AND2 I769 (rd_4r1[25:25], dt_0[25:25], rg_4r);
  AND2 I770 (rd_4r1[26:26], dt_0[26:26], rg_4r);
  AND2 I771 (rd_4r1[27:27], dt_0[27:27], rg_4r);
  AND2 I772 (rd_4r1[28:28], dt_0[28:28], rg_4r);
  AND2 I773 (rd_4r1[29:29], dt_0[29:29], rg_4r);
  AND2 I774 (rd_4r1[30:30], dt_0[30:30], rg_4r);
  AND2 I775 (rd_4r1[31:31], dt_0[31:31], rg_4r);
  AND2 I776 (rd_5r1[0:0], dt_0[0:0], rg_5r);
  AND2 I777 (rd_5r1[1:1], dt_0[1:1], rg_5r);
  AND2 I778 (rd_5r1[2:2], dt_0[2:2], rg_5r);
  AND2 I779 (rd_5r1[3:3], dt_0[3:3], rg_5r);
  AND2 I780 (rd_5r1[4:4], dt_0[4:4], rg_5r);
  AND2 I781 (rd_5r1[5:5], dt_0[5:5], rg_5r);
  AND2 I782 (rd_5r1[6:6], dt_0[6:6], rg_5r);
  AND2 I783 (rd_5r1[7:7], dt_0[7:7], rg_5r);
  AND2 I784 (rd_5r1[8:8], dt_0[8:8], rg_5r);
  AND2 I785 (rd_5r1[9:9], dt_0[9:9], rg_5r);
  AND2 I786 (rd_5r1[10:10], dt_0[10:10], rg_5r);
  AND2 I787 (rd_5r1[11:11], dt_0[11:11], rg_5r);
  AND2 I788 (rd_5r1[12:12], dt_0[12:12], rg_5r);
  AND2 I789 (rd_5r1[13:13], dt_0[13:13], rg_5r);
  AND2 I790 (rd_5r1[14:14], dt_0[14:14], rg_5r);
  AND2 I791 (rd_5r1[15:15], dt_0[15:15], rg_5r);
  AND2 I792 (rd_5r1[16:16], dt_0[16:16], rg_5r);
  AND2 I793 (rd_5r1[17:17], dt_0[17:17], rg_5r);
  AND2 I794 (rd_5r1[18:18], dt_0[18:18], rg_5r);
  AND2 I795 (rd_5r1[19:19], dt_0[19:19], rg_5r);
  AND2 I796 (rd_5r1[20:20], dt_0[20:20], rg_5r);
  AND2 I797 (rd_5r1[21:21], dt_0[21:21], rg_5r);
  AND2 I798 (rd_5r1[22:22], dt_0[22:22], rg_5r);
  AND2 I799 (rd_5r1[23:23], dt_0[23:23], rg_5r);
  AND2 I800 (rd_5r1[24:24], dt_0[24:24], rg_5r);
  AND2 I801 (rd_5r1[25:25], dt_0[25:25], rg_5r);
  AND2 I802 (rd_5r1[26:26], dt_0[26:26], rg_5r);
  AND2 I803 (rd_5r1[27:27], dt_0[27:27], rg_5r);
  AND2 I804 (rd_5r1[28:28], dt_0[28:28], rg_5r);
  AND2 I805 (rd_5r1[29:29], dt_0[29:29], rg_5r);
  AND2 I806 (rd_5r1[30:30], dt_0[30:30], rg_5r);
  AND2 I807 (rd_5r1[31:31], dt_0[31:31], rg_5r);
  NOR3 I808 (simp7921_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I809 (simp7921_0[1:1], rg_3r, rg_4r, rg_5r);
  NOR3 I810 (simp7921_0[2:2], rg_0a, rg_1a, rg_2a);
  NOR3 I811 (simp7921_0[3:3], rg_3a, rg_4a, rg_5a);
  NAND3 I812 (simp7922_0[0:0], simp7921_0[0:0], simp7921_0[1:1], simp7921_0[2:2]);
  INV I813 (simp7922_0[1:1], simp7921_0[3:3]);
  OR2 I814 (anyread_0, simp7922_0[0:0], simp7922_0[1:1]);
  BUFF I815 (wg_0a, wd_0a);
  BUFF I816 (rg_0a, rd_0a);
  BUFF I817 (rg_1a, rd_1a);
  BUFF I818 (rg_2a, rd_2a);
  BUFF I819 (rg_3a, rd_3a);
  BUFF I820 (rg_4a, rd_4a);
  BUFF I821 (rg_5a, rd_5a);
endmodule

// tkvinouts_19116032_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 TeakV "inouts[191:160]" 32 [] [0] [0,0,0,0
//   ,0,0] [Many [32],Many [0],Many [0,0,0,0,0,0],Many [32,32,32,32,32,32]]
module tkvinouts_19116032_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rg_5r, rg_5a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, rd_5r0, rd_5r1, rd_5a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  input rg_5r;
  output rg_5a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  output [31:0] rd_3r0;
  output [31:0] rd_3r1;
  input rd_3a;
  output [31:0] rd_4r0;
  output [31:0] rd_4r1;
  input rd_4a;
  output [31:0] rd_5r0;
  output [31:0] rd_5r1;
  input rd_5a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [3:0] simp7921_0;
  wire [1:0] simp7922_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_3r0[0:0], df_0[0:0], rg_3r);
  AND2 I521 (rd_3r0[1:1], df_0[1:1], rg_3r);
  AND2 I522 (rd_3r0[2:2], df_0[2:2], rg_3r);
  AND2 I523 (rd_3r0[3:3], df_0[3:3], rg_3r);
  AND2 I524 (rd_3r0[4:4], df_0[4:4], rg_3r);
  AND2 I525 (rd_3r0[5:5], df_0[5:5], rg_3r);
  AND2 I526 (rd_3r0[6:6], df_0[6:6], rg_3r);
  AND2 I527 (rd_3r0[7:7], df_0[7:7], rg_3r);
  AND2 I528 (rd_3r0[8:8], df_0[8:8], rg_3r);
  AND2 I529 (rd_3r0[9:9], df_0[9:9], rg_3r);
  AND2 I530 (rd_3r0[10:10], df_0[10:10], rg_3r);
  AND2 I531 (rd_3r0[11:11], df_0[11:11], rg_3r);
  AND2 I532 (rd_3r0[12:12], df_0[12:12], rg_3r);
  AND2 I533 (rd_3r0[13:13], df_0[13:13], rg_3r);
  AND2 I534 (rd_3r0[14:14], df_0[14:14], rg_3r);
  AND2 I535 (rd_3r0[15:15], df_0[15:15], rg_3r);
  AND2 I536 (rd_3r0[16:16], df_0[16:16], rg_3r);
  AND2 I537 (rd_3r0[17:17], df_0[17:17], rg_3r);
  AND2 I538 (rd_3r0[18:18], df_0[18:18], rg_3r);
  AND2 I539 (rd_3r0[19:19], df_0[19:19], rg_3r);
  AND2 I540 (rd_3r0[20:20], df_0[20:20], rg_3r);
  AND2 I541 (rd_3r0[21:21], df_0[21:21], rg_3r);
  AND2 I542 (rd_3r0[22:22], df_0[22:22], rg_3r);
  AND2 I543 (rd_3r0[23:23], df_0[23:23], rg_3r);
  AND2 I544 (rd_3r0[24:24], df_0[24:24], rg_3r);
  AND2 I545 (rd_3r0[25:25], df_0[25:25], rg_3r);
  AND2 I546 (rd_3r0[26:26], df_0[26:26], rg_3r);
  AND2 I547 (rd_3r0[27:27], df_0[27:27], rg_3r);
  AND2 I548 (rd_3r0[28:28], df_0[28:28], rg_3r);
  AND2 I549 (rd_3r0[29:29], df_0[29:29], rg_3r);
  AND2 I550 (rd_3r0[30:30], df_0[30:30], rg_3r);
  AND2 I551 (rd_3r0[31:31], df_0[31:31], rg_3r);
  AND2 I552 (rd_4r0[0:0], df_0[0:0], rg_4r);
  AND2 I553 (rd_4r0[1:1], df_0[1:1], rg_4r);
  AND2 I554 (rd_4r0[2:2], df_0[2:2], rg_4r);
  AND2 I555 (rd_4r0[3:3], df_0[3:3], rg_4r);
  AND2 I556 (rd_4r0[4:4], df_0[4:4], rg_4r);
  AND2 I557 (rd_4r0[5:5], df_0[5:5], rg_4r);
  AND2 I558 (rd_4r0[6:6], df_0[6:6], rg_4r);
  AND2 I559 (rd_4r0[7:7], df_0[7:7], rg_4r);
  AND2 I560 (rd_4r0[8:8], df_0[8:8], rg_4r);
  AND2 I561 (rd_4r0[9:9], df_0[9:9], rg_4r);
  AND2 I562 (rd_4r0[10:10], df_0[10:10], rg_4r);
  AND2 I563 (rd_4r0[11:11], df_0[11:11], rg_4r);
  AND2 I564 (rd_4r0[12:12], df_0[12:12], rg_4r);
  AND2 I565 (rd_4r0[13:13], df_0[13:13], rg_4r);
  AND2 I566 (rd_4r0[14:14], df_0[14:14], rg_4r);
  AND2 I567 (rd_4r0[15:15], df_0[15:15], rg_4r);
  AND2 I568 (rd_4r0[16:16], df_0[16:16], rg_4r);
  AND2 I569 (rd_4r0[17:17], df_0[17:17], rg_4r);
  AND2 I570 (rd_4r0[18:18], df_0[18:18], rg_4r);
  AND2 I571 (rd_4r0[19:19], df_0[19:19], rg_4r);
  AND2 I572 (rd_4r0[20:20], df_0[20:20], rg_4r);
  AND2 I573 (rd_4r0[21:21], df_0[21:21], rg_4r);
  AND2 I574 (rd_4r0[22:22], df_0[22:22], rg_4r);
  AND2 I575 (rd_4r0[23:23], df_0[23:23], rg_4r);
  AND2 I576 (rd_4r0[24:24], df_0[24:24], rg_4r);
  AND2 I577 (rd_4r0[25:25], df_0[25:25], rg_4r);
  AND2 I578 (rd_4r0[26:26], df_0[26:26], rg_4r);
  AND2 I579 (rd_4r0[27:27], df_0[27:27], rg_4r);
  AND2 I580 (rd_4r0[28:28], df_0[28:28], rg_4r);
  AND2 I581 (rd_4r0[29:29], df_0[29:29], rg_4r);
  AND2 I582 (rd_4r0[30:30], df_0[30:30], rg_4r);
  AND2 I583 (rd_4r0[31:31], df_0[31:31], rg_4r);
  AND2 I584 (rd_5r0[0:0], df_0[0:0], rg_5r);
  AND2 I585 (rd_5r0[1:1], df_0[1:1], rg_5r);
  AND2 I586 (rd_5r0[2:2], df_0[2:2], rg_5r);
  AND2 I587 (rd_5r0[3:3], df_0[3:3], rg_5r);
  AND2 I588 (rd_5r0[4:4], df_0[4:4], rg_5r);
  AND2 I589 (rd_5r0[5:5], df_0[5:5], rg_5r);
  AND2 I590 (rd_5r0[6:6], df_0[6:6], rg_5r);
  AND2 I591 (rd_5r0[7:7], df_0[7:7], rg_5r);
  AND2 I592 (rd_5r0[8:8], df_0[8:8], rg_5r);
  AND2 I593 (rd_5r0[9:9], df_0[9:9], rg_5r);
  AND2 I594 (rd_5r0[10:10], df_0[10:10], rg_5r);
  AND2 I595 (rd_5r0[11:11], df_0[11:11], rg_5r);
  AND2 I596 (rd_5r0[12:12], df_0[12:12], rg_5r);
  AND2 I597 (rd_5r0[13:13], df_0[13:13], rg_5r);
  AND2 I598 (rd_5r0[14:14], df_0[14:14], rg_5r);
  AND2 I599 (rd_5r0[15:15], df_0[15:15], rg_5r);
  AND2 I600 (rd_5r0[16:16], df_0[16:16], rg_5r);
  AND2 I601 (rd_5r0[17:17], df_0[17:17], rg_5r);
  AND2 I602 (rd_5r0[18:18], df_0[18:18], rg_5r);
  AND2 I603 (rd_5r0[19:19], df_0[19:19], rg_5r);
  AND2 I604 (rd_5r0[20:20], df_0[20:20], rg_5r);
  AND2 I605 (rd_5r0[21:21], df_0[21:21], rg_5r);
  AND2 I606 (rd_5r0[22:22], df_0[22:22], rg_5r);
  AND2 I607 (rd_5r0[23:23], df_0[23:23], rg_5r);
  AND2 I608 (rd_5r0[24:24], df_0[24:24], rg_5r);
  AND2 I609 (rd_5r0[25:25], df_0[25:25], rg_5r);
  AND2 I610 (rd_5r0[26:26], df_0[26:26], rg_5r);
  AND2 I611 (rd_5r0[27:27], df_0[27:27], rg_5r);
  AND2 I612 (rd_5r0[28:28], df_0[28:28], rg_5r);
  AND2 I613 (rd_5r0[29:29], df_0[29:29], rg_5r);
  AND2 I614 (rd_5r0[30:30], df_0[30:30], rg_5r);
  AND2 I615 (rd_5r0[31:31], df_0[31:31], rg_5r);
  AND2 I616 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I617 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I618 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I619 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I620 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I621 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I622 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I623 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I624 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I625 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I626 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I627 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I628 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I629 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I630 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I631 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I632 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I633 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I634 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I635 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I636 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I637 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I638 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I639 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I640 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I641 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I642 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I643 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I644 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I645 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I646 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I647 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I648 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I649 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I650 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I651 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I652 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I653 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I654 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I655 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I656 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I657 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I658 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I659 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I660 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I661 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I662 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I663 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I664 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I665 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I666 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I667 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I668 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I669 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I670 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I671 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I672 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I673 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I674 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I675 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I676 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I677 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I678 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I679 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I680 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I681 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I682 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I683 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I684 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I685 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I686 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I687 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I688 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I689 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I690 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I691 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I692 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I693 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I694 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I695 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I696 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I697 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I698 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I699 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I700 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I701 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I702 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I703 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I704 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I705 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I706 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I707 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I708 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I709 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I710 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I711 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  AND2 I712 (rd_3r1[0:0], dt_0[0:0], rg_3r);
  AND2 I713 (rd_3r1[1:1], dt_0[1:1], rg_3r);
  AND2 I714 (rd_3r1[2:2], dt_0[2:2], rg_3r);
  AND2 I715 (rd_3r1[3:3], dt_0[3:3], rg_3r);
  AND2 I716 (rd_3r1[4:4], dt_0[4:4], rg_3r);
  AND2 I717 (rd_3r1[5:5], dt_0[5:5], rg_3r);
  AND2 I718 (rd_3r1[6:6], dt_0[6:6], rg_3r);
  AND2 I719 (rd_3r1[7:7], dt_0[7:7], rg_3r);
  AND2 I720 (rd_3r1[8:8], dt_0[8:8], rg_3r);
  AND2 I721 (rd_3r1[9:9], dt_0[9:9], rg_3r);
  AND2 I722 (rd_3r1[10:10], dt_0[10:10], rg_3r);
  AND2 I723 (rd_3r1[11:11], dt_0[11:11], rg_3r);
  AND2 I724 (rd_3r1[12:12], dt_0[12:12], rg_3r);
  AND2 I725 (rd_3r1[13:13], dt_0[13:13], rg_3r);
  AND2 I726 (rd_3r1[14:14], dt_0[14:14], rg_3r);
  AND2 I727 (rd_3r1[15:15], dt_0[15:15], rg_3r);
  AND2 I728 (rd_3r1[16:16], dt_0[16:16], rg_3r);
  AND2 I729 (rd_3r1[17:17], dt_0[17:17], rg_3r);
  AND2 I730 (rd_3r1[18:18], dt_0[18:18], rg_3r);
  AND2 I731 (rd_3r1[19:19], dt_0[19:19], rg_3r);
  AND2 I732 (rd_3r1[20:20], dt_0[20:20], rg_3r);
  AND2 I733 (rd_3r1[21:21], dt_0[21:21], rg_3r);
  AND2 I734 (rd_3r1[22:22], dt_0[22:22], rg_3r);
  AND2 I735 (rd_3r1[23:23], dt_0[23:23], rg_3r);
  AND2 I736 (rd_3r1[24:24], dt_0[24:24], rg_3r);
  AND2 I737 (rd_3r1[25:25], dt_0[25:25], rg_3r);
  AND2 I738 (rd_3r1[26:26], dt_0[26:26], rg_3r);
  AND2 I739 (rd_3r1[27:27], dt_0[27:27], rg_3r);
  AND2 I740 (rd_3r1[28:28], dt_0[28:28], rg_3r);
  AND2 I741 (rd_3r1[29:29], dt_0[29:29], rg_3r);
  AND2 I742 (rd_3r1[30:30], dt_0[30:30], rg_3r);
  AND2 I743 (rd_3r1[31:31], dt_0[31:31], rg_3r);
  AND2 I744 (rd_4r1[0:0], dt_0[0:0], rg_4r);
  AND2 I745 (rd_4r1[1:1], dt_0[1:1], rg_4r);
  AND2 I746 (rd_4r1[2:2], dt_0[2:2], rg_4r);
  AND2 I747 (rd_4r1[3:3], dt_0[3:3], rg_4r);
  AND2 I748 (rd_4r1[4:4], dt_0[4:4], rg_4r);
  AND2 I749 (rd_4r1[5:5], dt_0[5:5], rg_4r);
  AND2 I750 (rd_4r1[6:6], dt_0[6:6], rg_4r);
  AND2 I751 (rd_4r1[7:7], dt_0[7:7], rg_4r);
  AND2 I752 (rd_4r1[8:8], dt_0[8:8], rg_4r);
  AND2 I753 (rd_4r1[9:9], dt_0[9:9], rg_4r);
  AND2 I754 (rd_4r1[10:10], dt_0[10:10], rg_4r);
  AND2 I755 (rd_4r1[11:11], dt_0[11:11], rg_4r);
  AND2 I756 (rd_4r1[12:12], dt_0[12:12], rg_4r);
  AND2 I757 (rd_4r1[13:13], dt_0[13:13], rg_4r);
  AND2 I758 (rd_4r1[14:14], dt_0[14:14], rg_4r);
  AND2 I759 (rd_4r1[15:15], dt_0[15:15], rg_4r);
  AND2 I760 (rd_4r1[16:16], dt_0[16:16], rg_4r);
  AND2 I761 (rd_4r1[17:17], dt_0[17:17], rg_4r);
  AND2 I762 (rd_4r1[18:18], dt_0[18:18], rg_4r);
  AND2 I763 (rd_4r1[19:19], dt_0[19:19], rg_4r);
  AND2 I764 (rd_4r1[20:20], dt_0[20:20], rg_4r);
  AND2 I765 (rd_4r1[21:21], dt_0[21:21], rg_4r);
  AND2 I766 (rd_4r1[22:22], dt_0[22:22], rg_4r);
  AND2 I767 (rd_4r1[23:23], dt_0[23:23], rg_4r);
  AND2 I768 (rd_4r1[24:24], dt_0[24:24], rg_4r);
  AND2 I769 (rd_4r1[25:25], dt_0[25:25], rg_4r);
  AND2 I770 (rd_4r1[26:26], dt_0[26:26], rg_4r);
  AND2 I771 (rd_4r1[27:27], dt_0[27:27], rg_4r);
  AND2 I772 (rd_4r1[28:28], dt_0[28:28], rg_4r);
  AND2 I773 (rd_4r1[29:29], dt_0[29:29], rg_4r);
  AND2 I774 (rd_4r1[30:30], dt_0[30:30], rg_4r);
  AND2 I775 (rd_4r1[31:31], dt_0[31:31], rg_4r);
  AND2 I776 (rd_5r1[0:0], dt_0[0:0], rg_5r);
  AND2 I777 (rd_5r1[1:1], dt_0[1:1], rg_5r);
  AND2 I778 (rd_5r1[2:2], dt_0[2:2], rg_5r);
  AND2 I779 (rd_5r1[3:3], dt_0[3:3], rg_5r);
  AND2 I780 (rd_5r1[4:4], dt_0[4:4], rg_5r);
  AND2 I781 (rd_5r1[5:5], dt_0[5:5], rg_5r);
  AND2 I782 (rd_5r1[6:6], dt_0[6:6], rg_5r);
  AND2 I783 (rd_5r1[7:7], dt_0[7:7], rg_5r);
  AND2 I784 (rd_5r1[8:8], dt_0[8:8], rg_5r);
  AND2 I785 (rd_5r1[9:9], dt_0[9:9], rg_5r);
  AND2 I786 (rd_5r1[10:10], dt_0[10:10], rg_5r);
  AND2 I787 (rd_5r1[11:11], dt_0[11:11], rg_5r);
  AND2 I788 (rd_5r1[12:12], dt_0[12:12], rg_5r);
  AND2 I789 (rd_5r1[13:13], dt_0[13:13], rg_5r);
  AND2 I790 (rd_5r1[14:14], dt_0[14:14], rg_5r);
  AND2 I791 (rd_5r1[15:15], dt_0[15:15], rg_5r);
  AND2 I792 (rd_5r1[16:16], dt_0[16:16], rg_5r);
  AND2 I793 (rd_5r1[17:17], dt_0[17:17], rg_5r);
  AND2 I794 (rd_5r1[18:18], dt_0[18:18], rg_5r);
  AND2 I795 (rd_5r1[19:19], dt_0[19:19], rg_5r);
  AND2 I796 (rd_5r1[20:20], dt_0[20:20], rg_5r);
  AND2 I797 (rd_5r1[21:21], dt_0[21:21], rg_5r);
  AND2 I798 (rd_5r1[22:22], dt_0[22:22], rg_5r);
  AND2 I799 (rd_5r1[23:23], dt_0[23:23], rg_5r);
  AND2 I800 (rd_5r1[24:24], dt_0[24:24], rg_5r);
  AND2 I801 (rd_5r1[25:25], dt_0[25:25], rg_5r);
  AND2 I802 (rd_5r1[26:26], dt_0[26:26], rg_5r);
  AND2 I803 (rd_5r1[27:27], dt_0[27:27], rg_5r);
  AND2 I804 (rd_5r1[28:28], dt_0[28:28], rg_5r);
  AND2 I805 (rd_5r1[29:29], dt_0[29:29], rg_5r);
  AND2 I806 (rd_5r1[30:30], dt_0[30:30], rg_5r);
  AND2 I807 (rd_5r1[31:31], dt_0[31:31], rg_5r);
  NOR3 I808 (simp7921_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I809 (simp7921_0[1:1], rg_3r, rg_4r, rg_5r);
  NOR3 I810 (simp7921_0[2:2], rg_0a, rg_1a, rg_2a);
  NOR3 I811 (simp7921_0[3:3], rg_3a, rg_4a, rg_5a);
  NAND3 I812 (simp7922_0[0:0], simp7921_0[0:0], simp7921_0[1:1], simp7921_0[2:2]);
  INV I813 (simp7922_0[1:1], simp7921_0[3:3]);
  OR2 I814 (anyread_0, simp7922_0[0:0], simp7922_0[1:1]);
  BUFF I815 (wg_0a, wd_0a);
  BUFF I816 (rg_0a, rd_0a);
  BUFF I817 (rg_1a, rd_1a);
  BUFF I818 (rg_2a, rd_2a);
  BUFF I819 (rg_3a, rd_3a);
  BUFF I820 (rg_4a, rd_4a);
  BUFF I821 (rg_5a, rd_5a);
endmodule

// tkvinouts_22319232_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 TeakV "inouts[223:192]" 32 [] [0] [0,0,0,0
//   ,0,0] [Many [32],Many [0],Many [0,0,0,0,0,0],Many [32,32,32,32,32,32]]
module tkvinouts_22319232_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rg_5r, rg_5a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, rd_5r0, rd_5r1, rd_5a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  input rg_5r;
  output rg_5a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  output [31:0] rd_3r0;
  output [31:0] rd_3r1;
  input rd_3a;
  output [31:0] rd_4r0;
  output [31:0] rd_4r1;
  input rd_4a;
  output [31:0] rd_5r0;
  output [31:0] rd_5r1;
  input rd_5a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [3:0] simp7921_0;
  wire [1:0] simp7922_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_3r0[0:0], df_0[0:0], rg_3r);
  AND2 I521 (rd_3r0[1:1], df_0[1:1], rg_3r);
  AND2 I522 (rd_3r0[2:2], df_0[2:2], rg_3r);
  AND2 I523 (rd_3r0[3:3], df_0[3:3], rg_3r);
  AND2 I524 (rd_3r0[4:4], df_0[4:4], rg_3r);
  AND2 I525 (rd_3r0[5:5], df_0[5:5], rg_3r);
  AND2 I526 (rd_3r0[6:6], df_0[6:6], rg_3r);
  AND2 I527 (rd_3r0[7:7], df_0[7:7], rg_3r);
  AND2 I528 (rd_3r0[8:8], df_0[8:8], rg_3r);
  AND2 I529 (rd_3r0[9:9], df_0[9:9], rg_3r);
  AND2 I530 (rd_3r0[10:10], df_0[10:10], rg_3r);
  AND2 I531 (rd_3r0[11:11], df_0[11:11], rg_3r);
  AND2 I532 (rd_3r0[12:12], df_0[12:12], rg_3r);
  AND2 I533 (rd_3r0[13:13], df_0[13:13], rg_3r);
  AND2 I534 (rd_3r0[14:14], df_0[14:14], rg_3r);
  AND2 I535 (rd_3r0[15:15], df_0[15:15], rg_3r);
  AND2 I536 (rd_3r0[16:16], df_0[16:16], rg_3r);
  AND2 I537 (rd_3r0[17:17], df_0[17:17], rg_3r);
  AND2 I538 (rd_3r0[18:18], df_0[18:18], rg_3r);
  AND2 I539 (rd_3r0[19:19], df_0[19:19], rg_3r);
  AND2 I540 (rd_3r0[20:20], df_0[20:20], rg_3r);
  AND2 I541 (rd_3r0[21:21], df_0[21:21], rg_3r);
  AND2 I542 (rd_3r0[22:22], df_0[22:22], rg_3r);
  AND2 I543 (rd_3r0[23:23], df_0[23:23], rg_3r);
  AND2 I544 (rd_3r0[24:24], df_0[24:24], rg_3r);
  AND2 I545 (rd_3r0[25:25], df_0[25:25], rg_3r);
  AND2 I546 (rd_3r0[26:26], df_0[26:26], rg_3r);
  AND2 I547 (rd_3r0[27:27], df_0[27:27], rg_3r);
  AND2 I548 (rd_3r0[28:28], df_0[28:28], rg_3r);
  AND2 I549 (rd_3r0[29:29], df_0[29:29], rg_3r);
  AND2 I550 (rd_3r0[30:30], df_0[30:30], rg_3r);
  AND2 I551 (rd_3r0[31:31], df_0[31:31], rg_3r);
  AND2 I552 (rd_4r0[0:0], df_0[0:0], rg_4r);
  AND2 I553 (rd_4r0[1:1], df_0[1:1], rg_4r);
  AND2 I554 (rd_4r0[2:2], df_0[2:2], rg_4r);
  AND2 I555 (rd_4r0[3:3], df_0[3:3], rg_4r);
  AND2 I556 (rd_4r0[4:4], df_0[4:4], rg_4r);
  AND2 I557 (rd_4r0[5:5], df_0[5:5], rg_4r);
  AND2 I558 (rd_4r0[6:6], df_0[6:6], rg_4r);
  AND2 I559 (rd_4r0[7:7], df_0[7:7], rg_4r);
  AND2 I560 (rd_4r0[8:8], df_0[8:8], rg_4r);
  AND2 I561 (rd_4r0[9:9], df_0[9:9], rg_4r);
  AND2 I562 (rd_4r0[10:10], df_0[10:10], rg_4r);
  AND2 I563 (rd_4r0[11:11], df_0[11:11], rg_4r);
  AND2 I564 (rd_4r0[12:12], df_0[12:12], rg_4r);
  AND2 I565 (rd_4r0[13:13], df_0[13:13], rg_4r);
  AND2 I566 (rd_4r0[14:14], df_0[14:14], rg_4r);
  AND2 I567 (rd_4r0[15:15], df_0[15:15], rg_4r);
  AND2 I568 (rd_4r0[16:16], df_0[16:16], rg_4r);
  AND2 I569 (rd_4r0[17:17], df_0[17:17], rg_4r);
  AND2 I570 (rd_4r0[18:18], df_0[18:18], rg_4r);
  AND2 I571 (rd_4r0[19:19], df_0[19:19], rg_4r);
  AND2 I572 (rd_4r0[20:20], df_0[20:20], rg_4r);
  AND2 I573 (rd_4r0[21:21], df_0[21:21], rg_4r);
  AND2 I574 (rd_4r0[22:22], df_0[22:22], rg_4r);
  AND2 I575 (rd_4r0[23:23], df_0[23:23], rg_4r);
  AND2 I576 (rd_4r0[24:24], df_0[24:24], rg_4r);
  AND2 I577 (rd_4r0[25:25], df_0[25:25], rg_4r);
  AND2 I578 (rd_4r0[26:26], df_0[26:26], rg_4r);
  AND2 I579 (rd_4r0[27:27], df_0[27:27], rg_4r);
  AND2 I580 (rd_4r0[28:28], df_0[28:28], rg_4r);
  AND2 I581 (rd_4r0[29:29], df_0[29:29], rg_4r);
  AND2 I582 (rd_4r0[30:30], df_0[30:30], rg_4r);
  AND2 I583 (rd_4r0[31:31], df_0[31:31], rg_4r);
  AND2 I584 (rd_5r0[0:0], df_0[0:0], rg_5r);
  AND2 I585 (rd_5r0[1:1], df_0[1:1], rg_5r);
  AND2 I586 (rd_5r0[2:2], df_0[2:2], rg_5r);
  AND2 I587 (rd_5r0[3:3], df_0[3:3], rg_5r);
  AND2 I588 (rd_5r0[4:4], df_0[4:4], rg_5r);
  AND2 I589 (rd_5r0[5:5], df_0[5:5], rg_5r);
  AND2 I590 (rd_5r0[6:6], df_0[6:6], rg_5r);
  AND2 I591 (rd_5r0[7:7], df_0[7:7], rg_5r);
  AND2 I592 (rd_5r0[8:8], df_0[8:8], rg_5r);
  AND2 I593 (rd_5r0[9:9], df_0[9:9], rg_5r);
  AND2 I594 (rd_5r0[10:10], df_0[10:10], rg_5r);
  AND2 I595 (rd_5r0[11:11], df_0[11:11], rg_5r);
  AND2 I596 (rd_5r0[12:12], df_0[12:12], rg_5r);
  AND2 I597 (rd_5r0[13:13], df_0[13:13], rg_5r);
  AND2 I598 (rd_5r0[14:14], df_0[14:14], rg_5r);
  AND2 I599 (rd_5r0[15:15], df_0[15:15], rg_5r);
  AND2 I600 (rd_5r0[16:16], df_0[16:16], rg_5r);
  AND2 I601 (rd_5r0[17:17], df_0[17:17], rg_5r);
  AND2 I602 (rd_5r0[18:18], df_0[18:18], rg_5r);
  AND2 I603 (rd_5r0[19:19], df_0[19:19], rg_5r);
  AND2 I604 (rd_5r0[20:20], df_0[20:20], rg_5r);
  AND2 I605 (rd_5r0[21:21], df_0[21:21], rg_5r);
  AND2 I606 (rd_5r0[22:22], df_0[22:22], rg_5r);
  AND2 I607 (rd_5r0[23:23], df_0[23:23], rg_5r);
  AND2 I608 (rd_5r0[24:24], df_0[24:24], rg_5r);
  AND2 I609 (rd_5r0[25:25], df_0[25:25], rg_5r);
  AND2 I610 (rd_5r0[26:26], df_0[26:26], rg_5r);
  AND2 I611 (rd_5r0[27:27], df_0[27:27], rg_5r);
  AND2 I612 (rd_5r0[28:28], df_0[28:28], rg_5r);
  AND2 I613 (rd_5r0[29:29], df_0[29:29], rg_5r);
  AND2 I614 (rd_5r0[30:30], df_0[30:30], rg_5r);
  AND2 I615 (rd_5r0[31:31], df_0[31:31], rg_5r);
  AND2 I616 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I617 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I618 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I619 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I620 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I621 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I622 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I623 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I624 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I625 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I626 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I627 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I628 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I629 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I630 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I631 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I632 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I633 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I634 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I635 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I636 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I637 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I638 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I639 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I640 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I641 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I642 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I643 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I644 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I645 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I646 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I647 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I648 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I649 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I650 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I651 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I652 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I653 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I654 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I655 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I656 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I657 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I658 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I659 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I660 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I661 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I662 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I663 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I664 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I665 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I666 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I667 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I668 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I669 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I670 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I671 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I672 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I673 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I674 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I675 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I676 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I677 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I678 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I679 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I680 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I681 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I682 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I683 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I684 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I685 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I686 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I687 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I688 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I689 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I690 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I691 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I692 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I693 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I694 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I695 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I696 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I697 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I698 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I699 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I700 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I701 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I702 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I703 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I704 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I705 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I706 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I707 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I708 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I709 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I710 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I711 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  AND2 I712 (rd_3r1[0:0], dt_0[0:0], rg_3r);
  AND2 I713 (rd_3r1[1:1], dt_0[1:1], rg_3r);
  AND2 I714 (rd_3r1[2:2], dt_0[2:2], rg_3r);
  AND2 I715 (rd_3r1[3:3], dt_0[3:3], rg_3r);
  AND2 I716 (rd_3r1[4:4], dt_0[4:4], rg_3r);
  AND2 I717 (rd_3r1[5:5], dt_0[5:5], rg_3r);
  AND2 I718 (rd_3r1[6:6], dt_0[6:6], rg_3r);
  AND2 I719 (rd_3r1[7:7], dt_0[7:7], rg_3r);
  AND2 I720 (rd_3r1[8:8], dt_0[8:8], rg_3r);
  AND2 I721 (rd_3r1[9:9], dt_0[9:9], rg_3r);
  AND2 I722 (rd_3r1[10:10], dt_0[10:10], rg_3r);
  AND2 I723 (rd_3r1[11:11], dt_0[11:11], rg_3r);
  AND2 I724 (rd_3r1[12:12], dt_0[12:12], rg_3r);
  AND2 I725 (rd_3r1[13:13], dt_0[13:13], rg_3r);
  AND2 I726 (rd_3r1[14:14], dt_0[14:14], rg_3r);
  AND2 I727 (rd_3r1[15:15], dt_0[15:15], rg_3r);
  AND2 I728 (rd_3r1[16:16], dt_0[16:16], rg_3r);
  AND2 I729 (rd_3r1[17:17], dt_0[17:17], rg_3r);
  AND2 I730 (rd_3r1[18:18], dt_0[18:18], rg_3r);
  AND2 I731 (rd_3r1[19:19], dt_0[19:19], rg_3r);
  AND2 I732 (rd_3r1[20:20], dt_0[20:20], rg_3r);
  AND2 I733 (rd_3r1[21:21], dt_0[21:21], rg_3r);
  AND2 I734 (rd_3r1[22:22], dt_0[22:22], rg_3r);
  AND2 I735 (rd_3r1[23:23], dt_0[23:23], rg_3r);
  AND2 I736 (rd_3r1[24:24], dt_0[24:24], rg_3r);
  AND2 I737 (rd_3r1[25:25], dt_0[25:25], rg_3r);
  AND2 I738 (rd_3r1[26:26], dt_0[26:26], rg_3r);
  AND2 I739 (rd_3r1[27:27], dt_0[27:27], rg_3r);
  AND2 I740 (rd_3r1[28:28], dt_0[28:28], rg_3r);
  AND2 I741 (rd_3r1[29:29], dt_0[29:29], rg_3r);
  AND2 I742 (rd_3r1[30:30], dt_0[30:30], rg_3r);
  AND2 I743 (rd_3r1[31:31], dt_0[31:31], rg_3r);
  AND2 I744 (rd_4r1[0:0], dt_0[0:0], rg_4r);
  AND2 I745 (rd_4r1[1:1], dt_0[1:1], rg_4r);
  AND2 I746 (rd_4r1[2:2], dt_0[2:2], rg_4r);
  AND2 I747 (rd_4r1[3:3], dt_0[3:3], rg_4r);
  AND2 I748 (rd_4r1[4:4], dt_0[4:4], rg_4r);
  AND2 I749 (rd_4r1[5:5], dt_0[5:5], rg_4r);
  AND2 I750 (rd_4r1[6:6], dt_0[6:6], rg_4r);
  AND2 I751 (rd_4r1[7:7], dt_0[7:7], rg_4r);
  AND2 I752 (rd_4r1[8:8], dt_0[8:8], rg_4r);
  AND2 I753 (rd_4r1[9:9], dt_0[9:9], rg_4r);
  AND2 I754 (rd_4r1[10:10], dt_0[10:10], rg_4r);
  AND2 I755 (rd_4r1[11:11], dt_0[11:11], rg_4r);
  AND2 I756 (rd_4r1[12:12], dt_0[12:12], rg_4r);
  AND2 I757 (rd_4r1[13:13], dt_0[13:13], rg_4r);
  AND2 I758 (rd_4r1[14:14], dt_0[14:14], rg_4r);
  AND2 I759 (rd_4r1[15:15], dt_0[15:15], rg_4r);
  AND2 I760 (rd_4r1[16:16], dt_0[16:16], rg_4r);
  AND2 I761 (rd_4r1[17:17], dt_0[17:17], rg_4r);
  AND2 I762 (rd_4r1[18:18], dt_0[18:18], rg_4r);
  AND2 I763 (rd_4r1[19:19], dt_0[19:19], rg_4r);
  AND2 I764 (rd_4r1[20:20], dt_0[20:20], rg_4r);
  AND2 I765 (rd_4r1[21:21], dt_0[21:21], rg_4r);
  AND2 I766 (rd_4r1[22:22], dt_0[22:22], rg_4r);
  AND2 I767 (rd_4r1[23:23], dt_0[23:23], rg_4r);
  AND2 I768 (rd_4r1[24:24], dt_0[24:24], rg_4r);
  AND2 I769 (rd_4r1[25:25], dt_0[25:25], rg_4r);
  AND2 I770 (rd_4r1[26:26], dt_0[26:26], rg_4r);
  AND2 I771 (rd_4r1[27:27], dt_0[27:27], rg_4r);
  AND2 I772 (rd_4r1[28:28], dt_0[28:28], rg_4r);
  AND2 I773 (rd_4r1[29:29], dt_0[29:29], rg_4r);
  AND2 I774 (rd_4r1[30:30], dt_0[30:30], rg_4r);
  AND2 I775 (rd_4r1[31:31], dt_0[31:31], rg_4r);
  AND2 I776 (rd_5r1[0:0], dt_0[0:0], rg_5r);
  AND2 I777 (rd_5r1[1:1], dt_0[1:1], rg_5r);
  AND2 I778 (rd_5r1[2:2], dt_0[2:2], rg_5r);
  AND2 I779 (rd_5r1[3:3], dt_0[3:3], rg_5r);
  AND2 I780 (rd_5r1[4:4], dt_0[4:4], rg_5r);
  AND2 I781 (rd_5r1[5:5], dt_0[5:5], rg_5r);
  AND2 I782 (rd_5r1[6:6], dt_0[6:6], rg_5r);
  AND2 I783 (rd_5r1[7:7], dt_0[7:7], rg_5r);
  AND2 I784 (rd_5r1[8:8], dt_0[8:8], rg_5r);
  AND2 I785 (rd_5r1[9:9], dt_0[9:9], rg_5r);
  AND2 I786 (rd_5r1[10:10], dt_0[10:10], rg_5r);
  AND2 I787 (rd_5r1[11:11], dt_0[11:11], rg_5r);
  AND2 I788 (rd_5r1[12:12], dt_0[12:12], rg_5r);
  AND2 I789 (rd_5r1[13:13], dt_0[13:13], rg_5r);
  AND2 I790 (rd_5r1[14:14], dt_0[14:14], rg_5r);
  AND2 I791 (rd_5r1[15:15], dt_0[15:15], rg_5r);
  AND2 I792 (rd_5r1[16:16], dt_0[16:16], rg_5r);
  AND2 I793 (rd_5r1[17:17], dt_0[17:17], rg_5r);
  AND2 I794 (rd_5r1[18:18], dt_0[18:18], rg_5r);
  AND2 I795 (rd_5r1[19:19], dt_0[19:19], rg_5r);
  AND2 I796 (rd_5r1[20:20], dt_0[20:20], rg_5r);
  AND2 I797 (rd_5r1[21:21], dt_0[21:21], rg_5r);
  AND2 I798 (rd_5r1[22:22], dt_0[22:22], rg_5r);
  AND2 I799 (rd_5r1[23:23], dt_0[23:23], rg_5r);
  AND2 I800 (rd_5r1[24:24], dt_0[24:24], rg_5r);
  AND2 I801 (rd_5r1[25:25], dt_0[25:25], rg_5r);
  AND2 I802 (rd_5r1[26:26], dt_0[26:26], rg_5r);
  AND2 I803 (rd_5r1[27:27], dt_0[27:27], rg_5r);
  AND2 I804 (rd_5r1[28:28], dt_0[28:28], rg_5r);
  AND2 I805 (rd_5r1[29:29], dt_0[29:29], rg_5r);
  AND2 I806 (rd_5r1[30:30], dt_0[30:30], rg_5r);
  AND2 I807 (rd_5r1[31:31], dt_0[31:31], rg_5r);
  NOR3 I808 (simp7921_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I809 (simp7921_0[1:1], rg_3r, rg_4r, rg_5r);
  NOR3 I810 (simp7921_0[2:2], rg_0a, rg_1a, rg_2a);
  NOR3 I811 (simp7921_0[3:3], rg_3a, rg_4a, rg_5a);
  NAND3 I812 (simp7922_0[0:0], simp7921_0[0:0], simp7921_0[1:1], simp7921_0[2:2]);
  INV I813 (simp7922_0[1:1], simp7921_0[3:3]);
  OR2 I814 (anyread_0, simp7922_0[0:0], simp7922_0[1:1]);
  BUFF I815 (wg_0a, wd_0a);
  BUFF I816 (rg_0a, rd_0a);
  BUFF I817 (rg_1a, rd_1a);
  BUFF I818 (rg_2a, rd_2a);
  BUFF I819 (rg_3a, rd_3a);
  BUFF I820 (rg_4a, rd_4a);
  BUFF I821 (rg_5a, rd_5a);
endmodule

// tkvinouts_25522432_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 TeakV "inouts[255:224]" 32 [] [0] [0,0,0,0
//   ,0,0] [Many [32],Many [0],Many [0,0,0,0,0,0],Many [32,32,32,32,32,32]]
module tkvinouts_25522432_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rg_5r, rg_5a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, rd_5r0, rd_5r1, rd_5a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  input rg_5r;
  output rg_5a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  output [31:0] rd_3r0;
  output [31:0] rd_3r1;
  input rd_3a;
  output [31:0] rd_4r0;
  output [31:0] rd_4r1;
  input rd_4a;
  output [31:0] rd_5r0;
  output [31:0] rd_5r1;
  input rd_5a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [3:0] simp7921_0;
  wire [1:0] simp7922_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_3r0[0:0], df_0[0:0], rg_3r);
  AND2 I521 (rd_3r0[1:1], df_0[1:1], rg_3r);
  AND2 I522 (rd_3r0[2:2], df_0[2:2], rg_3r);
  AND2 I523 (rd_3r0[3:3], df_0[3:3], rg_3r);
  AND2 I524 (rd_3r0[4:4], df_0[4:4], rg_3r);
  AND2 I525 (rd_3r0[5:5], df_0[5:5], rg_3r);
  AND2 I526 (rd_3r0[6:6], df_0[6:6], rg_3r);
  AND2 I527 (rd_3r0[7:7], df_0[7:7], rg_3r);
  AND2 I528 (rd_3r0[8:8], df_0[8:8], rg_3r);
  AND2 I529 (rd_3r0[9:9], df_0[9:9], rg_3r);
  AND2 I530 (rd_3r0[10:10], df_0[10:10], rg_3r);
  AND2 I531 (rd_3r0[11:11], df_0[11:11], rg_3r);
  AND2 I532 (rd_3r0[12:12], df_0[12:12], rg_3r);
  AND2 I533 (rd_3r0[13:13], df_0[13:13], rg_3r);
  AND2 I534 (rd_3r0[14:14], df_0[14:14], rg_3r);
  AND2 I535 (rd_3r0[15:15], df_0[15:15], rg_3r);
  AND2 I536 (rd_3r0[16:16], df_0[16:16], rg_3r);
  AND2 I537 (rd_3r0[17:17], df_0[17:17], rg_3r);
  AND2 I538 (rd_3r0[18:18], df_0[18:18], rg_3r);
  AND2 I539 (rd_3r0[19:19], df_0[19:19], rg_3r);
  AND2 I540 (rd_3r0[20:20], df_0[20:20], rg_3r);
  AND2 I541 (rd_3r0[21:21], df_0[21:21], rg_3r);
  AND2 I542 (rd_3r0[22:22], df_0[22:22], rg_3r);
  AND2 I543 (rd_3r0[23:23], df_0[23:23], rg_3r);
  AND2 I544 (rd_3r0[24:24], df_0[24:24], rg_3r);
  AND2 I545 (rd_3r0[25:25], df_0[25:25], rg_3r);
  AND2 I546 (rd_3r0[26:26], df_0[26:26], rg_3r);
  AND2 I547 (rd_3r0[27:27], df_0[27:27], rg_3r);
  AND2 I548 (rd_3r0[28:28], df_0[28:28], rg_3r);
  AND2 I549 (rd_3r0[29:29], df_0[29:29], rg_3r);
  AND2 I550 (rd_3r0[30:30], df_0[30:30], rg_3r);
  AND2 I551 (rd_3r0[31:31], df_0[31:31], rg_3r);
  AND2 I552 (rd_4r0[0:0], df_0[0:0], rg_4r);
  AND2 I553 (rd_4r0[1:1], df_0[1:1], rg_4r);
  AND2 I554 (rd_4r0[2:2], df_0[2:2], rg_4r);
  AND2 I555 (rd_4r0[3:3], df_0[3:3], rg_4r);
  AND2 I556 (rd_4r0[4:4], df_0[4:4], rg_4r);
  AND2 I557 (rd_4r0[5:5], df_0[5:5], rg_4r);
  AND2 I558 (rd_4r0[6:6], df_0[6:6], rg_4r);
  AND2 I559 (rd_4r0[7:7], df_0[7:7], rg_4r);
  AND2 I560 (rd_4r0[8:8], df_0[8:8], rg_4r);
  AND2 I561 (rd_4r0[9:9], df_0[9:9], rg_4r);
  AND2 I562 (rd_4r0[10:10], df_0[10:10], rg_4r);
  AND2 I563 (rd_4r0[11:11], df_0[11:11], rg_4r);
  AND2 I564 (rd_4r0[12:12], df_0[12:12], rg_4r);
  AND2 I565 (rd_4r0[13:13], df_0[13:13], rg_4r);
  AND2 I566 (rd_4r0[14:14], df_0[14:14], rg_4r);
  AND2 I567 (rd_4r0[15:15], df_0[15:15], rg_4r);
  AND2 I568 (rd_4r0[16:16], df_0[16:16], rg_4r);
  AND2 I569 (rd_4r0[17:17], df_0[17:17], rg_4r);
  AND2 I570 (rd_4r0[18:18], df_0[18:18], rg_4r);
  AND2 I571 (rd_4r0[19:19], df_0[19:19], rg_4r);
  AND2 I572 (rd_4r0[20:20], df_0[20:20], rg_4r);
  AND2 I573 (rd_4r0[21:21], df_0[21:21], rg_4r);
  AND2 I574 (rd_4r0[22:22], df_0[22:22], rg_4r);
  AND2 I575 (rd_4r0[23:23], df_0[23:23], rg_4r);
  AND2 I576 (rd_4r0[24:24], df_0[24:24], rg_4r);
  AND2 I577 (rd_4r0[25:25], df_0[25:25], rg_4r);
  AND2 I578 (rd_4r0[26:26], df_0[26:26], rg_4r);
  AND2 I579 (rd_4r0[27:27], df_0[27:27], rg_4r);
  AND2 I580 (rd_4r0[28:28], df_0[28:28], rg_4r);
  AND2 I581 (rd_4r0[29:29], df_0[29:29], rg_4r);
  AND2 I582 (rd_4r0[30:30], df_0[30:30], rg_4r);
  AND2 I583 (rd_4r0[31:31], df_0[31:31], rg_4r);
  AND2 I584 (rd_5r0[0:0], df_0[0:0], rg_5r);
  AND2 I585 (rd_5r0[1:1], df_0[1:1], rg_5r);
  AND2 I586 (rd_5r0[2:2], df_0[2:2], rg_5r);
  AND2 I587 (rd_5r0[3:3], df_0[3:3], rg_5r);
  AND2 I588 (rd_5r0[4:4], df_0[4:4], rg_5r);
  AND2 I589 (rd_5r0[5:5], df_0[5:5], rg_5r);
  AND2 I590 (rd_5r0[6:6], df_0[6:6], rg_5r);
  AND2 I591 (rd_5r0[7:7], df_0[7:7], rg_5r);
  AND2 I592 (rd_5r0[8:8], df_0[8:8], rg_5r);
  AND2 I593 (rd_5r0[9:9], df_0[9:9], rg_5r);
  AND2 I594 (rd_5r0[10:10], df_0[10:10], rg_5r);
  AND2 I595 (rd_5r0[11:11], df_0[11:11], rg_5r);
  AND2 I596 (rd_5r0[12:12], df_0[12:12], rg_5r);
  AND2 I597 (rd_5r0[13:13], df_0[13:13], rg_5r);
  AND2 I598 (rd_5r0[14:14], df_0[14:14], rg_5r);
  AND2 I599 (rd_5r0[15:15], df_0[15:15], rg_5r);
  AND2 I600 (rd_5r0[16:16], df_0[16:16], rg_5r);
  AND2 I601 (rd_5r0[17:17], df_0[17:17], rg_5r);
  AND2 I602 (rd_5r0[18:18], df_0[18:18], rg_5r);
  AND2 I603 (rd_5r0[19:19], df_0[19:19], rg_5r);
  AND2 I604 (rd_5r0[20:20], df_0[20:20], rg_5r);
  AND2 I605 (rd_5r0[21:21], df_0[21:21], rg_5r);
  AND2 I606 (rd_5r0[22:22], df_0[22:22], rg_5r);
  AND2 I607 (rd_5r0[23:23], df_0[23:23], rg_5r);
  AND2 I608 (rd_5r0[24:24], df_0[24:24], rg_5r);
  AND2 I609 (rd_5r0[25:25], df_0[25:25], rg_5r);
  AND2 I610 (rd_5r0[26:26], df_0[26:26], rg_5r);
  AND2 I611 (rd_5r0[27:27], df_0[27:27], rg_5r);
  AND2 I612 (rd_5r0[28:28], df_0[28:28], rg_5r);
  AND2 I613 (rd_5r0[29:29], df_0[29:29], rg_5r);
  AND2 I614 (rd_5r0[30:30], df_0[30:30], rg_5r);
  AND2 I615 (rd_5r0[31:31], df_0[31:31], rg_5r);
  AND2 I616 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I617 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I618 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I619 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I620 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I621 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I622 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I623 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I624 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I625 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I626 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I627 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I628 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I629 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I630 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I631 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I632 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I633 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I634 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I635 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I636 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I637 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I638 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I639 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I640 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I641 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I642 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I643 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I644 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I645 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I646 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I647 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I648 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I649 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I650 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I651 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I652 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I653 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I654 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I655 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I656 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I657 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I658 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I659 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I660 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I661 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I662 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I663 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I664 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I665 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I666 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I667 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I668 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I669 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I670 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I671 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I672 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I673 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I674 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I675 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I676 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I677 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I678 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I679 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I680 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I681 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I682 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I683 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I684 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I685 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I686 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I687 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I688 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I689 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I690 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I691 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I692 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I693 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I694 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I695 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I696 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I697 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I698 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I699 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I700 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I701 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I702 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I703 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I704 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I705 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I706 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I707 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I708 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I709 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I710 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I711 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  AND2 I712 (rd_3r1[0:0], dt_0[0:0], rg_3r);
  AND2 I713 (rd_3r1[1:1], dt_0[1:1], rg_3r);
  AND2 I714 (rd_3r1[2:2], dt_0[2:2], rg_3r);
  AND2 I715 (rd_3r1[3:3], dt_0[3:3], rg_3r);
  AND2 I716 (rd_3r1[4:4], dt_0[4:4], rg_3r);
  AND2 I717 (rd_3r1[5:5], dt_0[5:5], rg_3r);
  AND2 I718 (rd_3r1[6:6], dt_0[6:6], rg_3r);
  AND2 I719 (rd_3r1[7:7], dt_0[7:7], rg_3r);
  AND2 I720 (rd_3r1[8:8], dt_0[8:8], rg_3r);
  AND2 I721 (rd_3r1[9:9], dt_0[9:9], rg_3r);
  AND2 I722 (rd_3r1[10:10], dt_0[10:10], rg_3r);
  AND2 I723 (rd_3r1[11:11], dt_0[11:11], rg_3r);
  AND2 I724 (rd_3r1[12:12], dt_0[12:12], rg_3r);
  AND2 I725 (rd_3r1[13:13], dt_0[13:13], rg_3r);
  AND2 I726 (rd_3r1[14:14], dt_0[14:14], rg_3r);
  AND2 I727 (rd_3r1[15:15], dt_0[15:15], rg_3r);
  AND2 I728 (rd_3r1[16:16], dt_0[16:16], rg_3r);
  AND2 I729 (rd_3r1[17:17], dt_0[17:17], rg_3r);
  AND2 I730 (rd_3r1[18:18], dt_0[18:18], rg_3r);
  AND2 I731 (rd_3r1[19:19], dt_0[19:19], rg_3r);
  AND2 I732 (rd_3r1[20:20], dt_0[20:20], rg_3r);
  AND2 I733 (rd_3r1[21:21], dt_0[21:21], rg_3r);
  AND2 I734 (rd_3r1[22:22], dt_0[22:22], rg_3r);
  AND2 I735 (rd_3r1[23:23], dt_0[23:23], rg_3r);
  AND2 I736 (rd_3r1[24:24], dt_0[24:24], rg_3r);
  AND2 I737 (rd_3r1[25:25], dt_0[25:25], rg_3r);
  AND2 I738 (rd_3r1[26:26], dt_0[26:26], rg_3r);
  AND2 I739 (rd_3r1[27:27], dt_0[27:27], rg_3r);
  AND2 I740 (rd_3r1[28:28], dt_0[28:28], rg_3r);
  AND2 I741 (rd_3r1[29:29], dt_0[29:29], rg_3r);
  AND2 I742 (rd_3r1[30:30], dt_0[30:30], rg_3r);
  AND2 I743 (rd_3r1[31:31], dt_0[31:31], rg_3r);
  AND2 I744 (rd_4r1[0:0], dt_0[0:0], rg_4r);
  AND2 I745 (rd_4r1[1:1], dt_0[1:1], rg_4r);
  AND2 I746 (rd_4r1[2:2], dt_0[2:2], rg_4r);
  AND2 I747 (rd_4r1[3:3], dt_0[3:3], rg_4r);
  AND2 I748 (rd_4r1[4:4], dt_0[4:4], rg_4r);
  AND2 I749 (rd_4r1[5:5], dt_0[5:5], rg_4r);
  AND2 I750 (rd_4r1[6:6], dt_0[6:6], rg_4r);
  AND2 I751 (rd_4r1[7:7], dt_0[7:7], rg_4r);
  AND2 I752 (rd_4r1[8:8], dt_0[8:8], rg_4r);
  AND2 I753 (rd_4r1[9:9], dt_0[9:9], rg_4r);
  AND2 I754 (rd_4r1[10:10], dt_0[10:10], rg_4r);
  AND2 I755 (rd_4r1[11:11], dt_0[11:11], rg_4r);
  AND2 I756 (rd_4r1[12:12], dt_0[12:12], rg_4r);
  AND2 I757 (rd_4r1[13:13], dt_0[13:13], rg_4r);
  AND2 I758 (rd_4r1[14:14], dt_0[14:14], rg_4r);
  AND2 I759 (rd_4r1[15:15], dt_0[15:15], rg_4r);
  AND2 I760 (rd_4r1[16:16], dt_0[16:16], rg_4r);
  AND2 I761 (rd_4r1[17:17], dt_0[17:17], rg_4r);
  AND2 I762 (rd_4r1[18:18], dt_0[18:18], rg_4r);
  AND2 I763 (rd_4r1[19:19], dt_0[19:19], rg_4r);
  AND2 I764 (rd_4r1[20:20], dt_0[20:20], rg_4r);
  AND2 I765 (rd_4r1[21:21], dt_0[21:21], rg_4r);
  AND2 I766 (rd_4r1[22:22], dt_0[22:22], rg_4r);
  AND2 I767 (rd_4r1[23:23], dt_0[23:23], rg_4r);
  AND2 I768 (rd_4r1[24:24], dt_0[24:24], rg_4r);
  AND2 I769 (rd_4r1[25:25], dt_0[25:25], rg_4r);
  AND2 I770 (rd_4r1[26:26], dt_0[26:26], rg_4r);
  AND2 I771 (rd_4r1[27:27], dt_0[27:27], rg_4r);
  AND2 I772 (rd_4r1[28:28], dt_0[28:28], rg_4r);
  AND2 I773 (rd_4r1[29:29], dt_0[29:29], rg_4r);
  AND2 I774 (rd_4r1[30:30], dt_0[30:30], rg_4r);
  AND2 I775 (rd_4r1[31:31], dt_0[31:31], rg_4r);
  AND2 I776 (rd_5r1[0:0], dt_0[0:0], rg_5r);
  AND2 I777 (rd_5r1[1:1], dt_0[1:1], rg_5r);
  AND2 I778 (rd_5r1[2:2], dt_0[2:2], rg_5r);
  AND2 I779 (rd_5r1[3:3], dt_0[3:3], rg_5r);
  AND2 I780 (rd_5r1[4:4], dt_0[4:4], rg_5r);
  AND2 I781 (rd_5r1[5:5], dt_0[5:5], rg_5r);
  AND2 I782 (rd_5r1[6:6], dt_0[6:6], rg_5r);
  AND2 I783 (rd_5r1[7:7], dt_0[7:7], rg_5r);
  AND2 I784 (rd_5r1[8:8], dt_0[8:8], rg_5r);
  AND2 I785 (rd_5r1[9:9], dt_0[9:9], rg_5r);
  AND2 I786 (rd_5r1[10:10], dt_0[10:10], rg_5r);
  AND2 I787 (rd_5r1[11:11], dt_0[11:11], rg_5r);
  AND2 I788 (rd_5r1[12:12], dt_0[12:12], rg_5r);
  AND2 I789 (rd_5r1[13:13], dt_0[13:13], rg_5r);
  AND2 I790 (rd_5r1[14:14], dt_0[14:14], rg_5r);
  AND2 I791 (rd_5r1[15:15], dt_0[15:15], rg_5r);
  AND2 I792 (rd_5r1[16:16], dt_0[16:16], rg_5r);
  AND2 I793 (rd_5r1[17:17], dt_0[17:17], rg_5r);
  AND2 I794 (rd_5r1[18:18], dt_0[18:18], rg_5r);
  AND2 I795 (rd_5r1[19:19], dt_0[19:19], rg_5r);
  AND2 I796 (rd_5r1[20:20], dt_0[20:20], rg_5r);
  AND2 I797 (rd_5r1[21:21], dt_0[21:21], rg_5r);
  AND2 I798 (rd_5r1[22:22], dt_0[22:22], rg_5r);
  AND2 I799 (rd_5r1[23:23], dt_0[23:23], rg_5r);
  AND2 I800 (rd_5r1[24:24], dt_0[24:24], rg_5r);
  AND2 I801 (rd_5r1[25:25], dt_0[25:25], rg_5r);
  AND2 I802 (rd_5r1[26:26], dt_0[26:26], rg_5r);
  AND2 I803 (rd_5r1[27:27], dt_0[27:27], rg_5r);
  AND2 I804 (rd_5r1[28:28], dt_0[28:28], rg_5r);
  AND2 I805 (rd_5r1[29:29], dt_0[29:29], rg_5r);
  AND2 I806 (rd_5r1[30:30], dt_0[30:30], rg_5r);
  AND2 I807 (rd_5r1[31:31], dt_0[31:31], rg_5r);
  NOR3 I808 (simp7921_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I809 (simp7921_0[1:1], rg_3r, rg_4r, rg_5r);
  NOR3 I810 (simp7921_0[2:2], rg_0a, rg_1a, rg_2a);
  NOR3 I811 (simp7921_0[3:3], rg_3a, rg_4a, rg_5a);
  NAND3 I812 (simp7922_0[0:0], simp7921_0[0:0], simp7921_0[1:1], simp7921_0[2:2]);
  INV I813 (simp7922_0[1:1], simp7921_0[3:3]);
  OR2 I814 (anyread_0, simp7922_0[0:0], simp7922_0[1:1]);
  BUFF I815 (wg_0a, wd_0a);
  BUFF I816 (rg_0a, rd_0a);
  BUFF I817 (rg_1a, rd_1a);
  BUFF I818 (rg_2a, rd_2a);
  BUFF I819 (rg_3a, rd_3a);
  BUFF I820 (rg_4a, rd_4a);
  BUFF I821 (rg_5a, rd_5a);
endmodule

// tkvlocals_31032_wo0w32_ro0w32o0w32o0w32 TeakV "locals[31:0]" 32 [] [0] [0,0,0] [Many [32],Many [0],M
//   any [0,0,0],Many [32,32,32]]
module tkvlocals_31032_wo0w32_ro0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp6001_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I521 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I522 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I523 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I524 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I525 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I526 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I527 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I528 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I529 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I530 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I531 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I532 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I533 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I534 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I535 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I536 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I537 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I538 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I539 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I540 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I541 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I542 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I543 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I544 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I545 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I546 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I547 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I548 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I549 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I550 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I551 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I552 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I553 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I554 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I555 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I556 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I557 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I558 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I559 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I560 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I561 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I562 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I563 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I564 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I565 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I566 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I567 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I568 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I569 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I570 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I571 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I572 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I573 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I574 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I575 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I576 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I577 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I578 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I579 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I580 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I581 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I582 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I583 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I608 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I609 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I610 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I611 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I612 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I613 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I614 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I615 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  NOR3 I616 (simp6001_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I617 (simp6001_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I618 (anyread_0, simp6001_0[0:0], simp6001_0[1:1]);
  BUFF I619 (wg_0a, wd_0a);
  BUFF I620 (rg_0a, rd_0a);
  BUFF I621 (rg_1a, rd_1a);
  BUFF I622 (rg_2a, rd_2a);
endmodule

// tkvlocals_633232_wo0w32_ro0w32o0w32o0w32 TeakV "locals[63:32]" 32 [] [0] [0,0,0] [Many [32],Many [0]
//   ,Many [0,0,0],Many [32,32,32]]
module tkvlocals_633232_wo0w32_ro0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp6001_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I521 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I522 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I523 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I524 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I525 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I526 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I527 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I528 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I529 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I530 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I531 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I532 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I533 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I534 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I535 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I536 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I537 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I538 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I539 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I540 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I541 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I542 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I543 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I544 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I545 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I546 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I547 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I548 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I549 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I550 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I551 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I552 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I553 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I554 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I555 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I556 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I557 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I558 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I559 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I560 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I561 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I562 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I563 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I564 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I565 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I566 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I567 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I568 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I569 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I570 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I571 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I572 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I573 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I574 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I575 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I576 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I577 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I578 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I579 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I580 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I581 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I582 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I583 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I608 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I609 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I610 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I611 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I612 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I613 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I614 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I615 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  NOR3 I616 (simp6001_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I617 (simp6001_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I618 (anyread_0, simp6001_0[0:0], simp6001_0[1:1]);
  BUFF I619 (wg_0a, wd_0a);
  BUFF I620 (rg_0a, rd_0a);
  BUFF I621 (rg_1a, rd_1a);
  BUFF I622 (rg_2a, rd_2a);
endmodule

// tkvlocals_956432_wo0w32_ro0w32o0w32o0w32 TeakV "locals[95:64]" 32 [] [0] [0,0,0] [Many [32],Many [0]
//   ,Many [0,0,0],Many [32,32,32]]
module tkvlocals_956432_wo0w32_ro0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp6001_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I521 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I522 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I523 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I524 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I525 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I526 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I527 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I528 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I529 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I530 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I531 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I532 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I533 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I534 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I535 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I536 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I537 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I538 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I539 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I540 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I541 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I542 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I543 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I544 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I545 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I546 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I547 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I548 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I549 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I550 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I551 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I552 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I553 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I554 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I555 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I556 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I557 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I558 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I559 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I560 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I561 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I562 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I563 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I564 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I565 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I566 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I567 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I568 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I569 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I570 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I571 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I572 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I573 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I574 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I575 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I576 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I577 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I578 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I579 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I580 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I581 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I582 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I583 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I608 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I609 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I610 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I611 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I612 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I613 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I614 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I615 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  NOR3 I616 (simp6001_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I617 (simp6001_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I618 (anyread_0, simp6001_0[0:0], simp6001_0[1:1]);
  BUFF I619 (wg_0a, wd_0a);
  BUFF I620 (rg_0a, rd_0a);
  BUFF I621 (rg_1a, rd_1a);
  BUFF I622 (rg_2a, rd_2a);
endmodule

// tkvlocals_1279632_wo0w32_ro0w32o0w32o0w32 TeakV "locals[127:96]" 32 [] [0] [0,0,0] [Many [32],Many [
//   0],Many [0,0,0],Many [32,32,32]]
module tkvlocals_1279632_wo0w32_ro0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp6001_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I521 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I522 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I523 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I524 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I525 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I526 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I527 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I528 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I529 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I530 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I531 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I532 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I533 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I534 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I535 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I536 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I537 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I538 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I539 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I540 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I541 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I542 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I543 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I544 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I545 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I546 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I547 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I548 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I549 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I550 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I551 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I552 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I553 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I554 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I555 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I556 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I557 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I558 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I559 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I560 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I561 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I562 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I563 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I564 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I565 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I566 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I567 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I568 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I569 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I570 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I571 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I572 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I573 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I574 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I575 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I576 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I577 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I578 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I579 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I580 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I581 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I582 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I583 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I608 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I609 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I610 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I611 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I612 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I613 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I614 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I615 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  NOR3 I616 (simp6001_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I617 (simp6001_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I618 (anyread_0, simp6001_0[0:0], simp6001_0[1:1]);
  BUFF I619 (wg_0a, wd_0a);
  BUFF I620 (rg_0a, rd_0a);
  BUFF I621 (rg_1a, rd_1a);
  BUFF I622 (rg_2a, rd_2a);
endmodule

// tkvlocals_15912832_wo0w32_ro0w32o0w32o0w32 TeakV "locals[159:128]" 32 [] [0] [0,0,0] [Many [32],Many
//    [0],Many [0,0,0],Many [32,32,32]]
module tkvlocals_15912832_wo0w32_ro0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp6001_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I521 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I522 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I523 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I524 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I525 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I526 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I527 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I528 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I529 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I530 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I531 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I532 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I533 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I534 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I535 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I536 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I537 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I538 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I539 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I540 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I541 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I542 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I543 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I544 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I545 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I546 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I547 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I548 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I549 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I550 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I551 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I552 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I553 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I554 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I555 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I556 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I557 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I558 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I559 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I560 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I561 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I562 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I563 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I564 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I565 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I566 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I567 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I568 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I569 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I570 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I571 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I572 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I573 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I574 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I575 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I576 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I577 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I578 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I579 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I580 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I581 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I582 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I583 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I608 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I609 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I610 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I611 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I612 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I613 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I614 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I615 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  NOR3 I616 (simp6001_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I617 (simp6001_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I618 (anyread_0, simp6001_0[0:0], simp6001_0[1:1]);
  BUFF I619 (wg_0a, wd_0a);
  BUFF I620 (rg_0a, rd_0a);
  BUFF I621 (rg_1a, rd_1a);
  BUFF I622 (rg_2a, rd_2a);
endmodule

// tkvlocals_19116032_wo0w32_ro0w32o0w32o0w32 TeakV "locals[191:160]" 32 [] [0] [0,0,0] [Many [32],Many
//    [0],Many [0,0,0],Many [32,32,32]]
module tkvlocals_19116032_wo0w32_ro0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp6001_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I521 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I522 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I523 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I524 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I525 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I526 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I527 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I528 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I529 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I530 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I531 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I532 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I533 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I534 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I535 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I536 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I537 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I538 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I539 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I540 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I541 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I542 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I543 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I544 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I545 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I546 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I547 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I548 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I549 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I550 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I551 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I552 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I553 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I554 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I555 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I556 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I557 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I558 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I559 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I560 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I561 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I562 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I563 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I564 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I565 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I566 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I567 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I568 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I569 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I570 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I571 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I572 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I573 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I574 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I575 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I576 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I577 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I578 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I579 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I580 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I581 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I582 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I583 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I608 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I609 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I610 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I611 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I612 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I613 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I614 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I615 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  NOR3 I616 (simp6001_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I617 (simp6001_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I618 (anyread_0, simp6001_0[0:0], simp6001_0[1:1]);
  BUFF I619 (wg_0a, wd_0a);
  BUFF I620 (rg_0a, rd_0a);
  BUFF I621 (rg_1a, rd_1a);
  BUFF I622 (rg_2a, rd_2a);
endmodule

// tkvlocals_22319232_wo0w32_ro0w32o0w32o0w32 TeakV "locals[223:192]" 32 [] [0] [0,0,0] [Many [32],Many
//    [0],Many [0,0,0],Many [32,32,32]]
module tkvlocals_22319232_wo0w32_ro0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp6001_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I521 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I522 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I523 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I524 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I525 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I526 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I527 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I528 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I529 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I530 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I531 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I532 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I533 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I534 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I535 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I536 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I537 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I538 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I539 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I540 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I541 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I542 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I543 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I544 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I545 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I546 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I547 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I548 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I549 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I550 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I551 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I552 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I553 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I554 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I555 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I556 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I557 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I558 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I559 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I560 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I561 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I562 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I563 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I564 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I565 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I566 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I567 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I568 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I569 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I570 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I571 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I572 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I573 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I574 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I575 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I576 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I577 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I578 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I579 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I580 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I581 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I582 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I583 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I608 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I609 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I610 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I611 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I612 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I613 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I614 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I615 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  NOR3 I616 (simp6001_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I617 (simp6001_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I618 (anyread_0, simp6001_0[0:0], simp6001_0[1:1]);
  BUFF I619 (wg_0a, wd_0a);
  BUFF I620 (rg_0a, rd_0a);
  BUFF I621 (rg_1a, rd_1a);
  BUFF I622 (rg_2a, rd_2a);
endmodule

// tkvlocals_25522432_wo0w32_ro0w32o0w32o0w32 TeakV "locals[255:224]" 32 [] [0] [0,0,0] [Many [32],Many
//    [0],Many [0,0,0],Many [32,32,32]]
module tkvlocals_25522432_wo0w32_ro0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp6001_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I521 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I522 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I523 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I524 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I525 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I526 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I527 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I528 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I529 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I530 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I531 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I532 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I533 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I534 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I535 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I536 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I537 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I538 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I539 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I540 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I541 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I542 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I543 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I544 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I545 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I546 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I547 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I548 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I549 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I550 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I551 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I552 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I553 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I554 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I555 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I556 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I557 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I558 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I559 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I560 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I561 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I562 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I563 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I564 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I565 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I566 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I567 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I568 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I569 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I570 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I571 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I572 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I573 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I574 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I575 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I576 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I577 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I578 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I579 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I580 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I581 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I582 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I583 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I608 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I609 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I610 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I611 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I612 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I613 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I614 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I615 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  NOR3 I616 (simp6001_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I617 (simp6001_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I618 (anyread_0, simp6001_0[0:0], simp6001_0[1:1]);
  BUFF I619 (wg_0a, wd_0a);
  BUFF I620 (rg_0a, rd_0a);
  BUFF I621 (rg_1a, rd_1a);
  BUFF I622 (rg_2a, rd_2a);
endmodule

// tkvglobals_31032_wo0w32_ro0w32o0w32o0w32 TeakV "globals[31:0]" 32 [] [0] [0,0,0] [Many [32],Many [0]
//   ,Many [0,0,0],Many [32,32,32]]
module tkvglobals_31032_wo0w32_ro0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp6001_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I521 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I522 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I523 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I524 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I525 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I526 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I527 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I528 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I529 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I530 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I531 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I532 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I533 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I534 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I535 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I536 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I537 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I538 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I539 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I540 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I541 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I542 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I543 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I544 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I545 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I546 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I547 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I548 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I549 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I550 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I551 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I552 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I553 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I554 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I555 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I556 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I557 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I558 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I559 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I560 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I561 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I562 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I563 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I564 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I565 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I566 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I567 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I568 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I569 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I570 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I571 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I572 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I573 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I574 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I575 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I576 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I577 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I578 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I579 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I580 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I581 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I582 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I583 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I608 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I609 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I610 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I611 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I612 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I613 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I614 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I615 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  NOR3 I616 (simp6001_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I617 (simp6001_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I618 (anyread_0, simp6001_0[0:0], simp6001_0[1:1]);
  BUFF I619 (wg_0a, wd_0a);
  BUFF I620 (rg_0a, rd_0a);
  BUFF I621 (rg_1a, rd_1a);
  BUFF I622 (rg_2a, rd_2a);
endmodule

// tkvglobals_633232_wo0w32_ro0w32o0w32o0w32 TeakV "globals[63:32]" 32 [] [0] [0,0,0] [Many [32],Many [
//   0],Many [0,0,0],Many [32,32,32]]
module tkvglobals_633232_wo0w32_ro0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp6001_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I521 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I522 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I523 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I524 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I525 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I526 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I527 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I528 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I529 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I530 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I531 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I532 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I533 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I534 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I535 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I536 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I537 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I538 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I539 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I540 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I541 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I542 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I543 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I544 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I545 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I546 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I547 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I548 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I549 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I550 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I551 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I552 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I553 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I554 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I555 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I556 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I557 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I558 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I559 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I560 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I561 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I562 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I563 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I564 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I565 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I566 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I567 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I568 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I569 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I570 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I571 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I572 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I573 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I574 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I575 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I576 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I577 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I578 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I579 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I580 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I581 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I582 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I583 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I608 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I609 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I610 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I611 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I612 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I613 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I614 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I615 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  NOR3 I616 (simp6001_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I617 (simp6001_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I618 (anyread_0, simp6001_0[0:0], simp6001_0[1:1]);
  BUFF I619 (wg_0a, wd_0a);
  BUFF I620 (rg_0a, rd_0a);
  BUFF I621 (rg_1a, rd_1a);
  BUFF I622 (rg_2a, rd_2a);
endmodule

// tkvglobals_956432_wo0w32_ro0w32o0w32o0w32 TeakV "globals[95:64]" 32 [] [0] [0,0,0] [Many [32],Many [
//   0],Many [0,0,0],Many [32,32,32]]
module tkvglobals_956432_wo0w32_ro0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp6001_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I521 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I522 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I523 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I524 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I525 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I526 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I527 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I528 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I529 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I530 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I531 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I532 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I533 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I534 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I535 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I536 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I537 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I538 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I539 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I540 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I541 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I542 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I543 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I544 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I545 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I546 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I547 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I548 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I549 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I550 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I551 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I552 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I553 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I554 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I555 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I556 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I557 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I558 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I559 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I560 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I561 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I562 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I563 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I564 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I565 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I566 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I567 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I568 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I569 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I570 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I571 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I572 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I573 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I574 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I575 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I576 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I577 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I578 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I579 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I580 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I581 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I582 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I583 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I608 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I609 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I610 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I611 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I612 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I613 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I614 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I615 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  NOR3 I616 (simp6001_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I617 (simp6001_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I618 (anyread_0, simp6001_0[0:0], simp6001_0[1:1]);
  BUFF I619 (wg_0a, wd_0a);
  BUFF I620 (rg_0a, rd_0a);
  BUFF I621 (rg_1a, rd_1a);
  BUFF I622 (rg_2a, rd_2a);
endmodule

// tkvglobals_1279632_wo0w32_ro0w32o0w32o0w32 TeakV "globals[127:96]" 32 [] [0] [0,0,0] [Many [32],Many
//    [0],Many [0,0,0],Many [32,32,32]]
module tkvglobals_1279632_wo0w32_ro0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp6001_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I521 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I522 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I523 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I524 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I525 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I526 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I527 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I528 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I529 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I530 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I531 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I532 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I533 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I534 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I535 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I536 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I537 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I538 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I539 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I540 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I541 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I542 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I543 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I544 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I545 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I546 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I547 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I548 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I549 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I550 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I551 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I552 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I553 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I554 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I555 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I556 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I557 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I558 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I559 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I560 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I561 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I562 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I563 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I564 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I565 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I566 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I567 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I568 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I569 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I570 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I571 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I572 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I573 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I574 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I575 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I576 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I577 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I578 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I579 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I580 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I581 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I582 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I583 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I608 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I609 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I610 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I611 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I612 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I613 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I614 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I615 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  NOR3 I616 (simp6001_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I617 (simp6001_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I618 (anyread_0, simp6001_0[0:0], simp6001_0[1:1]);
  BUFF I619 (wg_0a, wd_0a);
  BUFF I620 (rg_0a, rd_0a);
  BUFF I621 (rg_1a, rd_1a);
  BUFF I622 (rg_2a, rd_2a);
endmodule

// tkvglobals_15912832_wo0w32_ro0w32o0w32o0w32 TeakV "globals[159:128]" 32 [] [0] [0,0,0] [Many [32],Ma
//   ny [0],Many [0,0,0],Many [32,32,32]]
module tkvglobals_15912832_wo0w32_ro0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp6001_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I521 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I522 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I523 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I524 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I525 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I526 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I527 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I528 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I529 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I530 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I531 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I532 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I533 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I534 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I535 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I536 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I537 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I538 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I539 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I540 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I541 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I542 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I543 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I544 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I545 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I546 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I547 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I548 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I549 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I550 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I551 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I552 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I553 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I554 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I555 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I556 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I557 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I558 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I559 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I560 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I561 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I562 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I563 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I564 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I565 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I566 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I567 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I568 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I569 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I570 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I571 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I572 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I573 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I574 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I575 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I576 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I577 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I578 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I579 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I580 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I581 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I582 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I583 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I608 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I609 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I610 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I611 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I612 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I613 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I614 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I615 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  NOR3 I616 (simp6001_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I617 (simp6001_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I618 (anyread_0, simp6001_0[0:0], simp6001_0[1:1]);
  BUFF I619 (wg_0a, wd_0a);
  BUFF I620 (rg_0a, rd_0a);
  BUFF I621 (rg_1a, rd_1a);
  BUFF I622 (rg_2a, rd_2a);
endmodule

// tkvglobals_19116032_wo0w32_ro0w32o0w32o0w32 TeakV "globals[191:160]" 32 [] [0] [0,0,0] [Many [32],Ma
//   ny [0],Many [0,0,0],Many [32,32,32]]
module tkvglobals_19116032_wo0w32_ro0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp6001_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I521 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I522 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I523 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I524 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I525 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I526 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I527 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I528 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I529 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I530 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I531 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I532 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I533 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I534 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I535 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I536 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I537 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I538 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I539 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I540 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I541 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I542 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I543 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I544 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I545 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I546 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I547 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I548 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I549 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I550 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I551 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I552 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I553 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I554 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I555 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I556 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I557 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I558 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I559 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I560 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I561 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I562 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I563 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I564 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I565 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I566 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I567 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I568 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I569 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I570 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I571 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I572 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I573 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I574 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I575 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I576 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I577 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I578 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I579 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I580 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I581 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I582 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I583 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I608 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I609 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I610 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I611 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I612 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I613 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I614 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I615 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  NOR3 I616 (simp6001_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I617 (simp6001_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I618 (anyread_0, simp6001_0[0:0], simp6001_0[1:1]);
  BUFF I619 (wg_0a, wd_0a);
  BUFF I620 (rg_0a, rd_0a);
  BUFF I621 (rg_1a, rd_1a);
  BUFF I622 (rg_2a, rd_2a);
endmodule

// tkvglobals_22319232_wo0w32_ro0w32o0w32o0w32 TeakV "globals[223:192]" 32 [] [0] [0,0,0] [Many [32],Ma
//   ny [0],Many [0,0,0],Many [32,32,32]]
module tkvglobals_22319232_wo0w32_ro0w32o0w32o0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output [31:0] rd_1r0;
  output [31:0] rd_1r1;
  input rd_1a;
  output [31:0] rd_2r0;
  output [31:0] rd_2r1;
  input rd_2a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  wire [1:0] simp6001_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_1r0[0:0], df_0[0:0], rg_1r);
  AND2 I457 (rd_1r0[1:1], df_0[1:1], rg_1r);
  AND2 I458 (rd_1r0[2:2], df_0[2:2], rg_1r);
  AND2 I459 (rd_1r0[3:3], df_0[3:3], rg_1r);
  AND2 I460 (rd_1r0[4:4], df_0[4:4], rg_1r);
  AND2 I461 (rd_1r0[5:5], df_0[5:5], rg_1r);
  AND2 I462 (rd_1r0[6:6], df_0[6:6], rg_1r);
  AND2 I463 (rd_1r0[7:7], df_0[7:7], rg_1r);
  AND2 I464 (rd_1r0[8:8], df_0[8:8], rg_1r);
  AND2 I465 (rd_1r0[9:9], df_0[9:9], rg_1r);
  AND2 I466 (rd_1r0[10:10], df_0[10:10], rg_1r);
  AND2 I467 (rd_1r0[11:11], df_0[11:11], rg_1r);
  AND2 I468 (rd_1r0[12:12], df_0[12:12], rg_1r);
  AND2 I469 (rd_1r0[13:13], df_0[13:13], rg_1r);
  AND2 I470 (rd_1r0[14:14], df_0[14:14], rg_1r);
  AND2 I471 (rd_1r0[15:15], df_0[15:15], rg_1r);
  AND2 I472 (rd_1r0[16:16], df_0[16:16], rg_1r);
  AND2 I473 (rd_1r0[17:17], df_0[17:17], rg_1r);
  AND2 I474 (rd_1r0[18:18], df_0[18:18], rg_1r);
  AND2 I475 (rd_1r0[19:19], df_0[19:19], rg_1r);
  AND2 I476 (rd_1r0[20:20], df_0[20:20], rg_1r);
  AND2 I477 (rd_1r0[21:21], df_0[21:21], rg_1r);
  AND2 I478 (rd_1r0[22:22], df_0[22:22], rg_1r);
  AND2 I479 (rd_1r0[23:23], df_0[23:23], rg_1r);
  AND2 I480 (rd_1r0[24:24], df_0[24:24], rg_1r);
  AND2 I481 (rd_1r0[25:25], df_0[25:25], rg_1r);
  AND2 I482 (rd_1r0[26:26], df_0[26:26], rg_1r);
  AND2 I483 (rd_1r0[27:27], df_0[27:27], rg_1r);
  AND2 I484 (rd_1r0[28:28], df_0[28:28], rg_1r);
  AND2 I485 (rd_1r0[29:29], df_0[29:29], rg_1r);
  AND2 I486 (rd_1r0[30:30], df_0[30:30], rg_1r);
  AND2 I487 (rd_1r0[31:31], df_0[31:31], rg_1r);
  AND2 I488 (rd_2r0[0:0], df_0[0:0], rg_2r);
  AND2 I489 (rd_2r0[1:1], df_0[1:1], rg_2r);
  AND2 I490 (rd_2r0[2:2], df_0[2:2], rg_2r);
  AND2 I491 (rd_2r0[3:3], df_0[3:3], rg_2r);
  AND2 I492 (rd_2r0[4:4], df_0[4:4], rg_2r);
  AND2 I493 (rd_2r0[5:5], df_0[5:5], rg_2r);
  AND2 I494 (rd_2r0[6:6], df_0[6:6], rg_2r);
  AND2 I495 (rd_2r0[7:7], df_0[7:7], rg_2r);
  AND2 I496 (rd_2r0[8:8], df_0[8:8], rg_2r);
  AND2 I497 (rd_2r0[9:9], df_0[9:9], rg_2r);
  AND2 I498 (rd_2r0[10:10], df_0[10:10], rg_2r);
  AND2 I499 (rd_2r0[11:11], df_0[11:11], rg_2r);
  AND2 I500 (rd_2r0[12:12], df_0[12:12], rg_2r);
  AND2 I501 (rd_2r0[13:13], df_0[13:13], rg_2r);
  AND2 I502 (rd_2r0[14:14], df_0[14:14], rg_2r);
  AND2 I503 (rd_2r0[15:15], df_0[15:15], rg_2r);
  AND2 I504 (rd_2r0[16:16], df_0[16:16], rg_2r);
  AND2 I505 (rd_2r0[17:17], df_0[17:17], rg_2r);
  AND2 I506 (rd_2r0[18:18], df_0[18:18], rg_2r);
  AND2 I507 (rd_2r0[19:19], df_0[19:19], rg_2r);
  AND2 I508 (rd_2r0[20:20], df_0[20:20], rg_2r);
  AND2 I509 (rd_2r0[21:21], df_0[21:21], rg_2r);
  AND2 I510 (rd_2r0[22:22], df_0[22:22], rg_2r);
  AND2 I511 (rd_2r0[23:23], df_0[23:23], rg_2r);
  AND2 I512 (rd_2r0[24:24], df_0[24:24], rg_2r);
  AND2 I513 (rd_2r0[25:25], df_0[25:25], rg_2r);
  AND2 I514 (rd_2r0[26:26], df_0[26:26], rg_2r);
  AND2 I515 (rd_2r0[27:27], df_0[27:27], rg_2r);
  AND2 I516 (rd_2r0[28:28], df_0[28:28], rg_2r);
  AND2 I517 (rd_2r0[29:29], df_0[29:29], rg_2r);
  AND2 I518 (rd_2r0[30:30], df_0[30:30], rg_2r);
  AND2 I519 (rd_2r0[31:31], df_0[31:31], rg_2r);
  AND2 I520 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I521 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I522 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I523 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I524 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I525 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I526 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I527 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I528 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I529 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I530 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I531 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I532 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I533 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I534 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I535 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I536 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I537 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I538 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I539 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I540 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I541 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I542 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I543 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I544 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I545 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I546 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I547 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I548 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I549 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I550 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I551 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I552 (rd_1r1[0:0], dt_0[0:0], rg_1r);
  AND2 I553 (rd_1r1[1:1], dt_0[1:1], rg_1r);
  AND2 I554 (rd_1r1[2:2], dt_0[2:2], rg_1r);
  AND2 I555 (rd_1r1[3:3], dt_0[3:3], rg_1r);
  AND2 I556 (rd_1r1[4:4], dt_0[4:4], rg_1r);
  AND2 I557 (rd_1r1[5:5], dt_0[5:5], rg_1r);
  AND2 I558 (rd_1r1[6:6], dt_0[6:6], rg_1r);
  AND2 I559 (rd_1r1[7:7], dt_0[7:7], rg_1r);
  AND2 I560 (rd_1r1[8:8], dt_0[8:8], rg_1r);
  AND2 I561 (rd_1r1[9:9], dt_0[9:9], rg_1r);
  AND2 I562 (rd_1r1[10:10], dt_0[10:10], rg_1r);
  AND2 I563 (rd_1r1[11:11], dt_0[11:11], rg_1r);
  AND2 I564 (rd_1r1[12:12], dt_0[12:12], rg_1r);
  AND2 I565 (rd_1r1[13:13], dt_0[13:13], rg_1r);
  AND2 I566 (rd_1r1[14:14], dt_0[14:14], rg_1r);
  AND2 I567 (rd_1r1[15:15], dt_0[15:15], rg_1r);
  AND2 I568 (rd_1r1[16:16], dt_0[16:16], rg_1r);
  AND2 I569 (rd_1r1[17:17], dt_0[17:17], rg_1r);
  AND2 I570 (rd_1r1[18:18], dt_0[18:18], rg_1r);
  AND2 I571 (rd_1r1[19:19], dt_0[19:19], rg_1r);
  AND2 I572 (rd_1r1[20:20], dt_0[20:20], rg_1r);
  AND2 I573 (rd_1r1[21:21], dt_0[21:21], rg_1r);
  AND2 I574 (rd_1r1[22:22], dt_0[22:22], rg_1r);
  AND2 I575 (rd_1r1[23:23], dt_0[23:23], rg_1r);
  AND2 I576 (rd_1r1[24:24], dt_0[24:24], rg_1r);
  AND2 I577 (rd_1r1[25:25], dt_0[25:25], rg_1r);
  AND2 I578 (rd_1r1[26:26], dt_0[26:26], rg_1r);
  AND2 I579 (rd_1r1[27:27], dt_0[27:27], rg_1r);
  AND2 I580 (rd_1r1[28:28], dt_0[28:28], rg_1r);
  AND2 I581 (rd_1r1[29:29], dt_0[29:29], rg_1r);
  AND2 I582 (rd_1r1[30:30], dt_0[30:30], rg_1r);
  AND2 I583 (rd_1r1[31:31], dt_0[31:31], rg_1r);
  AND2 I584 (rd_2r1[0:0], dt_0[0:0], rg_2r);
  AND2 I585 (rd_2r1[1:1], dt_0[1:1], rg_2r);
  AND2 I586 (rd_2r1[2:2], dt_0[2:2], rg_2r);
  AND2 I587 (rd_2r1[3:3], dt_0[3:3], rg_2r);
  AND2 I588 (rd_2r1[4:4], dt_0[4:4], rg_2r);
  AND2 I589 (rd_2r1[5:5], dt_0[5:5], rg_2r);
  AND2 I590 (rd_2r1[6:6], dt_0[6:6], rg_2r);
  AND2 I591 (rd_2r1[7:7], dt_0[7:7], rg_2r);
  AND2 I592 (rd_2r1[8:8], dt_0[8:8], rg_2r);
  AND2 I593 (rd_2r1[9:9], dt_0[9:9], rg_2r);
  AND2 I594 (rd_2r1[10:10], dt_0[10:10], rg_2r);
  AND2 I595 (rd_2r1[11:11], dt_0[11:11], rg_2r);
  AND2 I596 (rd_2r1[12:12], dt_0[12:12], rg_2r);
  AND2 I597 (rd_2r1[13:13], dt_0[13:13], rg_2r);
  AND2 I598 (rd_2r1[14:14], dt_0[14:14], rg_2r);
  AND2 I599 (rd_2r1[15:15], dt_0[15:15], rg_2r);
  AND2 I600 (rd_2r1[16:16], dt_0[16:16], rg_2r);
  AND2 I601 (rd_2r1[17:17], dt_0[17:17], rg_2r);
  AND2 I602 (rd_2r1[18:18], dt_0[18:18], rg_2r);
  AND2 I603 (rd_2r1[19:19], dt_0[19:19], rg_2r);
  AND2 I604 (rd_2r1[20:20], dt_0[20:20], rg_2r);
  AND2 I605 (rd_2r1[21:21], dt_0[21:21], rg_2r);
  AND2 I606 (rd_2r1[22:22], dt_0[22:22], rg_2r);
  AND2 I607 (rd_2r1[23:23], dt_0[23:23], rg_2r);
  AND2 I608 (rd_2r1[24:24], dt_0[24:24], rg_2r);
  AND2 I609 (rd_2r1[25:25], dt_0[25:25], rg_2r);
  AND2 I610 (rd_2r1[26:26], dt_0[26:26], rg_2r);
  AND2 I611 (rd_2r1[27:27], dt_0[27:27], rg_2r);
  AND2 I612 (rd_2r1[28:28], dt_0[28:28], rg_2r);
  AND2 I613 (rd_2r1[29:29], dt_0[29:29], rg_2r);
  AND2 I614 (rd_2r1[30:30], dt_0[30:30], rg_2r);
  AND2 I615 (rd_2r1[31:31], dt_0[31:31], rg_2r);
  NOR3 I616 (simp6001_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I617 (simp6001_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I618 (anyread_0, simp6001_0[0:0], simp6001_0[1:1]);
  BUFF I619 (wg_0a, wd_0a);
  BUFF I620 (rg_0a, rd_0a);
  BUFF I621 (rg_1a, rd_1a);
  BUFF I622 (rg_2a, rd_2a);
endmodule

// tkm5x32b TeakM [Many [32,32,32,32,32],One 32]
module tkm5x32b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, i_4r0, i_4r1, i_4a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [31:0] i_1r0;
  input [31:0] i_1r1;
  output i_1a;
  input [31:0] i_2r0;
  input [31:0] i_2r1;
  output i_2a;
  input [31:0] i_3r0;
  input [31:0] i_3r1;
  output i_3a;
  input [31:0] i_4r0;
  input [31:0] i_4r1;
  output i_4a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  input reset;
  wire [31:0] gfint_0;
  wire [31:0] gfint_1;
  wire [31:0] gfint_2;
  wire [31:0] gfint_3;
  wire [31:0] gfint_4;
  wire [31:0] gtint_0;
  wire [31:0] gtint_1;
  wire [31:0] gtint_2;
  wire [31:0] gtint_3;
  wire [31:0] gtint_4;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire choice_4;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire icomp_3;
  wire icomp_4;
  wire nchosen_0;
  wire [1:0] simp221_0;
  wire [1:0] simp231_0;
  wire [1:0] simp241_0;
  wire [1:0] simp251_0;
  wire [1:0] simp261_0;
  wire [1:0] simp271_0;
  wire [1:0] simp281_0;
  wire [1:0] simp291_0;
  wire [1:0] simp301_0;
  wire [1:0] simp311_0;
  wire [1:0] simp321_0;
  wire [1:0] simp331_0;
  wire [1:0] simp341_0;
  wire [1:0] simp351_0;
  wire [1:0] simp361_0;
  wire [1:0] simp371_0;
  wire [1:0] simp381_0;
  wire [1:0] simp391_0;
  wire [1:0] simp401_0;
  wire [1:0] simp411_0;
  wire [1:0] simp421_0;
  wire [1:0] simp431_0;
  wire [1:0] simp441_0;
  wire [1:0] simp451_0;
  wire [1:0] simp461_0;
  wire [1:0] simp471_0;
  wire [1:0] simp481_0;
  wire [1:0] simp491_0;
  wire [1:0] simp501_0;
  wire [1:0] simp511_0;
  wire [1:0] simp521_0;
  wire [1:0] simp531_0;
  wire [1:0] simp541_0;
  wire [1:0] simp551_0;
  wire [1:0] simp561_0;
  wire [1:0] simp571_0;
  wire [1:0] simp581_0;
  wire [1:0] simp591_0;
  wire [1:0] simp601_0;
  wire [1:0] simp611_0;
  wire [1:0] simp621_0;
  wire [1:0] simp631_0;
  wire [1:0] simp641_0;
  wire [1:0] simp651_0;
  wire [1:0] simp661_0;
  wire [1:0] simp671_0;
  wire [1:0] simp681_0;
  wire [1:0] simp691_0;
  wire [1:0] simp701_0;
  wire [1:0] simp711_0;
  wire [1:0] simp721_0;
  wire [1:0] simp731_0;
  wire [1:0] simp741_0;
  wire [1:0] simp751_0;
  wire [1:0] simp761_0;
  wire [1:0] simp771_0;
  wire [1:0] simp781_0;
  wire [1:0] simp791_0;
  wire [1:0] simp801_0;
  wire [1:0] simp811_0;
  wire [1:0] simp821_0;
  wire [1:0] simp831_0;
  wire [1:0] simp841_0;
  wire [1:0] simp851_0;
  wire [31:0] comp0_0;
  wire [10:0] simp4391_0;
  wire [3:0] simp4392_0;
  wire [1:0] simp4393_0;
  wire [31:0] comp1_0;
  wire [10:0] simp4731_0;
  wire [3:0] simp4732_0;
  wire [1:0] simp4733_0;
  wire [31:0] comp2_0;
  wire [10:0] simp5071_0;
  wire [3:0] simp5072_0;
  wire [1:0] simp5073_0;
  wire [31:0] comp3_0;
  wire [10:0] simp5411_0;
  wire [3:0] simp5412_0;
  wire [1:0] simp5413_0;
  wire [31:0] comp4_0;
  wire [10:0] simp5751_0;
  wire [3:0] simp5752_0;
  wire [1:0] simp5753_0;
  wire [1:0] simp5811_0;
  NOR3 I0 (simp221_0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  NOR2 I1 (simp221_0[1:1], gfint_3[0:0], gfint_4[0:0]);
  NAND2 I2 (o_0r0[0:0], simp221_0[0:0], simp221_0[1:1]);
  NOR3 I3 (simp231_0[0:0], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  NOR2 I4 (simp231_0[1:1], gfint_3[1:1], gfint_4[1:1]);
  NAND2 I5 (o_0r0[1:1], simp231_0[0:0], simp231_0[1:1]);
  NOR3 I6 (simp241_0[0:0], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  NOR2 I7 (simp241_0[1:1], gfint_3[2:2], gfint_4[2:2]);
  NAND2 I8 (o_0r0[2:2], simp241_0[0:0], simp241_0[1:1]);
  NOR3 I9 (simp251_0[0:0], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  NOR2 I10 (simp251_0[1:1], gfint_3[3:3], gfint_4[3:3]);
  NAND2 I11 (o_0r0[3:3], simp251_0[0:0], simp251_0[1:1]);
  NOR3 I12 (simp261_0[0:0], gfint_0[4:4], gfint_1[4:4], gfint_2[4:4]);
  NOR2 I13 (simp261_0[1:1], gfint_3[4:4], gfint_4[4:4]);
  NAND2 I14 (o_0r0[4:4], simp261_0[0:0], simp261_0[1:1]);
  NOR3 I15 (simp271_0[0:0], gfint_0[5:5], gfint_1[5:5], gfint_2[5:5]);
  NOR2 I16 (simp271_0[1:1], gfint_3[5:5], gfint_4[5:5]);
  NAND2 I17 (o_0r0[5:5], simp271_0[0:0], simp271_0[1:1]);
  NOR3 I18 (simp281_0[0:0], gfint_0[6:6], gfint_1[6:6], gfint_2[6:6]);
  NOR2 I19 (simp281_0[1:1], gfint_3[6:6], gfint_4[6:6]);
  NAND2 I20 (o_0r0[6:6], simp281_0[0:0], simp281_0[1:1]);
  NOR3 I21 (simp291_0[0:0], gfint_0[7:7], gfint_1[7:7], gfint_2[7:7]);
  NOR2 I22 (simp291_0[1:1], gfint_3[7:7], gfint_4[7:7]);
  NAND2 I23 (o_0r0[7:7], simp291_0[0:0], simp291_0[1:1]);
  NOR3 I24 (simp301_0[0:0], gfint_0[8:8], gfint_1[8:8], gfint_2[8:8]);
  NOR2 I25 (simp301_0[1:1], gfint_3[8:8], gfint_4[8:8]);
  NAND2 I26 (o_0r0[8:8], simp301_0[0:0], simp301_0[1:1]);
  NOR3 I27 (simp311_0[0:0], gfint_0[9:9], gfint_1[9:9], gfint_2[9:9]);
  NOR2 I28 (simp311_0[1:1], gfint_3[9:9], gfint_4[9:9]);
  NAND2 I29 (o_0r0[9:9], simp311_0[0:0], simp311_0[1:1]);
  NOR3 I30 (simp321_0[0:0], gfint_0[10:10], gfint_1[10:10], gfint_2[10:10]);
  NOR2 I31 (simp321_0[1:1], gfint_3[10:10], gfint_4[10:10]);
  NAND2 I32 (o_0r0[10:10], simp321_0[0:0], simp321_0[1:1]);
  NOR3 I33 (simp331_0[0:0], gfint_0[11:11], gfint_1[11:11], gfint_2[11:11]);
  NOR2 I34 (simp331_0[1:1], gfint_3[11:11], gfint_4[11:11]);
  NAND2 I35 (o_0r0[11:11], simp331_0[0:0], simp331_0[1:1]);
  NOR3 I36 (simp341_0[0:0], gfint_0[12:12], gfint_1[12:12], gfint_2[12:12]);
  NOR2 I37 (simp341_0[1:1], gfint_3[12:12], gfint_4[12:12]);
  NAND2 I38 (o_0r0[12:12], simp341_0[0:0], simp341_0[1:1]);
  NOR3 I39 (simp351_0[0:0], gfint_0[13:13], gfint_1[13:13], gfint_2[13:13]);
  NOR2 I40 (simp351_0[1:1], gfint_3[13:13], gfint_4[13:13]);
  NAND2 I41 (o_0r0[13:13], simp351_0[0:0], simp351_0[1:1]);
  NOR3 I42 (simp361_0[0:0], gfint_0[14:14], gfint_1[14:14], gfint_2[14:14]);
  NOR2 I43 (simp361_0[1:1], gfint_3[14:14], gfint_4[14:14]);
  NAND2 I44 (o_0r0[14:14], simp361_0[0:0], simp361_0[1:1]);
  NOR3 I45 (simp371_0[0:0], gfint_0[15:15], gfint_1[15:15], gfint_2[15:15]);
  NOR2 I46 (simp371_0[1:1], gfint_3[15:15], gfint_4[15:15]);
  NAND2 I47 (o_0r0[15:15], simp371_0[0:0], simp371_0[1:1]);
  NOR3 I48 (simp381_0[0:0], gfint_0[16:16], gfint_1[16:16], gfint_2[16:16]);
  NOR2 I49 (simp381_0[1:1], gfint_3[16:16], gfint_4[16:16]);
  NAND2 I50 (o_0r0[16:16], simp381_0[0:0], simp381_0[1:1]);
  NOR3 I51 (simp391_0[0:0], gfint_0[17:17], gfint_1[17:17], gfint_2[17:17]);
  NOR2 I52 (simp391_0[1:1], gfint_3[17:17], gfint_4[17:17]);
  NAND2 I53 (o_0r0[17:17], simp391_0[0:0], simp391_0[1:1]);
  NOR3 I54 (simp401_0[0:0], gfint_0[18:18], gfint_1[18:18], gfint_2[18:18]);
  NOR2 I55 (simp401_0[1:1], gfint_3[18:18], gfint_4[18:18]);
  NAND2 I56 (o_0r0[18:18], simp401_0[0:0], simp401_0[1:1]);
  NOR3 I57 (simp411_0[0:0], gfint_0[19:19], gfint_1[19:19], gfint_2[19:19]);
  NOR2 I58 (simp411_0[1:1], gfint_3[19:19], gfint_4[19:19]);
  NAND2 I59 (o_0r0[19:19], simp411_0[0:0], simp411_0[1:1]);
  NOR3 I60 (simp421_0[0:0], gfint_0[20:20], gfint_1[20:20], gfint_2[20:20]);
  NOR2 I61 (simp421_0[1:1], gfint_3[20:20], gfint_4[20:20]);
  NAND2 I62 (o_0r0[20:20], simp421_0[0:0], simp421_0[1:1]);
  NOR3 I63 (simp431_0[0:0], gfint_0[21:21], gfint_1[21:21], gfint_2[21:21]);
  NOR2 I64 (simp431_0[1:1], gfint_3[21:21], gfint_4[21:21]);
  NAND2 I65 (o_0r0[21:21], simp431_0[0:0], simp431_0[1:1]);
  NOR3 I66 (simp441_0[0:0], gfint_0[22:22], gfint_1[22:22], gfint_2[22:22]);
  NOR2 I67 (simp441_0[1:1], gfint_3[22:22], gfint_4[22:22]);
  NAND2 I68 (o_0r0[22:22], simp441_0[0:0], simp441_0[1:1]);
  NOR3 I69 (simp451_0[0:0], gfint_0[23:23], gfint_1[23:23], gfint_2[23:23]);
  NOR2 I70 (simp451_0[1:1], gfint_3[23:23], gfint_4[23:23]);
  NAND2 I71 (o_0r0[23:23], simp451_0[0:0], simp451_0[1:1]);
  NOR3 I72 (simp461_0[0:0], gfint_0[24:24], gfint_1[24:24], gfint_2[24:24]);
  NOR2 I73 (simp461_0[1:1], gfint_3[24:24], gfint_4[24:24]);
  NAND2 I74 (o_0r0[24:24], simp461_0[0:0], simp461_0[1:1]);
  NOR3 I75 (simp471_0[0:0], gfint_0[25:25], gfint_1[25:25], gfint_2[25:25]);
  NOR2 I76 (simp471_0[1:1], gfint_3[25:25], gfint_4[25:25]);
  NAND2 I77 (o_0r0[25:25], simp471_0[0:0], simp471_0[1:1]);
  NOR3 I78 (simp481_0[0:0], gfint_0[26:26], gfint_1[26:26], gfint_2[26:26]);
  NOR2 I79 (simp481_0[1:1], gfint_3[26:26], gfint_4[26:26]);
  NAND2 I80 (o_0r0[26:26], simp481_0[0:0], simp481_0[1:1]);
  NOR3 I81 (simp491_0[0:0], gfint_0[27:27], gfint_1[27:27], gfint_2[27:27]);
  NOR2 I82 (simp491_0[1:1], gfint_3[27:27], gfint_4[27:27]);
  NAND2 I83 (o_0r0[27:27], simp491_0[0:0], simp491_0[1:1]);
  NOR3 I84 (simp501_0[0:0], gfint_0[28:28], gfint_1[28:28], gfint_2[28:28]);
  NOR2 I85 (simp501_0[1:1], gfint_3[28:28], gfint_4[28:28]);
  NAND2 I86 (o_0r0[28:28], simp501_0[0:0], simp501_0[1:1]);
  NOR3 I87 (simp511_0[0:0], gfint_0[29:29], gfint_1[29:29], gfint_2[29:29]);
  NOR2 I88 (simp511_0[1:1], gfint_3[29:29], gfint_4[29:29]);
  NAND2 I89 (o_0r0[29:29], simp511_0[0:0], simp511_0[1:1]);
  NOR3 I90 (simp521_0[0:0], gfint_0[30:30], gfint_1[30:30], gfint_2[30:30]);
  NOR2 I91 (simp521_0[1:1], gfint_3[30:30], gfint_4[30:30]);
  NAND2 I92 (o_0r0[30:30], simp521_0[0:0], simp521_0[1:1]);
  NOR3 I93 (simp531_0[0:0], gfint_0[31:31], gfint_1[31:31], gfint_2[31:31]);
  NOR2 I94 (simp531_0[1:1], gfint_3[31:31], gfint_4[31:31]);
  NAND2 I95 (o_0r0[31:31], simp531_0[0:0], simp531_0[1:1]);
  NOR3 I96 (simp541_0[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  NOR2 I97 (simp541_0[1:1], gtint_3[0:0], gtint_4[0:0]);
  NAND2 I98 (o_0r1[0:0], simp541_0[0:0], simp541_0[1:1]);
  NOR3 I99 (simp551_0[0:0], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  NOR2 I100 (simp551_0[1:1], gtint_3[1:1], gtint_4[1:1]);
  NAND2 I101 (o_0r1[1:1], simp551_0[0:0], simp551_0[1:1]);
  NOR3 I102 (simp561_0[0:0], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  NOR2 I103 (simp561_0[1:1], gtint_3[2:2], gtint_4[2:2]);
  NAND2 I104 (o_0r1[2:2], simp561_0[0:0], simp561_0[1:1]);
  NOR3 I105 (simp571_0[0:0], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  NOR2 I106 (simp571_0[1:1], gtint_3[3:3], gtint_4[3:3]);
  NAND2 I107 (o_0r1[3:3], simp571_0[0:0], simp571_0[1:1]);
  NOR3 I108 (simp581_0[0:0], gtint_0[4:4], gtint_1[4:4], gtint_2[4:4]);
  NOR2 I109 (simp581_0[1:1], gtint_3[4:4], gtint_4[4:4]);
  NAND2 I110 (o_0r1[4:4], simp581_0[0:0], simp581_0[1:1]);
  NOR3 I111 (simp591_0[0:0], gtint_0[5:5], gtint_1[5:5], gtint_2[5:5]);
  NOR2 I112 (simp591_0[1:1], gtint_3[5:5], gtint_4[5:5]);
  NAND2 I113 (o_0r1[5:5], simp591_0[0:0], simp591_0[1:1]);
  NOR3 I114 (simp601_0[0:0], gtint_0[6:6], gtint_1[6:6], gtint_2[6:6]);
  NOR2 I115 (simp601_0[1:1], gtint_3[6:6], gtint_4[6:6]);
  NAND2 I116 (o_0r1[6:6], simp601_0[0:0], simp601_0[1:1]);
  NOR3 I117 (simp611_0[0:0], gtint_0[7:7], gtint_1[7:7], gtint_2[7:7]);
  NOR2 I118 (simp611_0[1:1], gtint_3[7:7], gtint_4[7:7]);
  NAND2 I119 (o_0r1[7:7], simp611_0[0:0], simp611_0[1:1]);
  NOR3 I120 (simp621_0[0:0], gtint_0[8:8], gtint_1[8:8], gtint_2[8:8]);
  NOR2 I121 (simp621_0[1:1], gtint_3[8:8], gtint_4[8:8]);
  NAND2 I122 (o_0r1[8:8], simp621_0[0:0], simp621_0[1:1]);
  NOR3 I123 (simp631_0[0:0], gtint_0[9:9], gtint_1[9:9], gtint_2[9:9]);
  NOR2 I124 (simp631_0[1:1], gtint_3[9:9], gtint_4[9:9]);
  NAND2 I125 (o_0r1[9:9], simp631_0[0:0], simp631_0[1:1]);
  NOR3 I126 (simp641_0[0:0], gtint_0[10:10], gtint_1[10:10], gtint_2[10:10]);
  NOR2 I127 (simp641_0[1:1], gtint_3[10:10], gtint_4[10:10]);
  NAND2 I128 (o_0r1[10:10], simp641_0[0:0], simp641_0[1:1]);
  NOR3 I129 (simp651_0[0:0], gtint_0[11:11], gtint_1[11:11], gtint_2[11:11]);
  NOR2 I130 (simp651_0[1:1], gtint_3[11:11], gtint_4[11:11]);
  NAND2 I131 (o_0r1[11:11], simp651_0[0:0], simp651_0[1:1]);
  NOR3 I132 (simp661_0[0:0], gtint_0[12:12], gtint_1[12:12], gtint_2[12:12]);
  NOR2 I133 (simp661_0[1:1], gtint_3[12:12], gtint_4[12:12]);
  NAND2 I134 (o_0r1[12:12], simp661_0[0:0], simp661_0[1:1]);
  NOR3 I135 (simp671_0[0:0], gtint_0[13:13], gtint_1[13:13], gtint_2[13:13]);
  NOR2 I136 (simp671_0[1:1], gtint_3[13:13], gtint_4[13:13]);
  NAND2 I137 (o_0r1[13:13], simp671_0[0:0], simp671_0[1:1]);
  NOR3 I138 (simp681_0[0:0], gtint_0[14:14], gtint_1[14:14], gtint_2[14:14]);
  NOR2 I139 (simp681_0[1:1], gtint_3[14:14], gtint_4[14:14]);
  NAND2 I140 (o_0r1[14:14], simp681_0[0:0], simp681_0[1:1]);
  NOR3 I141 (simp691_0[0:0], gtint_0[15:15], gtint_1[15:15], gtint_2[15:15]);
  NOR2 I142 (simp691_0[1:1], gtint_3[15:15], gtint_4[15:15]);
  NAND2 I143 (o_0r1[15:15], simp691_0[0:0], simp691_0[1:1]);
  NOR3 I144 (simp701_0[0:0], gtint_0[16:16], gtint_1[16:16], gtint_2[16:16]);
  NOR2 I145 (simp701_0[1:1], gtint_3[16:16], gtint_4[16:16]);
  NAND2 I146 (o_0r1[16:16], simp701_0[0:0], simp701_0[1:1]);
  NOR3 I147 (simp711_0[0:0], gtint_0[17:17], gtint_1[17:17], gtint_2[17:17]);
  NOR2 I148 (simp711_0[1:1], gtint_3[17:17], gtint_4[17:17]);
  NAND2 I149 (o_0r1[17:17], simp711_0[0:0], simp711_0[1:1]);
  NOR3 I150 (simp721_0[0:0], gtint_0[18:18], gtint_1[18:18], gtint_2[18:18]);
  NOR2 I151 (simp721_0[1:1], gtint_3[18:18], gtint_4[18:18]);
  NAND2 I152 (o_0r1[18:18], simp721_0[0:0], simp721_0[1:1]);
  NOR3 I153 (simp731_0[0:0], gtint_0[19:19], gtint_1[19:19], gtint_2[19:19]);
  NOR2 I154 (simp731_0[1:1], gtint_3[19:19], gtint_4[19:19]);
  NAND2 I155 (o_0r1[19:19], simp731_0[0:0], simp731_0[1:1]);
  NOR3 I156 (simp741_0[0:0], gtint_0[20:20], gtint_1[20:20], gtint_2[20:20]);
  NOR2 I157 (simp741_0[1:1], gtint_3[20:20], gtint_4[20:20]);
  NAND2 I158 (o_0r1[20:20], simp741_0[0:0], simp741_0[1:1]);
  NOR3 I159 (simp751_0[0:0], gtint_0[21:21], gtint_1[21:21], gtint_2[21:21]);
  NOR2 I160 (simp751_0[1:1], gtint_3[21:21], gtint_4[21:21]);
  NAND2 I161 (o_0r1[21:21], simp751_0[0:0], simp751_0[1:1]);
  NOR3 I162 (simp761_0[0:0], gtint_0[22:22], gtint_1[22:22], gtint_2[22:22]);
  NOR2 I163 (simp761_0[1:1], gtint_3[22:22], gtint_4[22:22]);
  NAND2 I164 (o_0r1[22:22], simp761_0[0:0], simp761_0[1:1]);
  NOR3 I165 (simp771_0[0:0], gtint_0[23:23], gtint_1[23:23], gtint_2[23:23]);
  NOR2 I166 (simp771_0[1:1], gtint_3[23:23], gtint_4[23:23]);
  NAND2 I167 (o_0r1[23:23], simp771_0[0:0], simp771_0[1:1]);
  NOR3 I168 (simp781_0[0:0], gtint_0[24:24], gtint_1[24:24], gtint_2[24:24]);
  NOR2 I169 (simp781_0[1:1], gtint_3[24:24], gtint_4[24:24]);
  NAND2 I170 (o_0r1[24:24], simp781_0[0:0], simp781_0[1:1]);
  NOR3 I171 (simp791_0[0:0], gtint_0[25:25], gtint_1[25:25], gtint_2[25:25]);
  NOR2 I172 (simp791_0[1:1], gtint_3[25:25], gtint_4[25:25]);
  NAND2 I173 (o_0r1[25:25], simp791_0[0:0], simp791_0[1:1]);
  NOR3 I174 (simp801_0[0:0], gtint_0[26:26], gtint_1[26:26], gtint_2[26:26]);
  NOR2 I175 (simp801_0[1:1], gtint_3[26:26], gtint_4[26:26]);
  NAND2 I176 (o_0r1[26:26], simp801_0[0:0], simp801_0[1:1]);
  NOR3 I177 (simp811_0[0:0], gtint_0[27:27], gtint_1[27:27], gtint_2[27:27]);
  NOR2 I178 (simp811_0[1:1], gtint_3[27:27], gtint_4[27:27]);
  NAND2 I179 (o_0r1[27:27], simp811_0[0:0], simp811_0[1:1]);
  NOR3 I180 (simp821_0[0:0], gtint_0[28:28], gtint_1[28:28], gtint_2[28:28]);
  NOR2 I181 (simp821_0[1:1], gtint_3[28:28], gtint_4[28:28]);
  NAND2 I182 (o_0r1[28:28], simp821_0[0:0], simp821_0[1:1]);
  NOR3 I183 (simp831_0[0:0], gtint_0[29:29], gtint_1[29:29], gtint_2[29:29]);
  NOR2 I184 (simp831_0[1:1], gtint_3[29:29], gtint_4[29:29]);
  NAND2 I185 (o_0r1[29:29], simp831_0[0:0], simp831_0[1:1]);
  NOR3 I186 (simp841_0[0:0], gtint_0[30:30], gtint_1[30:30], gtint_2[30:30]);
  NOR2 I187 (simp841_0[1:1], gtint_3[30:30], gtint_4[30:30]);
  NAND2 I188 (o_0r1[30:30], simp841_0[0:0], simp841_0[1:1]);
  NOR3 I189 (simp851_0[0:0], gtint_0[31:31], gtint_1[31:31], gtint_2[31:31]);
  NOR2 I190 (simp851_0[1:1], gtint_3[31:31], gtint_4[31:31]);
  NAND2 I191 (o_0r1[31:31], simp851_0[0:0], simp851_0[1:1]);
  AND2 I192 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I193 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I194 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I195 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I196 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I197 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I198 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I199 (gtint_0[7:7], choice_0, i_0r1[7:7]);
  AND2 I200 (gtint_0[8:8], choice_0, i_0r1[8:8]);
  AND2 I201 (gtint_0[9:9], choice_0, i_0r1[9:9]);
  AND2 I202 (gtint_0[10:10], choice_0, i_0r1[10:10]);
  AND2 I203 (gtint_0[11:11], choice_0, i_0r1[11:11]);
  AND2 I204 (gtint_0[12:12], choice_0, i_0r1[12:12]);
  AND2 I205 (gtint_0[13:13], choice_0, i_0r1[13:13]);
  AND2 I206 (gtint_0[14:14], choice_0, i_0r1[14:14]);
  AND2 I207 (gtint_0[15:15], choice_0, i_0r1[15:15]);
  AND2 I208 (gtint_0[16:16], choice_0, i_0r1[16:16]);
  AND2 I209 (gtint_0[17:17], choice_0, i_0r1[17:17]);
  AND2 I210 (gtint_0[18:18], choice_0, i_0r1[18:18]);
  AND2 I211 (gtint_0[19:19], choice_0, i_0r1[19:19]);
  AND2 I212 (gtint_0[20:20], choice_0, i_0r1[20:20]);
  AND2 I213 (gtint_0[21:21], choice_0, i_0r1[21:21]);
  AND2 I214 (gtint_0[22:22], choice_0, i_0r1[22:22]);
  AND2 I215 (gtint_0[23:23], choice_0, i_0r1[23:23]);
  AND2 I216 (gtint_0[24:24], choice_0, i_0r1[24:24]);
  AND2 I217 (gtint_0[25:25], choice_0, i_0r1[25:25]);
  AND2 I218 (gtint_0[26:26], choice_0, i_0r1[26:26]);
  AND2 I219 (gtint_0[27:27], choice_0, i_0r1[27:27]);
  AND2 I220 (gtint_0[28:28], choice_0, i_0r1[28:28]);
  AND2 I221 (gtint_0[29:29], choice_0, i_0r1[29:29]);
  AND2 I222 (gtint_0[30:30], choice_0, i_0r1[30:30]);
  AND2 I223 (gtint_0[31:31], choice_0, i_0r1[31:31]);
  AND2 I224 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I225 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I226 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I227 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I228 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I229 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I230 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I231 (gtint_1[7:7], choice_1, i_1r1[7:7]);
  AND2 I232 (gtint_1[8:8], choice_1, i_1r1[8:8]);
  AND2 I233 (gtint_1[9:9], choice_1, i_1r1[9:9]);
  AND2 I234 (gtint_1[10:10], choice_1, i_1r1[10:10]);
  AND2 I235 (gtint_1[11:11], choice_1, i_1r1[11:11]);
  AND2 I236 (gtint_1[12:12], choice_1, i_1r1[12:12]);
  AND2 I237 (gtint_1[13:13], choice_1, i_1r1[13:13]);
  AND2 I238 (gtint_1[14:14], choice_1, i_1r1[14:14]);
  AND2 I239 (gtint_1[15:15], choice_1, i_1r1[15:15]);
  AND2 I240 (gtint_1[16:16], choice_1, i_1r1[16:16]);
  AND2 I241 (gtint_1[17:17], choice_1, i_1r1[17:17]);
  AND2 I242 (gtint_1[18:18], choice_1, i_1r1[18:18]);
  AND2 I243 (gtint_1[19:19], choice_1, i_1r1[19:19]);
  AND2 I244 (gtint_1[20:20], choice_1, i_1r1[20:20]);
  AND2 I245 (gtint_1[21:21], choice_1, i_1r1[21:21]);
  AND2 I246 (gtint_1[22:22], choice_1, i_1r1[22:22]);
  AND2 I247 (gtint_1[23:23], choice_1, i_1r1[23:23]);
  AND2 I248 (gtint_1[24:24], choice_1, i_1r1[24:24]);
  AND2 I249 (gtint_1[25:25], choice_1, i_1r1[25:25]);
  AND2 I250 (gtint_1[26:26], choice_1, i_1r1[26:26]);
  AND2 I251 (gtint_1[27:27], choice_1, i_1r1[27:27]);
  AND2 I252 (gtint_1[28:28], choice_1, i_1r1[28:28]);
  AND2 I253 (gtint_1[29:29], choice_1, i_1r1[29:29]);
  AND2 I254 (gtint_1[30:30], choice_1, i_1r1[30:30]);
  AND2 I255 (gtint_1[31:31], choice_1, i_1r1[31:31]);
  AND2 I256 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I257 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I258 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I259 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AND2 I260 (gtint_2[4:4], choice_2, i_2r1[4:4]);
  AND2 I261 (gtint_2[5:5], choice_2, i_2r1[5:5]);
  AND2 I262 (gtint_2[6:6], choice_2, i_2r1[6:6]);
  AND2 I263 (gtint_2[7:7], choice_2, i_2r1[7:7]);
  AND2 I264 (gtint_2[8:8], choice_2, i_2r1[8:8]);
  AND2 I265 (gtint_2[9:9], choice_2, i_2r1[9:9]);
  AND2 I266 (gtint_2[10:10], choice_2, i_2r1[10:10]);
  AND2 I267 (gtint_2[11:11], choice_2, i_2r1[11:11]);
  AND2 I268 (gtint_2[12:12], choice_2, i_2r1[12:12]);
  AND2 I269 (gtint_2[13:13], choice_2, i_2r1[13:13]);
  AND2 I270 (gtint_2[14:14], choice_2, i_2r1[14:14]);
  AND2 I271 (gtint_2[15:15], choice_2, i_2r1[15:15]);
  AND2 I272 (gtint_2[16:16], choice_2, i_2r1[16:16]);
  AND2 I273 (gtint_2[17:17], choice_2, i_2r1[17:17]);
  AND2 I274 (gtint_2[18:18], choice_2, i_2r1[18:18]);
  AND2 I275 (gtint_2[19:19], choice_2, i_2r1[19:19]);
  AND2 I276 (gtint_2[20:20], choice_2, i_2r1[20:20]);
  AND2 I277 (gtint_2[21:21], choice_2, i_2r1[21:21]);
  AND2 I278 (gtint_2[22:22], choice_2, i_2r1[22:22]);
  AND2 I279 (gtint_2[23:23], choice_2, i_2r1[23:23]);
  AND2 I280 (gtint_2[24:24], choice_2, i_2r1[24:24]);
  AND2 I281 (gtint_2[25:25], choice_2, i_2r1[25:25]);
  AND2 I282 (gtint_2[26:26], choice_2, i_2r1[26:26]);
  AND2 I283 (gtint_2[27:27], choice_2, i_2r1[27:27]);
  AND2 I284 (gtint_2[28:28], choice_2, i_2r1[28:28]);
  AND2 I285 (gtint_2[29:29], choice_2, i_2r1[29:29]);
  AND2 I286 (gtint_2[30:30], choice_2, i_2r1[30:30]);
  AND2 I287 (gtint_2[31:31], choice_2, i_2r1[31:31]);
  AND2 I288 (gtint_3[0:0], choice_3, i_3r1[0:0]);
  AND2 I289 (gtint_3[1:1], choice_3, i_3r1[1:1]);
  AND2 I290 (gtint_3[2:2], choice_3, i_3r1[2:2]);
  AND2 I291 (gtint_3[3:3], choice_3, i_3r1[3:3]);
  AND2 I292 (gtint_3[4:4], choice_3, i_3r1[4:4]);
  AND2 I293 (gtint_3[5:5], choice_3, i_3r1[5:5]);
  AND2 I294 (gtint_3[6:6], choice_3, i_3r1[6:6]);
  AND2 I295 (gtint_3[7:7], choice_3, i_3r1[7:7]);
  AND2 I296 (gtint_3[8:8], choice_3, i_3r1[8:8]);
  AND2 I297 (gtint_3[9:9], choice_3, i_3r1[9:9]);
  AND2 I298 (gtint_3[10:10], choice_3, i_3r1[10:10]);
  AND2 I299 (gtint_3[11:11], choice_3, i_3r1[11:11]);
  AND2 I300 (gtint_3[12:12], choice_3, i_3r1[12:12]);
  AND2 I301 (gtint_3[13:13], choice_3, i_3r1[13:13]);
  AND2 I302 (gtint_3[14:14], choice_3, i_3r1[14:14]);
  AND2 I303 (gtint_3[15:15], choice_3, i_3r1[15:15]);
  AND2 I304 (gtint_3[16:16], choice_3, i_3r1[16:16]);
  AND2 I305 (gtint_3[17:17], choice_3, i_3r1[17:17]);
  AND2 I306 (gtint_3[18:18], choice_3, i_3r1[18:18]);
  AND2 I307 (gtint_3[19:19], choice_3, i_3r1[19:19]);
  AND2 I308 (gtint_3[20:20], choice_3, i_3r1[20:20]);
  AND2 I309 (gtint_3[21:21], choice_3, i_3r1[21:21]);
  AND2 I310 (gtint_3[22:22], choice_3, i_3r1[22:22]);
  AND2 I311 (gtint_3[23:23], choice_3, i_3r1[23:23]);
  AND2 I312 (gtint_3[24:24], choice_3, i_3r1[24:24]);
  AND2 I313 (gtint_3[25:25], choice_3, i_3r1[25:25]);
  AND2 I314 (gtint_3[26:26], choice_3, i_3r1[26:26]);
  AND2 I315 (gtint_3[27:27], choice_3, i_3r1[27:27]);
  AND2 I316 (gtint_3[28:28], choice_3, i_3r1[28:28]);
  AND2 I317 (gtint_3[29:29], choice_3, i_3r1[29:29]);
  AND2 I318 (gtint_3[30:30], choice_3, i_3r1[30:30]);
  AND2 I319 (gtint_3[31:31], choice_3, i_3r1[31:31]);
  AND2 I320 (gtint_4[0:0], choice_4, i_4r1[0:0]);
  AND2 I321 (gtint_4[1:1], choice_4, i_4r1[1:1]);
  AND2 I322 (gtint_4[2:2], choice_4, i_4r1[2:2]);
  AND2 I323 (gtint_4[3:3], choice_4, i_4r1[3:3]);
  AND2 I324 (gtint_4[4:4], choice_4, i_4r1[4:4]);
  AND2 I325 (gtint_4[5:5], choice_4, i_4r1[5:5]);
  AND2 I326 (gtint_4[6:6], choice_4, i_4r1[6:6]);
  AND2 I327 (gtint_4[7:7], choice_4, i_4r1[7:7]);
  AND2 I328 (gtint_4[8:8], choice_4, i_4r1[8:8]);
  AND2 I329 (gtint_4[9:9], choice_4, i_4r1[9:9]);
  AND2 I330 (gtint_4[10:10], choice_4, i_4r1[10:10]);
  AND2 I331 (gtint_4[11:11], choice_4, i_4r1[11:11]);
  AND2 I332 (gtint_4[12:12], choice_4, i_4r1[12:12]);
  AND2 I333 (gtint_4[13:13], choice_4, i_4r1[13:13]);
  AND2 I334 (gtint_4[14:14], choice_4, i_4r1[14:14]);
  AND2 I335 (gtint_4[15:15], choice_4, i_4r1[15:15]);
  AND2 I336 (gtint_4[16:16], choice_4, i_4r1[16:16]);
  AND2 I337 (gtint_4[17:17], choice_4, i_4r1[17:17]);
  AND2 I338 (gtint_4[18:18], choice_4, i_4r1[18:18]);
  AND2 I339 (gtint_4[19:19], choice_4, i_4r1[19:19]);
  AND2 I340 (gtint_4[20:20], choice_4, i_4r1[20:20]);
  AND2 I341 (gtint_4[21:21], choice_4, i_4r1[21:21]);
  AND2 I342 (gtint_4[22:22], choice_4, i_4r1[22:22]);
  AND2 I343 (gtint_4[23:23], choice_4, i_4r1[23:23]);
  AND2 I344 (gtint_4[24:24], choice_4, i_4r1[24:24]);
  AND2 I345 (gtint_4[25:25], choice_4, i_4r1[25:25]);
  AND2 I346 (gtint_4[26:26], choice_4, i_4r1[26:26]);
  AND2 I347 (gtint_4[27:27], choice_4, i_4r1[27:27]);
  AND2 I348 (gtint_4[28:28], choice_4, i_4r1[28:28]);
  AND2 I349 (gtint_4[29:29], choice_4, i_4r1[29:29]);
  AND2 I350 (gtint_4[30:30], choice_4, i_4r1[30:30]);
  AND2 I351 (gtint_4[31:31], choice_4, i_4r1[31:31]);
  AND2 I352 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I353 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I354 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I355 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I356 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I357 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I358 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I359 (gfint_0[7:7], choice_0, i_0r0[7:7]);
  AND2 I360 (gfint_0[8:8], choice_0, i_0r0[8:8]);
  AND2 I361 (gfint_0[9:9], choice_0, i_0r0[9:9]);
  AND2 I362 (gfint_0[10:10], choice_0, i_0r0[10:10]);
  AND2 I363 (gfint_0[11:11], choice_0, i_0r0[11:11]);
  AND2 I364 (gfint_0[12:12], choice_0, i_0r0[12:12]);
  AND2 I365 (gfint_0[13:13], choice_0, i_0r0[13:13]);
  AND2 I366 (gfint_0[14:14], choice_0, i_0r0[14:14]);
  AND2 I367 (gfint_0[15:15], choice_0, i_0r0[15:15]);
  AND2 I368 (gfint_0[16:16], choice_0, i_0r0[16:16]);
  AND2 I369 (gfint_0[17:17], choice_0, i_0r0[17:17]);
  AND2 I370 (gfint_0[18:18], choice_0, i_0r0[18:18]);
  AND2 I371 (gfint_0[19:19], choice_0, i_0r0[19:19]);
  AND2 I372 (gfint_0[20:20], choice_0, i_0r0[20:20]);
  AND2 I373 (gfint_0[21:21], choice_0, i_0r0[21:21]);
  AND2 I374 (gfint_0[22:22], choice_0, i_0r0[22:22]);
  AND2 I375 (gfint_0[23:23], choice_0, i_0r0[23:23]);
  AND2 I376 (gfint_0[24:24], choice_0, i_0r0[24:24]);
  AND2 I377 (gfint_0[25:25], choice_0, i_0r0[25:25]);
  AND2 I378 (gfint_0[26:26], choice_0, i_0r0[26:26]);
  AND2 I379 (gfint_0[27:27], choice_0, i_0r0[27:27]);
  AND2 I380 (gfint_0[28:28], choice_0, i_0r0[28:28]);
  AND2 I381 (gfint_0[29:29], choice_0, i_0r0[29:29]);
  AND2 I382 (gfint_0[30:30], choice_0, i_0r0[30:30]);
  AND2 I383 (gfint_0[31:31], choice_0, i_0r0[31:31]);
  AND2 I384 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I385 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I386 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I387 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I388 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I389 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I390 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I391 (gfint_1[7:7], choice_1, i_1r0[7:7]);
  AND2 I392 (gfint_1[8:8], choice_1, i_1r0[8:8]);
  AND2 I393 (gfint_1[9:9], choice_1, i_1r0[9:9]);
  AND2 I394 (gfint_1[10:10], choice_1, i_1r0[10:10]);
  AND2 I395 (gfint_1[11:11], choice_1, i_1r0[11:11]);
  AND2 I396 (gfint_1[12:12], choice_1, i_1r0[12:12]);
  AND2 I397 (gfint_1[13:13], choice_1, i_1r0[13:13]);
  AND2 I398 (gfint_1[14:14], choice_1, i_1r0[14:14]);
  AND2 I399 (gfint_1[15:15], choice_1, i_1r0[15:15]);
  AND2 I400 (gfint_1[16:16], choice_1, i_1r0[16:16]);
  AND2 I401 (gfint_1[17:17], choice_1, i_1r0[17:17]);
  AND2 I402 (gfint_1[18:18], choice_1, i_1r0[18:18]);
  AND2 I403 (gfint_1[19:19], choice_1, i_1r0[19:19]);
  AND2 I404 (gfint_1[20:20], choice_1, i_1r0[20:20]);
  AND2 I405 (gfint_1[21:21], choice_1, i_1r0[21:21]);
  AND2 I406 (gfint_1[22:22], choice_1, i_1r0[22:22]);
  AND2 I407 (gfint_1[23:23], choice_1, i_1r0[23:23]);
  AND2 I408 (gfint_1[24:24], choice_1, i_1r0[24:24]);
  AND2 I409 (gfint_1[25:25], choice_1, i_1r0[25:25]);
  AND2 I410 (gfint_1[26:26], choice_1, i_1r0[26:26]);
  AND2 I411 (gfint_1[27:27], choice_1, i_1r0[27:27]);
  AND2 I412 (gfint_1[28:28], choice_1, i_1r0[28:28]);
  AND2 I413 (gfint_1[29:29], choice_1, i_1r0[29:29]);
  AND2 I414 (gfint_1[30:30], choice_1, i_1r0[30:30]);
  AND2 I415 (gfint_1[31:31], choice_1, i_1r0[31:31]);
  AND2 I416 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I417 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I418 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I419 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AND2 I420 (gfint_2[4:4], choice_2, i_2r0[4:4]);
  AND2 I421 (gfint_2[5:5], choice_2, i_2r0[5:5]);
  AND2 I422 (gfint_2[6:6], choice_2, i_2r0[6:6]);
  AND2 I423 (gfint_2[7:7], choice_2, i_2r0[7:7]);
  AND2 I424 (gfint_2[8:8], choice_2, i_2r0[8:8]);
  AND2 I425 (gfint_2[9:9], choice_2, i_2r0[9:9]);
  AND2 I426 (gfint_2[10:10], choice_2, i_2r0[10:10]);
  AND2 I427 (gfint_2[11:11], choice_2, i_2r0[11:11]);
  AND2 I428 (gfint_2[12:12], choice_2, i_2r0[12:12]);
  AND2 I429 (gfint_2[13:13], choice_2, i_2r0[13:13]);
  AND2 I430 (gfint_2[14:14], choice_2, i_2r0[14:14]);
  AND2 I431 (gfint_2[15:15], choice_2, i_2r0[15:15]);
  AND2 I432 (gfint_2[16:16], choice_2, i_2r0[16:16]);
  AND2 I433 (gfint_2[17:17], choice_2, i_2r0[17:17]);
  AND2 I434 (gfint_2[18:18], choice_2, i_2r0[18:18]);
  AND2 I435 (gfint_2[19:19], choice_2, i_2r0[19:19]);
  AND2 I436 (gfint_2[20:20], choice_2, i_2r0[20:20]);
  AND2 I437 (gfint_2[21:21], choice_2, i_2r0[21:21]);
  AND2 I438 (gfint_2[22:22], choice_2, i_2r0[22:22]);
  AND2 I439 (gfint_2[23:23], choice_2, i_2r0[23:23]);
  AND2 I440 (gfint_2[24:24], choice_2, i_2r0[24:24]);
  AND2 I441 (gfint_2[25:25], choice_2, i_2r0[25:25]);
  AND2 I442 (gfint_2[26:26], choice_2, i_2r0[26:26]);
  AND2 I443 (gfint_2[27:27], choice_2, i_2r0[27:27]);
  AND2 I444 (gfint_2[28:28], choice_2, i_2r0[28:28]);
  AND2 I445 (gfint_2[29:29], choice_2, i_2r0[29:29]);
  AND2 I446 (gfint_2[30:30], choice_2, i_2r0[30:30]);
  AND2 I447 (gfint_2[31:31], choice_2, i_2r0[31:31]);
  AND2 I448 (gfint_3[0:0], choice_3, i_3r0[0:0]);
  AND2 I449 (gfint_3[1:1], choice_3, i_3r0[1:1]);
  AND2 I450 (gfint_3[2:2], choice_3, i_3r0[2:2]);
  AND2 I451 (gfint_3[3:3], choice_3, i_3r0[3:3]);
  AND2 I452 (gfint_3[4:4], choice_3, i_3r0[4:4]);
  AND2 I453 (gfint_3[5:5], choice_3, i_3r0[5:5]);
  AND2 I454 (gfint_3[6:6], choice_3, i_3r0[6:6]);
  AND2 I455 (gfint_3[7:7], choice_3, i_3r0[7:7]);
  AND2 I456 (gfint_3[8:8], choice_3, i_3r0[8:8]);
  AND2 I457 (gfint_3[9:9], choice_3, i_3r0[9:9]);
  AND2 I458 (gfint_3[10:10], choice_3, i_3r0[10:10]);
  AND2 I459 (gfint_3[11:11], choice_3, i_3r0[11:11]);
  AND2 I460 (gfint_3[12:12], choice_3, i_3r0[12:12]);
  AND2 I461 (gfint_3[13:13], choice_3, i_3r0[13:13]);
  AND2 I462 (gfint_3[14:14], choice_3, i_3r0[14:14]);
  AND2 I463 (gfint_3[15:15], choice_3, i_3r0[15:15]);
  AND2 I464 (gfint_3[16:16], choice_3, i_3r0[16:16]);
  AND2 I465 (gfint_3[17:17], choice_3, i_3r0[17:17]);
  AND2 I466 (gfint_3[18:18], choice_3, i_3r0[18:18]);
  AND2 I467 (gfint_3[19:19], choice_3, i_3r0[19:19]);
  AND2 I468 (gfint_3[20:20], choice_3, i_3r0[20:20]);
  AND2 I469 (gfint_3[21:21], choice_3, i_3r0[21:21]);
  AND2 I470 (gfint_3[22:22], choice_3, i_3r0[22:22]);
  AND2 I471 (gfint_3[23:23], choice_3, i_3r0[23:23]);
  AND2 I472 (gfint_3[24:24], choice_3, i_3r0[24:24]);
  AND2 I473 (gfint_3[25:25], choice_3, i_3r0[25:25]);
  AND2 I474 (gfint_3[26:26], choice_3, i_3r0[26:26]);
  AND2 I475 (gfint_3[27:27], choice_3, i_3r0[27:27]);
  AND2 I476 (gfint_3[28:28], choice_3, i_3r0[28:28]);
  AND2 I477 (gfint_3[29:29], choice_3, i_3r0[29:29]);
  AND2 I478 (gfint_3[30:30], choice_3, i_3r0[30:30]);
  AND2 I479 (gfint_3[31:31], choice_3, i_3r0[31:31]);
  AND2 I480 (gfint_4[0:0], choice_4, i_4r0[0:0]);
  AND2 I481 (gfint_4[1:1], choice_4, i_4r0[1:1]);
  AND2 I482 (gfint_4[2:2], choice_4, i_4r0[2:2]);
  AND2 I483 (gfint_4[3:3], choice_4, i_4r0[3:3]);
  AND2 I484 (gfint_4[4:4], choice_4, i_4r0[4:4]);
  AND2 I485 (gfint_4[5:5], choice_4, i_4r0[5:5]);
  AND2 I486 (gfint_4[6:6], choice_4, i_4r0[6:6]);
  AND2 I487 (gfint_4[7:7], choice_4, i_4r0[7:7]);
  AND2 I488 (gfint_4[8:8], choice_4, i_4r0[8:8]);
  AND2 I489 (gfint_4[9:9], choice_4, i_4r0[9:9]);
  AND2 I490 (gfint_4[10:10], choice_4, i_4r0[10:10]);
  AND2 I491 (gfint_4[11:11], choice_4, i_4r0[11:11]);
  AND2 I492 (gfint_4[12:12], choice_4, i_4r0[12:12]);
  AND2 I493 (gfint_4[13:13], choice_4, i_4r0[13:13]);
  AND2 I494 (gfint_4[14:14], choice_4, i_4r0[14:14]);
  AND2 I495 (gfint_4[15:15], choice_4, i_4r0[15:15]);
  AND2 I496 (gfint_4[16:16], choice_4, i_4r0[16:16]);
  AND2 I497 (gfint_4[17:17], choice_4, i_4r0[17:17]);
  AND2 I498 (gfint_4[18:18], choice_4, i_4r0[18:18]);
  AND2 I499 (gfint_4[19:19], choice_4, i_4r0[19:19]);
  AND2 I500 (gfint_4[20:20], choice_4, i_4r0[20:20]);
  AND2 I501 (gfint_4[21:21], choice_4, i_4r0[21:21]);
  AND2 I502 (gfint_4[22:22], choice_4, i_4r0[22:22]);
  AND2 I503 (gfint_4[23:23], choice_4, i_4r0[23:23]);
  AND2 I504 (gfint_4[24:24], choice_4, i_4r0[24:24]);
  AND2 I505 (gfint_4[25:25], choice_4, i_4r0[25:25]);
  AND2 I506 (gfint_4[26:26], choice_4, i_4r0[26:26]);
  AND2 I507 (gfint_4[27:27], choice_4, i_4r0[27:27]);
  AND2 I508 (gfint_4[28:28], choice_4, i_4r0[28:28]);
  AND2 I509 (gfint_4[29:29], choice_4, i_4r0[29:29]);
  AND2 I510 (gfint_4[30:30], choice_4, i_4r0[30:30]);
  AND2 I511 (gfint_4[31:31], choice_4, i_4r0[31:31]);
  OR2 I512 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I513 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I514 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I515 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I516 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I517 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I518 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I519 (comp0_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I520 (comp0_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I521 (comp0_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I522 (comp0_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I523 (comp0_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I524 (comp0_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I525 (comp0_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I526 (comp0_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I527 (comp0_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I528 (comp0_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I529 (comp0_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I530 (comp0_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I531 (comp0_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I532 (comp0_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I533 (comp0_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I534 (comp0_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I535 (comp0_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I536 (comp0_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I537 (comp0_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I538 (comp0_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I539 (comp0_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I540 (comp0_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I541 (comp0_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I542 (comp0_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I543 (comp0_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  C3 I544 (simp4391_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I545 (simp4391_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I546 (simp4391_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I547 (simp4391_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I548 (simp4391_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I549 (simp4391_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I550 (simp4391_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I551 (simp4391_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I552 (simp4391_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I553 (simp4391_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I554 (simp4391_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I555 (simp4392_0[0:0], simp4391_0[0:0], simp4391_0[1:1], simp4391_0[2:2]);
  C3 I556 (simp4392_0[1:1], simp4391_0[3:3], simp4391_0[4:4], simp4391_0[5:5]);
  C3 I557 (simp4392_0[2:2], simp4391_0[6:6], simp4391_0[7:7], simp4391_0[8:8]);
  C2 I558 (simp4392_0[3:3], simp4391_0[9:9], simp4391_0[10:10]);
  C3 I559 (simp4393_0[0:0], simp4392_0[0:0], simp4392_0[1:1], simp4392_0[2:2]);
  BUFF I560 (simp4393_0[1:1], simp4392_0[3:3]);
  C2 I561 (icomp_0, simp4393_0[0:0], simp4393_0[1:1]);
  OR2 I562 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I563 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I564 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I565 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I566 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I567 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I568 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  OR2 I569 (comp1_0[7:7], i_1r0[7:7], i_1r1[7:7]);
  OR2 I570 (comp1_0[8:8], i_1r0[8:8], i_1r1[8:8]);
  OR2 I571 (comp1_0[9:9], i_1r0[9:9], i_1r1[9:9]);
  OR2 I572 (comp1_0[10:10], i_1r0[10:10], i_1r1[10:10]);
  OR2 I573 (comp1_0[11:11], i_1r0[11:11], i_1r1[11:11]);
  OR2 I574 (comp1_0[12:12], i_1r0[12:12], i_1r1[12:12]);
  OR2 I575 (comp1_0[13:13], i_1r0[13:13], i_1r1[13:13]);
  OR2 I576 (comp1_0[14:14], i_1r0[14:14], i_1r1[14:14]);
  OR2 I577 (comp1_0[15:15], i_1r0[15:15], i_1r1[15:15]);
  OR2 I578 (comp1_0[16:16], i_1r0[16:16], i_1r1[16:16]);
  OR2 I579 (comp1_0[17:17], i_1r0[17:17], i_1r1[17:17]);
  OR2 I580 (comp1_0[18:18], i_1r0[18:18], i_1r1[18:18]);
  OR2 I581 (comp1_0[19:19], i_1r0[19:19], i_1r1[19:19]);
  OR2 I582 (comp1_0[20:20], i_1r0[20:20], i_1r1[20:20]);
  OR2 I583 (comp1_0[21:21], i_1r0[21:21], i_1r1[21:21]);
  OR2 I584 (comp1_0[22:22], i_1r0[22:22], i_1r1[22:22]);
  OR2 I585 (comp1_0[23:23], i_1r0[23:23], i_1r1[23:23]);
  OR2 I586 (comp1_0[24:24], i_1r0[24:24], i_1r1[24:24]);
  OR2 I587 (comp1_0[25:25], i_1r0[25:25], i_1r1[25:25]);
  OR2 I588 (comp1_0[26:26], i_1r0[26:26], i_1r1[26:26]);
  OR2 I589 (comp1_0[27:27], i_1r0[27:27], i_1r1[27:27]);
  OR2 I590 (comp1_0[28:28], i_1r0[28:28], i_1r1[28:28]);
  OR2 I591 (comp1_0[29:29], i_1r0[29:29], i_1r1[29:29]);
  OR2 I592 (comp1_0[30:30], i_1r0[30:30], i_1r1[30:30]);
  OR2 I593 (comp1_0[31:31], i_1r0[31:31], i_1r1[31:31]);
  C3 I594 (simp4731_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I595 (simp4731_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  C3 I596 (simp4731_0[2:2], comp1_0[6:6], comp1_0[7:7], comp1_0[8:8]);
  C3 I597 (simp4731_0[3:3], comp1_0[9:9], comp1_0[10:10], comp1_0[11:11]);
  C3 I598 (simp4731_0[4:4], comp1_0[12:12], comp1_0[13:13], comp1_0[14:14]);
  C3 I599 (simp4731_0[5:5], comp1_0[15:15], comp1_0[16:16], comp1_0[17:17]);
  C3 I600 (simp4731_0[6:6], comp1_0[18:18], comp1_0[19:19], comp1_0[20:20]);
  C3 I601 (simp4731_0[7:7], comp1_0[21:21], comp1_0[22:22], comp1_0[23:23]);
  C3 I602 (simp4731_0[8:8], comp1_0[24:24], comp1_0[25:25], comp1_0[26:26]);
  C3 I603 (simp4731_0[9:9], comp1_0[27:27], comp1_0[28:28], comp1_0[29:29]);
  C2 I604 (simp4731_0[10:10], comp1_0[30:30], comp1_0[31:31]);
  C3 I605 (simp4732_0[0:0], simp4731_0[0:0], simp4731_0[1:1], simp4731_0[2:2]);
  C3 I606 (simp4732_0[1:1], simp4731_0[3:3], simp4731_0[4:4], simp4731_0[5:5]);
  C3 I607 (simp4732_0[2:2], simp4731_0[6:6], simp4731_0[7:7], simp4731_0[8:8]);
  C2 I608 (simp4732_0[3:3], simp4731_0[9:9], simp4731_0[10:10]);
  C3 I609 (simp4733_0[0:0], simp4732_0[0:0], simp4732_0[1:1], simp4732_0[2:2]);
  BUFF I610 (simp4733_0[1:1], simp4732_0[3:3]);
  C2 I611 (icomp_1, simp4733_0[0:0], simp4733_0[1:1]);
  OR2 I612 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I613 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I614 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2 I615 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  OR2 I616 (comp2_0[4:4], i_2r0[4:4], i_2r1[4:4]);
  OR2 I617 (comp2_0[5:5], i_2r0[5:5], i_2r1[5:5]);
  OR2 I618 (comp2_0[6:6], i_2r0[6:6], i_2r1[6:6]);
  OR2 I619 (comp2_0[7:7], i_2r0[7:7], i_2r1[7:7]);
  OR2 I620 (comp2_0[8:8], i_2r0[8:8], i_2r1[8:8]);
  OR2 I621 (comp2_0[9:9], i_2r0[9:9], i_2r1[9:9]);
  OR2 I622 (comp2_0[10:10], i_2r0[10:10], i_2r1[10:10]);
  OR2 I623 (comp2_0[11:11], i_2r0[11:11], i_2r1[11:11]);
  OR2 I624 (comp2_0[12:12], i_2r0[12:12], i_2r1[12:12]);
  OR2 I625 (comp2_0[13:13], i_2r0[13:13], i_2r1[13:13]);
  OR2 I626 (comp2_0[14:14], i_2r0[14:14], i_2r1[14:14]);
  OR2 I627 (comp2_0[15:15], i_2r0[15:15], i_2r1[15:15]);
  OR2 I628 (comp2_0[16:16], i_2r0[16:16], i_2r1[16:16]);
  OR2 I629 (comp2_0[17:17], i_2r0[17:17], i_2r1[17:17]);
  OR2 I630 (comp2_0[18:18], i_2r0[18:18], i_2r1[18:18]);
  OR2 I631 (comp2_0[19:19], i_2r0[19:19], i_2r1[19:19]);
  OR2 I632 (comp2_0[20:20], i_2r0[20:20], i_2r1[20:20]);
  OR2 I633 (comp2_0[21:21], i_2r0[21:21], i_2r1[21:21]);
  OR2 I634 (comp2_0[22:22], i_2r0[22:22], i_2r1[22:22]);
  OR2 I635 (comp2_0[23:23], i_2r0[23:23], i_2r1[23:23]);
  OR2 I636 (comp2_0[24:24], i_2r0[24:24], i_2r1[24:24]);
  OR2 I637 (comp2_0[25:25], i_2r0[25:25], i_2r1[25:25]);
  OR2 I638 (comp2_0[26:26], i_2r0[26:26], i_2r1[26:26]);
  OR2 I639 (comp2_0[27:27], i_2r0[27:27], i_2r1[27:27]);
  OR2 I640 (comp2_0[28:28], i_2r0[28:28], i_2r1[28:28]);
  OR2 I641 (comp2_0[29:29], i_2r0[29:29], i_2r1[29:29]);
  OR2 I642 (comp2_0[30:30], i_2r0[30:30], i_2r1[30:30]);
  OR2 I643 (comp2_0[31:31], i_2r0[31:31], i_2r1[31:31]);
  C3 I644 (simp5071_0[0:0], comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C3 I645 (simp5071_0[1:1], comp2_0[3:3], comp2_0[4:4], comp2_0[5:5]);
  C3 I646 (simp5071_0[2:2], comp2_0[6:6], comp2_0[7:7], comp2_0[8:8]);
  C3 I647 (simp5071_0[3:3], comp2_0[9:9], comp2_0[10:10], comp2_0[11:11]);
  C3 I648 (simp5071_0[4:4], comp2_0[12:12], comp2_0[13:13], comp2_0[14:14]);
  C3 I649 (simp5071_0[5:5], comp2_0[15:15], comp2_0[16:16], comp2_0[17:17]);
  C3 I650 (simp5071_0[6:6], comp2_0[18:18], comp2_0[19:19], comp2_0[20:20]);
  C3 I651 (simp5071_0[7:7], comp2_0[21:21], comp2_0[22:22], comp2_0[23:23]);
  C3 I652 (simp5071_0[8:8], comp2_0[24:24], comp2_0[25:25], comp2_0[26:26]);
  C3 I653 (simp5071_0[9:9], comp2_0[27:27], comp2_0[28:28], comp2_0[29:29]);
  C2 I654 (simp5071_0[10:10], comp2_0[30:30], comp2_0[31:31]);
  C3 I655 (simp5072_0[0:0], simp5071_0[0:0], simp5071_0[1:1], simp5071_0[2:2]);
  C3 I656 (simp5072_0[1:1], simp5071_0[3:3], simp5071_0[4:4], simp5071_0[5:5]);
  C3 I657 (simp5072_0[2:2], simp5071_0[6:6], simp5071_0[7:7], simp5071_0[8:8]);
  C2 I658 (simp5072_0[3:3], simp5071_0[9:9], simp5071_0[10:10]);
  C3 I659 (simp5073_0[0:0], simp5072_0[0:0], simp5072_0[1:1], simp5072_0[2:2]);
  BUFF I660 (simp5073_0[1:1], simp5072_0[3:3]);
  C2 I661 (icomp_2, simp5073_0[0:0], simp5073_0[1:1]);
  OR2 I662 (comp3_0[0:0], i_3r0[0:0], i_3r1[0:0]);
  OR2 I663 (comp3_0[1:1], i_3r0[1:1], i_3r1[1:1]);
  OR2 I664 (comp3_0[2:2], i_3r0[2:2], i_3r1[2:2]);
  OR2 I665 (comp3_0[3:3], i_3r0[3:3], i_3r1[3:3]);
  OR2 I666 (comp3_0[4:4], i_3r0[4:4], i_3r1[4:4]);
  OR2 I667 (comp3_0[5:5], i_3r0[5:5], i_3r1[5:5]);
  OR2 I668 (comp3_0[6:6], i_3r0[6:6], i_3r1[6:6]);
  OR2 I669 (comp3_0[7:7], i_3r0[7:7], i_3r1[7:7]);
  OR2 I670 (comp3_0[8:8], i_3r0[8:8], i_3r1[8:8]);
  OR2 I671 (comp3_0[9:9], i_3r0[9:9], i_3r1[9:9]);
  OR2 I672 (comp3_0[10:10], i_3r0[10:10], i_3r1[10:10]);
  OR2 I673 (comp3_0[11:11], i_3r0[11:11], i_3r1[11:11]);
  OR2 I674 (comp3_0[12:12], i_3r0[12:12], i_3r1[12:12]);
  OR2 I675 (comp3_0[13:13], i_3r0[13:13], i_3r1[13:13]);
  OR2 I676 (comp3_0[14:14], i_3r0[14:14], i_3r1[14:14]);
  OR2 I677 (comp3_0[15:15], i_3r0[15:15], i_3r1[15:15]);
  OR2 I678 (comp3_0[16:16], i_3r0[16:16], i_3r1[16:16]);
  OR2 I679 (comp3_0[17:17], i_3r0[17:17], i_3r1[17:17]);
  OR2 I680 (comp3_0[18:18], i_3r0[18:18], i_3r1[18:18]);
  OR2 I681 (comp3_0[19:19], i_3r0[19:19], i_3r1[19:19]);
  OR2 I682 (comp3_0[20:20], i_3r0[20:20], i_3r1[20:20]);
  OR2 I683 (comp3_0[21:21], i_3r0[21:21], i_3r1[21:21]);
  OR2 I684 (comp3_0[22:22], i_3r0[22:22], i_3r1[22:22]);
  OR2 I685 (comp3_0[23:23], i_3r0[23:23], i_3r1[23:23]);
  OR2 I686 (comp3_0[24:24], i_3r0[24:24], i_3r1[24:24]);
  OR2 I687 (comp3_0[25:25], i_3r0[25:25], i_3r1[25:25]);
  OR2 I688 (comp3_0[26:26], i_3r0[26:26], i_3r1[26:26]);
  OR2 I689 (comp3_0[27:27], i_3r0[27:27], i_3r1[27:27]);
  OR2 I690 (comp3_0[28:28], i_3r0[28:28], i_3r1[28:28]);
  OR2 I691 (comp3_0[29:29], i_3r0[29:29], i_3r1[29:29]);
  OR2 I692 (comp3_0[30:30], i_3r0[30:30], i_3r1[30:30]);
  OR2 I693 (comp3_0[31:31], i_3r0[31:31], i_3r1[31:31]);
  C3 I694 (simp5411_0[0:0], comp3_0[0:0], comp3_0[1:1], comp3_0[2:2]);
  C3 I695 (simp5411_0[1:1], comp3_0[3:3], comp3_0[4:4], comp3_0[5:5]);
  C3 I696 (simp5411_0[2:2], comp3_0[6:6], comp3_0[7:7], comp3_0[8:8]);
  C3 I697 (simp5411_0[3:3], comp3_0[9:9], comp3_0[10:10], comp3_0[11:11]);
  C3 I698 (simp5411_0[4:4], comp3_0[12:12], comp3_0[13:13], comp3_0[14:14]);
  C3 I699 (simp5411_0[5:5], comp3_0[15:15], comp3_0[16:16], comp3_0[17:17]);
  C3 I700 (simp5411_0[6:6], comp3_0[18:18], comp3_0[19:19], comp3_0[20:20]);
  C3 I701 (simp5411_0[7:7], comp3_0[21:21], comp3_0[22:22], comp3_0[23:23]);
  C3 I702 (simp5411_0[8:8], comp3_0[24:24], comp3_0[25:25], comp3_0[26:26]);
  C3 I703 (simp5411_0[9:9], comp3_0[27:27], comp3_0[28:28], comp3_0[29:29]);
  C2 I704 (simp5411_0[10:10], comp3_0[30:30], comp3_0[31:31]);
  C3 I705 (simp5412_0[0:0], simp5411_0[0:0], simp5411_0[1:1], simp5411_0[2:2]);
  C3 I706 (simp5412_0[1:1], simp5411_0[3:3], simp5411_0[4:4], simp5411_0[5:5]);
  C3 I707 (simp5412_0[2:2], simp5411_0[6:6], simp5411_0[7:7], simp5411_0[8:8]);
  C2 I708 (simp5412_0[3:3], simp5411_0[9:9], simp5411_0[10:10]);
  C3 I709 (simp5413_0[0:0], simp5412_0[0:0], simp5412_0[1:1], simp5412_0[2:2]);
  BUFF I710 (simp5413_0[1:1], simp5412_0[3:3]);
  C2 I711 (icomp_3, simp5413_0[0:0], simp5413_0[1:1]);
  OR2 I712 (comp4_0[0:0], i_4r0[0:0], i_4r1[0:0]);
  OR2 I713 (comp4_0[1:1], i_4r0[1:1], i_4r1[1:1]);
  OR2 I714 (comp4_0[2:2], i_4r0[2:2], i_4r1[2:2]);
  OR2 I715 (comp4_0[3:3], i_4r0[3:3], i_4r1[3:3]);
  OR2 I716 (comp4_0[4:4], i_4r0[4:4], i_4r1[4:4]);
  OR2 I717 (comp4_0[5:5], i_4r0[5:5], i_4r1[5:5]);
  OR2 I718 (comp4_0[6:6], i_4r0[6:6], i_4r1[6:6]);
  OR2 I719 (comp4_0[7:7], i_4r0[7:7], i_4r1[7:7]);
  OR2 I720 (comp4_0[8:8], i_4r0[8:8], i_4r1[8:8]);
  OR2 I721 (comp4_0[9:9], i_4r0[9:9], i_4r1[9:9]);
  OR2 I722 (comp4_0[10:10], i_4r0[10:10], i_4r1[10:10]);
  OR2 I723 (comp4_0[11:11], i_4r0[11:11], i_4r1[11:11]);
  OR2 I724 (comp4_0[12:12], i_4r0[12:12], i_4r1[12:12]);
  OR2 I725 (comp4_0[13:13], i_4r0[13:13], i_4r1[13:13]);
  OR2 I726 (comp4_0[14:14], i_4r0[14:14], i_4r1[14:14]);
  OR2 I727 (comp4_0[15:15], i_4r0[15:15], i_4r1[15:15]);
  OR2 I728 (comp4_0[16:16], i_4r0[16:16], i_4r1[16:16]);
  OR2 I729 (comp4_0[17:17], i_4r0[17:17], i_4r1[17:17]);
  OR2 I730 (comp4_0[18:18], i_4r0[18:18], i_4r1[18:18]);
  OR2 I731 (comp4_0[19:19], i_4r0[19:19], i_4r1[19:19]);
  OR2 I732 (comp4_0[20:20], i_4r0[20:20], i_4r1[20:20]);
  OR2 I733 (comp4_0[21:21], i_4r0[21:21], i_4r1[21:21]);
  OR2 I734 (comp4_0[22:22], i_4r0[22:22], i_4r1[22:22]);
  OR2 I735 (comp4_0[23:23], i_4r0[23:23], i_4r1[23:23]);
  OR2 I736 (comp4_0[24:24], i_4r0[24:24], i_4r1[24:24]);
  OR2 I737 (comp4_0[25:25], i_4r0[25:25], i_4r1[25:25]);
  OR2 I738 (comp4_0[26:26], i_4r0[26:26], i_4r1[26:26]);
  OR2 I739 (comp4_0[27:27], i_4r0[27:27], i_4r1[27:27]);
  OR2 I740 (comp4_0[28:28], i_4r0[28:28], i_4r1[28:28]);
  OR2 I741 (comp4_0[29:29], i_4r0[29:29], i_4r1[29:29]);
  OR2 I742 (comp4_0[30:30], i_4r0[30:30], i_4r1[30:30]);
  OR2 I743 (comp4_0[31:31], i_4r0[31:31], i_4r1[31:31]);
  C3 I744 (simp5751_0[0:0], comp4_0[0:0], comp4_0[1:1], comp4_0[2:2]);
  C3 I745 (simp5751_0[1:1], comp4_0[3:3], comp4_0[4:4], comp4_0[5:5]);
  C3 I746 (simp5751_0[2:2], comp4_0[6:6], comp4_0[7:7], comp4_0[8:8]);
  C3 I747 (simp5751_0[3:3], comp4_0[9:9], comp4_0[10:10], comp4_0[11:11]);
  C3 I748 (simp5751_0[4:4], comp4_0[12:12], comp4_0[13:13], comp4_0[14:14]);
  C3 I749 (simp5751_0[5:5], comp4_0[15:15], comp4_0[16:16], comp4_0[17:17]);
  C3 I750 (simp5751_0[6:6], comp4_0[18:18], comp4_0[19:19], comp4_0[20:20]);
  C3 I751 (simp5751_0[7:7], comp4_0[21:21], comp4_0[22:22], comp4_0[23:23]);
  C3 I752 (simp5751_0[8:8], comp4_0[24:24], comp4_0[25:25], comp4_0[26:26]);
  C3 I753 (simp5751_0[9:9], comp4_0[27:27], comp4_0[28:28], comp4_0[29:29]);
  C2 I754 (simp5751_0[10:10], comp4_0[30:30], comp4_0[31:31]);
  C3 I755 (simp5752_0[0:0], simp5751_0[0:0], simp5751_0[1:1], simp5751_0[2:2]);
  C3 I756 (simp5752_0[1:1], simp5751_0[3:3], simp5751_0[4:4], simp5751_0[5:5]);
  C3 I757 (simp5752_0[2:2], simp5751_0[6:6], simp5751_0[7:7], simp5751_0[8:8]);
  C2 I758 (simp5752_0[3:3], simp5751_0[9:9], simp5751_0[10:10]);
  C3 I759 (simp5753_0[0:0], simp5752_0[0:0], simp5752_0[1:1], simp5752_0[2:2]);
  BUFF I760 (simp5753_0[1:1], simp5752_0[3:3]);
  C2 I761 (icomp_4, simp5753_0[0:0], simp5753_0[1:1]);
  C2R I762 (choice_0, icomp_0, nchosen_0, reset);
  C2R I763 (choice_1, icomp_1, nchosen_0, reset);
  C2R I764 (choice_2, icomp_2, nchosen_0, reset);
  C2R I765 (choice_3, icomp_3, nchosen_0, reset);
  C2R I766 (choice_4, icomp_4, nchosen_0, reset);
  NOR3 I767 (simp5811_0[0:0], choice_0, choice_1, choice_2);
  NOR2 I768 (simp5811_0[1:1], choice_3, choice_4);
  NAND2 I769 (anychoice_0, simp5811_0[0:0], simp5811_0[1:1]);
  NOR2 I770 (nchosen_0, anychoice_0, o_0a);
  C2R I771 (i_0a, choice_0, o_0a, reset);
  C2R I772 (i_1a, choice_1, o_0a, reset);
  C2R I773 (i_2a, choice_2, o_0a, reset);
  C2R I774 (i_3a, choice_3, o_0a, reset);
  C2R I775 (i_4a, choice_4, o_0a, reset);
endmodule

// tkj0m0_0_0_0 TeakJ [Many [0,0,0,0],One 0]
module tkj0m0_0_0_0 (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, i_3r, i_3a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  output o_0r;
  input o_0a;
  input reset;
  wire [1:0] simp01_0;
  C3 I0 (simp01_0[0:0], i_0r, i_1r, i_2r);
  BUFF I1 (simp01_0[1:1], i_3r);
  C2 I2 (o_0r, simp01_0[0:0], simp01_0[1:1]);
  BUFF I3 (i_0a, o_0a);
  BUFF I4 (i_1a, o_0a);
  BUFF I5 (i_2a, o_0a);
  BUFF I6 (i_3a, o_0a);
endmodule

// tko2m1_1api0w1b_2api1w1b_3andt1o0w1bt2o0w1b TeakO [
//     (1,TeakOAppend 1 [(0,0+:1)]),
//     (2,TeakOAppend 1 [(0,1+:1)]),
//     (3,TeakOp TeakOpAnd [(1,0+:1),(2,0+:1)])] [One 2,One 1]
module tko2m1_1api0w1b_2api1w1b_3andt1o0w1bt2o0w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire termf_1;
  wire termf_2;
  wire termt_1;
  wire termt_2;
  wire [3:0] op3_0_0;
  BUFF I0 (termf_1, i_0r0[0:0]);
  BUFF I1 (termt_1, i_0r1[0:0]);
  BUFF I2 (termf_2, i_0r0[1:1]);
  BUFF I3 (termt_2, i_0r1[1:1]);
  C2 I4 (op3_0_0[0:0], termf_2, termf_1);
  C2 I5 (op3_0_0[1:1], termf_2, termt_1);
  C2 I6 (op3_0_0[2:2], termt_2, termf_1);
  C2 I7 (op3_0_0[3:3], termt_2, termt_1);
  OR3 I8 (o_0r0, op3_0_0[0:0], op3_0_0[1:1], op3_0_0[2:2]);
  BUFF I9 (o_0r1, op3_0_0[3:3]);
  BUFF I10 (i_0a, o_0a);
endmodule

// tko2m1_1api0w1b_2api1w1b_3ort1o0w1bt2o0w1b TeakO [
//     (1,TeakOAppend 1 [(0,0+:1)]),
//     (2,TeakOAppend 1 [(0,1+:1)]),
//     (3,TeakOp TeakOpOr [(1,0+:1),(2,0+:1)])] [One 2,One 1]
module tko2m1_1api0w1b_2api1w1b_3ort1o0w1bt2o0w1b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire termf_1;
  wire termf_2;
  wire termt_1;
  wire termt_2;
  wire [3:0] op3_0_0;
  BUFF I0 (termf_1, i_0r0[0:0]);
  BUFF I1 (termt_1, i_0r1[0:0]);
  BUFF I2 (termf_2, i_0r0[1:1]);
  BUFF I3 (termt_2, i_0r1[1:1]);
  C2 I4 (op3_0_0[0:0], termf_2, termf_1);
  C2 I5 (op3_0_0[1:1], termf_2, termt_1);
  C2 I6 (op3_0_0[2:2], termt_2, termf_1);
  C2 I7 (op3_0_0[3:3], termt_2, termt_1);
  BUFF I8 (o_0r0, op3_0_0[0:0]);
  OR3 I9 (o_0r1, op3_0_0[1:1], op3_0_0[2:2], op3_0_0[3:3]);
  BUFF I10 (i_0a, o_0a);
endmodule

// tks4_o0w4_0m8o0w0_1m9o0w0_2mao0w0_3mbo0w0_4mco0w0_5mdo0w0_6meo0w0_7mfo0w0 TeakS (0+:4) [([Imp 0 0,Im
//   p 8 0],0),([Imp 1 0,Imp 9 0],0),([Imp 2 0,Imp 10 0],0),([Imp 3 0,Imp 11 0],0),([Imp 4 0,Imp 12 0],0)
//   ,([Imp 5 0,Imp 13 0],0),([Imp 6 0,Imp 14 0],0),([Imp 7 0,Imp 15 0],0)] [One 4,Many [0,0,0,0,0,0,0,0]
//   ]
module tks4_o0w4_0m8o0w0_1m9o0w0_2mao0w0_3mbo0w0_4mco0w0_5mdo0w0_6meo0w0_7mfo0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, o_5r, o_5a, o_6r, o_6a, o_7r, o_7a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  output o_7r;
  input o_7a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire sel_4;
  wire sel_5;
  wire sel_6;
  wire sel_7;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire gsel_4;
  wire gsel_5;
  wire gsel_6;
  wire gsel_7;
  wire oack_0;
  wire [1:0] match0_0;
  wire [1:0] simp201_0;
  wire [1:0] simp211_0;
  wire [1:0] match1_0;
  wire [1:0] simp241_0;
  wire [1:0] simp251_0;
  wire [1:0] match2_0;
  wire [1:0] simp281_0;
  wire [1:0] simp291_0;
  wire [1:0] match3_0;
  wire [1:0] simp321_0;
  wire [1:0] simp331_0;
  wire [1:0] match4_0;
  wire [1:0] simp361_0;
  wire [1:0] simp371_0;
  wire [1:0] match5_0;
  wire [1:0] simp401_0;
  wire [1:0] simp411_0;
  wire [1:0] match6_0;
  wire [1:0] simp441_0;
  wire [1:0] simp451_0;
  wire [1:0] match7_0;
  wire [1:0] simp481_0;
  wire [1:0] simp491_0;
  wire [3:0] comp_0;
  wire [1:0] simp631_0;
  wire [2:0] simp721_0;
  OR2 I0 (sel_0, match0_0[0:0], match0_0[1:1]);
  C3 I1 (simp201_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I2 (simp201_0[1:1], i_0r0[3:3]);
  C2 I3 (match0_0[0:0], simp201_0[0:0], simp201_0[1:1]);
  C3 I4 (simp211_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I5 (simp211_0[1:1], i_0r1[3:3]);
  C2 I6 (match0_0[1:1], simp211_0[0:0], simp211_0[1:1]);
  OR2 I7 (sel_1, match1_0[0:0], match1_0[1:1]);
  C3 I8 (simp241_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I9 (simp241_0[1:1], i_0r0[3:3]);
  C2 I10 (match1_0[0:0], simp241_0[0:0], simp241_0[1:1]);
  C3 I11 (simp251_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I12 (simp251_0[1:1], i_0r1[3:3]);
  C2 I13 (match1_0[1:1], simp251_0[0:0], simp251_0[1:1]);
  OR2 I14 (sel_2, match2_0[0:0], match2_0[1:1]);
  C3 I15 (simp281_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I16 (simp281_0[1:1], i_0r0[3:3]);
  C2 I17 (match2_0[0:0], simp281_0[0:0], simp281_0[1:1]);
  C3 I18 (simp291_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I19 (simp291_0[1:1], i_0r1[3:3]);
  C2 I20 (match2_0[1:1], simp291_0[0:0], simp291_0[1:1]);
  OR2 I21 (sel_3, match3_0[0:0], match3_0[1:1]);
  C3 I22 (simp321_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I23 (simp321_0[1:1], i_0r0[3:3]);
  C2 I24 (match3_0[0:0], simp321_0[0:0], simp321_0[1:1]);
  C3 I25 (simp331_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I26 (simp331_0[1:1], i_0r1[3:3]);
  C2 I27 (match3_0[1:1], simp331_0[0:0], simp331_0[1:1]);
  OR2 I28 (sel_4, match4_0[0:0], match4_0[1:1]);
  C3 I29 (simp361_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I30 (simp361_0[1:1], i_0r0[3:3]);
  C2 I31 (match4_0[0:0], simp361_0[0:0], simp361_0[1:1]);
  C3 I32 (simp371_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I33 (simp371_0[1:1], i_0r1[3:3]);
  C2 I34 (match4_0[1:1], simp371_0[0:0], simp371_0[1:1]);
  OR2 I35 (sel_5, match5_0[0:0], match5_0[1:1]);
  C3 I36 (simp401_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I37 (simp401_0[1:1], i_0r0[3:3]);
  C2 I38 (match5_0[0:0], simp401_0[0:0], simp401_0[1:1]);
  C3 I39 (simp411_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I40 (simp411_0[1:1], i_0r1[3:3]);
  C2 I41 (match5_0[1:1], simp411_0[0:0], simp411_0[1:1]);
  OR2 I42 (sel_6, match6_0[0:0], match6_0[1:1]);
  C3 I43 (simp441_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I44 (simp441_0[1:1], i_0r0[3:3]);
  C2 I45 (match6_0[0:0], simp441_0[0:0], simp441_0[1:1]);
  C3 I46 (simp451_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I47 (simp451_0[1:1], i_0r1[3:3]);
  C2 I48 (match6_0[1:1], simp451_0[0:0], simp451_0[1:1]);
  OR2 I49 (sel_7, match7_0[0:0], match7_0[1:1]);
  C3 I50 (simp481_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I51 (simp481_0[1:1], i_0r0[3:3]);
  C2 I52 (match7_0[0:0], simp481_0[0:0], simp481_0[1:1]);
  C3 I53 (simp491_0[0:0], i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I54 (simp491_0[1:1], i_0r1[3:3]);
  C2 I55 (match7_0[1:1], simp491_0[0:0], simp491_0[1:1]);
  C2 I56 (gsel_0, sel_0, icomplete_0);
  C2 I57 (gsel_1, sel_1, icomplete_0);
  C2 I58 (gsel_2, sel_2, icomplete_0);
  C2 I59 (gsel_3, sel_3, icomplete_0);
  C2 I60 (gsel_4, sel_4, icomplete_0);
  C2 I61 (gsel_5, sel_5, icomplete_0);
  C2 I62 (gsel_6, sel_6, icomplete_0);
  C2 I63 (gsel_7, sel_7, icomplete_0);
  OR2 I64 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I65 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I66 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I67 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  C3 I68 (simp631_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  BUFF I69 (simp631_0[1:1], comp_0[3:3]);
  C2 I70 (icomplete_0, simp631_0[0:0], simp631_0[1:1]);
  BUFF I71 (o_0r, gsel_0);
  BUFF I72 (o_1r, gsel_1);
  BUFF I73 (o_2r, gsel_2);
  BUFF I74 (o_3r, gsel_3);
  BUFF I75 (o_4r, gsel_4);
  BUFF I76 (o_5r, gsel_5);
  BUFF I77 (o_6r, gsel_6);
  BUFF I78 (o_7r, gsel_7);
  NOR3 I79 (simp721_0[0:0], o_0a, o_1a, o_2a);
  NOR3 I80 (simp721_0[1:1], o_3a, o_4a, o_5a);
  NOR2 I81 (simp721_0[2:2], o_6a, o_7a);
  NAND3 I82 (oack_0, simp721_0[0:0], simp721_0[1:1], simp721_0[2:2]);
  C2 I83 (i_0a, oack_0, icomplete_0);
endmodule

// tko64m33_1api0w32b_2api32w32b_3nm1b0_4apt1o0w32bt3o0w1b_5nm1b0_6apt2o0w32bt5o0w1b_7addt4o0w33bt6o0w3
//   3b TeakO [
//     (1,TeakOAppend 1 [(0,0+:32)]),
//     (2,TeakOAppend 1 [(0,32+:32)]),
//     (3,TeakOConstant 1 0),
//     (4,TeakOAppend 1 [(1,0+:32),(3,0+:1)]),
//     (5,TeakOConstant 1 0),
//     (6,TeakOAppend 1 [(2,0+:32),(5,0+:1)]),
//     (7,TeakOp TeakOpAdd [(4,0+:33),(6,0+:33)])] [One 64,One 33]
module tko64m33_1api0w32b_2api32w32b_3nm1b0_4apt1o0w32bt3o0w1b_5nm1b0_6apt2o0w32bt5o0w1b_7addt4o0w33bt6o0w33b (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, reset);
  input [63:0] i_0r0;
  input [63:0] i_0r1;
  output i_0a;
  output [32:0] o_0r0;
  output [32:0] o_0r1;
  input o_0a;
  input reset;
  wire go_0;
  wire [63:0] gocomp_0;
  wire [21:0] simp661_0;
  wire [7:0] simp662_0;
  wire [2:0] simp663_0;
  wire [31:0] termf_1;
  wire [31:0] termf_2;
  wire termf_3;
  wire [32:0] termf_4;
  wire termf_5;
  wire [32:0] termf_6;
  wire [31:0] termt_1;
  wire [31:0] termt_2;
  wire termt_3;
  wire [32:0] termt_4;
  wire termt_5;
  wire [32:0] termt_6;
  wire [32:0] cf7__0;
  wire [32:0] ct7__0;
  wire [3:0] ha7__0;
  wire [7:0] fa7_1min_0;
  wire [1:0] simp3651_0;
  wire [1:0] simp3661_0;
  wire [7:0] fa7_2min_0;
  wire [1:0] simp3781_0;
  wire [1:0] simp3791_0;
  wire [7:0] fa7_3min_0;
  wire [1:0] simp3911_0;
  wire [1:0] simp3921_0;
  wire [7:0] fa7_4min_0;
  wire [1:0] simp4041_0;
  wire [1:0] simp4051_0;
  wire [7:0] fa7_5min_0;
  wire [1:0] simp4171_0;
  wire [1:0] simp4181_0;
  wire [7:0] fa7_6min_0;
  wire [1:0] simp4301_0;
  wire [1:0] simp4311_0;
  wire [7:0] fa7_7min_0;
  wire [1:0] simp4431_0;
  wire [1:0] simp4441_0;
  wire [7:0] fa7_8min_0;
  wire [1:0] simp4561_0;
  wire [1:0] simp4571_0;
  wire [7:0] fa7_9min_0;
  wire [1:0] simp4691_0;
  wire [1:0] simp4701_0;
  wire [7:0] fa7_10min_0;
  wire [1:0] simp4821_0;
  wire [1:0] simp4831_0;
  wire [7:0] fa7_11min_0;
  wire [1:0] simp4951_0;
  wire [1:0] simp4961_0;
  wire [7:0] fa7_12min_0;
  wire [1:0] simp5081_0;
  wire [1:0] simp5091_0;
  wire [7:0] fa7_13min_0;
  wire [1:0] simp5211_0;
  wire [1:0] simp5221_0;
  wire [7:0] fa7_14min_0;
  wire [1:0] simp5341_0;
  wire [1:0] simp5351_0;
  wire [7:0] fa7_15min_0;
  wire [1:0] simp5471_0;
  wire [1:0] simp5481_0;
  wire [7:0] fa7_16min_0;
  wire [1:0] simp5601_0;
  wire [1:0] simp5611_0;
  wire [7:0] fa7_17min_0;
  wire [1:0] simp5731_0;
  wire [1:0] simp5741_0;
  wire [7:0] fa7_18min_0;
  wire [1:0] simp5861_0;
  wire [1:0] simp5871_0;
  wire [7:0] fa7_19min_0;
  wire [1:0] simp5991_0;
  wire [1:0] simp6001_0;
  wire [7:0] fa7_20min_0;
  wire [1:0] simp6121_0;
  wire [1:0] simp6131_0;
  wire [7:0] fa7_21min_0;
  wire [1:0] simp6251_0;
  wire [1:0] simp6261_0;
  wire [7:0] fa7_22min_0;
  wire [1:0] simp6381_0;
  wire [1:0] simp6391_0;
  wire [7:0] fa7_23min_0;
  wire [1:0] simp6511_0;
  wire [1:0] simp6521_0;
  wire [7:0] fa7_24min_0;
  wire [1:0] simp6641_0;
  wire [1:0] simp6651_0;
  wire [7:0] fa7_25min_0;
  wire [1:0] simp6771_0;
  wire [1:0] simp6781_0;
  wire [7:0] fa7_26min_0;
  wire [1:0] simp6901_0;
  wire [1:0] simp6911_0;
  wire [7:0] fa7_27min_0;
  wire [1:0] simp7031_0;
  wire [1:0] simp7041_0;
  wire [7:0] fa7_28min_0;
  wire [1:0] simp7161_0;
  wire [1:0] simp7171_0;
  wire [7:0] fa7_29min_0;
  wire [1:0] simp7291_0;
  wire [1:0] simp7301_0;
  wire [7:0] fa7_30min_0;
  wire [1:0] simp7421_0;
  wire [1:0] simp7431_0;
  wire [7:0] fa7_31min_0;
  wire [1:0] simp7551_0;
  wire [1:0] simp7561_0;
  wire [7:0] fa7_32min_0;
  wire [1:0] simp7681_0;
  wire [1:0] simp7691_0;
  OR2 I0 (gocomp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (gocomp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I2 (gocomp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I3 (gocomp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I4 (gocomp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I5 (gocomp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I6 (gocomp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I7 (gocomp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I8 (gocomp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I9 (gocomp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I10 (gocomp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I11 (gocomp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I12 (gocomp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I13 (gocomp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I14 (gocomp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I15 (gocomp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I16 (gocomp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I17 (gocomp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I18 (gocomp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I19 (gocomp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I20 (gocomp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I21 (gocomp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I22 (gocomp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I23 (gocomp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I24 (gocomp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I25 (gocomp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I26 (gocomp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I27 (gocomp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I28 (gocomp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I29 (gocomp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I30 (gocomp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I31 (gocomp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I32 (gocomp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  OR2 I33 (gocomp_0[33:33], i_0r0[33:33], i_0r1[33:33]);
  OR2 I34 (gocomp_0[34:34], i_0r0[34:34], i_0r1[34:34]);
  OR2 I35 (gocomp_0[35:35], i_0r0[35:35], i_0r1[35:35]);
  OR2 I36 (gocomp_0[36:36], i_0r0[36:36], i_0r1[36:36]);
  OR2 I37 (gocomp_0[37:37], i_0r0[37:37], i_0r1[37:37]);
  OR2 I38 (gocomp_0[38:38], i_0r0[38:38], i_0r1[38:38]);
  OR2 I39 (gocomp_0[39:39], i_0r0[39:39], i_0r1[39:39]);
  OR2 I40 (gocomp_0[40:40], i_0r0[40:40], i_0r1[40:40]);
  OR2 I41 (gocomp_0[41:41], i_0r0[41:41], i_0r1[41:41]);
  OR2 I42 (gocomp_0[42:42], i_0r0[42:42], i_0r1[42:42]);
  OR2 I43 (gocomp_0[43:43], i_0r0[43:43], i_0r1[43:43]);
  OR2 I44 (gocomp_0[44:44], i_0r0[44:44], i_0r1[44:44]);
  OR2 I45 (gocomp_0[45:45], i_0r0[45:45], i_0r1[45:45]);
  OR2 I46 (gocomp_0[46:46], i_0r0[46:46], i_0r1[46:46]);
  OR2 I47 (gocomp_0[47:47], i_0r0[47:47], i_0r1[47:47]);
  OR2 I48 (gocomp_0[48:48], i_0r0[48:48], i_0r1[48:48]);
  OR2 I49 (gocomp_0[49:49], i_0r0[49:49], i_0r1[49:49]);
  OR2 I50 (gocomp_0[50:50], i_0r0[50:50], i_0r1[50:50]);
  OR2 I51 (gocomp_0[51:51], i_0r0[51:51], i_0r1[51:51]);
  OR2 I52 (gocomp_0[52:52], i_0r0[52:52], i_0r1[52:52]);
  OR2 I53 (gocomp_0[53:53], i_0r0[53:53], i_0r1[53:53]);
  OR2 I54 (gocomp_0[54:54], i_0r0[54:54], i_0r1[54:54]);
  OR2 I55 (gocomp_0[55:55], i_0r0[55:55], i_0r1[55:55]);
  OR2 I56 (gocomp_0[56:56], i_0r0[56:56], i_0r1[56:56]);
  OR2 I57 (gocomp_0[57:57], i_0r0[57:57], i_0r1[57:57]);
  OR2 I58 (gocomp_0[58:58], i_0r0[58:58], i_0r1[58:58]);
  OR2 I59 (gocomp_0[59:59], i_0r0[59:59], i_0r1[59:59]);
  OR2 I60 (gocomp_0[60:60], i_0r0[60:60], i_0r1[60:60]);
  OR2 I61 (gocomp_0[61:61], i_0r0[61:61], i_0r1[61:61]);
  OR2 I62 (gocomp_0[62:62], i_0r0[62:62], i_0r1[62:62]);
  OR2 I63 (gocomp_0[63:63], i_0r0[63:63], i_0r1[63:63]);
  C3 I64 (simp661_0[0:0], gocomp_0[0:0], gocomp_0[1:1], gocomp_0[2:2]);
  C3 I65 (simp661_0[1:1], gocomp_0[3:3], gocomp_0[4:4], gocomp_0[5:5]);
  C3 I66 (simp661_0[2:2], gocomp_0[6:6], gocomp_0[7:7], gocomp_0[8:8]);
  C3 I67 (simp661_0[3:3], gocomp_0[9:9], gocomp_0[10:10], gocomp_0[11:11]);
  C3 I68 (simp661_0[4:4], gocomp_0[12:12], gocomp_0[13:13], gocomp_0[14:14]);
  C3 I69 (simp661_0[5:5], gocomp_0[15:15], gocomp_0[16:16], gocomp_0[17:17]);
  C3 I70 (simp661_0[6:6], gocomp_0[18:18], gocomp_0[19:19], gocomp_0[20:20]);
  C3 I71 (simp661_0[7:7], gocomp_0[21:21], gocomp_0[22:22], gocomp_0[23:23]);
  C3 I72 (simp661_0[8:8], gocomp_0[24:24], gocomp_0[25:25], gocomp_0[26:26]);
  C3 I73 (simp661_0[9:9], gocomp_0[27:27], gocomp_0[28:28], gocomp_0[29:29]);
  C3 I74 (simp661_0[10:10], gocomp_0[30:30], gocomp_0[31:31], gocomp_0[32:32]);
  C3 I75 (simp661_0[11:11], gocomp_0[33:33], gocomp_0[34:34], gocomp_0[35:35]);
  C3 I76 (simp661_0[12:12], gocomp_0[36:36], gocomp_0[37:37], gocomp_0[38:38]);
  C3 I77 (simp661_0[13:13], gocomp_0[39:39], gocomp_0[40:40], gocomp_0[41:41]);
  C3 I78 (simp661_0[14:14], gocomp_0[42:42], gocomp_0[43:43], gocomp_0[44:44]);
  C3 I79 (simp661_0[15:15], gocomp_0[45:45], gocomp_0[46:46], gocomp_0[47:47]);
  C3 I80 (simp661_0[16:16], gocomp_0[48:48], gocomp_0[49:49], gocomp_0[50:50]);
  C3 I81 (simp661_0[17:17], gocomp_0[51:51], gocomp_0[52:52], gocomp_0[53:53]);
  C3 I82 (simp661_0[18:18], gocomp_0[54:54], gocomp_0[55:55], gocomp_0[56:56]);
  C3 I83 (simp661_0[19:19], gocomp_0[57:57], gocomp_0[58:58], gocomp_0[59:59]);
  C3 I84 (simp661_0[20:20], gocomp_0[60:60], gocomp_0[61:61], gocomp_0[62:62]);
  BUFF I85 (simp661_0[21:21], gocomp_0[63:63]);
  C3 I86 (simp662_0[0:0], simp661_0[0:0], simp661_0[1:1], simp661_0[2:2]);
  C3 I87 (simp662_0[1:1], simp661_0[3:3], simp661_0[4:4], simp661_0[5:5]);
  C3 I88 (simp662_0[2:2], simp661_0[6:6], simp661_0[7:7], simp661_0[8:8]);
  C3 I89 (simp662_0[3:3], simp661_0[9:9], simp661_0[10:10], simp661_0[11:11]);
  C3 I90 (simp662_0[4:4], simp661_0[12:12], simp661_0[13:13], simp661_0[14:14]);
  C3 I91 (simp662_0[5:5], simp661_0[15:15], simp661_0[16:16], simp661_0[17:17]);
  C3 I92 (simp662_0[6:6], simp661_0[18:18], simp661_0[19:19], simp661_0[20:20]);
  BUFF I93 (simp662_0[7:7], simp661_0[21:21]);
  C3 I94 (simp663_0[0:0], simp662_0[0:0], simp662_0[1:1], simp662_0[2:2]);
  C3 I95 (simp663_0[1:1], simp662_0[3:3], simp662_0[4:4], simp662_0[5:5]);
  C2 I96 (simp663_0[2:2], simp662_0[6:6], simp662_0[7:7]);
  C3 I97 (go_0, simp663_0[0:0], simp663_0[1:1], simp663_0[2:2]);
  BUFF I98 (termf_1[0:0], i_0r0[0:0]);
  BUFF I99 (termf_1[1:1], i_0r0[1:1]);
  BUFF I100 (termf_1[2:2], i_0r0[2:2]);
  BUFF I101 (termf_1[3:3], i_0r0[3:3]);
  BUFF I102 (termf_1[4:4], i_0r0[4:4]);
  BUFF I103 (termf_1[5:5], i_0r0[5:5]);
  BUFF I104 (termf_1[6:6], i_0r0[6:6]);
  BUFF I105 (termf_1[7:7], i_0r0[7:7]);
  BUFF I106 (termf_1[8:8], i_0r0[8:8]);
  BUFF I107 (termf_1[9:9], i_0r0[9:9]);
  BUFF I108 (termf_1[10:10], i_0r0[10:10]);
  BUFF I109 (termf_1[11:11], i_0r0[11:11]);
  BUFF I110 (termf_1[12:12], i_0r0[12:12]);
  BUFF I111 (termf_1[13:13], i_0r0[13:13]);
  BUFF I112 (termf_1[14:14], i_0r0[14:14]);
  BUFF I113 (termf_1[15:15], i_0r0[15:15]);
  BUFF I114 (termf_1[16:16], i_0r0[16:16]);
  BUFF I115 (termf_1[17:17], i_0r0[17:17]);
  BUFF I116 (termf_1[18:18], i_0r0[18:18]);
  BUFF I117 (termf_1[19:19], i_0r0[19:19]);
  BUFF I118 (termf_1[20:20], i_0r0[20:20]);
  BUFF I119 (termf_1[21:21], i_0r0[21:21]);
  BUFF I120 (termf_1[22:22], i_0r0[22:22]);
  BUFF I121 (termf_1[23:23], i_0r0[23:23]);
  BUFF I122 (termf_1[24:24], i_0r0[24:24]);
  BUFF I123 (termf_1[25:25], i_0r0[25:25]);
  BUFF I124 (termf_1[26:26], i_0r0[26:26]);
  BUFF I125 (termf_1[27:27], i_0r0[27:27]);
  BUFF I126 (termf_1[28:28], i_0r0[28:28]);
  BUFF I127 (termf_1[29:29], i_0r0[29:29]);
  BUFF I128 (termf_1[30:30], i_0r0[30:30]);
  BUFF I129 (termf_1[31:31], i_0r0[31:31]);
  BUFF I130 (termt_1[0:0], i_0r1[0:0]);
  BUFF I131 (termt_1[1:1], i_0r1[1:1]);
  BUFF I132 (termt_1[2:2], i_0r1[2:2]);
  BUFF I133 (termt_1[3:3], i_0r1[3:3]);
  BUFF I134 (termt_1[4:4], i_0r1[4:4]);
  BUFF I135 (termt_1[5:5], i_0r1[5:5]);
  BUFF I136 (termt_1[6:6], i_0r1[6:6]);
  BUFF I137 (termt_1[7:7], i_0r1[7:7]);
  BUFF I138 (termt_1[8:8], i_0r1[8:8]);
  BUFF I139 (termt_1[9:9], i_0r1[9:9]);
  BUFF I140 (termt_1[10:10], i_0r1[10:10]);
  BUFF I141 (termt_1[11:11], i_0r1[11:11]);
  BUFF I142 (termt_1[12:12], i_0r1[12:12]);
  BUFF I143 (termt_1[13:13], i_0r1[13:13]);
  BUFF I144 (termt_1[14:14], i_0r1[14:14]);
  BUFF I145 (termt_1[15:15], i_0r1[15:15]);
  BUFF I146 (termt_1[16:16], i_0r1[16:16]);
  BUFF I147 (termt_1[17:17], i_0r1[17:17]);
  BUFF I148 (termt_1[18:18], i_0r1[18:18]);
  BUFF I149 (termt_1[19:19], i_0r1[19:19]);
  BUFF I150 (termt_1[20:20], i_0r1[20:20]);
  BUFF I151 (termt_1[21:21], i_0r1[21:21]);
  BUFF I152 (termt_1[22:22], i_0r1[22:22]);
  BUFF I153 (termt_1[23:23], i_0r1[23:23]);
  BUFF I154 (termt_1[24:24], i_0r1[24:24]);
  BUFF I155 (termt_1[25:25], i_0r1[25:25]);
  BUFF I156 (termt_1[26:26], i_0r1[26:26]);
  BUFF I157 (termt_1[27:27], i_0r1[27:27]);
  BUFF I158 (termt_1[28:28], i_0r1[28:28]);
  BUFF I159 (termt_1[29:29], i_0r1[29:29]);
  BUFF I160 (termt_1[30:30], i_0r1[30:30]);
  BUFF I161 (termt_1[31:31], i_0r1[31:31]);
  BUFF I162 (termf_2[0:0], i_0r0[32:32]);
  BUFF I163 (termf_2[1:1], i_0r0[33:33]);
  BUFF I164 (termf_2[2:2], i_0r0[34:34]);
  BUFF I165 (termf_2[3:3], i_0r0[35:35]);
  BUFF I166 (termf_2[4:4], i_0r0[36:36]);
  BUFF I167 (termf_2[5:5], i_0r0[37:37]);
  BUFF I168 (termf_2[6:6], i_0r0[38:38]);
  BUFF I169 (termf_2[7:7], i_0r0[39:39]);
  BUFF I170 (termf_2[8:8], i_0r0[40:40]);
  BUFF I171 (termf_2[9:9], i_0r0[41:41]);
  BUFF I172 (termf_2[10:10], i_0r0[42:42]);
  BUFF I173 (termf_2[11:11], i_0r0[43:43]);
  BUFF I174 (termf_2[12:12], i_0r0[44:44]);
  BUFF I175 (termf_2[13:13], i_0r0[45:45]);
  BUFF I176 (termf_2[14:14], i_0r0[46:46]);
  BUFF I177 (termf_2[15:15], i_0r0[47:47]);
  BUFF I178 (termf_2[16:16], i_0r0[48:48]);
  BUFF I179 (termf_2[17:17], i_0r0[49:49]);
  BUFF I180 (termf_2[18:18], i_0r0[50:50]);
  BUFF I181 (termf_2[19:19], i_0r0[51:51]);
  BUFF I182 (termf_2[20:20], i_0r0[52:52]);
  BUFF I183 (termf_2[21:21], i_0r0[53:53]);
  BUFF I184 (termf_2[22:22], i_0r0[54:54]);
  BUFF I185 (termf_2[23:23], i_0r0[55:55]);
  BUFF I186 (termf_2[24:24], i_0r0[56:56]);
  BUFF I187 (termf_2[25:25], i_0r0[57:57]);
  BUFF I188 (termf_2[26:26], i_0r0[58:58]);
  BUFF I189 (termf_2[27:27], i_0r0[59:59]);
  BUFF I190 (termf_2[28:28], i_0r0[60:60]);
  BUFF I191 (termf_2[29:29], i_0r0[61:61]);
  BUFF I192 (termf_2[30:30], i_0r0[62:62]);
  BUFF I193 (termf_2[31:31], i_0r0[63:63]);
  BUFF I194 (termt_2[0:0], i_0r1[32:32]);
  BUFF I195 (termt_2[1:1], i_0r1[33:33]);
  BUFF I196 (termt_2[2:2], i_0r1[34:34]);
  BUFF I197 (termt_2[3:3], i_0r1[35:35]);
  BUFF I198 (termt_2[4:4], i_0r1[36:36]);
  BUFF I199 (termt_2[5:5], i_0r1[37:37]);
  BUFF I200 (termt_2[6:6], i_0r1[38:38]);
  BUFF I201 (termt_2[7:7], i_0r1[39:39]);
  BUFF I202 (termt_2[8:8], i_0r1[40:40]);
  BUFF I203 (termt_2[9:9], i_0r1[41:41]);
  BUFF I204 (termt_2[10:10], i_0r1[42:42]);
  BUFF I205 (termt_2[11:11], i_0r1[43:43]);
  BUFF I206 (termt_2[12:12], i_0r1[44:44]);
  BUFF I207 (termt_2[13:13], i_0r1[45:45]);
  BUFF I208 (termt_2[14:14], i_0r1[46:46]);
  BUFF I209 (termt_2[15:15], i_0r1[47:47]);
  BUFF I210 (termt_2[16:16], i_0r1[48:48]);
  BUFF I211 (termt_2[17:17], i_0r1[49:49]);
  BUFF I212 (termt_2[18:18], i_0r1[50:50]);
  BUFF I213 (termt_2[19:19], i_0r1[51:51]);
  BUFF I214 (termt_2[20:20], i_0r1[52:52]);
  BUFF I215 (termt_2[21:21], i_0r1[53:53]);
  BUFF I216 (termt_2[22:22], i_0r1[54:54]);
  BUFF I217 (termt_2[23:23], i_0r1[55:55]);
  BUFF I218 (termt_2[24:24], i_0r1[56:56]);
  BUFF I219 (termt_2[25:25], i_0r1[57:57]);
  BUFF I220 (termt_2[26:26], i_0r1[58:58]);
  BUFF I221 (termt_2[27:27], i_0r1[59:59]);
  BUFF I222 (termt_2[28:28], i_0r1[60:60]);
  BUFF I223 (termt_2[29:29], i_0r1[61:61]);
  BUFF I224 (termt_2[30:30], i_0r1[62:62]);
  BUFF I225 (termt_2[31:31], i_0r1[63:63]);
  BUFF I226 (termf_3, go_0);
  GND I227 (termt_3);
  BUFF I228 (termf_4[0:0], termf_1[0:0]);
  BUFF I229 (termf_4[1:1], termf_1[1:1]);
  BUFF I230 (termf_4[2:2], termf_1[2:2]);
  BUFF I231 (termf_4[3:3], termf_1[3:3]);
  BUFF I232 (termf_4[4:4], termf_1[4:4]);
  BUFF I233 (termf_4[5:5], termf_1[5:5]);
  BUFF I234 (termf_4[6:6], termf_1[6:6]);
  BUFF I235 (termf_4[7:7], termf_1[7:7]);
  BUFF I236 (termf_4[8:8], termf_1[8:8]);
  BUFF I237 (termf_4[9:9], termf_1[9:9]);
  BUFF I238 (termf_4[10:10], termf_1[10:10]);
  BUFF I239 (termf_4[11:11], termf_1[11:11]);
  BUFF I240 (termf_4[12:12], termf_1[12:12]);
  BUFF I241 (termf_4[13:13], termf_1[13:13]);
  BUFF I242 (termf_4[14:14], termf_1[14:14]);
  BUFF I243 (termf_4[15:15], termf_1[15:15]);
  BUFF I244 (termf_4[16:16], termf_1[16:16]);
  BUFF I245 (termf_4[17:17], termf_1[17:17]);
  BUFF I246 (termf_4[18:18], termf_1[18:18]);
  BUFF I247 (termf_4[19:19], termf_1[19:19]);
  BUFF I248 (termf_4[20:20], termf_1[20:20]);
  BUFF I249 (termf_4[21:21], termf_1[21:21]);
  BUFF I250 (termf_4[22:22], termf_1[22:22]);
  BUFF I251 (termf_4[23:23], termf_1[23:23]);
  BUFF I252 (termf_4[24:24], termf_1[24:24]);
  BUFF I253 (termf_4[25:25], termf_1[25:25]);
  BUFF I254 (termf_4[26:26], termf_1[26:26]);
  BUFF I255 (termf_4[27:27], termf_1[27:27]);
  BUFF I256 (termf_4[28:28], termf_1[28:28]);
  BUFF I257 (termf_4[29:29], termf_1[29:29]);
  BUFF I258 (termf_4[30:30], termf_1[30:30]);
  BUFF I259 (termf_4[31:31], termf_1[31:31]);
  BUFF I260 (termf_4[32:32], termf_3);
  BUFF I261 (termt_4[0:0], termt_1[0:0]);
  BUFF I262 (termt_4[1:1], termt_1[1:1]);
  BUFF I263 (termt_4[2:2], termt_1[2:2]);
  BUFF I264 (termt_4[3:3], termt_1[3:3]);
  BUFF I265 (termt_4[4:4], termt_1[4:4]);
  BUFF I266 (termt_4[5:5], termt_1[5:5]);
  BUFF I267 (termt_4[6:6], termt_1[6:6]);
  BUFF I268 (termt_4[7:7], termt_1[7:7]);
  BUFF I269 (termt_4[8:8], termt_1[8:8]);
  BUFF I270 (termt_4[9:9], termt_1[9:9]);
  BUFF I271 (termt_4[10:10], termt_1[10:10]);
  BUFF I272 (termt_4[11:11], termt_1[11:11]);
  BUFF I273 (termt_4[12:12], termt_1[12:12]);
  BUFF I274 (termt_4[13:13], termt_1[13:13]);
  BUFF I275 (termt_4[14:14], termt_1[14:14]);
  BUFF I276 (termt_4[15:15], termt_1[15:15]);
  BUFF I277 (termt_4[16:16], termt_1[16:16]);
  BUFF I278 (termt_4[17:17], termt_1[17:17]);
  BUFF I279 (termt_4[18:18], termt_1[18:18]);
  BUFF I280 (termt_4[19:19], termt_1[19:19]);
  BUFF I281 (termt_4[20:20], termt_1[20:20]);
  BUFF I282 (termt_4[21:21], termt_1[21:21]);
  BUFF I283 (termt_4[22:22], termt_1[22:22]);
  BUFF I284 (termt_4[23:23], termt_1[23:23]);
  BUFF I285 (termt_4[24:24], termt_1[24:24]);
  BUFF I286 (termt_4[25:25], termt_1[25:25]);
  BUFF I287 (termt_4[26:26], termt_1[26:26]);
  BUFF I288 (termt_4[27:27], termt_1[27:27]);
  BUFF I289 (termt_4[28:28], termt_1[28:28]);
  BUFF I290 (termt_4[29:29], termt_1[29:29]);
  BUFF I291 (termt_4[30:30], termt_1[30:30]);
  BUFF I292 (termt_4[31:31], termt_1[31:31]);
  BUFF I293 (termt_4[32:32], termt_3);
  BUFF I294 (termf_5, go_0);
  GND I295 (termt_5);
  BUFF I296 (termf_6[0:0], termf_2[0:0]);
  BUFF I297 (termf_6[1:1], termf_2[1:1]);
  BUFF I298 (termf_6[2:2], termf_2[2:2]);
  BUFF I299 (termf_6[3:3], termf_2[3:3]);
  BUFF I300 (termf_6[4:4], termf_2[4:4]);
  BUFF I301 (termf_6[5:5], termf_2[5:5]);
  BUFF I302 (termf_6[6:6], termf_2[6:6]);
  BUFF I303 (termf_6[7:7], termf_2[7:7]);
  BUFF I304 (termf_6[8:8], termf_2[8:8]);
  BUFF I305 (termf_6[9:9], termf_2[9:9]);
  BUFF I306 (termf_6[10:10], termf_2[10:10]);
  BUFF I307 (termf_6[11:11], termf_2[11:11]);
  BUFF I308 (termf_6[12:12], termf_2[12:12]);
  BUFF I309 (termf_6[13:13], termf_2[13:13]);
  BUFF I310 (termf_6[14:14], termf_2[14:14]);
  BUFF I311 (termf_6[15:15], termf_2[15:15]);
  BUFF I312 (termf_6[16:16], termf_2[16:16]);
  BUFF I313 (termf_6[17:17], termf_2[17:17]);
  BUFF I314 (termf_6[18:18], termf_2[18:18]);
  BUFF I315 (termf_6[19:19], termf_2[19:19]);
  BUFF I316 (termf_6[20:20], termf_2[20:20]);
  BUFF I317 (termf_6[21:21], termf_2[21:21]);
  BUFF I318 (termf_6[22:22], termf_2[22:22]);
  BUFF I319 (termf_6[23:23], termf_2[23:23]);
  BUFF I320 (termf_6[24:24], termf_2[24:24]);
  BUFF I321 (termf_6[25:25], termf_2[25:25]);
  BUFF I322 (termf_6[26:26], termf_2[26:26]);
  BUFF I323 (termf_6[27:27], termf_2[27:27]);
  BUFF I324 (termf_6[28:28], termf_2[28:28]);
  BUFF I325 (termf_6[29:29], termf_2[29:29]);
  BUFF I326 (termf_6[30:30], termf_2[30:30]);
  BUFF I327 (termf_6[31:31], termf_2[31:31]);
  BUFF I328 (termf_6[32:32], termf_5);
  BUFF I329 (termt_6[0:0], termt_2[0:0]);
  BUFF I330 (termt_6[1:1], termt_2[1:1]);
  BUFF I331 (termt_6[2:2], termt_2[2:2]);
  BUFF I332 (termt_6[3:3], termt_2[3:3]);
  BUFF I333 (termt_6[4:4], termt_2[4:4]);
  BUFF I334 (termt_6[5:5], termt_2[5:5]);
  BUFF I335 (termt_6[6:6], termt_2[6:6]);
  BUFF I336 (termt_6[7:7], termt_2[7:7]);
  BUFF I337 (termt_6[8:8], termt_2[8:8]);
  BUFF I338 (termt_6[9:9], termt_2[9:9]);
  BUFF I339 (termt_6[10:10], termt_2[10:10]);
  BUFF I340 (termt_6[11:11], termt_2[11:11]);
  BUFF I341 (termt_6[12:12], termt_2[12:12]);
  BUFF I342 (termt_6[13:13], termt_2[13:13]);
  BUFF I343 (termt_6[14:14], termt_2[14:14]);
  BUFF I344 (termt_6[15:15], termt_2[15:15]);
  BUFF I345 (termt_6[16:16], termt_2[16:16]);
  BUFF I346 (termt_6[17:17], termt_2[17:17]);
  BUFF I347 (termt_6[18:18], termt_2[18:18]);
  BUFF I348 (termt_6[19:19], termt_2[19:19]);
  BUFF I349 (termt_6[20:20], termt_2[20:20]);
  BUFF I350 (termt_6[21:21], termt_2[21:21]);
  BUFF I351 (termt_6[22:22], termt_2[22:22]);
  BUFF I352 (termt_6[23:23], termt_2[23:23]);
  BUFF I353 (termt_6[24:24], termt_2[24:24]);
  BUFF I354 (termt_6[25:25], termt_2[25:25]);
  BUFF I355 (termt_6[26:26], termt_2[26:26]);
  BUFF I356 (termt_6[27:27], termt_2[27:27]);
  BUFF I357 (termt_6[28:28], termt_2[28:28]);
  BUFF I358 (termt_6[29:29], termt_2[29:29]);
  BUFF I359 (termt_6[30:30], termt_2[30:30]);
  BUFF I360 (termt_6[31:31], termt_2[31:31]);
  BUFF I361 (termt_6[32:32], termt_5);
  C2 I362 (ha7__0[0:0], termf_6[0:0], termf_4[0:0]);
  C2 I363 (ha7__0[1:1], termf_6[0:0], termt_4[0:0]);
  C2 I364 (ha7__0[2:2], termt_6[0:0], termf_4[0:0]);
  C2 I365 (ha7__0[3:3], termt_6[0:0], termt_4[0:0]);
  OR3 I366 (cf7__0[0:0], ha7__0[0:0], ha7__0[1:1], ha7__0[2:2]);
  BUFF I367 (ct7__0[0:0], ha7__0[3:3]);
  OR2 I368 (o_0r0[0:0], ha7__0[0:0], ha7__0[3:3]);
  OR2 I369 (o_0r1[0:0], ha7__0[1:1], ha7__0[2:2]);
  C3 I370 (fa7_1min_0[0:0], cf7__0[0:0], termf_6[1:1], termf_4[1:1]);
  C3 I371 (fa7_1min_0[1:1], cf7__0[0:0], termf_6[1:1], termt_4[1:1]);
  C3 I372 (fa7_1min_0[2:2], cf7__0[0:0], termt_6[1:1], termf_4[1:1]);
  C3 I373 (fa7_1min_0[3:3], cf7__0[0:0], termt_6[1:1], termt_4[1:1]);
  C3 I374 (fa7_1min_0[4:4], ct7__0[0:0], termf_6[1:1], termf_4[1:1]);
  C3 I375 (fa7_1min_0[5:5], ct7__0[0:0], termf_6[1:1], termt_4[1:1]);
  C3 I376 (fa7_1min_0[6:6], ct7__0[0:0], termt_6[1:1], termf_4[1:1]);
  C3 I377 (fa7_1min_0[7:7], ct7__0[0:0], termt_6[1:1], termt_4[1:1]);
  NOR3 I378 (simp3651_0[0:0], fa7_1min_0[0:0], fa7_1min_0[3:3], fa7_1min_0[5:5]);
  INV I379 (simp3651_0[1:1], fa7_1min_0[6:6]);
  NAND2 I380 (o_0r0[1:1], simp3651_0[0:0], simp3651_0[1:1]);
  NOR3 I381 (simp3661_0[0:0], fa7_1min_0[1:1], fa7_1min_0[2:2], fa7_1min_0[4:4]);
  INV I382 (simp3661_0[1:1], fa7_1min_0[7:7]);
  NAND2 I383 (o_0r1[1:1], simp3661_0[0:0], simp3661_0[1:1]);
  AO222 I384 (ct7__0[1:1], termt_4[1:1], termt_6[1:1], termt_4[1:1], ct7__0[0:0], termt_6[1:1], ct7__0[0:0]);
  AO222 I385 (cf7__0[1:1], termf_4[1:1], termf_6[1:1], termf_4[1:1], cf7__0[0:0], termf_6[1:1], cf7__0[0:0]);
  C3 I386 (fa7_2min_0[0:0], cf7__0[1:1], termf_6[2:2], termf_4[2:2]);
  C3 I387 (fa7_2min_0[1:1], cf7__0[1:1], termf_6[2:2], termt_4[2:2]);
  C3 I388 (fa7_2min_0[2:2], cf7__0[1:1], termt_6[2:2], termf_4[2:2]);
  C3 I389 (fa7_2min_0[3:3], cf7__0[1:1], termt_6[2:2], termt_4[2:2]);
  C3 I390 (fa7_2min_0[4:4], ct7__0[1:1], termf_6[2:2], termf_4[2:2]);
  C3 I391 (fa7_2min_0[5:5], ct7__0[1:1], termf_6[2:2], termt_4[2:2]);
  C3 I392 (fa7_2min_0[6:6], ct7__0[1:1], termt_6[2:2], termf_4[2:2]);
  C3 I393 (fa7_2min_0[7:7], ct7__0[1:1], termt_6[2:2], termt_4[2:2]);
  NOR3 I394 (simp3781_0[0:0], fa7_2min_0[0:0], fa7_2min_0[3:3], fa7_2min_0[5:5]);
  INV I395 (simp3781_0[1:1], fa7_2min_0[6:6]);
  NAND2 I396 (o_0r0[2:2], simp3781_0[0:0], simp3781_0[1:1]);
  NOR3 I397 (simp3791_0[0:0], fa7_2min_0[1:1], fa7_2min_0[2:2], fa7_2min_0[4:4]);
  INV I398 (simp3791_0[1:1], fa7_2min_0[7:7]);
  NAND2 I399 (o_0r1[2:2], simp3791_0[0:0], simp3791_0[1:1]);
  AO222 I400 (ct7__0[2:2], termt_4[2:2], termt_6[2:2], termt_4[2:2], ct7__0[1:1], termt_6[2:2], ct7__0[1:1]);
  AO222 I401 (cf7__0[2:2], termf_4[2:2], termf_6[2:2], termf_4[2:2], cf7__0[1:1], termf_6[2:2], cf7__0[1:1]);
  C3 I402 (fa7_3min_0[0:0], cf7__0[2:2], termf_6[3:3], termf_4[3:3]);
  C3 I403 (fa7_3min_0[1:1], cf7__0[2:2], termf_6[3:3], termt_4[3:3]);
  C3 I404 (fa7_3min_0[2:2], cf7__0[2:2], termt_6[3:3], termf_4[3:3]);
  C3 I405 (fa7_3min_0[3:3], cf7__0[2:2], termt_6[3:3], termt_4[3:3]);
  C3 I406 (fa7_3min_0[4:4], ct7__0[2:2], termf_6[3:3], termf_4[3:3]);
  C3 I407 (fa7_3min_0[5:5], ct7__0[2:2], termf_6[3:3], termt_4[3:3]);
  C3 I408 (fa7_3min_0[6:6], ct7__0[2:2], termt_6[3:3], termf_4[3:3]);
  C3 I409 (fa7_3min_0[7:7], ct7__0[2:2], termt_6[3:3], termt_4[3:3]);
  NOR3 I410 (simp3911_0[0:0], fa7_3min_0[0:0], fa7_3min_0[3:3], fa7_3min_0[5:5]);
  INV I411 (simp3911_0[1:1], fa7_3min_0[6:6]);
  NAND2 I412 (o_0r0[3:3], simp3911_0[0:0], simp3911_0[1:1]);
  NOR3 I413 (simp3921_0[0:0], fa7_3min_0[1:1], fa7_3min_0[2:2], fa7_3min_0[4:4]);
  INV I414 (simp3921_0[1:1], fa7_3min_0[7:7]);
  NAND2 I415 (o_0r1[3:3], simp3921_0[0:0], simp3921_0[1:1]);
  AO222 I416 (ct7__0[3:3], termt_4[3:3], termt_6[3:3], termt_4[3:3], ct7__0[2:2], termt_6[3:3], ct7__0[2:2]);
  AO222 I417 (cf7__0[3:3], termf_4[3:3], termf_6[3:3], termf_4[3:3], cf7__0[2:2], termf_6[3:3], cf7__0[2:2]);
  C3 I418 (fa7_4min_0[0:0], cf7__0[3:3], termf_6[4:4], termf_4[4:4]);
  C3 I419 (fa7_4min_0[1:1], cf7__0[3:3], termf_6[4:4], termt_4[4:4]);
  C3 I420 (fa7_4min_0[2:2], cf7__0[3:3], termt_6[4:4], termf_4[4:4]);
  C3 I421 (fa7_4min_0[3:3], cf7__0[3:3], termt_6[4:4], termt_4[4:4]);
  C3 I422 (fa7_4min_0[4:4], ct7__0[3:3], termf_6[4:4], termf_4[4:4]);
  C3 I423 (fa7_4min_0[5:5], ct7__0[3:3], termf_6[4:4], termt_4[4:4]);
  C3 I424 (fa7_4min_0[6:6], ct7__0[3:3], termt_6[4:4], termf_4[4:4]);
  C3 I425 (fa7_4min_0[7:7], ct7__0[3:3], termt_6[4:4], termt_4[4:4]);
  NOR3 I426 (simp4041_0[0:0], fa7_4min_0[0:0], fa7_4min_0[3:3], fa7_4min_0[5:5]);
  INV I427 (simp4041_0[1:1], fa7_4min_0[6:6]);
  NAND2 I428 (o_0r0[4:4], simp4041_0[0:0], simp4041_0[1:1]);
  NOR3 I429 (simp4051_0[0:0], fa7_4min_0[1:1], fa7_4min_0[2:2], fa7_4min_0[4:4]);
  INV I430 (simp4051_0[1:1], fa7_4min_0[7:7]);
  NAND2 I431 (o_0r1[4:4], simp4051_0[0:0], simp4051_0[1:1]);
  AO222 I432 (ct7__0[4:4], termt_4[4:4], termt_6[4:4], termt_4[4:4], ct7__0[3:3], termt_6[4:4], ct7__0[3:3]);
  AO222 I433 (cf7__0[4:4], termf_4[4:4], termf_6[4:4], termf_4[4:4], cf7__0[3:3], termf_6[4:4], cf7__0[3:3]);
  C3 I434 (fa7_5min_0[0:0], cf7__0[4:4], termf_6[5:5], termf_4[5:5]);
  C3 I435 (fa7_5min_0[1:1], cf7__0[4:4], termf_6[5:5], termt_4[5:5]);
  C3 I436 (fa7_5min_0[2:2], cf7__0[4:4], termt_6[5:5], termf_4[5:5]);
  C3 I437 (fa7_5min_0[3:3], cf7__0[4:4], termt_6[5:5], termt_4[5:5]);
  C3 I438 (fa7_5min_0[4:4], ct7__0[4:4], termf_6[5:5], termf_4[5:5]);
  C3 I439 (fa7_5min_0[5:5], ct7__0[4:4], termf_6[5:5], termt_4[5:5]);
  C3 I440 (fa7_5min_0[6:6], ct7__0[4:4], termt_6[5:5], termf_4[5:5]);
  C3 I441 (fa7_5min_0[7:7], ct7__0[4:4], termt_6[5:5], termt_4[5:5]);
  NOR3 I442 (simp4171_0[0:0], fa7_5min_0[0:0], fa7_5min_0[3:3], fa7_5min_0[5:5]);
  INV I443 (simp4171_0[1:1], fa7_5min_0[6:6]);
  NAND2 I444 (o_0r0[5:5], simp4171_0[0:0], simp4171_0[1:1]);
  NOR3 I445 (simp4181_0[0:0], fa7_5min_0[1:1], fa7_5min_0[2:2], fa7_5min_0[4:4]);
  INV I446 (simp4181_0[1:1], fa7_5min_0[7:7]);
  NAND2 I447 (o_0r1[5:5], simp4181_0[0:0], simp4181_0[1:1]);
  AO222 I448 (ct7__0[5:5], termt_4[5:5], termt_6[5:5], termt_4[5:5], ct7__0[4:4], termt_6[5:5], ct7__0[4:4]);
  AO222 I449 (cf7__0[5:5], termf_4[5:5], termf_6[5:5], termf_4[5:5], cf7__0[4:4], termf_6[5:5], cf7__0[4:4]);
  C3 I450 (fa7_6min_0[0:0], cf7__0[5:5], termf_6[6:6], termf_4[6:6]);
  C3 I451 (fa7_6min_0[1:1], cf7__0[5:5], termf_6[6:6], termt_4[6:6]);
  C3 I452 (fa7_6min_0[2:2], cf7__0[5:5], termt_6[6:6], termf_4[6:6]);
  C3 I453 (fa7_6min_0[3:3], cf7__0[5:5], termt_6[6:6], termt_4[6:6]);
  C3 I454 (fa7_6min_0[4:4], ct7__0[5:5], termf_6[6:6], termf_4[6:6]);
  C3 I455 (fa7_6min_0[5:5], ct7__0[5:5], termf_6[6:6], termt_4[6:6]);
  C3 I456 (fa7_6min_0[6:6], ct7__0[5:5], termt_6[6:6], termf_4[6:6]);
  C3 I457 (fa7_6min_0[7:7], ct7__0[5:5], termt_6[6:6], termt_4[6:6]);
  NOR3 I458 (simp4301_0[0:0], fa7_6min_0[0:0], fa7_6min_0[3:3], fa7_6min_0[5:5]);
  INV I459 (simp4301_0[1:1], fa7_6min_0[6:6]);
  NAND2 I460 (o_0r0[6:6], simp4301_0[0:0], simp4301_0[1:1]);
  NOR3 I461 (simp4311_0[0:0], fa7_6min_0[1:1], fa7_6min_0[2:2], fa7_6min_0[4:4]);
  INV I462 (simp4311_0[1:1], fa7_6min_0[7:7]);
  NAND2 I463 (o_0r1[6:6], simp4311_0[0:0], simp4311_0[1:1]);
  AO222 I464 (ct7__0[6:6], termt_4[6:6], termt_6[6:6], termt_4[6:6], ct7__0[5:5], termt_6[6:6], ct7__0[5:5]);
  AO222 I465 (cf7__0[6:6], termf_4[6:6], termf_6[6:6], termf_4[6:6], cf7__0[5:5], termf_6[6:6], cf7__0[5:5]);
  C3 I466 (fa7_7min_0[0:0], cf7__0[6:6], termf_6[7:7], termf_4[7:7]);
  C3 I467 (fa7_7min_0[1:1], cf7__0[6:6], termf_6[7:7], termt_4[7:7]);
  C3 I468 (fa7_7min_0[2:2], cf7__0[6:6], termt_6[7:7], termf_4[7:7]);
  C3 I469 (fa7_7min_0[3:3], cf7__0[6:6], termt_6[7:7], termt_4[7:7]);
  C3 I470 (fa7_7min_0[4:4], ct7__0[6:6], termf_6[7:7], termf_4[7:7]);
  C3 I471 (fa7_7min_0[5:5], ct7__0[6:6], termf_6[7:7], termt_4[7:7]);
  C3 I472 (fa7_7min_0[6:6], ct7__0[6:6], termt_6[7:7], termf_4[7:7]);
  C3 I473 (fa7_7min_0[7:7], ct7__0[6:6], termt_6[7:7], termt_4[7:7]);
  NOR3 I474 (simp4431_0[0:0], fa7_7min_0[0:0], fa7_7min_0[3:3], fa7_7min_0[5:5]);
  INV I475 (simp4431_0[1:1], fa7_7min_0[6:6]);
  NAND2 I476 (o_0r0[7:7], simp4431_0[0:0], simp4431_0[1:1]);
  NOR3 I477 (simp4441_0[0:0], fa7_7min_0[1:1], fa7_7min_0[2:2], fa7_7min_0[4:4]);
  INV I478 (simp4441_0[1:1], fa7_7min_0[7:7]);
  NAND2 I479 (o_0r1[7:7], simp4441_0[0:0], simp4441_0[1:1]);
  AO222 I480 (ct7__0[7:7], termt_4[7:7], termt_6[7:7], termt_4[7:7], ct7__0[6:6], termt_6[7:7], ct7__0[6:6]);
  AO222 I481 (cf7__0[7:7], termf_4[7:7], termf_6[7:7], termf_4[7:7], cf7__0[6:6], termf_6[7:7], cf7__0[6:6]);
  C3 I482 (fa7_8min_0[0:0], cf7__0[7:7], termf_6[8:8], termf_4[8:8]);
  C3 I483 (fa7_8min_0[1:1], cf7__0[7:7], termf_6[8:8], termt_4[8:8]);
  C3 I484 (fa7_8min_0[2:2], cf7__0[7:7], termt_6[8:8], termf_4[8:8]);
  C3 I485 (fa7_8min_0[3:3], cf7__0[7:7], termt_6[8:8], termt_4[8:8]);
  C3 I486 (fa7_8min_0[4:4], ct7__0[7:7], termf_6[8:8], termf_4[8:8]);
  C3 I487 (fa7_8min_0[5:5], ct7__0[7:7], termf_6[8:8], termt_4[8:8]);
  C3 I488 (fa7_8min_0[6:6], ct7__0[7:7], termt_6[8:8], termf_4[8:8]);
  C3 I489 (fa7_8min_0[7:7], ct7__0[7:7], termt_6[8:8], termt_4[8:8]);
  NOR3 I490 (simp4561_0[0:0], fa7_8min_0[0:0], fa7_8min_0[3:3], fa7_8min_0[5:5]);
  INV I491 (simp4561_0[1:1], fa7_8min_0[6:6]);
  NAND2 I492 (o_0r0[8:8], simp4561_0[0:0], simp4561_0[1:1]);
  NOR3 I493 (simp4571_0[0:0], fa7_8min_0[1:1], fa7_8min_0[2:2], fa7_8min_0[4:4]);
  INV I494 (simp4571_0[1:1], fa7_8min_0[7:7]);
  NAND2 I495 (o_0r1[8:8], simp4571_0[0:0], simp4571_0[1:1]);
  AO222 I496 (ct7__0[8:8], termt_4[8:8], termt_6[8:8], termt_4[8:8], ct7__0[7:7], termt_6[8:8], ct7__0[7:7]);
  AO222 I497 (cf7__0[8:8], termf_4[8:8], termf_6[8:8], termf_4[8:8], cf7__0[7:7], termf_6[8:8], cf7__0[7:7]);
  C3 I498 (fa7_9min_0[0:0], cf7__0[8:8], termf_6[9:9], termf_4[9:9]);
  C3 I499 (fa7_9min_0[1:1], cf7__0[8:8], termf_6[9:9], termt_4[9:9]);
  C3 I500 (fa7_9min_0[2:2], cf7__0[8:8], termt_6[9:9], termf_4[9:9]);
  C3 I501 (fa7_9min_0[3:3], cf7__0[8:8], termt_6[9:9], termt_4[9:9]);
  C3 I502 (fa7_9min_0[4:4], ct7__0[8:8], termf_6[9:9], termf_4[9:9]);
  C3 I503 (fa7_9min_0[5:5], ct7__0[8:8], termf_6[9:9], termt_4[9:9]);
  C3 I504 (fa7_9min_0[6:6], ct7__0[8:8], termt_6[9:9], termf_4[9:9]);
  C3 I505 (fa7_9min_0[7:7], ct7__0[8:8], termt_6[9:9], termt_4[9:9]);
  NOR3 I506 (simp4691_0[0:0], fa7_9min_0[0:0], fa7_9min_0[3:3], fa7_9min_0[5:5]);
  INV I507 (simp4691_0[1:1], fa7_9min_0[6:6]);
  NAND2 I508 (o_0r0[9:9], simp4691_0[0:0], simp4691_0[1:1]);
  NOR3 I509 (simp4701_0[0:0], fa7_9min_0[1:1], fa7_9min_0[2:2], fa7_9min_0[4:4]);
  INV I510 (simp4701_0[1:1], fa7_9min_0[7:7]);
  NAND2 I511 (o_0r1[9:9], simp4701_0[0:0], simp4701_0[1:1]);
  AO222 I512 (ct7__0[9:9], termt_4[9:9], termt_6[9:9], termt_4[9:9], ct7__0[8:8], termt_6[9:9], ct7__0[8:8]);
  AO222 I513 (cf7__0[9:9], termf_4[9:9], termf_6[9:9], termf_4[9:9], cf7__0[8:8], termf_6[9:9], cf7__0[8:8]);
  C3 I514 (fa7_10min_0[0:0], cf7__0[9:9], termf_6[10:10], termf_4[10:10]);
  C3 I515 (fa7_10min_0[1:1], cf7__0[9:9], termf_6[10:10], termt_4[10:10]);
  C3 I516 (fa7_10min_0[2:2], cf7__0[9:9], termt_6[10:10], termf_4[10:10]);
  C3 I517 (fa7_10min_0[3:3], cf7__0[9:9], termt_6[10:10], termt_4[10:10]);
  C3 I518 (fa7_10min_0[4:4], ct7__0[9:9], termf_6[10:10], termf_4[10:10]);
  C3 I519 (fa7_10min_0[5:5], ct7__0[9:9], termf_6[10:10], termt_4[10:10]);
  C3 I520 (fa7_10min_0[6:6], ct7__0[9:9], termt_6[10:10], termf_4[10:10]);
  C3 I521 (fa7_10min_0[7:7], ct7__0[9:9], termt_6[10:10], termt_4[10:10]);
  NOR3 I522 (simp4821_0[0:0], fa7_10min_0[0:0], fa7_10min_0[3:3], fa7_10min_0[5:5]);
  INV I523 (simp4821_0[1:1], fa7_10min_0[6:6]);
  NAND2 I524 (o_0r0[10:10], simp4821_0[0:0], simp4821_0[1:1]);
  NOR3 I525 (simp4831_0[0:0], fa7_10min_0[1:1], fa7_10min_0[2:2], fa7_10min_0[4:4]);
  INV I526 (simp4831_0[1:1], fa7_10min_0[7:7]);
  NAND2 I527 (o_0r1[10:10], simp4831_0[0:0], simp4831_0[1:1]);
  AO222 I528 (ct7__0[10:10], termt_4[10:10], termt_6[10:10], termt_4[10:10], ct7__0[9:9], termt_6[10:10], ct7__0[9:9]);
  AO222 I529 (cf7__0[10:10], termf_4[10:10], termf_6[10:10], termf_4[10:10], cf7__0[9:9], termf_6[10:10], cf7__0[9:9]);
  C3 I530 (fa7_11min_0[0:0], cf7__0[10:10], termf_6[11:11], termf_4[11:11]);
  C3 I531 (fa7_11min_0[1:1], cf7__0[10:10], termf_6[11:11], termt_4[11:11]);
  C3 I532 (fa7_11min_0[2:2], cf7__0[10:10], termt_6[11:11], termf_4[11:11]);
  C3 I533 (fa7_11min_0[3:3], cf7__0[10:10], termt_6[11:11], termt_4[11:11]);
  C3 I534 (fa7_11min_0[4:4], ct7__0[10:10], termf_6[11:11], termf_4[11:11]);
  C3 I535 (fa7_11min_0[5:5], ct7__0[10:10], termf_6[11:11], termt_4[11:11]);
  C3 I536 (fa7_11min_0[6:6], ct7__0[10:10], termt_6[11:11], termf_4[11:11]);
  C3 I537 (fa7_11min_0[7:7], ct7__0[10:10], termt_6[11:11], termt_4[11:11]);
  NOR3 I538 (simp4951_0[0:0], fa7_11min_0[0:0], fa7_11min_0[3:3], fa7_11min_0[5:5]);
  INV I539 (simp4951_0[1:1], fa7_11min_0[6:6]);
  NAND2 I540 (o_0r0[11:11], simp4951_0[0:0], simp4951_0[1:1]);
  NOR3 I541 (simp4961_0[0:0], fa7_11min_0[1:1], fa7_11min_0[2:2], fa7_11min_0[4:4]);
  INV I542 (simp4961_0[1:1], fa7_11min_0[7:7]);
  NAND2 I543 (o_0r1[11:11], simp4961_0[0:0], simp4961_0[1:1]);
  AO222 I544 (ct7__0[11:11], termt_4[11:11], termt_6[11:11], termt_4[11:11], ct7__0[10:10], termt_6[11:11], ct7__0[10:10]);
  AO222 I545 (cf7__0[11:11], termf_4[11:11], termf_6[11:11], termf_4[11:11], cf7__0[10:10], termf_6[11:11], cf7__0[10:10]);
  C3 I546 (fa7_12min_0[0:0], cf7__0[11:11], termf_6[12:12], termf_4[12:12]);
  C3 I547 (fa7_12min_0[1:1], cf7__0[11:11], termf_6[12:12], termt_4[12:12]);
  C3 I548 (fa7_12min_0[2:2], cf7__0[11:11], termt_6[12:12], termf_4[12:12]);
  C3 I549 (fa7_12min_0[3:3], cf7__0[11:11], termt_6[12:12], termt_4[12:12]);
  C3 I550 (fa7_12min_0[4:4], ct7__0[11:11], termf_6[12:12], termf_4[12:12]);
  C3 I551 (fa7_12min_0[5:5], ct7__0[11:11], termf_6[12:12], termt_4[12:12]);
  C3 I552 (fa7_12min_0[6:6], ct7__0[11:11], termt_6[12:12], termf_4[12:12]);
  C3 I553 (fa7_12min_0[7:7], ct7__0[11:11], termt_6[12:12], termt_4[12:12]);
  NOR3 I554 (simp5081_0[0:0], fa7_12min_0[0:0], fa7_12min_0[3:3], fa7_12min_0[5:5]);
  INV I555 (simp5081_0[1:1], fa7_12min_0[6:6]);
  NAND2 I556 (o_0r0[12:12], simp5081_0[0:0], simp5081_0[1:1]);
  NOR3 I557 (simp5091_0[0:0], fa7_12min_0[1:1], fa7_12min_0[2:2], fa7_12min_0[4:4]);
  INV I558 (simp5091_0[1:1], fa7_12min_0[7:7]);
  NAND2 I559 (o_0r1[12:12], simp5091_0[0:0], simp5091_0[1:1]);
  AO222 I560 (ct7__0[12:12], termt_4[12:12], termt_6[12:12], termt_4[12:12], ct7__0[11:11], termt_6[12:12], ct7__0[11:11]);
  AO222 I561 (cf7__0[12:12], termf_4[12:12], termf_6[12:12], termf_4[12:12], cf7__0[11:11], termf_6[12:12], cf7__0[11:11]);
  C3 I562 (fa7_13min_0[0:0], cf7__0[12:12], termf_6[13:13], termf_4[13:13]);
  C3 I563 (fa7_13min_0[1:1], cf7__0[12:12], termf_6[13:13], termt_4[13:13]);
  C3 I564 (fa7_13min_0[2:2], cf7__0[12:12], termt_6[13:13], termf_4[13:13]);
  C3 I565 (fa7_13min_0[3:3], cf7__0[12:12], termt_6[13:13], termt_4[13:13]);
  C3 I566 (fa7_13min_0[4:4], ct7__0[12:12], termf_6[13:13], termf_4[13:13]);
  C3 I567 (fa7_13min_0[5:5], ct7__0[12:12], termf_6[13:13], termt_4[13:13]);
  C3 I568 (fa7_13min_0[6:6], ct7__0[12:12], termt_6[13:13], termf_4[13:13]);
  C3 I569 (fa7_13min_0[7:7], ct7__0[12:12], termt_6[13:13], termt_4[13:13]);
  NOR3 I570 (simp5211_0[0:0], fa7_13min_0[0:0], fa7_13min_0[3:3], fa7_13min_0[5:5]);
  INV I571 (simp5211_0[1:1], fa7_13min_0[6:6]);
  NAND2 I572 (o_0r0[13:13], simp5211_0[0:0], simp5211_0[1:1]);
  NOR3 I573 (simp5221_0[0:0], fa7_13min_0[1:1], fa7_13min_0[2:2], fa7_13min_0[4:4]);
  INV I574 (simp5221_0[1:1], fa7_13min_0[7:7]);
  NAND2 I575 (o_0r1[13:13], simp5221_0[0:0], simp5221_0[1:1]);
  AO222 I576 (ct7__0[13:13], termt_4[13:13], termt_6[13:13], termt_4[13:13], ct7__0[12:12], termt_6[13:13], ct7__0[12:12]);
  AO222 I577 (cf7__0[13:13], termf_4[13:13], termf_6[13:13], termf_4[13:13], cf7__0[12:12], termf_6[13:13], cf7__0[12:12]);
  C3 I578 (fa7_14min_0[0:0], cf7__0[13:13], termf_6[14:14], termf_4[14:14]);
  C3 I579 (fa7_14min_0[1:1], cf7__0[13:13], termf_6[14:14], termt_4[14:14]);
  C3 I580 (fa7_14min_0[2:2], cf7__0[13:13], termt_6[14:14], termf_4[14:14]);
  C3 I581 (fa7_14min_0[3:3], cf7__0[13:13], termt_6[14:14], termt_4[14:14]);
  C3 I582 (fa7_14min_0[4:4], ct7__0[13:13], termf_6[14:14], termf_4[14:14]);
  C3 I583 (fa7_14min_0[5:5], ct7__0[13:13], termf_6[14:14], termt_4[14:14]);
  C3 I584 (fa7_14min_0[6:6], ct7__0[13:13], termt_6[14:14], termf_4[14:14]);
  C3 I585 (fa7_14min_0[7:7], ct7__0[13:13], termt_6[14:14], termt_4[14:14]);
  NOR3 I586 (simp5341_0[0:0], fa7_14min_0[0:0], fa7_14min_0[3:3], fa7_14min_0[5:5]);
  INV I587 (simp5341_0[1:1], fa7_14min_0[6:6]);
  NAND2 I588 (o_0r0[14:14], simp5341_0[0:0], simp5341_0[1:1]);
  NOR3 I589 (simp5351_0[0:0], fa7_14min_0[1:1], fa7_14min_0[2:2], fa7_14min_0[4:4]);
  INV I590 (simp5351_0[1:1], fa7_14min_0[7:7]);
  NAND2 I591 (o_0r1[14:14], simp5351_0[0:0], simp5351_0[1:1]);
  AO222 I592 (ct7__0[14:14], termt_4[14:14], termt_6[14:14], termt_4[14:14], ct7__0[13:13], termt_6[14:14], ct7__0[13:13]);
  AO222 I593 (cf7__0[14:14], termf_4[14:14], termf_6[14:14], termf_4[14:14], cf7__0[13:13], termf_6[14:14], cf7__0[13:13]);
  C3 I594 (fa7_15min_0[0:0], cf7__0[14:14], termf_6[15:15], termf_4[15:15]);
  C3 I595 (fa7_15min_0[1:1], cf7__0[14:14], termf_6[15:15], termt_4[15:15]);
  C3 I596 (fa7_15min_0[2:2], cf7__0[14:14], termt_6[15:15], termf_4[15:15]);
  C3 I597 (fa7_15min_0[3:3], cf7__0[14:14], termt_6[15:15], termt_4[15:15]);
  C3 I598 (fa7_15min_0[4:4], ct7__0[14:14], termf_6[15:15], termf_4[15:15]);
  C3 I599 (fa7_15min_0[5:5], ct7__0[14:14], termf_6[15:15], termt_4[15:15]);
  C3 I600 (fa7_15min_0[6:6], ct7__0[14:14], termt_6[15:15], termf_4[15:15]);
  C3 I601 (fa7_15min_0[7:7], ct7__0[14:14], termt_6[15:15], termt_4[15:15]);
  NOR3 I602 (simp5471_0[0:0], fa7_15min_0[0:0], fa7_15min_0[3:3], fa7_15min_0[5:5]);
  INV I603 (simp5471_0[1:1], fa7_15min_0[6:6]);
  NAND2 I604 (o_0r0[15:15], simp5471_0[0:0], simp5471_0[1:1]);
  NOR3 I605 (simp5481_0[0:0], fa7_15min_0[1:1], fa7_15min_0[2:2], fa7_15min_0[4:4]);
  INV I606 (simp5481_0[1:1], fa7_15min_0[7:7]);
  NAND2 I607 (o_0r1[15:15], simp5481_0[0:0], simp5481_0[1:1]);
  AO222 I608 (ct7__0[15:15], termt_4[15:15], termt_6[15:15], termt_4[15:15], ct7__0[14:14], termt_6[15:15], ct7__0[14:14]);
  AO222 I609 (cf7__0[15:15], termf_4[15:15], termf_6[15:15], termf_4[15:15], cf7__0[14:14], termf_6[15:15], cf7__0[14:14]);
  C3 I610 (fa7_16min_0[0:0], cf7__0[15:15], termf_6[16:16], termf_4[16:16]);
  C3 I611 (fa7_16min_0[1:1], cf7__0[15:15], termf_6[16:16], termt_4[16:16]);
  C3 I612 (fa7_16min_0[2:2], cf7__0[15:15], termt_6[16:16], termf_4[16:16]);
  C3 I613 (fa7_16min_0[3:3], cf7__0[15:15], termt_6[16:16], termt_4[16:16]);
  C3 I614 (fa7_16min_0[4:4], ct7__0[15:15], termf_6[16:16], termf_4[16:16]);
  C3 I615 (fa7_16min_0[5:5], ct7__0[15:15], termf_6[16:16], termt_4[16:16]);
  C3 I616 (fa7_16min_0[6:6], ct7__0[15:15], termt_6[16:16], termf_4[16:16]);
  C3 I617 (fa7_16min_0[7:7], ct7__0[15:15], termt_6[16:16], termt_4[16:16]);
  NOR3 I618 (simp5601_0[0:0], fa7_16min_0[0:0], fa7_16min_0[3:3], fa7_16min_0[5:5]);
  INV I619 (simp5601_0[1:1], fa7_16min_0[6:6]);
  NAND2 I620 (o_0r0[16:16], simp5601_0[0:0], simp5601_0[1:1]);
  NOR3 I621 (simp5611_0[0:0], fa7_16min_0[1:1], fa7_16min_0[2:2], fa7_16min_0[4:4]);
  INV I622 (simp5611_0[1:1], fa7_16min_0[7:7]);
  NAND2 I623 (o_0r1[16:16], simp5611_0[0:0], simp5611_0[1:1]);
  AO222 I624 (ct7__0[16:16], termt_4[16:16], termt_6[16:16], termt_4[16:16], ct7__0[15:15], termt_6[16:16], ct7__0[15:15]);
  AO222 I625 (cf7__0[16:16], termf_4[16:16], termf_6[16:16], termf_4[16:16], cf7__0[15:15], termf_6[16:16], cf7__0[15:15]);
  C3 I626 (fa7_17min_0[0:0], cf7__0[16:16], termf_6[17:17], termf_4[17:17]);
  C3 I627 (fa7_17min_0[1:1], cf7__0[16:16], termf_6[17:17], termt_4[17:17]);
  C3 I628 (fa7_17min_0[2:2], cf7__0[16:16], termt_6[17:17], termf_4[17:17]);
  C3 I629 (fa7_17min_0[3:3], cf7__0[16:16], termt_6[17:17], termt_4[17:17]);
  C3 I630 (fa7_17min_0[4:4], ct7__0[16:16], termf_6[17:17], termf_4[17:17]);
  C3 I631 (fa7_17min_0[5:5], ct7__0[16:16], termf_6[17:17], termt_4[17:17]);
  C3 I632 (fa7_17min_0[6:6], ct7__0[16:16], termt_6[17:17], termf_4[17:17]);
  C3 I633 (fa7_17min_0[7:7], ct7__0[16:16], termt_6[17:17], termt_4[17:17]);
  NOR3 I634 (simp5731_0[0:0], fa7_17min_0[0:0], fa7_17min_0[3:3], fa7_17min_0[5:5]);
  INV I635 (simp5731_0[1:1], fa7_17min_0[6:6]);
  NAND2 I636 (o_0r0[17:17], simp5731_0[0:0], simp5731_0[1:1]);
  NOR3 I637 (simp5741_0[0:0], fa7_17min_0[1:1], fa7_17min_0[2:2], fa7_17min_0[4:4]);
  INV I638 (simp5741_0[1:1], fa7_17min_0[7:7]);
  NAND2 I639 (o_0r1[17:17], simp5741_0[0:0], simp5741_0[1:1]);
  AO222 I640 (ct7__0[17:17], termt_4[17:17], termt_6[17:17], termt_4[17:17], ct7__0[16:16], termt_6[17:17], ct7__0[16:16]);
  AO222 I641 (cf7__0[17:17], termf_4[17:17], termf_6[17:17], termf_4[17:17], cf7__0[16:16], termf_6[17:17], cf7__0[16:16]);
  C3 I642 (fa7_18min_0[0:0], cf7__0[17:17], termf_6[18:18], termf_4[18:18]);
  C3 I643 (fa7_18min_0[1:1], cf7__0[17:17], termf_6[18:18], termt_4[18:18]);
  C3 I644 (fa7_18min_0[2:2], cf7__0[17:17], termt_6[18:18], termf_4[18:18]);
  C3 I645 (fa7_18min_0[3:3], cf7__0[17:17], termt_6[18:18], termt_4[18:18]);
  C3 I646 (fa7_18min_0[4:4], ct7__0[17:17], termf_6[18:18], termf_4[18:18]);
  C3 I647 (fa7_18min_0[5:5], ct7__0[17:17], termf_6[18:18], termt_4[18:18]);
  C3 I648 (fa7_18min_0[6:6], ct7__0[17:17], termt_6[18:18], termf_4[18:18]);
  C3 I649 (fa7_18min_0[7:7], ct7__0[17:17], termt_6[18:18], termt_4[18:18]);
  NOR3 I650 (simp5861_0[0:0], fa7_18min_0[0:0], fa7_18min_0[3:3], fa7_18min_0[5:5]);
  INV I651 (simp5861_0[1:1], fa7_18min_0[6:6]);
  NAND2 I652 (o_0r0[18:18], simp5861_0[0:0], simp5861_0[1:1]);
  NOR3 I653 (simp5871_0[0:0], fa7_18min_0[1:1], fa7_18min_0[2:2], fa7_18min_0[4:4]);
  INV I654 (simp5871_0[1:1], fa7_18min_0[7:7]);
  NAND2 I655 (o_0r1[18:18], simp5871_0[0:0], simp5871_0[1:1]);
  AO222 I656 (ct7__0[18:18], termt_4[18:18], termt_6[18:18], termt_4[18:18], ct7__0[17:17], termt_6[18:18], ct7__0[17:17]);
  AO222 I657 (cf7__0[18:18], termf_4[18:18], termf_6[18:18], termf_4[18:18], cf7__0[17:17], termf_6[18:18], cf7__0[17:17]);
  C3 I658 (fa7_19min_0[0:0], cf7__0[18:18], termf_6[19:19], termf_4[19:19]);
  C3 I659 (fa7_19min_0[1:1], cf7__0[18:18], termf_6[19:19], termt_4[19:19]);
  C3 I660 (fa7_19min_0[2:2], cf7__0[18:18], termt_6[19:19], termf_4[19:19]);
  C3 I661 (fa7_19min_0[3:3], cf7__0[18:18], termt_6[19:19], termt_4[19:19]);
  C3 I662 (fa7_19min_0[4:4], ct7__0[18:18], termf_6[19:19], termf_4[19:19]);
  C3 I663 (fa7_19min_0[5:5], ct7__0[18:18], termf_6[19:19], termt_4[19:19]);
  C3 I664 (fa7_19min_0[6:6], ct7__0[18:18], termt_6[19:19], termf_4[19:19]);
  C3 I665 (fa7_19min_0[7:7], ct7__0[18:18], termt_6[19:19], termt_4[19:19]);
  NOR3 I666 (simp5991_0[0:0], fa7_19min_0[0:0], fa7_19min_0[3:3], fa7_19min_0[5:5]);
  INV I667 (simp5991_0[1:1], fa7_19min_0[6:6]);
  NAND2 I668 (o_0r0[19:19], simp5991_0[0:0], simp5991_0[1:1]);
  NOR3 I669 (simp6001_0[0:0], fa7_19min_0[1:1], fa7_19min_0[2:2], fa7_19min_0[4:4]);
  INV I670 (simp6001_0[1:1], fa7_19min_0[7:7]);
  NAND2 I671 (o_0r1[19:19], simp6001_0[0:0], simp6001_0[1:1]);
  AO222 I672 (ct7__0[19:19], termt_4[19:19], termt_6[19:19], termt_4[19:19], ct7__0[18:18], termt_6[19:19], ct7__0[18:18]);
  AO222 I673 (cf7__0[19:19], termf_4[19:19], termf_6[19:19], termf_4[19:19], cf7__0[18:18], termf_6[19:19], cf7__0[18:18]);
  C3 I674 (fa7_20min_0[0:0], cf7__0[19:19], termf_6[20:20], termf_4[20:20]);
  C3 I675 (fa7_20min_0[1:1], cf7__0[19:19], termf_6[20:20], termt_4[20:20]);
  C3 I676 (fa7_20min_0[2:2], cf7__0[19:19], termt_6[20:20], termf_4[20:20]);
  C3 I677 (fa7_20min_0[3:3], cf7__0[19:19], termt_6[20:20], termt_4[20:20]);
  C3 I678 (fa7_20min_0[4:4], ct7__0[19:19], termf_6[20:20], termf_4[20:20]);
  C3 I679 (fa7_20min_0[5:5], ct7__0[19:19], termf_6[20:20], termt_4[20:20]);
  C3 I680 (fa7_20min_0[6:6], ct7__0[19:19], termt_6[20:20], termf_4[20:20]);
  C3 I681 (fa7_20min_0[7:7], ct7__0[19:19], termt_6[20:20], termt_4[20:20]);
  NOR3 I682 (simp6121_0[0:0], fa7_20min_0[0:0], fa7_20min_0[3:3], fa7_20min_0[5:5]);
  INV I683 (simp6121_0[1:1], fa7_20min_0[6:6]);
  NAND2 I684 (o_0r0[20:20], simp6121_0[0:0], simp6121_0[1:1]);
  NOR3 I685 (simp6131_0[0:0], fa7_20min_0[1:1], fa7_20min_0[2:2], fa7_20min_0[4:4]);
  INV I686 (simp6131_0[1:1], fa7_20min_0[7:7]);
  NAND2 I687 (o_0r1[20:20], simp6131_0[0:0], simp6131_0[1:1]);
  AO222 I688 (ct7__0[20:20], termt_4[20:20], termt_6[20:20], termt_4[20:20], ct7__0[19:19], termt_6[20:20], ct7__0[19:19]);
  AO222 I689 (cf7__0[20:20], termf_4[20:20], termf_6[20:20], termf_4[20:20], cf7__0[19:19], termf_6[20:20], cf7__0[19:19]);
  C3 I690 (fa7_21min_0[0:0], cf7__0[20:20], termf_6[21:21], termf_4[21:21]);
  C3 I691 (fa7_21min_0[1:1], cf7__0[20:20], termf_6[21:21], termt_4[21:21]);
  C3 I692 (fa7_21min_0[2:2], cf7__0[20:20], termt_6[21:21], termf_4[21:21]);
  C3 I693 (fa7_21min_0[3:3], cf7__0[20:20], termt_6[21:21], termt_4[21:21]);
  C3 I694 (fa7_21min_0[4:4], ct7__0[20:20], termf_6[21:21], termf_4[21:21]);
  C3 I695 (fa7_21min_0[5:5], ct7__0[20:20], termf_6[21:21], termt_4[21:21]);
  C3 I696 (fa7_21min_0[6:6], ct7__0[20:20], termt_6[21:21], termf_4[21:21]);
  C3 I697 (fa7_21min_0[7:7], ct7__0[20:20], termt_6[21:21], termt_4[21:21]);
  NOR3 I698 (simp6251_0[0:0], fa7_21min_0[0:0], fa7_21min_0[3:3], fa7_21min_0[5:5]);
  INV I699 (simp6251_0[1:1], fa7_21min_0[6:6]);
  NAND2 I700 (o_0r0[21:21], simp6251_0[0:0], simp6251_0[1:1]);
  NOR3 I701 (simp6261_0[0:0], fa7_21min_0[1:1], fa7_21min_0[2:2], fa7_21min_0[4:4]);
  INV I702 (simp6261_0[1:1], fa7_21min_0[7:7]);
  NAND2 I703 (o_0r1[21:21], simp6261_0[0:0], simp6261_0[1:1]);
  AO222 I704 (ct7__0[21:21], termt_4[21:21], termt_6[21:21], termt_4[21:21], ct7__0[20:20], termt_6[21:21], ct7__0[20:20]);
  AO222 I705 (cf7__0[21:21], termf_4[21:21], termf_6[21:21], termf_4[21:21], cf7__0[20:20], termf_6[21:21], cf7__0[20:20]);
  C3 I706 (fa7_22min_0[0:0], cf7__0[21:21], termf_6[22:22], termf_4[22:22]);
  C3 I707 (fa7_22min_0[1:1], cf7__0[21:21], termf_6[22:22], termt_4[22:22]);
  C3 I708 (fa7_22min_0[2:2], cf7__0[21:21], termt_6[22:22], termf_4[22:22]);
  C3 I709 (fa7_22min_0[3:3], cf7__0[21:21], termt_6[22:22], termt_4[22:22]);
  C3 I710 (fa7_22min_0[4:4], ct7__0[21:21], termf_6[22:22], termf_4[22:22]);
  C3 I711 (fa7_22min_0[5:5], ct7__0[21:21], termf_6[22:22], termt_4[22:22]);
  C3 I712 (fa7_22min_0[6:6], ct7__0[21:21], termt_6[22:22], termf_4[22:22]);
  C3 I713 (fa7_22min_0[7:7], ct7__0[21:21], termt_6[22:22], termt_4[22:22]);
  NOR3 I714 (simp6381_0[0:0], fa7_22min_0[0:0], fa7_22min_0[3:3], fa7_22min_0[5:5]);
  INV I715 (simp6381_0[1:1], fa7_22min_0[6:6]);
  NAND2 I716 (o_0r0[22:22], simp6381_0[0:0], simp6381_0[1:1]);
  NOR3 I717 (simp6391_0[0:0], fa7_22min_0[1:1], fa7_22min_0[2:2], fa7_22min_0[4:4]);
  INV I718 (simp6391_0[1:1], fa7_22min_0[7:7]);
  NAND2 I719 (o_0r1[22:22], simp6391_0[0:0], simp6391_0[1:1]);
  AO222 I720 (ct7__0[22:22], termt_4[22:22], termt_6[22:22], termt_4[22:22], ct7__0[21:21], termt_6[22:22], ct7__0[21:21]);
  AO222 I721 (cf7__0[22:22], termf_4[22:22], termf_6[22:22], termf_4[22:22], cf7__0[21:21], termf_6[22:22], cf7__0[21:21]);
  C3 I722 (fa7_23min_0[0:0], cf7__0[22:22], termf_6[23:23], termf_4[23:23]);
  C3 I723 (fa7_23min_0[1:1], cf7__0[22:22], termf_6[23:23], termt_4[23:23]);
  C3 I724 (fa7_23min_0[2:2], cf7__0[22:22], termt_6[23:23], termf_4[23:23]);
  C3 I725 (fa7_23min_0[3:3], cf7__0[22:22], termt_6[23:23], termt_4[23:23]);
  C3 I726 (fa7_23min_0[4:4], ct7__0[22:22], termf_6[23:23], termf_4[23:23]);
  C3 I727 (fa7_23min_0[5:5], ct7__0[22:22], termf_6[23:23], termt_4[23:23]);
  C3 I728 (fa7_23min_0[6:6], ct7__0[22:22], termt_6[23:23], termf_4[23:23]);
  C3 I729 (fa7_23min_0[7:7], ct7__0[22:22], termt_6[23:23], termt_4[23:23]);
  NOR3 I730 (simp6511_0[0:0], fa7_23min_0[0:0], fa7_23min_0[3:3], fa7_23min_0[5:5]);
  INV I731 (simp6511_0[1:1], fa7_23min_0[6:6]);
  NAND2 I732 (o_0r0[23:23], simp6511_0[0:0], simp6511_0[1:1]);
  NOR3 I733 (simp6521_0[0:0], fa7_23min_0[1:1], fa7_23min_0[2:2], fa7_23min_0[4:4]);
  INV I734 (simp6521_0[1:1], fa7_23min_0[7:7]);
  NAND2 I735 (o_0r1[23:23], simp6521_0[0:0], simp6521_0[1:1]);
  AO222 I736 (ct7__0[23:23], termt_4[23:23], termt_6[23:23], termt_4[23:23], ct7__0[22:22], termt_6[23:23], ct7__0[22:22]);
  AO222 I737 (cf7__0[23:23], termf_4[23:23], termf_6[23:23], termf_4[23:23], cf7__0[22:22], termf_6[23:23], cf7__0[22:22]);
  C3 I738 (fa7_24min_0[0:0], cf7__0[23:23], termf_6[24:24], termf_4[24:24]);
  C3 I739 (fa7_24min_0[1:1], cf7__0[23:23], termf_6[24:24], termt_4[24:24]);
  C3 I740 (fa7_24min_0[2:2], cf7__0[23:23], termt_6[24:24], termf_4[24:24]);
  C3 I741 (fa7_24min_0[3:3], cf7__0[23:23], termt_6[24:24], termt_4[24:24]);
  C3 I742 (fa7_24min_0[4:4], ct7__0[23:23], termf_6[24:24], termf_4[24:24]);
  C3 I743 (fa7_24min_0[5:5], ct7__0[23:23], termf_6[24:24], termt_4[24:24]);
  C3 I744 (fa7_24min_0[6:6], ct7__0[23:23], termt_6[24:24], termf_4[24:24]);
  C3 I745 (fa7_24min_0[7:7], ct7__0[23:23], termt_6[24:24], termt_4[24:24]);
  NOR3 I746 (simp6641_0[0:0], fa7_24min_0[0:0], fa7_24min_0[3:3], fa7_24min_0[5:5]);
  INV I747 (simp6641_0[1:1], fa7_24min_0[6:6]);
  NAND2 I748 (o_0r0[24:24], simp6641_0[0:0], simp6641_0[1:1]);
  NOR3 I749 (simp6651_0[0:0], fa7_24min_0[1:1], fa7_24min_0[2:2], fa7_24min_0[4:4]);
  INV I750 (simp6651_0[1:1], fa7_24min_0[7:7]);
  NAND2 I751 (o_0r1[24:24], simp6651_0[0:0], simp6651_0[1:1]);
  AO222 I752 (ct7__0[24:24], termt_4[24:24], termt_6[24:24], termt_4[24:24], ct7__0[23:23], termt_6[24:24], ct7__0[23:23]);
  AO222 I753 (cf7__0[24:24], termf_4[24:24], termf_6[24:24], termf_4[24:24], cf7__0[23:23], termf_6[24:24], cf7__0[23:23]);
  C3 I754 (fa7_25min_0[0:0], cf7__0[24:24], termf_6[25:25], termf_4[25:25]);
  C3 I755 (fa7_25min_0[1:1], cf7__0[24:24], termf_6[25:25], termt_4[25:25]);
  C3 I756 (fa7_25min_0[2:2], cf7__0[24:24], termt_6[25:25], termf_4[25:25]);
  C3 I757 (fa7_25min_0[3:3], cf7__0[24:24], termt_6[25:25], termt_4[25:25]);
  C3 I758 (fa7_25min_0[4:4], ct7__0[24:24], termf_6[25:25], termf_4[25:25]);
  C3 I759 (fa7_25min_0[5:5], ct7__0[24:24], termf_6[25:25], termt_4[25:25]);
  C3 I760 (fa7_25min_0[6:6], ct7__0[24:24], termt_6[25:25], termf_4[25:25]);
  C3 I761 (fa7_25min_0[7:7], ct7__0[24:24], termt_6[25:25], termt_4[25:25]);
  NOR3 I762 (simp6771_0[0:0], fa7_25min_0[0:0], fa7_25min_0[3:3], fa7_25min_0[5:5]);
  INV I763 (simp6771_0[1:1], fa7_25min_0[6:6]);
  NAND2 I764 (o_0r0[25:25], simp6771_0[0:0], simp6771_0[1:1]);
  NOR3 I765 (simp6781_0[0:0], fa7_25min_0[1:1], fa7_25min_0[2:2], fa7_25min_0[4:4]);
  INV I766 (simp6781_0[1:1], fa7_25min_0[7:7]);
  NAND2 I767 (o_0r1[25:25], simp6781_0[0:0], simp6781_0[1:1]);
  AO222 I768 (ct7__0[25:25], termt_4[25:25], termt_6[25:25], termt_4[25:25], ct7__0[24:24], termt_6[25:25], ct7__0[24:24]);
  AO222 I769 (cf7__0[25:25], termf_4[25:25], termf_6[25:25], termf_4[25:25], cf7__0[24:24], termf_6[25:25], cf7__0[24:24]);
  C3 I770 (fa7_26min_0[0:0], cf7__0[25:25], termf_6[26:26], termf_4[26:26]);
  C3 I771 (fa7_26min_0[1:1], cf7__0[25:25], termf_6[26:26], termt_4[26:26]);
  C3 I772 (fa7_26min_0[2:2], cf7__0[25:25], termt_6[26:26], termf_4[26:26]);
  C3 I773 (fa7_26min_0[3:3], cf7__0[25:25], termt_6[26:26], termt_4[26:26]);
  C3 I774 (fa7_26min_0[4:4], ct7__0[25:25], termf_6[26:26], termf_4[26:26]);
  C3 I775 (fa7_26min_0[5:5], ct7__0[25:25], termf_6[26:26], termt_4[26:26]);
  C3 I776 (fa7_26min_0[6:6], ct7__0[25:25], termt_6[26:26], termf_4[26:26]);
  C3 I777 (fa7_26min_0[7:7], ct7__0[25:25], termt_6[26:26], termt_4[26:26]);
  NOR3 I778 (simp6901_0[0:0], fa7_26min_0[0:0], fa7_26min_0[3:3], fa7_26min_0[5:5]);
  INV I779 (simp6901_0[1:1], fa7_26min_0[6:6]);
  NAND2 I780 (o_0r0[26:26], simp6901_0[0:0], simp6901_0[1:1]);
  NOR3 I781 (simp6911_0[0:0], fa7_26min_0[1:1], fa7_26min_0[2:2], fa7_26min_0[4:4]);
  INV I782 (simp6911_0[1:1], fa7_26min_0[7:7]);
  NAND2 I783 (o_0r1[26:26], simp6911_0[0:0], simp6911_0[1:1]);
  AO222 I784 (ct7__0[26:26], termt_4[26:26], termt_6[26:26], termt_4[26:26], ct7__0[25:25], termt_6[26:26], ct7__0[25:25]);
  AO222 I785 (cf7__0[26:26], termf_4[26:26], termf_6[26:26], termf_4[26:26], cf7__0[25:25], termf_6[26:26], cf7__0[25:25]);
  C3 I786 (fa7_27min_0[0:0], cf7__0[26:26], termf_6[27:27], termf_4[27:27]);
  C3 I787 (fa7_27min_0[1:1], cf7__0[26:26], termf_6[27:27], termt_4[27:27]);
  C3 I788 (fa7_27min_0[2:2], cf7__0[26:26], termt_6[27:27], termf_4[27:27]);
  C3 I789 (fa7_27min_0[3:3], cf7__0[26:26], termt_6[27:27], termt_4[27:27]);
  C3 I790 (fa7_27min_0[4:4], ct7__0[26:26], termf_6[27:27], termf_4[27:27]);
  C3 I791 (fa7_27min_0[5:5], ct7__0[26:26], termf_6[27:27], termt_4[27:27]);
  C3 I792 (fa7_27min_0[6:6], ct7__0[26:26], termt_6[27:27], termf_4[27:27]);
  C3 I793 (fa7_27min_0[7:7], ct7__0[26:26], termt_6[27:27], termt_4[27:27]);
  NOR3 I794 (simp7031_0[0:0], fa7_27min_0[0:0], fa7_27min_0[3:3], fa7_27min_0[5:5]);
  INV I795 (simp7031_0[1:1], fa7_27min_0[6:6]);
  NAND2 I796 (o_0r0[27:27], simp7031_0[0:0], simp7031_0[1:1]);
  NOR3 I797 (simp7041_0[0:0], fa7_27min_0[1:1], fa7_27min_0[2:2], fa7_27min_0[4:4]);
  INV I798 (simp7041_0[1:1], fa7_27min_0[7:7]);
  NAND2 I799 (o_0r1[27:27], simp7041_0[0:0], simp7041_0[1:1]);
  AO222 I800 (ct7__0[27:27], termt_4[27:27], termt_6[27:27], termt_4[27:27], ct7__0[26:26], termt_6[27:27], ct7__0[26:26]);
  AO222 I801 (cf7__0[27:27], termf_4[27:27], termf_6[27:27], termf_4[27:27], cf7__0[26:26], termf_6[27:27], cf7__0[26:26]);
  C3 I802 (fa7_28min_0[0:0], cf7__0[27:27], termf_6[28:28], termf_4[28:28]);
  C3 I803 (fa7_28min_0[1:1], cf7__0[27:27], termf_6[28:28], termt_4[28:28]);
  C3 I804 (fa7_28min_0[2:2], cf7__0[27:27], termt_6[28:28], termf_4[28:28]);
  C3 I805 (fa7_28min_0[3:3], cf7__0[27:27], termt_6[28:28], termt_4[28:28]);
  C3 I806 (fa7_28min_0[4:4], ct7__0[27:27], termf_6[28:28], termf_4[28:28]);
  C3 I807 (fa7_28min_0[5:5], ct7__0[27:27], termf_6[28:28], termt_4[28:28]);
  C3 I808 (fa7_28min_0[6:6], ct7__0[27:27], termt_6[28:28], termf_4[28:28]);
  C3 I809 (fa7_28min_0[7:7], ct7__0[27:27], termt_6[28:28], termt_4[28:28]);
  NOR3 I810 (simp7161_0[0:0], fa7_28min_0[0:0], fa7_28min_0[3:3], fa7_28min_0[5:5]);
  INV I811 (simp7161_0[1:1], fa7_28min_0[6:6]);
  NAND2 I812 (o_0r0[28:28], simp7161_0[0:0], simp7161_0[1:1]);
  NOR3 I813 (simp7171_0[0:0], fa7_28min_0[1:1], fa7_28min_0[2:2], fa7_28min_0[4:4]);
  INV I814 (simp7171_0[1:1], fa7_28min_0[7:7]);
  NAND2 I815 (o_0r1[28:28], simp7171_0[0:0], simp7171_0[1:1]);
  AO222 I816 (ct7__0[28:28], termt_4[28:28], termt_6[28:28], termt_4[28:28], ct7__0[27:27], termt_6[28:28], ct7__0[27:27]);
  AO222 I817 (cf7__0[28:28], termf_4[28:28], termf_6[28:28], termf_4[28:28], cf7__0[27:27], termf_6[28:28], cf7__0[27:27]);
  C3 I818 (fa7_29min_0[0:0], cf7__0[28:28], termf_6[29:29], termf_4[29:29]);
  C3 I819 (fa7_29min_0[1:1], cf7__0[28:28], termf_6[29:29], termt_4[29:29]);
  C3 I820 (fa7_29min_0[2:2], cf7__0[28:28], termt_6[29:29], termf_4[29:29]);
  C3 I821 (fa7_29min_0[3:3], cf7__0[28:28], termt_6[29:29], termt_4[29:29]);
  C3 I822 (fa7_29min_0[4:4], ct7__0[28:28], termf_6[29:29], termf_4[29:29]);
  C3 I823 (fa7_29min_0[5:5], ct7__0[28:28], termf_6[29:29], termt_4[29:29]);
  C3 I824 (fa7_29min_0[6:6], ct7__0[28:28], termt_6[29:29], termf_4[29:29]);
  C3 I825 (fa7_29min_0[7:7], ct7__0[28:28], termt_6[29:29], termt_4[29:29]);
  NOR3 I826 (simp7291_0[0:0], fa7_29min_0[0:0], fa7_29min_0[3:3], fa7_29min_0[5:5]);
  INV I827 (simp7291_0[1:1], fa7_29min_0[6:6]);
  NAND2 I828 (o_0r0[29:29], simp7291_0[0:0], simp7291_0[1:1]);
  NOR3 I829 (simp7301_0[0:0], fa7_29min_0[1:1], fa7_29min_0[2:2], fa7_29min_0[4:4]);
  INV I830 (simp7301_0[1:1], fa7_29min_0[7:7]);
  NAND2 I831 (o_0r1[29:29], simp7301_0[0:0], simp7301_0[1:1]);
  AO222 I832 (ct7__0[29:29], termt_4[29:29], termt_6[29:29], termt_4[29:29], ct7__0[28:28], termt_6[29:29], ct7__0[28:28]);
  AO222 I833 (cf7__0[29:29], termf_4[29:29], termf_6[29:29], termf_4[29:29], cf7__0[28:28], termf_6[29:29], cf7__0[28:28]);
  C3 I834 (fa7_30min_0[0:0], cf7__0[29:29], termf_6[30:30], termf_4[30:30]);
  C3 I835 (fa7_30min_0[1:1], cf7__0[29:29], termf_6[30:30], termt_4[30:30]);
  C3 I836 (fa7_30min_0[2:2], cf7__0[29:29], termt_6[30:30], termf_4[30:30]);
  C3 I837 (fa7_30min_0[3:3], cf7__0[29:29], termt_6[30:30], termt_4[30:30]);
  C3 I838 (fa7_30min_0[4:4], ct7__0[29:29], termf_6[30:30], termf_4[30:30]);
  C3 I839 (fa7_30min_0[5:5], ct7__0[29:29], termf_6[30:30], termt_4[30:30]);
  C3 I840 (fa7_30min_0[6:6], ct7__0[29:29], termt_6[30:30], termf_4[30:30]);
  C3 I841 (fa7_30min_0[7:7], ct7__0[29:29], termt_6[30:30], termt_4[30:30]);
  NOR3 I842 (simp7421_0[0:0], fa7_30min_0[0:0], fa7_30min_0[3:3], fa7_30min_0[5:5]);
  INV I843 (simp7421_0[1:1], fa7_30min_0[6:6]);
  NAND2 I844 (o_0r0[30:30], simp7421_0[0:0], simp7421_0[1:1]);
  NOR3 I845 (simp7431_0[0:0], fa7_30min_0[1:1], fa7_30min_0[2:2], fa7_30min_0[4:4]);
  INV I846 (simp7431_0[1:1], fa7_30min_0[7:7]);
  NAND2 I847 (o_0r1[30:30], simp7431_0[0:0], simp7431_0[1:1]);
  AO222 I848 (ct7__0[30:30], termt_4[30:30], termt_6[30:30], termt_4[30:30], ct7__0[29:29], termt_6[30:30], ct7__0[29:29]);
  AO222 I849 (cf7__0[30:30], termf_4[30:30], termf_6[30:30], termf_4[30:30], cf7__0[29:29], termf_6[30:30], cf7__0[29:29]);
  C3 I850 (fa7_31min_0[0:0], cf7__0[30:30], termf_6[31:31], termf_4[31:31]);
  C3 I851 (fa7_31min_0[1:1], cf7__0[30:30], termf_6[31:31], termt_4[31:31]);
  C3 I852 (fa7_31min_0[2:2], cf7__0[30:30], termt_6[31:31], termf_4[31:31]);
  C3 I853 (fa7_31min_0[3:3], cf7__0[30:30], termt_6[31:31], termt_4[31:31]);
  C3 I854 (fa7_31min_0[4:4], ct7__0[30:30], termf_6[31:31], termf_4[31:31]);
  C3 I855 (fa7_31min_0[5:5], ct7__0[30:30], termf_6[31:31], termt_4[31:31]);
  C3 I856 (fa7_31min_0[6:6], ct7__0[30:30], termt_6[31:31], termf_4[31:31]);
  C3 I857 (fa7_31min_0[7:7], ct7__0[30:30], termt_6[31:31], termt_4[31:31]);
  NOR3 I858 (simp7551_0[0:0], fa7_31min_0[0:0], fa7_31min_0[3:3], fa7_31min_0[5:5]);
  INV I859 (simp7551_0[1:1], fa7_31min_0[6:6]);
  NAND2 I860 (o_0r0[31:31], simp7551_0[0:0], simp7551_0[1:1]);
  NOR3 I861 (simp7561_0[0:0], fa7_31min_0[1:1], fa7_31min_0[2:2], fa7_31min_0[4:4]);
  INV I862 (simp7561_0[1:1], fa7_31min_0[7:7]);
  NAND2 I863 (o_0r1[31:31], simp7561_0[0:0], simp7561_0[1:1]);
  AO222 I864 (ct7__0[31:31], termt_4[31:31], termt_6[31:31], termt_4[31:31], ct7__0[30:30], termt_6[31:31], ct7__0[30:30]);
  AO222 I865 (cf7__0[31:31], termf_4[31:31], termf_6[31:31], termf_4[31:31], cf7__0[30:30], termf_6[31:31], cf7__0[30:30]);
  C3 I866 (fa7_32min_0[0:0], cf7__0[31:31], termf_6[32:32], termf_4[32:32]);
  C3 I867 (fa7_32min_0[1:1], cf7__0[31:31], termf_6[32:32], termt_4[32:32]);
  C3 I868 (fa7_32min_0[2:2], cf7__0[31:31], termt_6[32:32], termf_4[32:32]);
  C3 I869 (fa7_32min_0[3:3], cf7__0[31:31], termt_6[32:32], termt_4[32:32]);
  C3 I870 (fa7_32min_0[4:4], ct7__0[31:31], termf_6[32:32], termf_4[32:32]);
  C3 I871 (fa7_32min_0[5:5], ct7__0[31:31], termf_6[32:32], termt_4[32:32]);
  C3 I872 (fa7_32min_0[6:6], ct7__0[31:31], termt_6[32:32], termf_4[32:32]);
  C3 I873 (fa7_32min_0[7:7], ct7__0[31:31], termt_6[32:32], termt_4[32:32]);
  NOR3 I874 (simp7681_0[0:0], fa7_32min_0[0:0], fa7_32min_0[3:3], fa7_32min_0[5:5]);
  INV I875 (simp7681_0[1:1], fa7_32min_0[6:6]);
  NAND2 I876 (o_0r0[32:32], simp7681_0[0:0], simp7681_0[1:1]);
  NOR3 I877 (simp7691_0[0:0], fa7_32min_0[1:1], fa7_32min_0[2:2], fa7_32min_0[4:4]);
  INV I878 (simp7691_0[1:1], fa7_32min_0[7:7]);
  NAND2 I879 (o_0r1[32:32], simp7691_0[0:0], simp7691_0[1:1]);
  AO222 I880 (ct7__0[32:32], termt_4[32:32], termt_6[32:32], termt_4[32:32], ct7__0[31:31], termt_6[32:32], ct7__0[31:31]);
  AO222 I881 (cf7__0[32:32], termf_4[32:32], termf_6[32:32], termf_4[32:32], cf7__0[31:31], termf_6[32:32], cf7__0[31:31]);
  BUFF I882 (i_0a, o_0a);
endmodule

// tkvtake1_wo0w1_ro0w1 TeakV "take" 1 [] [0] [0] [Many [1],Many [0],Many [0],Many [1]]
module tkvtake1_wo0w1_ro0w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input wg_0r0;
  input wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  input reset;
  wire wf_0;
  wire wt_0;
  wire df_0;
  wire dt_0;
  wire wc_0;
  wire wacks_0;
  wire wenr_0;
  wire wen_0;
  wire anyread_0;
  wire nreset_0;
  wire drlgf_0;
  wire drlgt_0;
  wire comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire conwgit_0;
  wire conwgif_0;
  wire conwig_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0, wenr_0, nreset_0);
  AND2 I2 (drlgf_0, wf_0, wen_0);
  AND2 I3 (drlgt_0, wt_0, wen_0);
  NOR2 I4 (df_0, dt_0, drlgt_0);
  NOR3 I5 (dt_0, df_0, drlgf_0, reset);
  AO22 I6 (wacks_0, drlgf_0, df_0, drlgt_0, dt_0);
  OR2 I7 (comp0_0, wg_0r0, wg_0r1);
  BUFF I8 (wc_0, comp0_0);
  AND2 I9 (conwgif_0, wg_0r0, conwig_0);
  AND2 I10 (conwgit_0, wg_0r1, conwig_0);
  BUFF I11 (conwigc_0, wc_0);
  AO22 I12 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I13 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I14 (wf_0, conwgif_0);
  BUFF I15 (wt_0, conwgit_0);
  BUFF I16 (wenr_0, wc_0);
  C2 I17 (wd_0r, conwig_0, wacks_0);
  AND2 I18 (rd_0r0, df_0, rg_0r);
  AND2 I19 (rd_0r1, dt_0, rg_0r);
  OR2 I20 (anyread_0, rg_0r, rg_0a);
  BUFF I21 (wg_0a, wd_0a);
  BUFF I22 (rg_0a, rd_0a);
endmodule

// tkm8x1b TeakM [Many [1,1,1,1,1,1,1,1],One 1]
module tkm8x1b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, i_4r0, i_4r1, i_4a, i_5r0, i_5r1, i_5a, i_6r0, i_6r1, i_6a, i_7r0, i_7r1, i_7a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input i_1r0;
  input i_1r1;
  output i_1a;
  input i_2r0;
  input i_2r1;
  output i_2a;
  input i_3r0;
  input i_3r1;
  output i_3a;
  input i_4r0;
  input i_4r1;
  output i_4a;
  input i_5r0;
  input i_5r1;
  output i_5a;
  input i_6r0;
  input i_6r1;
  output i_6a;
  input i_7r0;
  input i_7r1;
  output i_7a;
  output o_0r0;
  output o_0r1;
  input o_0a;
  input reset;
  wire gfint_0;
  wire gfint_1;
  wire gfint_2;
  wire gfint_3;
  wire gfint_4;
  wire gfint_5;
  wire gfint_6;
  wire gfint_7;
  wire gtint_0;
  wire gtint_1;
  wire gtint_2;
  wire gtint_3;
  wire gtint_4;
  wire gtint_5;
  wire gtint_6;
  wire gtint_7;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire choice_4;
  wire choice_5;
  wire choice_6;
  wire choice_7;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire icomp_3;
  wire icomp_4;
  wire icomp_5;
  wire icomp_6;
  wire icomp_7;
  wire nchosen_0;
  wire [2:0] simp341_0;
  wire [2:0] simp351_0;
  wire comp0_0;
  wire comp1_0;
  wire comp2_0;
  wire comp3_0;
  wire comp4_0;
  wire comp5_0;
  wire comp6_0;
  wire comp7_0;
  wire [2:0] simp841_0;
  NOR3 I0 (simp341_0[0:0], gfint_0, gfint_1, gfint_2);
  NOR3 I1 (simp341_0[1:1], gfint_3, gfint_4, gfint_5);
  NOR2 I2 (simp341_0[2:2], gfint_6, gfint_7);
  NAND3 I3 (o_0r0, simp341_0[0:0], simp341_0[1:1], simp341_0[2:2]);
  NOR3 I4 (simp351_0[0:0], gtint_0, gtint_1, gtint_2);
  NOR3 I5 (simp351_0[1:1], gtint_3, gtint_4, gtint_5);
  NOR2 I6 (simp351_0[2:2], gtint_6, gtint_7);
  NAND3 I7 (o_0r1, simp351_0[0:0], simp351_0[1:1], simp351_0[2:2]);
  AND2 I8 (gtint_0, choice_0, i_0r1);
  AND2 I9 (gtint_1, choice_1, i_1r1);
  AND2 I10 (gtint_2, choice_2, i_2r1);
  AND2 I11 (gtint_3, choice_3, i_3r1);
  AND2 I12 (gtint_4, choice_4, i_4r1);
  AND2 I13 (gtint_5, choice_5, i_5r1);
  AND2 I14 (gtint_6, choice_6, i_6r1);
  AND2 I15 (gtint_7, choice_7, i_7r1);
  AND2 I16 (gfint_0, choice_0, i_0r0);
  AND2 I17 (gfint_1, choice_1, i_1r0);
  AND2 I18 (gfint_2, choice_2, i_2r0);
  AND2 I19 (gfint_3, choice_3, i_3r0);
  AND2 I20 (gfint_4, choice_4, i_4r0);
  AND2 I21 (gfint_5, choice_5, i_5r0);
  AND2 I22 (gfint_6, choice_6, i_6r0);
  AND2 I23 (gfint_7, choice_7, i_7r0);
  OR2 I24 (comp0_0, i_0r0, i_0r1);
  BUFF I25 (icomp_0, comp0_0);
  OR2 I26 (comp1_0, i_1r0, i_1r1);
  BUFF I27 (icomp_1, comp1_0);
  OR2 I28 (comp2_0, i_2r0, i_2r1);
  BUFF I29 (icomp_2, comp2_0);
  OR2 I30 (comp3_0, i_3r0, i_3r1);
  BUFF I31 (icomp_3, comp3_0);
  OR2 I32 (comp4_0, i_4r0, i_4r1);
  BUFF I33 (icomp_4, comp4_0);
  OR2 I34 (comp5_0, i_5r0, i_5r1);
  BUFF I35 (icomp_5, comp5_0);
  OR2 I36 (comp6_0, i_6r0, i_6r1);
  BUFF I37 (icomp_6, comp6_0);
  OR2 I38 (comp7_0, i_7r0, i_7r1);
  BUFF I39 (icomp_7, comp7_0);
  C2R I40 (choice_0, icomp_0, nchosen_0, reset);
  C2R I41 (choice_1, icomp_1, nchosen_0, reset);
  C2R I42 (choice_2, icomp_2, nchosen_0, reset);
  C2R I43 (choice_3, icomp_3, nchosen_0, reset);
  C2R I44 (choice_4, icomp_4, nchosen_0, reset);
  C2R I45 (choice_5, icomp_5, nchosen_0, reset);
  C2R I46 (choice_6, icomp_6, nchosen_0, reset);
  C2R I47 (choice_7, icomp_7, nchosen_0, reset);
  NOR3 I48 (simp841_0[0:0], choice_0, choice_1, choice_2);
  NOR3 I49 (simp841_0[1:1], choice_3, choice_4, choice_5);
  NOR2 I50 (simp841_0[2:2], choice_6, choice_7);
  NAND3 I51 (anychoice_0, simp841_0[0:0], simp841_0[1:1], simp841_0[2:2]);
  NOR2 I52 (nchosen_0, anychoice_0, o_0a);
  C2R I53 (i_0a, choice_0, o_0a, reset);
  C2R I54 (i_1a, choice_1, o_0a, reset);
  C2R I55 (i_2a, choice_2, o_0a, reset);
  C2R I56 (i_3a, choice_3, o_0a, reset);
  C2R I57 (i_4a, choice_4, o_0a, reset);
  C2R I58 (i_5a, choice_5, o_0a, reset);
  C2R I59 (i_6a, choice_6, o_0a, reset);
  C2R I60 (i_7a, choice_7, o_0a, reset);
endmodule

// tko0m8_1nm8b1 TeakO [
//     (1,TeakOConstant 8 1)] [One 0,One 8]
module tko0m8_1nm8b1 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [7:0] o_0r0;
  output [7:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  GND I1 (o_0r0[0:0]);
  BUFF I2 (o_0r0[1:1], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  BUFF I6 (o_0r0[5:5], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  BUFF I8 (o_0r0[7:7], i_0r);
  GND I9 (o_0r1[1:1]);
  GND I10 (o_0r1[2:2]);
  GND I11 (o_0r1[3:3]);
  GND I12 (o_0r1[4:4]);
  GND I13 (o_0r1[5:5]);
  GND I14 (o_0r1[6:6]);
  GND I15 (o_0r1[7:7]);
  BUFF I16 (i_0a, o_0a);
endmodule

// tko0m8_1nm8b2 TeakO [
//     (1,TeakOConstant 8 2)] [One 0,One 8]
module tko0m8_1nm8b2 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [7:0] o_0r0;
  output [7:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[1:1], i_0r);
  GND I1 (o_0r0[1:1]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  BUFF I6 (o_0r0[5:5], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  BUFF I8 (o_0r0[7:7], i_0r);
  GND I9 (o_0r1[0:0]);
  GND I10 (o_0r1[2:2]);
  GND I11 (o_0r1[3:3]);
  GND I12 (o_0r1[4:4]);
  GND I13 (o_0r1[5:5]);
  GND I14 (o_0r1[6:6]);
  GND I15 (o_0r1[7:7]);
  BUFF I16 (i_0a, o_0a);
endmodule

// tko0m8_1nm8b4 TeakO [
//     (1,TeakOConstant 8 4)] [One 0,One 8]
module tko0m8_1nm8b4 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [7:0] o_0r0;
  output [7:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[2:2], i_0r);
  GND I1 (o_0r0[2:2]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  BUFF I6 (o_0r0[5:5], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  BUFF I8 (o_0r0[7:7], i_0r);
  GND I9 (o_0r1[0:0]);
  GND I10 (o_0r1[1:1]);
  GND I11 (o_0r1[3:3]);
  GND I12 (o_0r1[4:4]);
  GND I13 (o_0r1[5:5]);
  GND I14 (o_0r1[6:6]);
  GND I15 (o_0r1[7:7]);
  BUFF I16 (i_0a, o_0a);
endmodule

// tko0m8_1nm8b8 TeakO [
//     (1,TeakOConstant 8 8)] [One 0,One 8]
module tko0m8_1nm8b8 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [7:0] o_0r0;
  output [7:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[3:3], i_0r);
  GND I1 (o_0r0[3:3]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  BUFF I6 (o_0r0[5:5], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  BUFF I8 (o_0r0[7:7], i_0r);
  GND I9 (o_0r1[0:0]);
  GND I10 (o_0r1[1:1]);
  GND I11 (o_0r1[2:2]);
  GND I12 (o_0r1[4:4]);
  GND I13 (o_0r1[5:5]);
  GND I14 (o_0r1[6:6]);
  GND I15 (o_0r1[7:7]);
  BUFF I16 (i_0a, o_0a);
endmodule

// tko0m8_1nm8b10 TeakO [
//     (1,TeakOConstant 8 16)] [One 0,One 8]
module tko0m8_1nm8b10 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [7:0] o_0r0;
  output [7:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[4:4], i_0r);
  GND I1 (o_0r0[4:4]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  BUFF I6 (o_0r0[5:5], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  BUFF I8 (o_0r0[7:7], i_0r);
  GND I9 (o_0r1[0:0]);
  GND I10 (o_0r1[1:1]);
  GND I11 (o_0r1[2:2]);
  GND I12 (o_0r1[3:3]);
  GND I13 (o_0r1[5:5]);
  GND I14 (o_0r1[6:6]);
  GND I15 (o_0r1[7:7]);
  BUFF I16 (i_0a, o_0a);
endmodule

// tko0m8_1nm8b20 TeakO [
//     (1,TeakOConstant 8 32)] [One 0,One 8]
module tko0m8_1nm8b20 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [7:0] o_0r0;
  output [7:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[5:5], i_0r);
  GND I1 (o_0r0[5:5]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  BUFF I6 (o_0r0[4:4], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  BUFF I8 (o_0r0[7:7], i_0r);
  GND I9 (o_0r1[0:0]);
  GND I10 (o_0r1[1:1]);
  GND I11 (o_0r1[2:2]);
  GND I12 (o_0r1[3:3]);
  GND I13 (o_0r1[4:4]);
  GND I14 (o_0r1[6:6]);
  GND I15 (o_0r1[7:7]);
  BUFF I16 (i_0a, o_0a);
endmodule

// tko0m8_1nm8b40 TeakO [
//     (1,TeakOConstant 8 64)] [One 0,One 8]
module tko0m8_1nm8b40 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [7:0] o_0r0;
  output [7:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[6:6], i_0r);
  GND I1 (o_0r0[6:6]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  BUFF I6 (o_0r0[4:4], i_0r);
  BUFF I7 (o_0r0[5:5], i_0r);
  BUFF I8 (o_0r0[7:7], i_0r);
  GND I9 (o_0r1[0:0]);
  GND I10 (o_0r1[1:1]);
  GND I11 (o_0r1[2:2]);
  GND I12 (o_0r1[3:3]);
  GND I13 (o_0r1[4:4]);
  GND I14 (o_0r1[5:5]);
  GND I15 (o_0r1[7:7]);
  BUFF I16 (i_0a, o_0a);
endmodule

// tko0m8_1nm8b80 TeakO [
//     (1,TeakOConstant 8 128)] [One 0,One 8]
module tko0m8_1nm8b80 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [7:0] o_0r0;
  output [7:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[7:7], i_0r);
  GND I1 (o_0r0[7:7]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  BUFF I6 (o_0r0[4:4], i_0r);
  BUFF I7 (o_0r0[5:5], i_0r);
  BUFF I8 (o_0r0[6:6], i_0r);
  GND I9 (o_0r1[0:0]);
  GND I10 (o_0r1[1:1]);
  GND I11 (o_0r1[2:2]);
  GND I12 (o_0r1[3:3]);
  GND I13 (o_0r1[4:4]);
  GND I14 (o_0r1[5:5]);
  GND I15 (o_0r1[6:6]);
  BUFF I16 (i_0a, o_0a);
endmodule

// tkm8x8b TeakM [Many [8,8,8,8,8,8,8,8],One 8]
module tkm8x8b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, i_4r0, i_4r1, i_4a, i_5r0, i_5r1, i_5a, i_6r0, i_6r1, i_6a, i_7r0, i_7r1, i_7a, o_0r0, o_0r1, o_0a, reset);
  input [7:0] i_0r0;
  input [7:0] i_0r1;
  output i_0a;
  input [7:0] i_1r0;
  input [7:0] i_1r1;
  output i_1a;
  input [7:0] i_2r0;
  input [7:0] i_2r1;
  output i_2a;
  input [7:0] i_3r0;
  input [7:0] i_3r1;
  output i_3a;
  input [7:0] i_4r0;
  input [7:0] i_4r1;
  output i_4a;
  input [7:0] i_5r0;
  input [7:0] i_5r1;
  output i_5a;
  input [7:0] i_6r0;
  input [7:0] i_6r1;
  output i_6a;
  input [7:0] i_7r0;
  input [7:0] i_7r1;
  output i_7a;
  output [7:0] o_0r0;
  output [7:0] o_0r1;
  input o_0a;
  input reset;
  wire [7:0] gfint_0;
  wire [7:0] gfint_1;
  wire [7:0] gfint_2;
  wire [7:0] gfint_3;
  wire [7:0] gfint_4;
  wire [7:0] gfint_5;
  wire [7:0] gfint_6;
  wire [7:0] gfint_7;
  wire [7:0] gtint_0;
  wire [7:0] gtint_1;
  wire [7:0] gtint_2;
  wire [7:0] gtint_3;
  wire [7:0] gtint_4;
  wire [7:0] gtint_5;
  wire [7:0] gtint_6;
  wire [7:0] gtint_7;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire choice_4;
  wire choice_5;
  wire choice_6;
  wire choice_7;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire icomp_3;
  wire icomp_4;
  wire icomp_5;
  wire icomp_6;
  wire icomp_7;
  wire nchosen_0;
  wire [2:0] simp341_0;
  wire [2:0] simp351_0;
  wire [2:0] simp361_0;
  wire [2:0] simp371_0;
  wire [2:0] simp381_0;
  wire [2:0] simp391_0;
  wire [2:0] simp401_0;
  wire [2:0] simp411_0;
  wire [2:0] simp421_0;
  wire [2:0] simp431_0;
  wire [2:0] simp441_0;
  wire [2:0] simp451_0;
  wire [2:0] simp461_0;
  wire [2:0] simp471_0;
  wire [2:0] simp481_0;
  wire [2:0] simp491_0;
  wire [7:0] comp0_0;
  wire [2:0] simp1871_0;
  wire [7:0] comp1_0;
  wire [2:0] simp1971_0;
  wire [7:0] comp2_0;
  wire [2:0] simp2071_0;
  wire [7:0] comp3_0;
  wire [2:0] simp2171_0;
  wire [7:0] comp4_0;
  wire [2:0] simp2271_0;
  wire [7:0] comp5_0;
  wire [2:0] simp2371_0;
  wire [7:0] comp6_0;
  wire [2:0] simp2471_0;
  wire [7:0] comp7_0;
  wire [2:0] simp2571_0;
  wire [2:0] simp2661_0;
  NOR3 I0 (simp341_0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  NOR3 I1 (simp341_0[1:1], gfint_3[0:0], gfint_4[0:0], gfint_5[0:0]);
  NOR2 I2 (simp341_0[2:2], gfint_6[0:0], gfint_7[0:0]);
  NAND3 I3 (o_0r0[0:0], simp341_0[0:0], simp341_0[1:1], simp341_0[2:2]);
  NOR3 I4 (simp351_0[0:0], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  NOR3 I5 (simp351_0[1:1], gfint_3[1:1], gfint_4[1:1], gfint_5[1:1]);
  NOR2 I6 (simp351_0[2:2], gfint_6[1:1], gfint_7[1:1]);
  NAND3 I7 (o_0r0[1:1], simp351_0[0:0], simp351_0[1:1], simp351_0[2:2]);
  NOR3 I8 (simp361_0[0:0], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  NOR3 I9 (simp361_0[1:1], gfint_3[2:2], gfint_4[2:2], gfint_5[2:2]);
  NOR2 I10 (simp361_0[2:2], gfint_6[2:2], gfint_7[2:2]);
  NAND3 I11 (o_0r0[2:2], simp361_0[0:0], simp361_0[1:1], simp361_0[2:2]);
  NOR3 I12 (simp371_0[0:0], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  NOR3 I13 (simp371_0[1:1], gfint_3[3:3], gfint_4[3:3], gfint_5[3:3]);
  NOR2 I14 (simp371_0[2:2], gfint_6[3:3], gfint_7[3:3]);
  NAND3 I15 (o_0r0[3:3], simp371_0[0:0], simp371_0[1:1], simp371_0[2:2]);
  NOR3 I16 (simp381_0[0:0], gfint_0[4:4], gfint_1[4:4], gfint_2[4:4]);
  NOR3 I17 (simp381_0[1:1], gfint_3[4:4], gfint_4[4:4], gfint_5[4:4]);
  NOR2 I18 (simp381_0[2:2], gfint_6[4:4], gfint_7[4:4]);
  NAND3 I19 (o_0r0[4:4], simp381_0[0:0], simp381_0[1:1], simp381_0[2:2]);
  NOR3 I20 (simp391_0[0:0], gfint_0[5:5], gfint_1[5:5], gfint_2[5:5]);
  NOR3 I21 (simp391_0[1:1], gfint_3[5:5], gfint_4[5:5], gfint_5[5:5]);
  NOR2 I22 (simp391_0[2:2], gfint_6[5:5], gfint_7[5:5]);
  NAND3 I23 (o_0r0[5:5], simp391_0[0:0], simp391_0[1:1], simp391_0[2:2]);
  NOR3 I24 (simp401_0[0:0], gfint_0[6:6], gfint_1[6:6], gfint_2[6:6]);
  NOR3 I25 (simp401_0[1:1], gfint_3[6:6], gfint_4[6:6], gfint_5[6:6]);
  NOR2 I26 (simp401_0[2:2], gfint_6[6:6], gfint_7[6:6]);
  NAND3 I27 (o_0r0[6:6], simp401_0[0:0], simp401_0[1:1], simp401_0[2:2]);
  NOR3 I28 (simp411_0[0:0], gfint_0[7:7], gfint_1[7:7], gfint_2[7:7]);
  NOR3 I29 (simp411_0[1:1], gfint_3[7:7], gfint_4[7:7], gfint_5[7:7]);
  NOR2 I30 (simp411_0[2:2], gfint_6[7:7], gfint_7[7:7]);
  NAND3 I31 (o_0r0[7:7], simp411_0[0:0], simp411_0[1:1], simp411_0[2:2]);
  NOR3 I32 (simp421_0[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  NOR3 I33 (simp421_0[1:1], gtint_3[0:0], gtint_4[0:0], gtint_5[0:0]);
  NOR2 I34 (simp421_0[2:2], gtint_6[0:0], gtint_7[0:0]);
  NAND3 I35 (o_0r1[0:0], simp421_0[0:0], simp421_0[1:1], simp421_0[2:2]);
  NOR3 I36 (simp431_0[0:0], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  NOR3 I37 (simp431_0[1:1], gtint_3[1:1], gtint_4[1:1], gtint_5[1:1]);
  NOR2 I38 (simp431_0[2:2], gtint_6[1:1], gtint_7[1:1]);
  NAND3 I39 (o_0r1[1:1], simp431_0[0:0], simp431_0[1:1], simp431_0[2:2]);
  NOR3 I40 (simp441_0[0:0], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  NOR3 I41 (simp441_0[1:1], gtint_3[2:2], gtint_4[2:2], gtint_5[2:2]);
  NOR2 I42 (simp441_0[2:2], gtint_6[2:2], gtint_7[2:2]);
  NAND3 I43 (o_0r1[2:2], simp441_0[0:0], simp441_0[1:1], simp441_0[2:2]);
  NOR3 I44 (simp451_0[0:0], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  NOR3 I45 (simp451_0[1:1], gtint_3[3:3], gtint_4[3:3], gtint_5[3:3]);
  NOR2 I46 (simp451_0[2:2], gtint_6[3:3], gtint_7[3:3]);
  NAND3 I47 (o_0r1[3:3], simp451_0[0:0], simp451_0[1:1], simp451_0[2:2]);
  NOR3 I48 (simp461_0[0:0], gtint_0[4:4], gtint_1[4:4], gtint_2[4:4]);
  NOR3 I49 (simp461_0[1:1], gtint_3[4:4], gtint_4[4:4], gtint_5[4:4]);
  NOR2 I50 (simp461_0[2:2], gtint_6[4:4], gtint_7[4:4]);
  NAND3 I51 (o_0r1[4:4], simp461_0[0:0], simp461_0[1:1], simp461_0[2:2]);
  NOR3 I52 (simp471_0[0:0], gtint_0[5:5], gtint_1[5:5], gtint_2[5:5]);
  NOR3 I53 (simp471_0[1:1], gtint_3[5:5], gtint_4[5:5], gtint_5[5:5]);
  NOR2 I54 (simp471_0[2:2], gtint_6[5:5], gtint_7[5:5]);
  NAND3 I55 (o_0r1[5:5], simp471_0[0:0], simp471_0[1:1], simp471_0[2:2]);
  NOR3 I56 (simp481_0[0:0], gtint_0[6:6], gtint_1[6:6], gtint_2[6:6]);
  NOR3 I57 (simp481_0[1:1], gtint_3[6:6], gtint_4[6:6], gtint_5[6:6]);
  NOR2 I58 (simp481_0[2:2], gtint_6[6:6], gtint_7[6:6]);
  NAND3 I59 (o_0r1[6:6], simp481_0[0:0], simp481_0[1:1], simp481_0[2:2]);
  NOR3 I60 (simp491_0[0:0], gtint_0[7:7], gtint_1[7:7], gtint_2[7:7]);
  NOR3 I61 (simp491_0[1:1], gtint_3[7:7], gtint_4[7:7], gtint_5[7:7]);
  NOR2 I62 (simp491_0[2:2], gtint_6[7:7], gtint_7[7:7]);
  NAND3 I63 (o_0r1[7:7], simp491_0[0:0], simp491_0[1:1], simp491_0[2:2]);
  AND2 I64 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I65 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I66 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I67 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I68 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I69 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I70 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I71 (gtint_0[7:7], choice_0, i_0r1[7:7]);
  AND2 I72 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I73 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I74 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I75 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I76 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I77 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I78 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I79 (gtint_1[7:7], choice_1, i_1r1[7:7]);
  AND2 I80 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I81 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I82 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I83 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AND2 I84 (gtint_2[4:4], choice_2, i_2r1[4:4]);
  AND2 I85 (gtint_2[5:5], choice_2, i_2r1[5:5]);
  AND2 I86 (gtint_2[6:6], choice_2, i_2r1[6:6]);
  AND2 I87 (gtint_2[7:7], choice_2, i_2r1[7:7]);
  AND2 I88 (gtint_3[0:0], choice_3, i_3r1[0:0]);
  AND2 I89 (gtint_3[1:1], choice_3, i_3r1[1:1]);
  AND2 I90 (gtint_3[2:2], choice_3, i_3r1[2:2]);
  AND2 I91 (gtint_3[3:3], choice_3, i_3r1[3:3]);
  AND2 I92 (gtint_3[4:4], choice_3, i_3r1[4:4]);
  AND2 I93 (gtint_3[5:5], choice_3, i_3r1[5:5]);
  AND2 I94 (gtint_3[6:6], choice_3, i_3r1[6:6]);
  AND2 I95 (gtint_3[7:7], choice_3, i_3r1[7:7]);
  AND2 I96 (gtint_4[0:0], choice_4, i_4r1[0:0]);
  AND2 I97 (gtint_4[1:1], choice_4, i_4r1[1:1]);
  AND2 I98 (gtint_4[2:2], choice_4, i_4r1[2:2]);
  AND2 I99 (gtint_4[3:3], choice_4, i_4r1[3:3]);
  AND2 I100 (gtint_4[4:4], choice_4, i_4r1[4:4]);
  AND2 I101 (gtint_4[5:5], choice_4, i_4r1[5:5]);
  AND2 I102 (gtint_4[6:6], choice_4, i_4r1[6:6]);
  AND2 I103 (gtint_4[7:7], choice_4, i_4r1[7:7]);
  AND2 I104 (gtint_5[0:0], choice_5, i_5r1[0:0]);
  AND2 I105 (gtint_5[1:1], choice_5, i_5r1[1:1]);
  AND2 I106 (gtint_5[2:2], choice_5, i_5r1[2:2]);
  AND2 I107 (gtint_5[3:3], choice_5, i_5r1[3:3]);
  AND2 I108 (gtint_5[4:4], choice_5, i_5r1[4:4]);
  AND2 I109 (gtint_5[5:5], choice_5, i_5r1[5:5]);
  AND2 I110 (gtint_5[6:6], choice_5, i_5r1[6:6]);
  AND2 I111 (gtint_5[7:7], choice_5, i_5r1[7:7]);
  AND2 I112 (gtint_6[0:0], choice_6, i_6r1[0:0]);
  AND2 I113 (gtint_6[1:1], choice_6, i_6r1[1:1]);
  AND2 I114 (gtint_6[2:2], choice_6, i_6r1[2:2]);
  AND2 I115 (gtint_6[3:3], choice_6, i_6r1[3:3]);
  AND2 I116 (gtint_6[4:4], choice_6, i_6r1[4:4]);
  AND2 I117 (gtint_6[5:5], choice_6, i_6r1[5:5]);
  AND2 I118 (gtint_6[6:6], choice_6, i_6r1[6:6]);
  AND2 I119 (gtint_6[7:7], choice_6, i_6r1[7:7]);
  AND2 I120 (gtint_7[0:0], choice_7, i_7r1[0:0]);
  AND2 I121 (gtint_7[1:1], choice_7, i_7r1[1:1]);
  AND2 I122 (gtint_7[2:2], choice_7, i_7r1[2:2]);
  AND2 I123 (gtint_7[3:3], choice_7, i_7r1[3:3]);
  AND2 I124 (gtint_7[4:4], choice_7, i_7r1[4:4]);
  AND2 I125 (gtint_7[5:5], choice_7, i_7r1[5:5]);
  AND2 I126 (gtint_7[6:6], choice_7, i_7r1[6:6]);
  AND2 I127 (gtint_7[7:7], choice_7, i_7r1[7:7]);
  AND2 I128 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I129 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I130 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I131 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I132 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I133 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I134 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I135 (gfint_0[7:7], choice_0, i_0r0[7:7]);
  AND2 I136 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I137 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I138 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I139 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I140 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I141 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I142 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I143 (gfint_1[7:7], choice_1, i_1r0[7:7]);
  AND2 I144 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I145 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I146 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I147 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AND2 I148 (gfint_2[4:4], choice_2, i_2r0[4:4]);
  AND2 I149 (gfint_2[5:5], choice_2, i_2r0[5:5]);
  AND2 I150 (gfint_2[6:6], choice_2, i_2r0[6:6]);
  AND2 I151 (gfint_2[7:7], choice_2, i_2r0[7:7]);
  AND2 I152 (gfint_3[0:0], choice_3, i_3r0[0:0]);
  AND2 I153 (gfint_3[1:1], choice_3, i_3r0[1:1]);
  AND2 I154 (gfint_3[2:2], choice_3, i_3r0[2:2]);
  AND2 I155 (gfint_3[3:3], choice_3, i_3r0[3:3]);
  AND2 I156 (gfint_3[4:4], choice_3, i_3r0[4:4]);
  AND2 I157 (gfint_3[5:5], choice_3, i_3r0[5:5]);
  AND2 I158 (gfint_3[6:6], choice_3, i_3r0[6:6]);
  AND2 I159 (gfint_3[7:7], choice_3, i_3r0[7:7]);
  AND2 I160 (gfint_4[0:0], choice_4, i_4r0[0:0]);
  AND2 I161 (gfint_4[1:1], choice_4, i_4r0[1:1]);
  AND2 I162 (gfint_4[2:2], choice_4, i_4r0[2:2]);
  AND2 I163 (gfint_4[3:3], choice_4, i_4r0[3:3]);
  AND2 I164 (gfint_4[4:4], choice_4, i_4r0[4:4]);
  AND2 I165 (gfint_4[5:5], choice_4, i_4r0[5:5]);
  AND2 I166 (gfint_4[6:6], choice_4, i_4r0[6:6]);
  AND2 I167 (gfint_4[7:7], choice_4, i_4r0[7:7]);
  AND2 I168 (gfint_5[0:0], choice_5, i_5r0[0:0]);
  AND2 I169 (gfint_5[1:1], choice_5, i_5r0[1:1]);
  AND2 I170 (gfint_5[2:2], choice_5, i_5r0[2:2]);
  AND2 I171 (gfint_5[3:3], choice_5, i_5r0[3:3]);
  AND2 I172 (gfint_5[4:4], choice_5, i_5r0[4:4]);
  AND2 I173 (gfint_5[5:5], choice_5, i_5r0[5:5]);
  AND2 I174 (gfint_5[6:6], choice_5, i_5r0[6:6]);
  AND2 I175 (gfint_5[7:7], choice_5, i_5r0[7:7]);
  AND2 I176 (gfint_6[0:0], choice_6, i_6r0[0:0]);
  AND2 I177 (gfint_6[1:1], choice_6, i_6r0[1:1]);
  AND2 I178 (gfint_6[2:2], choice_6, i_6r0[2:2]);
  AND2 I179 (gfint_6[3:3], choice_6, i_6r0[3:3]);
  AND2 I180 (gfint_6[4:4], choice_6, i_6r0[4:4]);
  AND2 I181 (gfint_6[5:5], choice_6, i_6r0[5:5]);
  AND2 I182 (gfint_6[6:6], choice_6, i_6r0[6:6]);
  AND2 I183 (gfint_6[7:7], choice_6, i_6r0[7:7]);
  AND2 I184 (gfint_7[0:0], choice_7, i_7r0[0:0]);
  AND2 I185 (gfint_7[1:1], choice_7, i_7r0[1:1]);
  AND2 I186 (gfint_7[2:2], choice_7, i_7r0[2:2]);
  AND2 I187 (gfint_7[3:3], choice_7, i_7r0[3:3]);
  AND2 I188 (gfint_7[4:4], choice_7, i_7r0[4:4]);
  AND2 I189 (gfint_7[5:5], choice_7, i_7r0[5:5]);
  AND2 I190 (gfint_7[6:6], choice_7, i_7r0[6:6]);
  AND2 I191 (gfint_7[7:7], choice_7, i_7r0[7:7]);
  OR2 I192 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I193 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I194 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I195 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I196 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I197 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I198 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I199 (comp0_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  C3 I200 (simp1871_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I201 (simp1871_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C2 I202 (simp1871_0[2:2], comp0_0[6:6], comp0_0[7:7]);
  C3 I203 (icomp_0, simp1871_0[0:0], simp1871_0[1:1], simp1871_0[2:2]);
  OR2 I204 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I205 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I206 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I207 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I208 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I209 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I210 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  OR2 I211 (comp1_0[7:7], i_1r0[7:7], i_1r1[7:7]);
  C3 I212 (simp1971_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I213 (simp1971_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  C2 I214 (simp1971_0[2:2], comp1_0[6:6], comp1_0[7:7]);
  C3 I215 (icomp_1, simp1971_0[0:0], simp1971_0[1:1], simp1971_0[2:2]);
  OR2 I216 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I217 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I218 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2 I219 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  OR2 I220 (comp2_0[4:4], i_2r0[4:4], i_2r1[4:4]);
  OR2 I221 (comp2_0[5:5], i_2r0[5:5], i_2r1[5:5]);
  OR2 I222 (comp2_0[6:6], i_2r0[6:6], i_2r1[6:6]);
  OR2 I223 (comp2_0[7:7], i_2r0[7:7], i_2r1[7:7]);
  C3 I224 (simp2071_0[0:0], comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C3 I225 (simp2071_0[1:1], comp2_0[3:3], comp2_0[4:4], comp2_0[5:5]);
  C2 I226 (simp2071_0[2:2], comp2_0[6:6], comp2_0[7:7]);
  C3 I227 (icomp_2, simp2071_0[0:0], simp2071_0[1:1], simp2071_0[2:2]);
  OR2 I228 (comp3_0[0:0], i_3r0[0:0], i_3r1[0:0]);
  OR2 I229 (comp3_0[1:1], i_3r0[1:1], i_3r1[1:1]);
  OR2 I230 (comp3_0[2:2], i_3r0[2:2], i_3r1[2:2]);
  OR2 I231 (comp3_0[3:3], i_3r0[3:3], i_3r1[3:3]);
  OR2 I232 (comp3_0[4:4], i_3r0[4:4], i_3r1[4:4]);
  OR2 I233 (comp3_0[5:5], i_3r0[5:5], i_3r1[5:5]);
  OR2 I234 (comp3_0[6:6], i_3r0[6:6], i_3r1[6:6]);
  OR2 I235 (comp3_0[7:7], i_3r0[7:7], i_3r1[7:7]);
  C3 I236 (simp2171_0[0:0], comp3_0[0:0], comp3_0[1:1], comp3_0[2:2]);
  C3 I237 (simp2171_0[1:1], comp3_0[3:3], comp3_0[4:4], comp3_0[5:5]);
  C2 I238 (simp2171_0[2:2], comp3_0[6:6], comp3_0[7:7]);
  C3 I239 (icomp_3, simp2171_0[0:0], simp2171_0[1:1], simp2171_0[2:2]);
  OR2 I240 (comp4_0[0:0], i_4r0[0:0], i_4r1[0:0]);
  OR2 I241 (comp4_0[1:1], i_4r0[1:1], i_4r1[1:1]);
  OR2 I242 (comp4_0[2:2], i_4r0[2:2], i_4r1[2:2]);
  OR2 I243 (comp4_0[3:3], i_4r0[3:3], i_4r1[3:3]);
  OR2 I244 (comp4_0[4:4], i_4r0[4:4], i_4r1[4:4]);
  OR2 I245 (comp4_0[5:5], i_4r0[5:5], i_4r1[5:5]);
  OR2 I246 (comp4_0[6:6], i_4r0[6:6], i_4r1[6:6]);
  OR2 I247 (comp4_0[7:7], i_4r0[7:7], i_4r1[7:7]);
  C3 I248 (simp2271_0[0:0], comp4_0[0:0], comp4_0[1:1], comp4_0[2:2]);
  C3 I249 (simp2271_0[1:1], comp4_0[3:3], comp4_0[4:4], comp4_0[5:5]);
  C2 I250 (simp2271_0[2:2], comp4_0[6:6], comp4_0[7:7]);
  C3 I251 (icomp_4, simp2271_0[0:0], simp2271_0[1:1], simp2271_0[2:2]);
  OR2 I252 (comp5_0[0:0], i_5r0[0:0], i_5r1[0:0]);
  OR2 I253 (comp5_0[1:1], i_5r0[1:1], i_5r1[1:1]);
  OR2 I254 (comp5_0[2:2], i_5r0[2:2], i_5r1[2:2]);
  OR2 I255 (comp5_0[3:3], i_5r0[3:3], i_5r1[3:3]);
  OR2 I256 (comp5_0[4:4], i_5r0[4:4], i_5r1[4:4]);
  OR2 I257 (comp5_0[5:5], i_5r0[5:5], i_5r1[5:5]);
  OR2 I258 (comp5_0[6:6], i_5r0[6:6], i_5r1[6:6]);
  OR2 I259 (comp5_0[7:7], i_5r0[7:7], i_5r1[7:7]);
  C3 I260 (simp2371_0[0:0], comp5_0[0:0], comp5_0[1:1], comp5_0[2:2]);
  C3 I261 (simp2371_0[1:1], comp5_0[3:3], comp5_0[4:4], comp5_0[5:5]);
  C2 I262 (simp2371_0[2:2], comp5_0[6:6], comp5_0[7:7]);
  C3 I263 (icomp_5, simp2371_0[0:0], simp2371_0[1:1], simp2371_0[2:2]);
  OR2 I264 (comp6_0[0:0], i_6r0[0:0], i_6r1[0:0]);
  OR2 I265 (comp6_0[1:1], i_6r0[1:1], i_6r1[1:1]);
  OR2 I266 (comp6_0[2:2], i_6r0[2:2], i_6r1[2:2]);
  OR2 I267 (comp6_0[3:3], i_6r0[3:3], i_6r1[3:3]);
  OR2 I268 (comp6_0[4:4], i_6r0[4:4], i_6r1[4:4]);
  OR2 I269 (comp6_0[5:5], i_6r0[5:5], i_6r1[5:5]);
  OR2 I270 (comp6_0[6:6], i_6r0[6:6], i_6r1[6:6]);
  OR2 I271 (comp6_0[7:7], i_6r0[7:7], i_6r1[7:7]);
  C3 I272 (simp2471_0[0:0], comp6_0[0:0], comp6_0[1:1], comp6_0[2:2]);
  C3 I273 (simp2471_0[1:1], comp6_0[3:3], comp6_0[4:4], comp6_0[5:5]);
  C2 I274 (simp2471_0[2:2], comp6_0[6:6], comp6_0[7:7]);
  C3 I275 (icomp_6, simp2471_0[0:0], simp2471_0[1:1], simp2471_0[2:2]);
  OR2 I276 (comp7_0[0:0], i_7r0[0:0], i_7r1[0:0]);
  OR2 I277 (comp7_0[1:1], i_7r0[1:1], i_7r1[1:1]);
  OR2 I278 (comp7_0[2:2], i_7r0[2:2], i_7r1[2:2]);
  OR2 I279 (comp7_0[3:3], i_7r0[3:3], i_7r1[3:3]);
  OR2 I280 (comp7_0[4:4], i_7r0[4:4], i_7r1[4:4]);
  OR2 I281 (comp7_0[5:5], i_7r0[5:5], i_7r1[5:5]);
  OR2 I282 (comp7_0[6:6], i_7r0[6:6], i_7r1[6:6]);
  OR2 I283 (comp7_0[7:7], i_7r0[7:7], i_7r1[7:7]);
  C3 I284 (simp2571_0[0:0], comp7_0[0:0], comp7_0[1:1], comp7_0[2:2]);
  C3 I285 (simp2571_0[1:1], comp7_0[3:3], comp7_0[4:4], comp7_0[5:5]);
  C2 I286 (simp2571_0[2:2], comp7_0[6:6], comp7_0[7:7]);
  C3 I287 (icomp_7, simp2571_0[0:0], simp2571_0[1:1], simp2571_0[2:2]);
  C2R I288 (choice_0, icomp_0, nchosen_0, reset);
  C2R I289 (choice_1, icomp_1, nchosen_0, reset);
  C2R I290 (choice_2, icomp_2, nchosen_0, reset);
  C2R I291 (choice_3, icomp_3, nchosen_0, reset);
  C2R I292 (choice_4, icomp_4, nchosen_0, reset);
  C2R I293 (choice_5, icomp_5, nchosen_0, reset);
  C2R I294 (choice_6, icomp_6, nchosen_0, reset);
  C2R I295 (choice_7, icomp_7, nchosen_0, reset);
  NOR3 I296 (simp2661_0[0:0], choice_0, choice_1, choice_2);
  NOR3 I297 (simp2661_0[1:1], choice_3, choice_4, choice_5);
  NOR2 I298 (simp2661_0[2:2], choice_6, choice_7);
  NAND3 I299 (anychoice_0, simp2661_0[0:0], simp2661_0[1:1], simp2661_0[2:2]);
  NOR2 I300 (nchosen_0, anychoice_0, o_0a);
  C2R I301 (i_0a, choice_0, o_0a, reset);
  C2R I302 (i_1a, choice_1, o_0a, reset);
  C2R I303 (i_2a, choice_2, o_0a, reset);
  C2R I304 (i_3a, choice_3, o_0a, reset);
  C2R I305 (i_4a, choice_4, o_0a, reset);
  C2R I306 (i_5a, choice_5, o_0a, reset);
  C2R I307 (i_6a, choice_6, o_0a, reset);
  C2R I308 (i_7a, choice_7, o_0a, reset);
endmodule

// tkj8m0_8 TeakJ [Many [0,8],One 8]
module tkj8m0_8 (i_0r, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  input [7:0] i_1r0;
  input [7:0] i_1r1;
  output i_1a;
  output [7:0] o_0r0;
  output [7:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [7:0] joinf_0;
  wire [7:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_1r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_1r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_1r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_1r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_1r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_1r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_1r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_1r0[7:7]);
  BUFF I8 (joint_0[0:0], i_1r1[0:0]);
  BUFF I9 (joint_0[1:1], i_1r1[1:1]);
  BUFF I10 (joint_0[2:2], i_1r1[2:2]);
  BUFF I11 (joint_0[3:3], i_1r1[3:3]);
  BUFF I12 (joint_0[4:4], i_1r1[4:4]);
  BUFF I13 (joint_0[5:5], i_1r1[5:5]);
  BUFF I14 (joint_0[6:6], i_1r1[6:6]);
  BUFF I15 (joint_0[7:7], i_1r1[7:7]);
  BUFF I16 (icomplete_0, i_0r);
  C2 I17 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I18 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I19 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I20 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I21 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I22 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I23 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I24 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I25 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I26 (o_0r1[1:1], joint_0[1:1]);
  BUFF I27 (o_0r1[2:2], joint_0[2:2]);
  BUFF I28 (o_0r1[3:3], joint_0[3:3]);
  BUFF I29 (o_0r1[4:4], joint_0[4:4]);
  BUFF I30 (o_0r1[5:5], joint_0[5:5]);
  BUFF I31 (o_0r1[6:6], joint_0[6:6]);
  BUFF I32 (o_0r1[7:7], joint_0[7:7]);
  BUFF I33 (i_0a, o_0a);
  BUFF I34 (i_1a, o_0a);
endmodule

// tks8_o0w8_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0_20o0w0_40o0w0_80o0w0 TeakS (0+:8) [([Imp 1 0],0),([Imp 2 0]
//   ,0),([Imp 4 0],0),([Imp 8 0],0),([Imp 16 0],0),([Imp 32 0],0),([Imp 64 0],0),([Imp 128 0],0)] [One 8
//   ,Many [0,0,0,0,0,0,0,0]]
module tks8_o0w8_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0_20o0w0_40o0w0_80o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, o_5r, o_5a, o_6r, o_6a, o_7r, o_7a, reset);
  input [7:0] i_0r0;
  input [7:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  output o_7r;
  input o_7a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire sel_4;
  wire sel_5;
  wire sel_6;
  wire sel_7;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire gsel_4;
  wire gsel_5;
  wire gsel_6;
  wire gsel_7;
  wire oack_0;
  wire match0_0;
  wire [2:0] simp201_0;
  wire match1_0;
  wire [2:0] simp231_0;
  wire match2_0;
  wire [2:0] simp261_0;
  wire match3_0;
  wire [2:0] simp291_0;
  wire match4_0;
  wire [2:0] simp321_0;
  wire match5_0;
  wire [2:0] simp351_0;
  wire match6_0;
  wire [2:0] simp381_0;
  wire match7_0;
  wire [2:0] simp411_0;
  wire [7:0] comp_0;
  wire [2:0] simp591_0;
  wire [2:0] simp681_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (simp201_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I2 (simp201_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I3 (simp201_0[2:2], i_0r0[6:6], i_0r0[7:7]);
  C3 I4 (match0_0, simp201_0[0:0], simp201_0[1:1], simp201_0[2:2]);
  BUFF I5 (sel_1, match1_0);
  C3 I6 (simp231_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I7 (simp231_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I8 (simp231_0[2:2], i_0r0[6:6], i_0r0[7:7]);
  C3 I9 (match1_0, simp231_0[0:0], simp231_0[1:1], simp231_0[2:2]);
  BUFF I10 (sel_2, match2_0);
  C3 I11 (simp261_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I12 (simp261_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I13 (simp261_0[2:2], i_0r0[6:6], i_0r0[7:7]);
  C3 I14 (match2_0, simp261_0[0:0], simp261_0[1:1], simp261_0[2:2]);
  BUFF I15 (sel_3, match3_0);
  C3 I16 (simp291_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I17 (simp291_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I18 (simp291_0[2:2], i_0r0[6:6], i_0r0[7:7]);
  C3 I19 (match3_0, simp291_0[0:0], simp291_0[1:1], simp291_0[2:2]);
  BUFF I20 (sel_4, match4_0);
  C3 I21 (simp321_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I22 (simp321_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  C2 I23 (simp321_0[2:2], i_0r0[6:6], i_0r0[7:7]);
  C3 I24 (match4_0, simp321_0[0:0], simp321_0[1:1], simp321_0[2:2]);
  BUFF I25 (sel_5, match5_0);
  C3 I26 (simp351_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I27 (simp351_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  C2 I28 (simp351_0[2:2], i_0r0[6:6], i_0r0[7:7]);
  C3 I29 (match5_0, simp351_0[0:0], simp351_0[1:1], simp351_0[2:2]);
  BUFF I30 (sel_6, match6_0);
  C3 I31 (simp381_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I32 (simp381_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I33 (simp381_0[2:2], i_0r1[6:6], i_0r0[7:7]);
  C3 I34 (match6_0, simp381_0[0:0], simp381_0[1:1], simp381_0[2:2]);
  BUFF I35 (sel_7, match7_0);
  C3 I36 (simp411_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I37 (simp411_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  C2 I38 (simp411_0[2:2], i_0r0[6:6], i_0r1[7:7]);
  C3 I39 (match7_0, simp411_0[0:0], simp411_0[1:1], simp411_0[2:2]);
  C2 I40 (gsel_0, sel_0, icomplete_0);
  C2 I41 (gsel_1, sel_1, icomplete_0);
  C2 I42 (gsel_2, sel_2, icomplete_0);
  C2 I43 (gsel_3, sel_3, icomplete_0);
  C2 I44 (gsel_4, sel_4, icomplete_0);
  C2 I45 (gsel_5, sel_5, icomplete_0);
  C2 I46 (gsel_6, sel_6, icomplete_0);
  C2 I47 (gsel_7, sel_7, icomplete_0);
  OR2 I48 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I49 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I50 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I51 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I52 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I53 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I54 (comp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I55 (comp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  C3 I56 (simp591_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I57 (simp591_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C2 I58 (simp591_0[2:2], comp_0[6:6], comp_0[7:7]);
  C3 I59 (icomplete_0, simp591_0[0:0], simp591_0[1:1], simp591_0[2:2]);
  BUFF I60 (o_0r, gsel_0);
  BUFF I61 (o_1r, gsel_1);
  BUFF I62 (o_2r, gsel_2);
  BUFF I63 (o_3r, gsel_3);
  BUFF I64 (o_4r, gsel_4);
  BUFF I65 (o_5r, gsel_5);
  BUFF I66 (o_6r, gsel_6);
  BUFF I67 (o_7r, gsel_7);
  NOR3 I68 (simp681_0[0:0], o_0a, o_1a, o_2a);
  NOR3 I69 (simp681_0[1:1], o_3a, o_4a, o_5a);
  NOR2 I70 (simp681_0[2:2], o_6a, o_7a);
  NAND3 I71 (oack_0, simp681_0[0:0], simp681_0[1:1], simp681_0[2:2]);
  C2 I72 (i_0a, oack_0, icomplete_0);
endmodule

// tkj7m6_1 TeakJ [Many [6,1],One 7]
module tkj7m6_1 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [5:0] i_0r0;
  input [5:0] i_0r1;
  output i_0a;
  input i_1r0;
  input i_1r1;
  output i_1a;
  output [6:0] o_0r0;
  output [6:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [6:0] joinf_0;
  wire [6:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_1r0);
  BUFF I7 (joint_0[0:0], i_0r1[0:0]);
  BUFF I8 (joint_0[1:1], i_0r1[1:1]);
  BUFF I9 (joint_0[2:2], i_0r1[2:2]);
  BUFF I10 (joint_0[3:3], i_0r1[3:3]);
  BUFF I11 (joint_0[4:4], i_0r1[4:4]);
  BUFF I12 (joint_0[5:5], i_0r1[5:5]);
  BUFF I13 (joint_0[6:6], i_1r1);
  OR2 I14 (dcomplete_0, i_1r0, i_1r1);
  BUFF I15 (icomplete_0, dcomplete_0);
  C2 I16 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I17 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I18 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I19 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I20 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I21 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I22 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I23 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I24 (o_0r1[1:1], joint_0[1:1]);
  BUFF I25 (o_0r1[2:2], joint_0[2:2]);
  BUFF I26 (o_0r1[3:3], joint_0[3:3]);
  BUFF I27 (o_0r1[4:4], joint_0[4:4]);
  BUFF I28 (o_0r1[5:5], joint_0[5:5]);
  BUFF I29 (o_0r1[6:6], joint_0[6:6]);
  BUFF I30 (i_0a, o_0a);
  BUFF I31 (i_1a, o_0a);
endmodule

// tkvaluResult32_wo0w32_ro0w32 TeakV "aluResult" 32 [] [0] [0] [Many [32],Many [0],Many [0],Many [32]]
module tkvaluResult32_wo0w32_ro0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I457 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I458 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I459 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I460 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I461 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I462 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I463 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I464 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I465 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I466 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I467 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I468 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I469 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I470 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I471 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I472 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I473 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I474 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I475 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I476 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I477 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I478 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I479 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I480 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I481 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I482 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I483 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I484 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I485 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I486 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I487 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  OR2 I488 (anyread_0, rg_0r, rg_0a);
  BUFF I489 (wg_0a, wd_0a);
  BUFF I490 (rg_0a, rd_0a);
endmodule

// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0 TeakF [0,0,0,0,0,0] [One 0,Many [0,0,0,0,0,0]]
module tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, o_5r, o_5a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  input reset;
  wire [1:0] simp11_0;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  BUFF I2 (o_2r, i_0r);
  BUFF I3 (o_3r, i_0r);
  BUFF I4 (o_4r, i_0r);
  BUFF I5 (o_5r, i_0r);
  C3 I6 (simp11_0[0:0], o_0a, o_1a, o_2a);
  C3 I7 (simp11_0[1:1], o_3a, o_4a, o_5a);
  C2 I8 (i_0a, simp11_0[0:0], simp11_0[1:1]);
endmodule

// tkj0m0_0_0_0_0_0 TeakJ [Many [0,0,0,0,0,0],One 0]
module tkj0m0_0_0_0_0_0 (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, i_3r, i_3a, i_4r, i_4a, i_5r, i_5a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  input i_4r;
  output i_4a;
  input i_5r;
  output i_5a;
  output o_0r;
  input o_0a;
  input reset;
  wire [1:0] simp01_0;
  C3 I0 (simp01_0[0:0], i_0r, i_1r, i_2r);
  C3 I1 (simp01_0[1:1], i_3r, i_4r, i_5r);
  C2 I2 (o_0r, simp01_0[0:0], simp01_0[1:1]);
  BUFF I3 (i_0a, o_0a);
  BUFF I4 (i_1a, o_0a);
  BUFF I5 (i_2a, o_0a);
  BUFF I6 (i_3a, o_0a);
  BUFF I7 (i_4a, o_0a);
  BUFF I8 (i_5a, o_0a);
endmodule

// tkj3m1_2 TeakJ [Many [1,2],One 3]
module tkj3m1_2 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r0;
  input i_0r1;
  output i_0a;
  input [1:0] i_1r0;
  input [1:0] i_1r1;
  output i_1a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [2:0] joinf_0;
  wire [2:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0);
  BUFF I1 (joinf_0[1:1], i_1r0[0:0]);
  BUFF I2 (joinf_0[2:2], i_1r0[1:1]);
  BUFF I3 (joint_0[0:0], i_0r1);
  BUFF I4 (joint_0[1:1], i_1r1[0:0]);
  BUFF I5 (joint_0[2:2], i_1r1[1:1]);
  OR2 I6 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I7 (icomplete_0, dcomplete_0);
  C2 I8 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I9 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I10 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I11 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I12 (o_0r1[1:1], joint_0[1:1]);
  BUFF I13 (o_0r1[2:2], joint_0[2:2]);
  BUFF I14 (i_0a, o_0a);
  BUFF I15 (i_1a, o_0a);
endmodule

// tkf4mo0w0 TeakF [0] [One 4,Many [0]]
module tkf4mo0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  wire ucomplete_0;
  wire [3:0] comp_0;
  wire [1:0] simp91_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I2 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I3 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I4 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  C3 I5 (simp91_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  BUFF I6 (simp91_0[1:1], comp_0[3:3]);
  C2 I7 (ucomplete_0, simp91_0[0:0], simp91_0[1:1]);
  C2 I8 (acomplete_0, ucomplete_0, icomplete_0);
  BUFF I9 (o_0r, icomplete_0);
  C2 I10 (i_0a, acomplete_0, o_0a);
endmodule

// tkvdread32_wo0w32_ro0w32 TeakV "dread" 32 [] [0] [0] [Many [32],Many [0],Many [0],Many [32]]
module tkvdread32_wo0w32_ro0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I457 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I458 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I459 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I460 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I461 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I462 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I463 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I464 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I465 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I466 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I467 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I468 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I469 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I470 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I471 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I472 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I473 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I474 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I475 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I476 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I477 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I478 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I479 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I480 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I481 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I482 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I483 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I484 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I485 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I486 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I487 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  OR2 I488 (anyread_0, rg_0r, rg_0a);
  BUFF I489 (wg_0a, wd_0a);
  BUFF I490 (rg_0a, rd_0a);
endmodule

// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 TeakF [0,0,0,0,0,0,0,0] [One 0,Many [0,0,0,0,0,0,0,0]]
module tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, o_5r, o_5a, o_6r, o_6a, o_7r, o_7a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  output o_7r;
  input o_7a;
  input reset;
  wire [2:0] simp11_0;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  BUFF I2 (o_2r, i_0r);
  BUFF I3 (o_3r, i_0r);
  BUFF I4 (o_4r, i_0r);
  BUFF I5 (o_5r, i_0r);
  BUFF I6 (o_6r, i_0r);
  BUFF I7 (o_7r, i_0r);
  C3 I8 (simp11_0[0:0], o_0a, o_1a, o_2a);
  C3 I9 (simp11_0[1:1], o_3a, o_4a, o_5a);
  C2 I10 (simp11_0[2:2], o_6a, o_7a);
  C3 I11 (i_0a, simp11_0[0:0], simp11_0[1:1], simp11_0[2:2]);
endmodule

// tkj0m0_0_0_0_0_0_0_0 TeakJ [Many [0,0,0,0,0,0,0,0],One 0]
module tkj0m0_0_0_0_0_0_0_0 (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, i_3r, i_3a, i_4r, i_4a, i_5r, i_5a, i_6r, i_6a, i_7r, i_7a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  input i_4r;
  output i_4a;
  input i_5r;
  output i_5a;
  input i_6r;
  output i_6a;
  input i_7r;
  output i_7a;
  output o_0r;
  input o_0a;
  input reset;
  wire [2:0] simp01_0;
  C3 I0 (simp01_0[0:0], i_0r, i_1r, i_2r);
  C3 I1 (simp01_0[1:1], i_3r, i_4r, i_5r);
  C2 I2 (simp01_0[2:2], i_6r, i_7r);
  C3 I3 (o_0r, simp01_0[0:0], simp01_0[1:1], simp01_0[2:2]);
  BUFF I4 (i_0a, o_0a);
  BUFF I5 (i_1a, o_0a);
  BUFF I6 (i_2a, o_0a);
  BUFF I7 (i_3a, o_0a);
  BUFF I8 (i_4a, o_0a);
  BUFF I9 (i_5a, o_0a);
  BUFF I10 (i_6a, o_0a);
  BUFF I11 (i_7a, o_0a);
endmodule

// tkvr232_wo0w32_ro0w32 TeakV "r2" 32 [] [0] [0] [Many [32],Many [0],Many [0],Many [32]]
module tkvr232_wo0w32_ro0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I457 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I458 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I459 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I460 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I461 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I462 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I463 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I464 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I465 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I466 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I467 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I468 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I469 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I470 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I471 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I472 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I473 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I474 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I475 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I476 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I477 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I478 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I479 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I480 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I481 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I482 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I483 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I484 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I485 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I486 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I487 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  OR2 I488 (anyread_0, rg_0r, rg_0a);
  BUFF I489 (wg_0a, wd_0a);
  BUFF I490 (rg_0a, rd_0a);
endmodule

// tks3_o0w3_7o0w0_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0 TeakS (0+:3) [([Imp 7 0],0),([Imp 0 0],0),
//   ([Imp 1 0],0),([Imp 2 0],0),([Imp 3 0],0),([Imp 4 0],0),([Imp 5 0],0),([Imp 6 0],0)] [One 3,Many [0,
//   0,0,0,0,0,0,0]]
module tks3_o0w3_7o0w0_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, o_5r, o_5a, o_6r, o_6a, o_7r, o_7a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  output o_7r;
  input o_7a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire sel_4;
  wire sel_5;
  wire sel_6;
  wire sel_7;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire gsel_4;
  wire gsel_5;
  wire gsel_6;
  wire gsel_7;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire match2_0;
  wire match3_0;
  wire match4_0;
  wire match5_0;
  wire match6_0;
  wire match7_0;
  wire [2:0] comp_0;
  wire [2:0] simp631_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (match0_0, i_0r1[0:0], i_0r1[1:1], i_0r1[2:2]);
  BUFF I2 (sel_1, match1_0);
  C3 I3 (match1_0, i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I4 (sel_2, match2_0);
  C3 I5 (match2_0, i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  BUFF I6 (sel_3, match3_0);
  C3 I7 (match3_0, i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I8 (sel_4, match4_0);
  C3 I9 (match4_0, i_0r1[0:0], i_0r1[1:1], i_0r0[2:2]);
  BUFF I10 (sel_5, match5_0);
  C3 I11 (match5_0, i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I12 (sel_6, match6_0);
  C3 I13 (match6_0, i_0r1[0:0], i_0r0[1:1], i_0r1[2:2]);
  BUFF I14 (sel_7, match7_0);
  C3 I15 (match7_0, i_0r0[0:0], i_0r1[1:1], i_0r1[2:2]);
  C2 I16 (gsel_0, sel_0, icomplete_0);
  C2 I17 (gsel_1, sel_1, icomplete_0);
  C2 I18 (gsel_2, sel_2, icomplete_0);
  C2 I19 (gsel_3, sel_3, icomplete_0);
  C2 I20 (gsel_4, sel_4, icomplete_0);
  C2 I21 (gsel_5, sel_5, icomplete_0);
  C2 I22 (gsel_6, sel_6, icomplete_0);
  C2 I23 (gsel_7, sel_7, icomplete_0);
  OR2 I24 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I25 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I26 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I27 (icomplete_0, comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  BUFF I28 (o_0r, gsel_0);
  BUFF I29 (o_1r, gsel_1);
  BUFF I30 (o_2r, gsel_2);
  BUFF I31 (o_3r, gsel_3);
  BUFF I32 (o_4r, gsel_4);
  BUFF I33 (o_5r, gsel_5);
  BUFF I34 (o_6r, gsel_6);
  BUFF I35 (o_7r, gsel_7);
  NOR3 I36 (simp631_0[0:0], o_0a, o_1a, o_2a);
  NOR3 I37 (simp631_0[1:1], o_3a, o_4a, o_5a);
  NOR2 I38 (simp631_0[2:2], o_6a, o_7a);
  NAND3 I39 (oack_0, simp631_0[0:0], simp631_0[1:1], simp631_0[2:2]);
  C2 I40 (i_0a, oack_0, icomplete_0);
endmodule

// tko0m7_1nm7b1 TeakO [
//     (1,TeakOConstant 7 1)] [One 0,One 7]
module tko0m7_1nm7b1 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [6:0] o_0r0;
  output [6:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[0:0], i_0r);
  GND I1 (o_0r0[0:0]);
  BUFF I2 (o_0r0[1:1], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  BUFF I6 (o_0r0[5:5], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  GND I8 (o_0r1[1:1]);
  GND I9 (o_0r1[2:2]);
  GND I10 (o_0r1[3:3]);
  GND I11 (o_0r1[4:4]);
  GND I12 (o_0r1[5:5]);
  GND I13 (o_0r1[6:6]);
  BUFF I14 (i_0a, o_0a);
endmodule

// tko0m7_1nm7b2 TeakO [
//     (1,TeakOConstant 7 2)] [One 0,One 7]
module tko0m7_1nm7b2 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [6:0] o_0r0;
  output [6:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[1:1], i_0r);
  GND I1 (o_0r0[1:1]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[2:2], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  BUFF I6 (o_0r0[5:5], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  GND I8 (o_0r1[0:0]);
  GND I9 (o_0r1[2:2]);
  GND I10 (o_0r1[3:3]);
  GND I11 (o_0r1[4:4]);
  GND I12 (o_0r1[5:5]);
  GND I13 (o_0r1[6:6]);
  BUFF I14 (i_0a, o_0a);
endmodule

// tko0m7_1nm7b4 TeakO [
//     (1,TeakOConstant 7 4)] [One 0,One 7]
module tko0m7_1nm7b4 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [6:0] o_0r0;
  output [6:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[2:2], i_0r);
  GND I1 (o_0r0[2:2]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[3:3], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  BUFF I6 (o_0r0[5:5], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  GND I8 (o_0r1[0:0]);
  GND I9 (o_0r1[1:1]);
  GND I10 (o_0r1[3:3]);
  GND I11 (o_0r1[4:4]);
  GND I12 (o_0r1[5:5]);
  GND I13 (o_0r1[6:6]);
  BUFF I14 (i_0a, o_0a);
endmodule

// tko0m7_1nm7b8 TeakO [
//     (1,TeakOConstant 7 8)] [One 0,One 7]
module tko0m7_1nm7b8 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [6:0] o_0r0;
  output [6:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[3:3], i_0r);
  GND I1 (o_0r0[3:3]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[4:4], i_0r);
  BUFF I6 (o_0r0[5:5], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  GND I8 (o_0r1[0:0]);
  GND I9 (o_0r1[1:1]);
  GND I10 (o_0r1[2:2]);
  GND I11 (o_0r1[4:4]);
  GND I12 (o_0r1[5:5]);
  GND I13 (o_0r1[6:6]);
  BUFF I14 (i_0a, o_0a);
endmodule

// tko0m7_1nm7b10 TeakO [
//     (1,TeakOConstant 7 16)] [One 0,One 7]
module tko0m7_1nm7b10 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [6:0] o_0r0;
  output [6:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[4:4], i_0r);
  GND I1 (o_0r0[4:4]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  BUFF I6 (o_0r0[5:5], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  GND I8 (o_0r1[0:0]);
  GND I9 (o_0r1[1:1]);
  GND I10 (o_0r1[2:2]);
  GND I11 (o_0r1[3:3]);
  GND I12 (o_0r1[5:5]);
  GND I13 (o_0r1[6:6]);
  BUFF I14 (i_0a, o_0a);
endmodule

// tko0m7_1nm7b20 TeakO [
//     (1,TeakOConstant 7 32)] [One 0,One 7]
module tko0m7_1nm7b20 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [6:0] o_0r0;
  output [6:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[5:5], i_0r);
  GND I1 (o_0r0[5:5]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  BUFF I6 (o_0r0[4:4], i_0r);
  BUFF I7 (o_0r0[6:6], i_0r);
  GND I8 (o_0r1[0:0]);
  GND I9 (o_0r1[1:1]);
  GND I10 (o_0r1[2:2]);
  GND I11 (o_0r1[3:3]);
  GND I12 (o_0r1[4:4]);
  GND I13 (o_0r1[6:6]);
  BUFF I14 (i_0a, o_0a);
endmodule

// tko0m7_1nm7b40 TeakO [
//     (1,TeakOConstant 7 64)] [One 0,One 7]
module tko0m7_1nm7b40 (i_0r, i_0a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  output [6:0] o_0r0;
  output [6:0] o_0r1;
  input o_0a;
  input reset;
  BUFF I0 (o_0r1[6:6], i_0r);
  GND I1 (o_0r0[6:6]);
  BUFF I2 (o_0r0[0:0], i_0r);
  BUFF I3 (o_0r0[1:1], i_0r);
  BUFF I4 (o_0r0[2:2], i_0r);
  BUFF I5 (o_0r0[3:3], i_0r);
  BUFF I6 (o_0r0[4:4], i_0r);
  BUFF I7 (o_0r0[5:5], i_0r);
  GND I8 (o_0r1[0:0]);
  GND I9 (o_0r1[1:1]);
  GND I10 (o_0r1[2:2]);
  GND I11 (o_0r1[3:3]);
  GND I12 (o_0r1[4:4]);
  GND I13 (o_0r1[5:5]);
  BUFF I14 (i_0a, o_0a);
endmodule

// tkm7x7b TeakM [Many [7,7,7,7,7,7,7],One 7]
module tkm7x7b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, i_3r0, i_3r1, i_3a, i_4r0, i_4r1, i_4a, i_5r0, i_5r1, i_5a, i_6r0, i_6r1, i_6a, o_0r0, o_0r1, o_0a, reset);
  input [6:0] i_0r0;
  input [6:0] i_0r1;
  output i_0a;
  input [6:0] i_1r0;
  input [6:0] i_1r1;
  output i_1a;
  input [6:0] i_2r0;
  input [6:0] i_2r1;
  output i_2a;
  input [6:0] i_3r0;
  input [6:0] i_3r1;
  output i_3a;
  input [6:0] i_4r0;
  input [6:0] i_4r1;
  output i_4a;
  input [6:0] i_5r0;
  input [6:0] i_5r1;
  output i_5a;
  input [6:0] i_6r0;
  input [6:0] i_6r1;
  output i_6a;
  output [6:0] o_0r0;
  output [6:0] o_0r1;
  input o_0a;
  input reset;
  wire [6:0] gfint_0;
  wire [6:0] gfint_1;
  wire [6:0] gfint_2;
  wire [6:0] gfint_3;
  wire [6:0] gfint_4;
  wire [6:0] gfint_5;
  wire [6:0] gfint_6;
  wire [6:0] gtint_0;
  wire [6:0] gtint_1;
  wire [6:0] gtint_2;
  wire [6:0] gtint_3;
  wire [6:0] gtint_4;
  wire [6:0] gtint_5;
  wire [6:0] gtint_6;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire choice_3;
  wire choice_4;
  wire choice_5;
  wire choice_6;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire icomp_3;
  wire icomp_4;
  wire icomp_5;
  wire icomp_6;
  wire nchosen_0;
  wire [2:0] simp301_0;
  wire [2:0] simp311_0;
  wire [2:0] simp321_0;
  wire [2:0] simp331_0;
  wire [2:0] simp341_0;
  wire [2:0] simp351_0;
  wire [2:0] simp361_0;
  wire [2:0] simp371_0;
  wire [2:0] simp381_0;
  wire [2:0] simp391_0;
  wire [2:0] simp401_0;
  wire [2:0] simp411_0;
  wire [2:0] simp421_0;
  wire [2:0] simp431_0;
  wire [6:0] comp0_0;
  wire [2:0] simp1501_0;
  wire [6:0] comp1_0;
  wire [2:0] simp1591_0;
  wire [6:0] comp2_0;
  wire [2:0] simp1681_0;
  wire [6:0] comp3_0;
  wire [2:0] simp1771_0;
  wire [6:0] comp4_0;
  wire [2:0] simp1861_0;
  wire [6:0] comp5_0;
  wire [2:0] simp1951_0;
  wire [6:0] comp6_0;
  wire [2:0] simp2041_0;
  wire [2:0] simp2121_0;
  NOR3 I0 (simp301_0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  NOR3 I1 (simp301_0[1:1], gfint_3[0:0], gfint_4[0:0], gfint_5[0:0]);
  INV I2 (simp301_0[2:2], gfint_6[0:0]);
  NAND3 I3 (o_0r0[0:0], simp301_0[0:0], simp301_0[1:1], simp301_0[2:2]);
  NOR3 I4 (simp311_0[0:0], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  NOR3 I5 (simp311_0[1:1], gfint_3[1:1], gfint_4[1:1], gfint_5[1:1]);
  INV I6 (simp311_0[2:2], gfint_6[1:1]);
  NAND3 I7 (o_0r0[1:1], simp311_0[0:0], simp311_0[1:1], simp311_0[2:2]);
  NOR3 I8 (simp321_0[0:0], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  NOR3 I9 (simp321_0[1:1], gfint_3[2:2], gfint_4[2:2], gfint_5[2:2]);
  INV I10 (simp321_0[2:2], gfint_6[2:2]);
  NAND3 I11 (o_0r0[2:2], simp321_0[0:0], simp321_0[1:1], simp321_0[2:2]);
  NOR3 I12 (simp331_0[0:0], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  NOR3 I13 (simp331_0[1:1], gfint_3[3:3], gfint_4[3:3], gfint_5[3:3]);
  INV I14 (simp331_0[2:2], gfint_6[3:3]);
  NAND3 I15 (o_0r0[3:3], simp331_0[0:0], simp331_0[1:1], simp331_0[2:2]);
  NOR3 I16 (simp341_0[0:0], gfint_0[4:4], gfint_1[4:4], gfint_2[4:4]);
  NOR3 I17 (simp341_0[1:1], gfint_3[4:4], gfint_4[4:4], gfint_5[4:4]);
  INV I18 (simp341_0[2:2], gfint_6[4:4]);
  NAND3 I19 (o_0r0[4:4], simp341_0[0:0], simp341_0[1:1], simp341_0[2:2]);
  NOR3 I20 (simp351_0[0:0], gfint_0[5:5], gfint_1[5:5], gfint_2[5:5]);
  NOR3 I21 (simp351_0[1:1], gfint_3[5:5], gfint_4[5:5], gfint_5[5:5]);
  INV I22 (simp351_0[2:2], gfint_6[5:5]);
  NAND3 I23 (o_0r0[5:5], simp351_0[0:0], simp351_0[1:1], simp351_0[2:2]);
  NOR3 I24 (simp361_0[0:0], gfint_0[6:6], gfint_1[6:6], gfint_2[6:6]);
  NOR3 I25 (simp361_0[1:1], gfint_3[6:6], gfint_4[6:6], gfint_5[6:6]);
  INV I26 (simp361_0[2:2], gfint_6[6:6]);
  NAND3 I27 (o_0r0[6:6], simp361_0[0:0], simp361_0[1:1], simp361_0[2:2]);
  NOR3 I28 (simp371_0[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  NOR3 I29 (simp371_0[1:1], gtint_3[0:0], gtint_4[0:0], gtint_5[0:0]);
  INV I30 (simp371_0[2:2], gtint_6[0:0]);
  NAND3 I31 (o_0r1[0:0], simp371_0[0:0], simp371_0[1:1], simp371_0[2:2]);
  NOR3 I32 (simp381_0[0:0], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  NOR3 I33 (simp381_0[1:1], gtint_3[1:1], gtint_4[1:1], gtint_5[1:1]);
  INV I34 (simp381_0[2:2], gtint_6[1:1]);
  NAND3 I35 (o_0r1[1:1], simp381_0[0:0], simp381_0[1:1], simp381_0[2:2]);
  NOR3 I36 (simp391_0[0:0], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  NOR3 I37 (simp391_0[1:1], gtint_3[2:2], gtint_4[2:2], gtint_5[2:2]);
  INV I38 (simp391_0[2:2], gtint_6[2:2]);
  NAND3 I39 (o_0r1[2:2], simp391_0[0:0], simp391_0[1:1], simp391_0[2:2]);
  NOR3 I40 (simp401_0[0:0], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  NOR3 I41 (simp401_0[1:1], gtint_3[3:3], gtint_4[3:3], gtint_5[3:3]);
  INV I42 (simp401_0[2:2], gtint_6[3:3]);
  NAND3 I43 (o_0r1[3:3], simp401_0[0:0], simp401_0[1:1], simp401_0[2:2]);
  NOR3 I44 (simp411_0[0:0], gtint_0[4:4], gtint_1[4:4], gtint_2[4:4]);
  NOR3 I45 (simp411_0[1:1], gtint_3[4:4], gtint_4[4:4], gtint_5[4:4]);
  INV I46 (simp411_0[2:2], gtint_6[4:4]);
  NAND3 I47 (o_0r1[4:4], simp411_0[0:0], simp411_0[1:1], simp411_0[2:2]);
  NOR3 I48 (simp421_0[0:0], gtint_0[5:5], gtint_1[5:5], gtint_2[5:5]);
  NOR3 I49 (simp421_0[1:1], gtint_3[5:5], gtint_4[5:5], gtint_5[5:5]);
  INV I50 (simp421_0[2:2], gtint_6[5:5]);
  NAND3 I51 (o_0r1[5:5], simp421_0[0:0], simp421_0[1:1], simp421_0[2:2]);
  NOR3 I52 (simp431_0[0:0], gtint_0[6:6], gtint_1[6:6], gtint_2[6:6]);
  NOR3 I53 (simp431_0[1:1], gtint_3[6:6], gtint_4[6:6], gtint_5[6:6]);
  INV I54 (simp431_0[2:2], gtint_6[6:6]);
  NAND3 I55 (o_0r1[6:6], simp431_0[0:0], simp431_0[1:1], simp431_0[2:2]);
  AND2 I56 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I57 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I58 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I59 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I60 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I61 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I62 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I63 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I64 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I65 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I66 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I67 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I68 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I69 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I70 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I71 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I72 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I73 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AND2 I74 (gtint_2[4:4], choice_2, i_2r1[4:4]);
  AND2 I75 (gtint_2[5:5], choice_2, i_2r1[5:5]);
  AND2 I76 (gtint_2[6:6], choice_2, i_2r1[6:6]);
  AND2 I77 (gtint_3[0:0], choice_3, i_3r1[0:0]);
  AND2 I78 (gtint_3[1:1], choice_3, i_3r1[1:1]);
  AND2 I79 (gtint_3[2:2], choice_3, i_3r1[2:2]);
  AND2 I80 (gtint_3[3:3], choice_3, i_3r1[3:3]);
  AND2 I81 (gtint_3[4:4], choice_3, i_3r1[4:4]);
  AND2 I82 (gtint_3[5:5], choice_3, i_3r1[5:5]);
  AND2 I83 (gtint_3[6:6], choice_3, i_3r1[6:6]);
  AND2 I84 (gtint_4[0:0], choice_4, i_4r1[0:0]);
  AND2 I85 (gtint_4[1:1], choice_4, i_4r1[1:1]);
  AND2 I86 (gtint_4[2:2], choice_4, i_4r1[2:2]);
  AND2 I87 (gtint_4[3:3], choice_4, i_4r1[3:3]);
  AND2 I88 (gtint_4[4:4], choice_4, i_4r1[4:4]);
  AND2 I89 (gtint_4[5:5], choice_4, i_4r1[5:5]);
  AND2 I90 (gtint_4[6:6], choice_4, i_4r1[6:6]);
  AND2 I91 (gtint_5[0:0], choice_5, i_5r1[0:0]);
  AND2 I92 (gtint_5[1:1], choice_5, i_5r1[1:1]);
  AND2 I93 (gtint_5[2:2], choice_5, i_5r1[2:2]);
  AND2 I94 (gtint_5[3:3], choice_5, i_5r1[3:3]);
  AND2 I95 (gtint_5[4:4], choice_5, i_5r1[4:4]);
  AND2 I96 (gtint_5[5:5], choice_5, i_5r1[5:5]);
  AND2 I97 (gtint_5[6:6], choice_5, i_5r1[6:6]);
  AND2 I98 (gtint_6[0:0], choice_6, i_6r1[0:0]);
  AND2 I99 (gtint_6[1:1], choice_6, i_6r1[1:1]);
  AND2 I100 (gtint_6[2:2], choice_6, i_6r1[2:2]);
  AND2 I101 (gtint_6[3:3], choice_6, i_6r1[3:3]);
  AND2 I102 (gtint_6[4:4], choice_6, i_6r1[4:4]);
  AND2 I103 (gtint_6[5:5], choice_6, i_6r1[5:5]);
  AND2 I104 (gtint_6[6:6], choice_6, i_6r1[6:6]);
  AND2 I105 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I106 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I107 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I108 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I109 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I110 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I111 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I112 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I113 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I114 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I115 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I116 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I117 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I118 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I119 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I120 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I121 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I122 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AND2 I123 (gfint_2[4:4], choice_2, i_2r0[4:4]);
  AND2 I124 (gfint_2[5:5], choice_2, i_2r0[5:5]);
  AND2 I125 (gfint_2[6:6], choice_2, i_2r0[6:6]);
  AND2 I126 (gfint_3[0:0], choice_3, i_3r0[0:0]);
  AND2 I127 (gfint_3[1:1], choice_3, i_3r0[1:1]);
  AND2 I128 (gfint_3[2:2], choice_3, i_3r0[2:2]);
  AND2 I129 (gfint_3[3:3], choice_3, i_3r0[3:3]);
  AND2 I130 (gfint_3[4:4], choice_3, i_3r0[4:4]);
  AND2 I131 (gfint_3[5:5], choice_3, i_3r0[5:5]);
  AND2 I132 (gfint_3[6:6], choice_3, i_3r0[6:6]);
  AND2 I133 (gfint_4[0:0], choice_4, i_4r0[0:0]);
  AND2 I134 (gfint_4[1:1], choice_4, i_4r0[1:1]);
  AND2 I135 (gfint_4[2:2], choice_4, i_4r0[2:2]);
  AND2 I136 (gfint_4[3:3], choice_4, i_4r0[3:3]);
  AND2 I137 (gfint_4[4:4], choice_4, i_4r0[4:4]);
  AND2 I138 (gfint_4[5:5], choice_4, i_4r0[5:5]);
  AND2 I139 (gfint_4[6:6], choice_4, i_4r0[6:6]);
  AND2 I140 (gfint_5[0:0], choice_5, i_5r0[0:0]);
  AND2 I141 (gfint_5[1:1], choice_5, i_5r0[1:1]);
  AND2 I142 (gfint_5[2:2], choice_5, i_5r0[2:2]);
  AND2 I143 (gfint_5[3:3], choice_5, i_5r0[3:3]);
  AND2 I144 (gfint_5[4:4], choice_5, i_5r0[4:4]);
  AND2 I145 (gfint_5[5:5], choice_5, i_5r0[5:5]);
  AND2 I146 (gfint_5[6:6], choice_5, i_5r0[6:6]);
  AND2 I147 (gfint_6[0:0], choice_6, i_6r0[0:0]);
  AND2 I148 (gfint_6[1:1], choice_6, i_6r0[1:1]);
  AND2 I149 (gfint_6[2:2], choice_6, i_6r0[2:2]);
  AND2 I150 (gfint_6[3:3], choice_6, i_6r0[3:3]);
  AND2 I151 (gfint_6[4:4], choice_6, i_6r0[4:4]);
  AND2 I152 (gfint_6[5:5], choice_6, i_6r0[5:5]);
  AND2 I153 (gfint_6[6:6], choice_6, i_6r0[6:6]);
  OR2 I154 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I155 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I156 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I157 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I158 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I159 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I160 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  C3 I161 (simp1501_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I162 (simp1501_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  BUFF I163 (simp1501_0[2:2], comp0_0[6:6]);
  C3 I164 (icomp_0, simp1501_0[0:0], simp1501_0[1:1], simp1501_0[2:2]);
  OR2 I165 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I166 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I167 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I168 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I169 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I170 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I171 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  C3 I172 (simp1591_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I173 (simp1591_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  BUFF I174 (simp1591_0[2:2], comp1_0[6:6]);
  C3 I175 (icomp_1, simp1591_0[0:0], simp1591_0[1:1], simp1591_0[2:2]);
  OR2 I176 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I177 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I178 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2 I179 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  OR2 I180 (comp2_0[4:4], i_2r0[4:4], i_2r1[4:4]);
  OR2 I181 (comp2_0[5:5], i_2r0[5:5], i_2r1[5:5]);
  OR2 I182 (comp2_0[6:6], i_2r0[6:6], i_2r1[6:6]);
  C3 I183 (simp1681_0[0:0], comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C3 I184 (simp1681_0[1:1], comp2_0[3:3], comp2_0[4:4], comp2_0[5:5]);
  BUFF I185 (simp1681_0[2:2], comp2_0[6:6]);
  C3 I186 (icomp_2, simp1681_0[0:0], simp1681_0[1:1], simp1681_0[2:2]);
  OR2 I187 (comp3_0[0:0], i_3r0[0:0], i_3r1[0:0]);
  OR2 I188 (comp3_0[1:1], i_3r0[1:1], i_3r1[1:1]);
  OR2 I189 (comp3_0[2:2], i_3r0[2:2], i_3r1[2:2]);
  OR2 I190 (comp3_0[3:3], i_3r0[3:3], i_3r1[3:3]);
  OR2 I191 (comp3_0[4:4], i_3r0[4:4], i_3r1[4:4]);
  OR2 I192 (comp3_0[5:5], i_3r0[5:5], i_3r1[5:5]);
  OR2 I193 (comp3_0[6:6], i_3r0[6:6], i_3r1[6:6]);
  C3 I194 (simp1771_0[0:0], comp3_0[0:0], comp3_0[1:1], comp3_0[2:2]);
  C3 I195 (simp1771_0[1:1], comp3_0[3:3], comp3_0[4:4], comp3_0[5:5]);
  BUFF I196 (simp1771_0[2:2], comp3_0[6:6]);
  C3 I197 (icomp_3, simp1771_0[0:0], simp1771_0[1:1], simp1771_0[2:2]);
  OR2 I198 (comp4_0[0:0], i_4r0[0:0], i_4r1[0:0]);
  OR2 I199 (comp4_0[1:1], i_4r0[1:1], i_4r1[1:1]);
  OR2 I200 (comp4_0[2:2], i_4r0[2:2], i_4r1[2:2]);
  OR2 I201 (comp4_0[3:3], i_4r0[3:3], i_4r1[3:3]);
  OR2 I202 (comp4_0[4:4], i_4r0[4:4], i_4r1[4:4]);
  OR2 I203 (comp4_0[5:5], i_4r0[5:5], i_4r1[5:5]);
  OR2 I204 (comp4_0[6:6], i_4r0[6:6], i_4r1[6:6]);
  C3 I205 (simp1861_0[0:0], comp4_0[0:0], comp4_0[1:1], comp4_0[2:2]);
  C3 I206 (simp1861_0[1:1], comp4_0[3:3], comp4_0[4:4], comp4_0[5:5]);
  BUFF I207 (simp1861_0[2:2], comp4_0[6:6]);
  C3 I208 (icomp_4, simp1861_0[0:0], simp1861_0[1:1], simp1861_0[2:2]);
  OR2 I209 (comp5_0[0:0], i_5r0[0:0], i_5r1[0:0]);
  OR2 I210 (comp5_0[1:1], i_5r0[1:1], i_5r1[1:1]);
  OR2 I211 (comp5_0[2:2], i_5r0[2:2], i_5r1[2:2]);
  OR2 I212 (comp5_0[3:3], i_5r0[3:3], i_5r1[3:3]);
  OR2 I213 (comp5_0[4:4], i_5r0[4:4], i_5r1[4:4]);
  OR2 I214 (comp5_0[5:5], i_5r0[5:5], i_5r1[5:5]);
  OR2 I215 (comp5_0[6:6], i_5r0[6:6], i_5r1[6:6]);
  C3 I216 (simp1951_0[0:0], comp5_0[0:0], comp5_0[1:1], comp5_0[2:2]);
  C3 I217 (simp1951_0[1:1], comp5_0[3:3], comp5_0[4:4], comp5_0[5:5]);
  BUFF I218 (simp1951_0[2:2], comp5_0[6:6]);
  C3 I219 (icomp_5, simp1951_0[0:0], simp1951_0[1:1], simp1951_0[2:2]);
  OR2 I220 (comp6_0[0:0], i_6r0[0:0], i_6r1[0:0]);
  OR2 I221 (comp6_0[1:1], i_6r0[1:1], i_6r1[1:1]);
  OR2 I222 (comp6_0[2:2], i_6r0[2:2], i_6r1[2:2]);
  OR2 I223 (comp6_0[3:3], i_6r0[3:3], i_6r1[3:3]);
  OR2 I224 (comp6_0[4:4], i_6r0[4:4], i_6r1[4:4]);
  OR2 I225 (comp6_0[5:5], i_6r0[5:5], i_6r1[5:5]);
  OR2 I226 (comp6_0[6:6], i_6r0[6:6], i_6r1[6:6]);
  C3 I227 (simp2041_0[0:0], comp6_0[0:0], comp6_0[1:1], comp6_0[2:2]);
  C3 I228 (simp2041_0[1:1], comp6_0[3:3], comp6_0[4:4], comp6_0[5:5]);
  BUFF I229 (simp2041_0[2:2], comp6_0[6:6]);
  C3 I230 (icomp_6, simp2041_0[0:0], simp2041_0[1:1], simp2041_0[2:2]);
  C2R I231 (choice_0, icomp_0, nchosen_0, reset);
  C2R I232 (choice_1, icomp_1, nchosen_0, reset);
  C2R I233 (choice_2, icomp_2, nchosen_0, reset);
  C2R I234 (choice_3, icomp_3, nchosen_0, reset);
  C2R I235 (choice_4, icomp_4, nchosen_0, reset);
  C2R I236 (choice_5, icomp_5, nchosen_0, reset);
  C2R I237 (choice_6, icomp_6, nchosen_0, reset);
  NOR3 I238 (simp2121_0[0:0], choice_0, choice_1, choice_2);
  NOR3 I239 (simp2121_0[1:1], choice_3, choice_4, choice_5);
  INV I240 (simp2121_0[2:2], choice_6);
  NAND3 I241 (anychoice_0, simp2121_0[0:0], simp2121_0[1:1], simp2121_0[2:2]);
  NOR2 I242 (nchosen_0, anychoice_0, o_0a);
  C2R I243 (i_0a, choice_0, o_0a, reset);
  C2R I244 (i_1a, choice_1, o_0a, reset);
  C2R I245 (i_2a, choice_2, o_0a, reset);
  C2R I246 (i_3a, choice_3, o_0a, reset);
  C2R I247 (i_4a, choice_4, o_0a, reset);
  C2R I248 (i_5a, choice_5, o_0a, reset);
  C2R I249 (i_6a, choice_6, o_0a, reset);
endmodule

// tkj7m0_7 TeakJ [Many [0,7],One 7]
module tkj7m0_7 (i_0r, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input i_0r;
  output i_0a;
  input [6:0] i_1r0;
  input [6:0] i_1r1;
  output i_1a;
  output [6:0] o_0r0;
  output [6:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [6:0] joinf_0;
  wire [6:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_1r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_1r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_1r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_1r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_1r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_1r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_1r0[6:6]);
  BUFF I7 (joint_0[0:0], i_1r1[0:0]);
  BUFF I8 (joint_0[1:1], i_1r1[1:1]);
  BUFF I9 (joint_0[2:2], i_1r1[2:2]);
  BUFF I10 (joint_0[3:3], i_1r1[3:3]);
  BUFF I11 (joint_0[4:4], i_1r1[4:4]);
  BUFF I12 (joint_0[5:5], i_1r1[5:5]);
  BUFF I13 (joint_0[6:6], i_1r1[6:6]);
  BUFF I14 (icomplete_0, i_0r);
  C2 I15 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I16 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I17 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I18 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I19 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I20 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I21 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I22 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I23 (o_0r1[1:1], joint_0[1:1]);
  BUFF I24 (o_0r1[2:2], joint_0[2:2]);
  BUFF I25 (o_0r1[3:3], joint_0[3:3]);
  BUFF I26 (o_0r1[4:4], joint_0[4:4]);
  BUFF I27 (o_0r1[5:5], joint_0[5:5]);
  BUFF I28 (o_0r1[6:6], joint_0[6:6]);
  BUFF I29 (i_0a, o_0a);
  BUFF I30 (i_1a, o_0a);
endmodule

// tks7_o0w7_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0_20o0w0_40o0w0 TeakS (0+:7) [([Imp 1 0],0),([Imp 2 0],0),([I
//   mp 4 0],0),([Imp 8 0],0),([Imp 16 0],0),([Imp 32 0],0),([Imp 64 0],0)] [One 7,Many [0,0,0,0,0,0,0]]
module tks7_o0w7_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0_20o0w0_40o0w0 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, o_5r, o_5a, o_6r, o_6a, reset);
  input [6:0] i_0r0;
  input [6:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire sel_3;
  wire sel_4;
  wire sel_5;
  wire sel_6;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire gsel_3;
  wire gsel_4;
  wire gsel_5;
  wire gsel_6;
  wire oack_0;
  wire match0_0;
  wire [2:0] simp181_0;
  wire match1_0;
  wire [2:0] simp211_0;
  wire match2_0;
  wire [2:0] simp241_0;
  wire match3_0;
  wire [2:0] simp271_0;
  wire match4_0;
  wire [2:0] simp301_0;
  wire match5_0;
  wire [2:0] simp331_0;
  wire match6_0;
  wire [2:0] simp361_0;
  wire [6:0] comp_0;
  wire [2:0] simp521_0;
  wire [2:0] simp601_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (simp181_0[0:0], i_0r1[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I2 (simp181_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  BUFF I3 (simp181_0[2:2], i_0r0[6:6]);
  C3 I4 (match0_0, simp181_0[0:0], simp181_0[1:1], simp181_0[2:2]);
  BUFF I5 (sel_1, match1_0);
  C3 I6 (simp211_0[0:0], i_0r0[0:0], i_0r1[1:1], i_0r0[2:2]);
  C3 I7 (simp211_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  BUFF I8 (simp211_0[2:2], i_0r0[6:6]);
  C3 I9 (match1_0, simp211_0[0:0], simp211_0[1:1], simp211_0[2:2]);
  BUFF I10 (sel_2, match2_0);
  C3 I11 (simp241_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r1[2:2]);
  C3 I12 (simp241_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  BUFF I13 (simp241_0[2:2], i_0r0[6:6]);
  C3 I14 (match2_0, simp241_0[0:0], simp241_0[1:1], simp241_0[2:2]);
  BUFF I15 (sel_3, match3_0);
  C3 I16 (simp271_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I17 (simp271_0[1:1], i_0r1[3:3], i_0r0[4:4], i_0r0[5:5]);
  BUFF I18 (simp271_0[2:2], i_0r0[6:6]);
  C3 I19 (match3_0, simp271_0[0:0], simp271_0[1:1], simp271_0[2:2]);
  BUFF I20 (sel_4, match4_0);
  C3 I21 (simp301_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I22 (simp301_0[1:1], i_0r0[3:3], i_0r1[4:4], i_0r0[5:5]);
  BUFF I23 (simp301_0[2:2], i_0r0[6:6]);
  C3 I24 (match4_0, simp301_0[0:0], simp301_0[1:1], simp301_0[2:2]);
  BUFF I25 (sel_5, match5_0);
  C3 I26 (simp331_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I27 (simp331_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r1[5:5]);
  BUFF I28 (simp331_0[2:2], i_0r0[6:6]);
  C3 I29 (match5_0, simp331_0[0:0], simp331_0[1:1], simp331_0[2:2]);
  BUFF I30 (sel_6, match6_0);
  C3 I31 (simp361_0[0:0], i_0r0[0:0], i_0r0[1:1], i_0r0[2:2]);
  C3 I32 (simp361_0[1:1], i_0r0[3:3], i_0r0[4:4], i_0r0[5:5]);
  BUFF I33 (simp361_0[2:2], i_0r1[6:6]);
  C3 I34 (match6_0, simp361_0[0:0], simp361_0[1:1], simp361_0[2:2]);
  C2 I35 (gsel_0, sel_0, icomplete_0);
  C2 I36 (gsel_1, sel_1, icomplete_0);
  C2 I37 (gsel_2, sel_2, icomplete_0);
  C2 I38 (gsel_3, sel_3, icomplete_0);
  C2 I39 (gsel_4, sel_4, icomplete_0);
  C2 I40 (gsel_5, sel_5, icomplete_0);
  C2 I41 (gsel_6, sel_6, icomplete_0);
  OR2 I42 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I43 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I44 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I45 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I46 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I47 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I48 (comp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  C3 I49 (simp521_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I50 (simp521_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  BUFF I51 (simp521_0[2:2], comp_0[6:6]);
  C3 I52 (icomplete_0, simp521_0[0:0], simp521_0[1:1], simp521_0[2:2]);
  BUFF I53 (o_0r, gsel_0);
  BUFF I54 (o_1r, gsel_1);
  BUFF I55 (o_2r, gsel_2);
  BUFF I56 (o_3r, gsel_3);
  BUFF I57 (o_4r, gsel_4);
  BUFF I58 (o_5r, gsel_5);
  BUFF I59 (o_6r, gsel_6);
  NOR3 I60 (simp601_0[0:0], o_0a, o_1a, o_2a);
  NOR3 I61 (simp601_0[1:1], o_3a, o_4a, o_5a);
  INV I62 (simp601_0[2:2], o_6a);
  NAND3 I63 (oack_0, simp601_0[0:0], simp601_0[1:1], simp601_0[2:2]);
  C2 I64 (i_0a, oack_0, icomplete_0);
endmodule

// tkvr132_wo0w32_ro0w32 TeakV "r1" 32 [] [0] [0] [Many [32],Many [0],Many [0],Many [32]]
module tkvr132_wo0w32_ro0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I457 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I458 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I459 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I460 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I461 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I462 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I463 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I464 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I465 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I466 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I467 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I468 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I469 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I470 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I471 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I472 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I473 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I474 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I475 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I476 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I477 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I478 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I479 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I480 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I481 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I482 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I483 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I484 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I485 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I486 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I487 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  OR2 I488 (anyread_0, rg_0r, rg_0a);
  BUFF I489 (wg_0a, wd_0a);
  BUFF I490 (rg_0a, rd_0a);
endmodule

// tkvr032_wo0w32_ro0w32 TeakV "r0" 32 [] [0] [0] [Many [32],Many [0],Many [0],Many [32]]
module tkvr032_wo0w32_ro0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I457 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I458 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I459 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I460 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I461 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I462 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I463 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I464 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I465 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I466 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I467 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I468 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I469 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I470 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I471 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I472 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I473 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I474 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I475 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I476 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I477 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I478 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I479 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I480 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I481 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I482 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I483 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I484 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I485 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I486 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I487 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  OR2 I488 (anyread_0, rg_0r, rg_0a);
  BUFF I489 (wg_0a, wd_0a);
  BUFF I490 (rg_0a, rd_0a);
endmodule

// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 TeakF [0,0,0,0,0,0,0] [One 0,Many [0,0,0,0,0,0,0]]
module tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 (i_0r, i_0a, o_0r, o_0a, o_1r, o_1a, o_2r, o_2a, o_3r, o_3a, o_4r, o_4a, o_5r, o_5a, o_6r, o_6a, reset);
  input i_0r;
  output i_0a;
  output o_0r;
  input o_0a;
  output o_1r;
  input o_1a;
  output o_2r;
  input o_2a;
  output o_3r;
  input o_3a;
  output o_4r;
  input o_4a;
  output o_5r;
  input o_5a;
  output o_6r;
  input o_6a;
  input reset;
  wire [2:0] simp11_0;
  BUFF I0 (o_0r, i_0r);
  BUFF I1 (o_1r, i_0r);
  BUFF I2 (o_2r, i_0r);
  BUFF I3 (o_3r, i_0r);
  BUFF I4 (o_4r, i_0r);
  BUFF I5 (o_5r, i_0r);
  BUFF I6 (o_6r, i_0r);
  C3 I7 (simp11_0[0:0], o_0a, o_1a, o_2a);
  C3 I8 (simp11_0[1:1], o_3a, o_4a, o_5a);
  BUFF I9 (simp11_0[2:2], o_6a);
  C3 I10 (i_0a, simp11_0[0:0], simp11_0[1:1], simp11_0[2:2]);
endmodule

// tkj0m0_0_0_0_0_0_0 TeakJ [Many [0,0,0,0,0,0,0],One 0]
module tkj0m0_0_0_0_0_0_0 (i_0r, i_0a, i_1r, i_1a, i_2r, i_2a, i_3r, i_3a, i_4r, i_4a, i_5r, i_5a, i_6r, i_6a, o_0r, o_0a, reset);
  input i_0r;
  output i_0a;
  input i_1r;
  output i_1a;
  input i_2r;
  output i_2a;
  input i_3r;
  output i_3a;
  input i_4r;
  output i_4a;
  input i_5r;
  output i_5a;
  input i_6r;
  output i_6a;
  output o_0r;
  input o_0a;
  input reset;
  wire [2:0] simp01_0;
  C3 I0 (simp01_0[0:0], i_0r, i_1r, i_2r);
  C3 I1 (simp01_0[1:1], i_3r, i_4r, i_5r);
  BUFF I2 (simp01_0[2:2], i_6r);
  C3 I3 (o_0r, simp01_0[0:0], simp01_0[1:1], simp01_0[2:2]);
  BUFF I4 (i_0a, o_0a);
  BUFF I5 (i_1a, o_0a);
  BUFF I6 (i_2a, o_0a);
  BUFF I7 (i_3a, o_0a);
  BUFF I8 (i_4a, o_0a);
  BUFF I9 (i_5a, o_0a);
  BUFF I10 (i_6a, o_0a);
endmodule

// tkvtakeBranch21_wo0w1_ro0w1 TeakV "takeBranch2" 1 [] [0] [0] [Many [1],Many [0],Many [0],Many [1]]
module tkvtakeBranch21_wo0w1_ro0w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input wg_0r0;
  input wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  input reset;
  wire wf_0;
  wire wt_0;
  wire df_0;
  wire dt_0;
  wire wc_0;
  wire wacks_0;
  wire wenr_0;
  wire wen_0;
  wire anyread_0;
  wire nreset_0;
  wire drlgf_0;
  wire drlgt_0;
  wire comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire conwgit_0;
  wire conwgif_0;
  wire conwig_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0, wenr_0, nreset_0);
  AND2 I2 (drlgf_0, wf_0, wen_0);
  AND2 I3 (drlgt_0, wt_0, wen_0);
  NOR2 I4 (df_0, dt_0, drlgt_0);
  NOR3 I5 (dt_0, df_0, drlgf_0, reset);
  AO22 I6 (wacks_0, drlgf_0, df_0, drlgt_0, dt_0);
  OR2 I7 (comp0_0, wg_0r0, wg_0r1);
  BUFF I8 (wc_0, comp0_0);
  AND2 I9 (conwgif_0, wg_0r0, conwig_0);
  AND2 I10 (conwgit_0, wg_0r1, conwig_0);
  BUFF I11 (conwigc_0, wc_0);
  AO22 I12 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I13 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I14 (wf_0, conwgif_0);
  BUFF I15 (wt_0, conwgit_0);
  BUFF I16 (wenr_0, wc_0);
  C2 I17 (wd_0r, conwig_0, wacks_0);
  AND2 I18 (rd_0r0, df_0, rg_0r);
  AND2 I19 (rd_0r1, dt_0, rg_0r);
  OR2 I20 (anyread_0, rg_0r, rg_0a);
  BUFF I21 (wg_0a, wd_0a);
  BUFF I22 (rg_0a, rd_0a);
endmodule

// tkvtakeBranch1_wo0w1_ro0w1o0w1 TeakV "takeBranch" 1 [] [0] [0,0] [Many [1],Many [0],Many [0,0],Many 
//   [1,1]]
module tkvtakeBranch1_wo0w1_ro0w1o0w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, reset);
  input wg_0r0;
  input wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  output rd_1r0;
  output rd_1r1;
  input rd_1a;
  input reset;
  wire wf_0;
  wire wt_0;
  wire df_0;
  wire dt_0;
  wire wc_0;
  wire wacks_0;
  wire wenr_0;
  wire wen_0;
  wire anyread_0;
  wire nreset_0;
  wire drlgf_0;
  wire drlgt_0;
  wire comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire conwgit_0;
  wire conwgif_0;
  wire conwig_0;
  wire [1:0] simp401_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0, wenr_0, nreset_0);
  AND2 I2 (drlgf_0, wf_0, wen_0);
  AND2 I3 (drlgt_0, wt_0, wen_0);
  NOR2 I4 (df_0, dt_0, drlgt_0);
  NOR3 I5 (dt_0, df_0, drlgf_0, reset);
  AO22 I6 (wacks_0, drlgf_0, df_0, drlgt_0, dt_0);
  OR2 I7 (comp0_0, wg_0r0, wg_0r1);
  BUFF I8 (wc_0, comp0_0);
  AND2 I9 (conwgif_0, wg_0r0, conwig_0);
  AND2 I10 (conwgit_0, wg_0r1, conwig_0);
  BUFF I11 (conwigc_0, wc_0);
  AO22 I12 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I13 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I14 (wf_0, conwgif_0);
  BUFF I15 (wt_0, conwgit_0);
  BUFF I16 (wenr_0, wc_0);
  C2 I17 (wd_0r, conwig_0, wacks_0);
  AND2 I18 (rd_0r0, df_0, rg_0r);
  AND2 I19 (rd_1r0, df_0, rg_1r);
  AND2 I20 (rd_0r1, dt_0, rg_0r);
  AND2 I21 (rd_1r1, dt_0, rg_1r);
  NOR3 I22 (simp401_0[0:0], rg_0r, rg_1r, rg_0a);
  INV I23 (simp401_0[1:1], rg_1a);
  NAND2 I24 (anyread_0, simp401_0[0:0], simp401_0[1:1]);
  BUFF I25 (wg_0a, wd_0a);
  BUFF I26 (rg_0a, rd_0a);
  BUFF I27 (rg_1a, rd_1a);
endmodule

// tkvcwp1_wo0w1_ro0w1 TeakV "cwp" 1 [] [0] [0] [Many [1],Many [0],Many [0],Many [1]]
module tkvcwp1_wo0w1_ro0w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input wg_0r0;
  input wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  input reset;
  wire wf_0;
  wire wt_0;
  wire df_0;
  wire dt_0;
  wire wc_0;
  wire wacks_0;
  wire wenr_0;
  wire wen_0;
  wire anyread_0;
  wire nreset_0;
  wire drlgf_0;
  wire drlgt_0;
  wire comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire conwgit_0;
  wire conwgif_0;
  wire conwig_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0, wenr_0, nreset_0);
  AND2 I2 (drlgf_0, wf_0, wen_0);
  AND2 I3 (drlgt_0, wt_0, wen_0);
  NOR2 I4 (df_0, dt_0, drlgt_0);
  NOR3 I5 (dt_0, df_0, drlgf_0, reset);
  AO22 I6 (wacks_0, drlgf_0, df_0, drlgt_0, dt_0);
  OR2 I7 (comp0_0, wg_0r0, wg_0r1);
  BUFF I8 (wc_0, comp0_0);
  AND2 I9 (conwgif_0, wg_0r0, conwig_0);
  AND2 I10 (conwgit_0, wg_0r1, conwig_0);
  BUFF I11 (conwigc_0, wc_0);
  AO22 I12 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I13 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I14 (wf_0, conwgif_0);
  BUFF I15 (wt_0, conwgit_0);
  BUFF I16 (wenr_0, wc_0);
  C2 I17 (wd_0r, conwig_0, wacks_0);
  AND2 I18 (rd_0r0, df_0, rg_0r);
  AND2 I19 (rd_0r1, dt_0, rg_0r);
  OR2 I20 (anyread_0, rg_0r, rg_0a);
  BUFF I21 (wg_0a, wd_0a);
  BUFF I22 (rg_0a, rd_0a);
endmodule

// tkvpreCarry1_wo0w1_ro0w1o0w1o0w1 TeakV "preCarry" 1 [] [0] [0,0,0] [Many [1],Many [0],Many [0,0,0],M
//   any [1,1,1]]
module tkvpreCarry1_wo0w1_ro0w1o0w1o0w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, reset);
  input wg_0r0;
  input wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  output rd_1r0;
  output rd_1r1;
  input rd_1a;
  output rd_2r0;
  output rd_2r1;
  input rd_2a;
  input reset;
  wire wf_0;
  wire wt_0;
  wire df_0;
  wire dt_0;
  wire wc_0;
  wire wacks_0;
  wire wenr_0;
  wire wen_0;
  wire anyread_0;
  wire nreset_0;
  wire drlgf_0;
  wire drlgt_0;
  wire comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire conwgit_0;
  wire conwgif_0;
  wire conwig_0;
  wire [1:0] simp421_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0, wenr_0, nreset_0);
  AND2 I2 (drlgf_0, wf_0, wen_0);
  AND2 I3 (drlgt_0, wt_0, wen_0);
  NOR2 I4 (df_0, dt_0, drlgt_0);
  NOR3 I5 (dt_0, df_0, drlgf_0, reset);
  AO22 I6 (wacks_0, drlgf_0, df_0, drlgt_0, dt_0);
  OR2 I7 (comp0_0, wg_0r0, wg_0r1);
  BUFF I8 (wc_0, comp0_0);
  AND2 I9 (conwgif_0, wg_0r0, conwig_0);
  AND2 I10 (conwgit_0, wg_0r1, conwig_0);
  BUFF I11 (conwigc_0, wc_0);
  AO22 I12 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I13 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I14 (wf_0, conwgif_0);
  BUFF I15 (wt_0, conwgit_0);
  BUFF I16 (wenr_0, wc_0);
  C2 I17 (wd_0r, conwig_0, wacks_0);
  AND2 I18 (rd_0r0, df_0, rg_0r);
  AND2 I19 (rd_1r0, df_0, rg_1r);
  AND2 I20 (rd_2r0, df_0, rg_2r);
  AND2 I21 (rd_0r1, dt_0, rg_0r);
  AND2 I22 (rd_1r1, dt_0, rg_1r);
  AND2 I23 (rd_2r1, dt_0, rg_2r);
  NOR3 I24 (simp421_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I25 (simp421_0[1:1], rg_0a, rg_1a, rg_2a);
  NAND2 I26 (anyread_0, simp421_0[0:0], simp421_0[1:1]);
  BUFF I27 (wg_0a, wd_0a);
  BUFF I28 (rg_0a, rd_0a);
  BUFF I29 (rg_1a, rd_1a);
  BUFF I30 (rg_2a, rd_2a);
endmodule

// tkm2x4b TeakM [Many [4,4],One 4]
module tkm2x4b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  input [3:0] i_1r0;
  input [3:0] i_1r1;
  output i_1a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  input reset;
  wire [3:0] gfint_0;
  wire [3:0] gfint_1;
  wire [3:0] gtint_0;
  wire [3:0] gtint_1;
  wire choice_0;
  wire choice_1;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire nchosen_0;
  wire [3:0] comp0_0;
  wire [1:0] simp391_0;
  wire [3:0] comp1_0;
  wire [1:0] simp451_0;
  OR2 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0]);
  OR2 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1]);
  OR2 I2 (o_0r0[2:2], gfint_0[2:2], gfint_1[2:2]);
  OR2 I3 (o_0r0[3:3], gfint_0[3:3], gfint_1[3:3]);
  OR2 I4 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0]);
  OR2 I5 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1]);
  OR2 I6 (o_0r1[2:2], gtint_0[2:2], gtint_1[2:2]);
  OR2 I7 (o_0r1[3:3], gtint_0[3:3], gtint_1[3:3]);
  AND2 I8 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I9 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I10 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I11 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I12 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I13 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I14 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I15 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I16 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I17 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I18 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I19 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I20 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I21 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I22 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I23 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  OR2 I24 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I25 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I26 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I27 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  C3 I28 (simp391_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  BUFF I29 (simp391_0[1:1], comp0_0[3:3]);
  C2 I30 (icomp_0, simp391_0[0:0], simp391_0[1:1]);
  OR2 I31 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I32 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I33 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I34 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  C3 I35 (simp451_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  BUFF I36 (simp451_0[1:1], comp1_0[3:3]);
  C2 I37 (icomp_1, simp451_0[0:0], simp451_0[1:1]);
  C2R I38 (choice_0, icomp_0, nchosen_0, reset);
  C2R I39 (choice_1, icomp_1, nchosen_0, reset);
  OR2 I40 (anychoice_0, choice_0, choice_1);
  NOR2 I41 (nchosen_0, anychoice_0, o_0a);
  C2R I42 (i_0a, choice_0, o_0a, reset);
  C2R I43 (i_1a, choice_1, o_0a, reset);
endmodule

// tkvflags4_wo0w4_ro2w1o1w1o3w1o0w1o3w1o2w1o1w1o2w1o1w1o0w1o0w1o3w1 TeakV "flags" 4 [] [0] [2,1,3,0,3,
//   2,1,2,1,0,0,3] [Many [4],Many [0],Many [0,0,0,0,0,0,0,0,0,0,0,0],Many [1,1,1,1,1,1,1,1,1,1,1,1]]
module tkvflags4_wo0w4_ro2w1o1w1o3w1o0w1o3w1o2w1o1w1o2w1o1w1o0w1o0w1o3w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rg_5r, rg_5a, rg_6r, rg_6a, rg_7r, rg_7a, rg_8r, rg_8a, rg_9r, rg_9a, rg_10r, rg_10a, rg_11r, rg_11a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, rd_5r0, rd_5r1, rd_5a, rd_6r0, rd_6r1, rd_6a, rd_7r0, rd_7r1, rd_7a, rd_8r0, rd_8r1, rd_8a, rd_9r0, rd_9r1, rd_9a, rd_10r0, rd_10r1, rd_10a, rd_11r0, rd_11r1, rd_11a, reset);
  input [3:0] wg_0r0;
  input [3:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  input rg_5r;
  output rg_5a;
  input rg_6r;
  output rg_6a;
  input rg_7r;
  output rg_7a;
  input rg_8r;
  output rg_8a;
  input rg_9r;
  output rg_9a;
  input rg_10r;
  output rg_10a;
  input rg_11r;
  output rg_11a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  output rd_1r0;
  output rd_1r1;
  input rd_1a;
  output rd_2r0;
  output rd_2r1;
  input rd_2a;
  output rd_3r0;
  output rd_3r1;
  input rd_3a;
  output rd_4r0;
  output rd_4r1;
  input rd_4a;
  output rd_5r0;
  output rd_5r1;
  input rd_5a;
  output rd_6r0;
  output rd_6r1;
  input rd_6a;
  output rd_7r0;
  output rd_7r1;
  input rd_7a;
  output rd_8r0;
  output rd_8r1;
  input rd_8a;
  output rd_9r0;
  output rd_9r1;
  input rd_9a;
  output rd_10r0;
  output rd_10r1;
  input rd_10a;
  output rd_11r0;
  output rd_11r1;
  input rd_11a;
  input reset;
  wire [3:0] wf_0;
  wire [3:0] wt_0;
  wire [3:0] df_0;
  wire [3:0] dt_0;
  wire wc_0;
  wire [3:0] wacks_0;
  wire [3:0] wenr_0;
  wire [3:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [3:0] drlgf_0;
  wire [3:0] drlgt_0;
  wire [3:0] comp0_0;
  wire [1:0] simp421_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [3:0] conwgit_0;
  wire [3:0] conwgif_0;
  wire conwig_0;
  wire [1:0] simp711_0;
  wire [7:0] simp961_0;
  wire [2:0] simp962_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I6 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I7 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I8 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I9 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I10 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I11 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I12 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  NOR2 I13 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I14 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I15 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I16 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR3 I17 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I18 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I19 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I20 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  AO22 I21 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I22 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I23 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I24 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  OR2 I25 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I26 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I27 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I28 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  C3 I29 (simp421_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  BUFF I30 (simp421_0[1:1], comp0_0[3:3]);
  C2 I31 (wc_0, simp421_0[0:0], simp421_0[1:1]);
  AND2 I32 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I33 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I34 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I35 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I36 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I37 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I38 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I39 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  BUFF I40 (conwigc_0, wc_0);
  AO22 I41 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I42 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I43 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I44 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I45 (wenr_0[0:0], wc_0);
  BUFF I46 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I47 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I48 (wenr_0[1:1], wc_0);
  BUFF I49 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I50 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I51 (wenr_0[2:2], wc_0);
  BUFF I52 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I53 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I54 (wenr_0[3:3], wc_0);
  C3 I55 (simp711_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C2 I56 (simp711_0[1:1], wacks_0[2:2], wacks_0[3:3]);
  C2 I57 (wd_0r, simp711_0[0:0], simp711_0[1:1]);
  AND2 I58 (rd_0r0, df_0[2:2], rg_0r);
  AND2 I59 (rd_1r0, df_0[1:1], rg_1r);
  AND2 I60 (rd_2r0, df_0[3:3], rg_2r);
  AND2 I61 (rd_3r0, df_0[0:0], rg_3r);
  AND2 I62 (rd_4r0, df_0[3:3], rg_4r);
  AND2 I63 (rd_5r0, df_0[2:2], rg_5r);
  AND2 I64 (rd_6r0, df_0[1:1], rg_6r);
  AND2 I65 (rd_7r0, df_0[2:2], rg_7r);
  AND2 I66 (rd_8r0, df_0[1:1], rg_8r);
  AND2 I67 (rd_9r0, df_0[0:0], rg_9r);
  AND2 I68 (rd_10r0, df_0[0:0], rg_10r);
  AND2 I69 (rd_11r0, df_0[3:3], rg_11r);
  AND2 I70 (rd_0r1, dt_0[2:2], rg_0r);
  AND2 I71 (rd_1r1, dt_0[1:1], rg_1r);
  AND2 I72 (rd_2r1, dt_0[3:3], rg_2r);
  AND2 I73 (rd_3r1, dt_0[0:0], rg_3r);
  AND2 I74 (rd_4r1, dt_0[3:3], rg_4r);
  AND2 I75 (rd_5r1, dt_0[2:2], rg_5r);
  AND2 I76 (rd_6r1, dt_0[1:1], rg_6r);
  AND2 I77 (rd_7r1, dt_0[2:2], rg_7r);
  AND2 I78 (rd_8r1, dt_0[1:1], rg_8r);
  AND2 I79 (rd_9r1, dt_0[0:0], rg_9r);
  AND2 I80 (rd_10r1, dt_0[0:0], rg_10r);
  AND2 I81 (rd_11r1, dt_0[3:3], rg_11r);
  NOR3 I82 (simp961_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I83 (simp961_0[1:1], rg_3r, rg_4r, rg_5r);
  NOR3 I84 (simp961_0[2:2], rg_6r, rg_7r, rg_8r);
  NOR3 I85 (simp961_0[3:3], rg_9r, rg_10r, rg_11r);
  NOR3 I86 (simp961_0[4:4], rg_0a, rg_1a, rg_2a);
  NOR3 I87 (simp961_0[5:5], rg_3a, rg_4a, rg_5a);
  NOR3 I88 (simp961_0[6:6], rg_6a, rg_7a, rg_8a);
  NOR3 I89 (simp961_0[7:7], rg_9a, rg_10a, rg_11a);
  NAND3 I90 (simp962_0[0:0], simp961_0[0:0], simp961_0[1:1], simp961_0[2:2]);
  NAND3 I91 (simp962_0[1:1], simp961_0[3:3], simp961_0[4:4], simp961_0[5:5]);
  NAND2 I92 (simp962_0[2:2], simp961_0[6:6], simp961_0[7:7]);
  OR3 I93 (anyread_0, simp962_0[0:0], simp962_0[1:1], simp962_0[2:2]);
  BUFF I94 (wg_0a, wd_0a);
  BUFF I95 (rg_0a, rd_0a);
  BUFF I96 (rg_1a, rd_1a);
  BUFF I97 (rg_2a, rd_2a);
  BUFF I98 (rg_3a, rd_3a);
  BUFF I99 (rg_4a, rd_4a);
  BUFF I100 (rg_5a, rd_5a);
  BUFF I101 (rg_6a, rd_6a);
  BUFF I102 (rg_7a, rd_7a);
  BUFF I103 (rg_8a, rd_8a);
  BUFF I104 (rg_9a, rd_9a);
  BUFF I105 (rg_10a, rd_10a);
  BUFF I106 (rg_11a, rd_11a);
endmodule

// tkvpcr33_wo0w33_ro0w32o32w1 TeakV "pcr" 33 [] [0] [0,32] [Many [33],Many [0],Many [0,0],Many [32,1]]
module tkvpcr33_wo0w33_ro0w32o32w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, reset);
  input [32:0] wg_0r0;
  input [32:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  output rd_1r0;
  output rd_1r1;
  input rd_1a;
  input reset;
  wire [32:0] wf_0;
  wire [32:0] wt_0;
  wire [32:0] df_0;
  wire [32:0] dt_0;
  wire wc_0;
  wire [32:0] wacks_0;
  wire [32:0] wenr_0;
  wire [32:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [32:0] drlgf_0;
  wire [32:0] drlgt_0;
  wire [32:0] comp0_0;
  wire [10:0] simp2451_0;
  wire [3:0] simp2452_0;
  wire [1:0] simp2453_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [32:0] conwgit_0;
  wire [32:0] conwgif_0;
  wire conwig_0;
  wire [11:0] simp4191_0;
  wire [3:0] simp4192_0;
  wire [1:0] simp4193_0;
  wire [1:0] simp4861_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (wen_0[32:32], wenr_0[32:32], nreset_0);
  AND2 I34 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I35 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I36 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I37 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I38 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I39 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I40 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I41 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I42 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I43 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I44 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I45 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I46 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I47 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I48 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I49 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I50 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I51 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I52 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I53 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I54 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I55 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I56 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I57 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I58 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I59 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I60 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I61 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I62 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I63 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I64 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I65 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I66 (drlgf_0[32:32], wf_0[32:32], wen_0[32:32]);
  AND2 I67 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I68 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I69 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I70 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I71 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I72 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I73 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I74 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I75 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I76 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I77 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I78 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I79 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I80 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I81 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I82 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I83 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I84 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I85 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I86 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I87 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I88 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I89 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I90 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I91 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I92 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I93 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I94 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I95 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I96 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I97 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I98 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  AND2 I99 (drlgt_0[32:32], wt_0[32:32], wen_0[32:32]);
  NOR2 I100 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I101 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I102 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I103 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I104 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I105 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I106 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I107 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I108 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I109 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I110 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I111 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I112 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I113 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I114 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I115 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I116 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I117 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I118 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I119 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I120 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I121 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I122 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I123 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I124 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I125 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I126 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I127 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I128 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I129 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I130 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I131 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR2 I132 (df_0[32:32], dt_0[32:32], drlgt_0[32:32]);
  NOR3 I133 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I134 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I135 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I136 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I137 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I138 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I139 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I140 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I141 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I142 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I143 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I144 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I145 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I146 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I147 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I148 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I149 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I150 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I151 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I152 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I153 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I154 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I155 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I156 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I157 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I158 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I159 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I160 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I161 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I162 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I163 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I164 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  NOR3 I165 (dt_0[32:32], df_0[32:32], drlgf_0[32:32], reset);
  AO22 I166 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I167 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I168 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I169 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I170 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I171 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I172 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I173 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I174 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I175 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I176 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I177 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I178 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I179 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I180 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I181 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I182 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I183 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I184 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I185 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I186 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I187 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I188 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I189 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I190 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I191 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I192 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I193 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I194 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I195 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I196 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I197 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  AO22 I198 (wacks_0[32:32], drlgf_0[32:32], df_0[32:32], drlgt_0[32:32], dt_0[32:32]);
  OR2 I199 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I200 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I201 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I202 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I203 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I204 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I205 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I206 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I207 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I208 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I209 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I210 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I211 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I212 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I213 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I214 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I215 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I216 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I217 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I218 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I219 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I220 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I221 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I222 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I223 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I224 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I225 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I226 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I227 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I228 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I229 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I230 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  OR2 I231 (comp0_0[32:32], wg_0r0[32:32], wg_0r1[32:32]);
  C3 I232 (simp2451_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I233 (simp2451_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I234 (simp2451_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I235 (simp2451_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I236 (simp2451_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I237 (simp2451_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I238 (simp2451_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I239 (simp2451_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I240 (simp2451_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I241 (simp2451_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C3 I242 (simp2451_0[10:10], comp0_0[30:30], comp0_0[31:31], comp0_0[32:32]);
  C3 I243 (simp2452_0[0:0], simp2451_0[0:0], simp2451_0[1:1], simp2451_0[2:2]);
  C3 I244 (simp2452_0[1:1], simp2451_0[3:3], simp2451_0[4:4], simp2451_0[5:5]);
  C3 I245 (simp2452_0[2:2], simp2451_0[6:6], simp2451_0[7:7], simp2451_0[8:8]);
  C2 I246 (simp2452_0[3:3], simp2451_0[9:9], simp2451_0[10:10]);
  C3 I247 (simp2453_0[0:0], simp2452_0[0:0], simp2452_0[1:1], simp2452_0[2:2]);
  BUFF I248 (simp2453_0[1:1], simp2452_0[3:3]);
  C2 I249 (wc_0, simp2453_0[0:0], simp2453_0[1:1]);
  AND2 I250 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I251 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I252 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I253 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I254 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I255 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I256 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I257 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I258 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I259 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I260 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I261 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I262 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I263 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I264 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I265 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I266 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I267 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I268 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I269 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I270 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I271 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I272 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I273 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I274 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I275 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I276 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I277 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I278 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I279 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I280 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I281 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I282 (conwgif_0[32:32], wg_0r0[32:32], conwig_0);
  AND2 I283 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I284 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I285 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I286 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I287 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I288 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I289 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I290 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I291 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I292 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I293 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I294 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I295 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I296 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I297 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I298 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I299 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I300 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I301 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I302 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I303 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I304 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I305 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I306 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I307 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I308 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I309 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I310 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I311 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I312 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I313 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I314 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  AND2 I315 (conwgit_0[32:32], wg_0r1[32:32], conwig_0);
  BUFF I316 (conwigc_0, wc_0);
  AO22 I317 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I318 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I319 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I320 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I321 (wenr_0[0:0], wc_0);
  BUFF I322 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I323 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I324 (wenr_0[1:1], wc_0);
  BUFF I325 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I326 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I327 (wenr_0[2:2], wc_0);
  BUFF I328 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I329 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I330 (wenr_0[3:3], wc_0);
  BUFF I331 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I332 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I333 (wenr_0[4:4], wc_0);
  BUFF I334 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I335 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I336 (wenr_0[5:5], wc_0);
  BUFF I337 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I338 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I339 (wenr_0[6:6], wc_0);
  BUFF I340 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I341 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I342 (wenr_0[7:7], wc_0);
  BUFF I343 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I344 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I345 (wenr_0[8:8], wc_0);
  BUFF I346 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I347 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I348 (wenr_0[9:9], wc_0);
  BUFF I349 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I350 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I351 (wenr_0[10:10], wc_0);
  BUFF I352 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I353 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I354 (wenr_0[11:11], wc_0);
  BUFF I355 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I356 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I357 (wenr_0[12:12], wc_0);
  BUFF I358 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I359 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I360 (wenr_0[13:13], wc_0);
  BUFF I361 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I362 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I363 (wenr_0[14:14], wc_0);
  BUFF I364 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I365 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I366 (wenr_0[15:15], wc_0);
  BUFF I367 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I368 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I369 (wenr_0[16:16], wc_0);
  BUFF I370 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I371 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I372 (wenr_0[17:17], wc_0);
  BUFF I373 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I374 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I375 (wenr_0[18:18], wc_0);
  BUFF I376 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I377 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I378 (wenr_0[19:19], wc_0);
  BUFF I379 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I380 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I381 (wenr_0[20:20], wc_0);
  BUFF I382 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I383 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I384 (wenr_0[21:21], wc_0);
  BUFF I385 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I386 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I387 (wenr_0[22:22], wc_0);
  BUFF I388 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I389 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I390 (wenr_0[23:23], wc_0);
  BUFF I391 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I392 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I393 (wenr_0[24:24], wc_0);
  BUFF I394 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I395 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I396 (wenr_0[25:25], wc_0);
  BUFF I397 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I398 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I399 (wenr_0[26:26], wc_0);
  BUFF I400 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I401 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I402 (wenr_0[27:27], wc_0);
  BUFF I403 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I404 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I405 (wenr_0[28:28], wc_0);
  BUFF I406 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I407 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I408 (wenr_0[29:29], wc_0);
  BUFF I409 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I410 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I411 (wenr_0[30:30], wc_0);
  BUFF I412 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I413 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I414 (wenr_0[31:31], wc_0);
  BUFF I415 (wf_0[32:32], conwgif_0[32:32]);
  BUFF I416 (wt_0[32:32], conwgit_0[32:32]);
  BUFF I417 (wenr_0[32:32], wc_0);
  C3 I418 (simp4191_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I419 (simp4191_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I420 (simp4191_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I421 (simp4191_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I422 (simp4191_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I423 (simp4191_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I424 (simp4191_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I425 (simp4191_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I426 (simp4191_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I427 (simp4191_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I428 (simp4191_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  BUFF I429 (simp4191_0[11:11], wacks_0[32:32]);
  C3 I430 (simp4192_0[0:0], simp4191_0[0:0], simp4191_0[1:1], simp4191_0[2:2]);
  C3 I431 (simp4192_0[1:1], simp4191_0[3:3], simp4191_0[4:4], simp4191_0[5:5]);
  C3 I432 (simp4192_0[2:2], simp4191_0[6:6], simp4191_0[7:7], simp4191_0[8:8]);
  C3 I433 (simp4192_0[3:3], simp4191_0[9:9], simp4191_0[10:10], simp4191_0[11:11]);
  C3 I434 (simp4193_0[0:0], simp4192_0[0:0], simp4192_0[1:1], simp4192_0[2:2]);
  BUFF I435 (simp4193_0[1:1], simp4192_0[3:3]);
  C2 I436 (wd_0r, simp4193_0[0:0], simp4193_0[1:1]);
  AND2 I437 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I438 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I439 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I440 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I441 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I442 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I443 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I444 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I445 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I446 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I447 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I448 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I449 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I450 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I451 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I452 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I453 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I454 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I455 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I456 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I457 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I458 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I459 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I460 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I461 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I462 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I463 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I464 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I465 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I466 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I467 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I468 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I469 (rd_1r0, df_0[32:32], rg_1r);
  AND2 I470 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I471 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I472 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I473 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I474 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I475 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I476 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I477 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I478 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I479 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I480 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I481 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I482 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I483 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I484 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I485 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I486 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I487 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I488 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I489 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I490 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I491 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I492 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I493 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I494 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I495 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I496 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I497 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I498 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I499 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I500 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I501 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I502 (rd_1r1, dt_0[32:32], rg_1r);
  NOR3 I503 (simp4861_0[0:0], rg_0r, rg_1r, rg_0a);
  INV I504 (simp4861_0[1:1], rg_1a);
  NAND2 I505 (anyread_0, simp4861_0[0:0], simp4861_0[1:1]);
  BUFF I506 (wg_0a, wd_0a);
  BUFF I507 (rg_0a, rd_0a);
  BUFF I508 (rg_1a, rd_1a);
endmodule

// tkvopr74_wo0w74_ro26w5o25w1o25w1o20w5o9w1o15w5o8w1o10w5o7w1o7w3o38w32o37w1o71w2o71w2o25w1o31w6o38w32
//   o6w1o3w4o0w3 TeakV "opr" 74 [] [0] [26,25,25,20,9,15,8,10,7,7,38,37,71,71,25,31,38,6,3,0] [Many [74]
//   ,Many [0],Many [0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0],Many [5,1,1,5,1,5,1,5,1,3,32,1,2,2,1,6,32,1
//   ,4,3]]
module tkvopr74_wo0w74_ro26w5o25w1o25w1o20w5o9w1o15w5o8w1o10w5o7w1o7w3o38w32o37w1o71w2o71w2o25w1o31w6o38w32o6w1o3w4o0w3 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rg_2r, rg_2a, rg_3r, rg_3a, rg_4r, rg_4a, rg_5r, rg_5a, rg_6r, rg_6a, rg_7r, rg_7a, rg_8r, rg_8a, rg_9r, rg_9a, rg_10r, rg_10a, rg_11r, rg_11a, rg_12r, rg_12a, rg_13r, rg_13a, rg_14r, rg_14a, rg_15r, rg_15a, rg_16r, rg_16a, rg_17r, rg_17a, rg_18r, rg_18a, rg_19r, rg_19a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, rd_2r0, rd_2r1, rd_2a, rd_3r0, rd_3r1, rd_3a, rd_4r0, rd_4r1, rd_4a, rd_5r0, rd_5r1, rd_5a, rd_6r0, rd_6r1, rd_6a, rd_7r0, rd_7r1, rd_7a, rd_8r0, rd_8r1, rd_8a, rd_9r0, rd_9r1, rd_9a, rd_10r0, rd_10r1, rd_10a, rd_11r0, rd_11r1, rd_11a, rd_12r0, rd_12r1, rd_12a, rd_13r0, rd_13r1, rd_13a, rd_14r0, rd_14r1, rd_14a, rd_15r0, rd_15r1, rd_15a, rd_16r0, rd_16r1, rd_16a, rd_17r0, rd_17r1, rd_17a, rd_18r0, rd_18r1, rd_18a, rd_19r0, rd_19r1, rd_19a, reset);
  input [73:0] wg_0r0;
  input [73:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  input rg_2r;
  output rg_2a;
  input rg_3r;
  output rg_3a;
  input rg_4r;
  output rg_4a;
  input rg_5r;
  output rg_5a;
  input rg_6r;
  output rg_6a;
  input rg_7r;
  output rg_7a;
  input rg_8r;
  output rg_8a;
  input rg_9r;
  output rg_9a;
  input rg_10r;
  output rg_10a;
  input rg_11r;
  output rg_11a;
  input rg_12r;
  output rg_12a;
  input rg_13r;
  output rg_13a;
  input rg_14r;
  output rg_14a;
  input rg_15r;
  output rg_15a;
  input rg_16r;
  output rg_16a;
  input rg_17r;
  output rg_17a;
  input rg_18r;
  output rg_18a;
  input rg_19r;
  output rg_19a;
  output [4:0] rd_0r0;
  output [4:0] rd_0r1;
  input rd_0a;
  output rd_1r0;
  output rd_1r1;
  input rd_1a;
  output rd_2r0;
  output rd_2r1;
  input rd_2a;
  output [4:0] rd_3r0;
  output [4:0] rd_3r1;
  input rd_3a;
  output rd_4r0;
  output rd_4r1;
  input rd_4a;
  output [4:0] rd_5r0;
  output [4:0] rd_5r1;
  input rd_5a;
  output rd_6r0;
  output rd_6r1;
  input rd_6a;
  output [4:0] rd_7r0;
  output [4:0] rd_7r1;
  input rd_7a;
  output rd_8r0;
  output rd_8r1;
  input rd_8a;
  output [2:0] rd_9r0;
  output [2:0] rd_9r1;
  input rd_9a;
  output [31:0] rd_10r0;
  output [31:0] rd_10r1;
  input rd_10a;
  output rd_11r0;
  output rd_11r1;
  input rd_11a;
  output [1:0] rd_12r0;
  output [1:0] rd_12r1;
  input rd_12a;
  output [1:0] rd_13r0;
  output [1:0] rd_13r1;
  input rd_13a;
  output rd_14r0;
  output rd_14r1;
  input rd_14a;
  output [5:0] rd_15r0;
  output [5:0] rd_15r1;
  input rd_15a;
  output [31:0] rd_16r0;
  output [31:0] rd_16r1;
  input rd_16a;
  output rd_17r0;
  output rd_17r1;
  input rd_17a;
  output [3:0] rd_18r0;
  output [3:0] rd_18r1;
  input rd_18a;
  output [2:0] rd_19r0;
  output [2:0] rd_19r1;
  input rd_19a;
  input reset;
  wire [73:0] wf_0;
  wire [73:0] wt_0;
  wire [73:0] df_0;
  wire [73:0] dt_0;
  wire wc_0;
  wire [73:0] wacks_0;
  wire [73:0] wenr_0;
  wire [73:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [73:0] drlgf_0;
  wire [73:0] drlgt_0;
  wire [73:0] comp0_0;
  wire [24:0] simp5321_0;
  wire [8:0] simp5322_0;
  wire [2:0] simp5323_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [73:0] conwgit_0;
  wire [73:0] conwgif_0;
  wire conwig_0;
  wire [24:0] simp9111_0;
  wire [8:0] simp9112_0;
  wire [2:0] simp9113_0;
  wire [13:0] simp11361_0;
  wire [4:0] simp11362_0;
  wire [1:0] simp11363_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (wen_0[32:32], wenr_0[32:32], nreset_0);
  AND2 I34 (wen_0[33:33], wenr_0[33:33], nreset_0);
  AND2 I35 (wen_0[34:34], wenr_0[34:34], nreset_0);
  AND2 I36 (wen_0[35:35], wenr_0[35:35], nreset_0);
  AND2 I37 (wen_0[36:36], wenr_0[36:36], nreset_0);
  AND2 I38 (wen_0[37:37], wenr_0[37:37], nreset_0);
  AND2 I39 (wen_0[38:38], wenr_0[38:38], nreset_0);
  AND2 I40 (wen_0[39:39], wenr_0[39:39], nreset_0);
  AND2 I41 (wen_0[40:40], wenr_0[40:40], nreset_0);
  AND2 I42 (wen_0[41:41], wenr_0[41:41], nreset_0);
  AND2 I43 (wen_0[42:42], wenr_0[42:42], nreset_0);
  AND2 I44 (wen_0[43:43], wenr_0[43:43], nreset_0);
  AND2 I45 (wen_0[44:44], wenr_0[44:44], nreset_0);
  AND2 I46 (wen_0[45:45], wenr_0[45:45], nreset_0);
  AND2 I47 (wen_0[46:46], wenr_0[46:46], nreset_0);
  AND2 I48 (wen_0[47:47], wenr_0[47:47], nreset_0);
  AND2 I49 (wen_0[48:48], wenr_0[48:48], nreset_0);
  AND2 I50 (wen_0[49:49], wenr_0[49:49], nreset_0);
  AND2 I51 (wen_0[50:50], wenr_0[50:50], nreset_0);
  AND2 I52 (wen_0[51:51], wenr_0[51:51], nreset_0);
  AND2 I53 (wen_0[52:52], wenr_0[52:52], nreset_0);
  AND2 I54 (wen_0[53:53], wenr_0[53:53], nreset_0);
  AND2 I55 (wen_0[54:54], wenr_0[54:54], nreset_0);
  AND2 I56 (wen_0[55:55], wenr_0[55:55], nreset_0);
  AND2 I57 (wen_0[56:56], wenr_0[56:56], nreset_0);
  AND2 I58 (wen_0[57:57], wenr_0[57:57], nreset_0);
  AND2 I59 (wen_0[58:58], wenr_0[58:58], nreset_0);
  AND2 I60 (wen_0[59:59], wenr_0[59:59], nreset_0);
  AND2 I61 (wen_0[60:60], wenr_0[60:60], nreset_0);
  AND2 I62 (wen_0[61:61], wenr_0[61:61], nreset_0);
  AND2 I63 (wen_0[62:62], wenr_0[62:62], nreset_0);
  AND2 I64 (wen_0[63:63], wenr_0[63:63], nreset_0);
  AND2 I65 (wen_0[64:64], wenr_0[64:64], nreset_0);
  AND2 I66 (wen_0[65:65], wenr_0[65:65], nreset_0);
  AND2 I67 (wen_0[66:66], wenr_0[66:66], nreset_0);
  AND2 I68 (wen_0[67:67], wenr_0[67:67], nreset_0);
  AND2 I69 (wen_0[68:68], wenr_0[68:68], nreset_0);
  AND2 I70 (wen_0[69:69], wenr_0[69:69], nreset_0);
  AND2 I71 (wen_0[70:70], wenr_0[70:70], nreset_0);
  AND2 I72 (wen_0[71:71], wenr_0[71:71], nreset_0);
  AND2 I73 (wen_0[72:72], wenr_0[72:72], nreset_0);
  AND2 I74 (wen_0[73:73], wenr_0[73:73], nreset_0);
  AND2 I75 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I76 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I77 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I78 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I79 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I80 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I81 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I82 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I83 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I84 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I85 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I86 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I87 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I88 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I89 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I90 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I91 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I92 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I93 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I94 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I95 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I96 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I97 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I98 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I99 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I100 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I101 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I102 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I103 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I104 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I105 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I106 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I107 (drlgf_0[32:32], wf_0[32:32], wen_0[32:32]);
  AND2 I108 (drlgf_0[33:33], wf_0[33:33], wen_0[33:33]);
  AND2 I109 (drlgf_0[34:34], wf_0[34:34], wen_0[34:34]);
  AND2 I110 (drlgf_0[35:35], wf_0[35:35], wen_0[35:35]);
  AND2 I111 (drlgf_0[36:36], wf_0[36:36], wen_0[36:36]);
  AND2 I112 (drlgf_0[37:37], wf_0[37:37], wen_0[37:37]);
  AND2 I113 (drlgf_0[38:38], wf_0[38:38], wen_0[38:38]);
  AND2 I114 (drlgf_0[39:39], wf_0[39:39], wen_0[39:39]);
  AND2 I115 (drlgf_0[40:40], wf_0[40:40], wen_0[40:40]);
  AND2 I116 (drlgf_0[41:41], wf_0[41:41], wen_0[41:41]);
  AND2 I117 (drlgf_0[42:42], wf_0[42:42], wen_0[42:42]);
  AND2 I118 (drlgf_0[43:43], wf_0[43:43], wen_0[43:43]);
  AND2 I119 (drlgf_0[44:44], wf_0[44:44], wen_0[44:44]);
  AND2 I120 (drlgf_0[45:45], wf_0[45:45], wen_0[45:45]);
  AND2 I121 (drlgf_0[46:46], wf_0[46:46], wen_0[46:46]);
  AND2 I122 (drlgf_0[47:47], wf_0[47:47], wen_0[47:47]);
  AND2 I123 (drlgf_0[48:48], wf_0[48:48], wen_0[48:48]);
  AND2 I124 (drlgf_0[49:49], wf_0[49:49], wen_0[49:49]);
  AND2 I125 (drlgf_0[50:50], wf_0[50:50], wen_0[50:50]);
  AND2 I126 (drlgf_0[51:51], wf_0[51:51], wen_0[51:51]);
  AND2 I127 (drlgf_0[52:52], wf_0[52:52], wen_0[52:52]);
  AND2 I128 (drlgf_0[53:53], wf_0[53:53], wen_0[53:53]);
  AND2 I129 (drlgf_0[54:54], wf_0[54:54], wen_0[54:54]);
  AND2 I130 (drlgf_0[55:55], wf_0[55:55], wen_0[55:55]);
  AND2 I131 (drlgf_0[56:56], wf_0[56:56], wen_0[56:56]);
  AND2 I132 (drlgf_0[57:57], wf_0[57:57], wen_0[57:57]);
  AND2 I133 (drlgf_0[58:58], wf_0[58:58], wen_0[58:58]);
  AND2 I134 (drlgf_0[59:59], wf_0[59:59], wen_0[59:59]);
  AND2 I135 (drlgf_0[60:60], wf_0[60:60], wen_0[60:60]);
  AND2 I136 (drlgf_0[61:61], wf_0[61:61], wen_0[61:61]);
  AND2 I137 (drlgf_0[62:62], wf_0[62:62], wen_0[62:62]);
  AND2 I138 (drlgf_0[63:63], wf_0[63:63], wen_0[63:63]);
  AND2 I139 (drlgf_0[64:64], wf_0[64:64], wen_0[64:64]);
  AND2 I140 (drlgf_0[65:65], wf_0[65:65], wen_0[65:65]);
  AND2 I141 (drlgf_0[66:66], wf_0[66:66], wen_0[66:66]);
  AND2 I142 (drlgf_0[67:67], wf_0[67:67], wen_0[67:67]);
  AND2 I143 (drlgf_0[68:68], wf_0[68:68], wen_0[68:68]);
  AND2 I144 (drlgf_0[69:69], wf_0[69:69], wen_0[69:69]);
  AND2 I145 (drlgf_0[70:70], wf_0[70:70], wen_0[70:70]);
  AND2 I146 (drlgf_0[71:71], wf_0[71:71], wen_0[71:71]);
  AND2 I147 (drlgf_0[72:72], wf_0[72:72], wen_0[72:72]);
  AND2 I148 (drlgf_0[73:73], wf_0[73:73], wen_0[73:73]);
  AND2 I149 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I150 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I151 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I152 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I153 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I154 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I155 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I156 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I157 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I158 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I159 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I160 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I161 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I162 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I163 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I164 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I165 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I166 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I167 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I168 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I169 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I170 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I171 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I172 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I173 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I174 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I175 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I176 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I177 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I178 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I179 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I180 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  AND2 I181 (drlgt_0[32:32], wt_0[32:32], wen_0[32:32]);
  AND2 I182 (drlgt_0[33:33], wt_0[33:33], wen_0[33:33]);
  AND2 I183 (drlgt_0[34:34], wt_0[34:34], wen_0[34:34]);
  AND2 I184 (drlgt_0[35:35], wt_0[35:35], wen_0[35:35]);
  AND2 I185 (drlgt_0[36:36], wt_0[36:36], wen_0[36:36]);
  AND2 I186 (drlgt_0[37:37], wt_0[37:37], wen_0[37:37]);
  AND2 I187 (drlgt_0[38:38], wt_0[38:38], wen_0[38:38]);
  AND2 I188 (drlgt_0[39:39], wt_0[39:39], wen_0[39:39]);
  AND2 I189 (drlgt_0[40:40], wt_0[40:40], wen_0[40:40]);
  AND2 I190 (drlgt_0[41:41], wt_0[41:41], wen_0[41:41]);
  AND2 I191 (drlgt_0[42:42], wt_0[42:42], wen_0[42:42]);
  AND2 I192 (drlgt_0[43:43], wt_0[43:43], wen_0[43:43]);
  AND2 I193 (drlgt_0[44:44], wt_0[44:44], wen_0[44:44]);
  AND2 I194 (drlgt_0[45:45], wt_0[45:45], wen_0[45:45]);
  AND2 I195 (drlgt_0[46:46], wt_0[46:46], wen_0[46:46]);
  AND2 I196 (drlgt_0[47:47], wt_0[47:47], wen_0[47:47]);
  AND2 I197 (drlgt_0[48:48], wt_0[48:48], wen_0[48:48]);
  AND2 I198 (drlgt_0[49:49], wt_0[49:49], wen_0[49:49]);
  AND2 I199 (drlgt_0[50:50], wt_0[50:50], wen_0[50:50]);
  AND2 I200 (drlgt_0[51:51], wt_0[51:51], wen_0[51:51]);
  AND2 I201 (drlgt_0[52:52], wt_0[52:52], wen_0[52:52]);
  AND2 I202 (drlgt_0[53:53], wt_0[53:53], wen_0[53:53]);
  AND2 I203 (drlgt_0[54:54], wt_0[54:54], wen_0[54:54]);
  AND2 I204 (drlgt_0[55:55], wt_0[55:55], wen_0[55:55]);
  AND2 I205 (drlgt_0[56:56], wt_0[56:56], wen_0[56:56]);
  AND2 I206 (drlgt_0[57:57], wt_0[57:57], wen_0[57:57]);
  AND2 I207 (drlgt_0[58:58], wt_0[58:58], wen_0[58:58]);
  AND2 I208 (drlgt_0[59:59], wt_0[59:59], wen_0[59:59]);
  AND2 I209 (drlgt_0[60:60], wt_0[60:60], wen_0[60:60]);
  AND2 I210 (drlgt_0[61:61], wt_0[61:61], wen_0[61:61]);
  AND2 I211 (drlgt_0[62:62], wt_0[62:62], wen_0[62:62]);
  AND2 I212 (drlgt_0[63:63], wt_0[63:63], wen_0[63:63]);
  AND2 I213 (drlgt_0[64:64], wt_0[64:64], wen_0[64:64]);
  AND2 I214 (drlgt_0[65:65], wt_0[65:65], wen_0[65:65]);
  AND2 I215 (drlgt_0[66:66], wt_0[66:66], wen_0[66:66]);
  AND2 I216 (drlgt_0[67:67], wt_0[67:67], wen_0[67:67]);
  AND2 I217 (drlgt_0[68:68], wt_0[68:68], wen_0[68:68]);
  AND2 I218 (drlgt_0[69:69], wt_0[69:69], wen_0[69:69]);
  AND2 I219 (drlgt_0[70:70], wt_0[70:70], wen_0[70:70]);
  AND2 I220 (drlgt_0[71:71], wt_0[71:71], wen_0[71:71]);
  AND2 I221 (drlgt_0[72:72], wt_0[72:72], wen_0[72:72]);
  AND2 I222 (drlgt_0[73:73], wt_0[73:73], wen_0[73:73]);
  NOR2 I223 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I224 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I225 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I226 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I227 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I228 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I229 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I230 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I231 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I232 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I233 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I234 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I235 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I236 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I237 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I238 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I239 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I240 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I241 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I242 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I243 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I244 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I245 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I246 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I247 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I248 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I249 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I250 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I251 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I252 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I253 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I254 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR2 I255 (df_0[32:32], dt_0[32:32], drlgt_0[32:32]);
  NOR2 I256 (df_0[33:33], dt_0[33:33], drlgt_0[33:33]);
  NOR2 I257 (df_0[34:34], dt_0[34:34], drlgt_0[34:34]);
  NOR2 I258 (df_0[35:35], dt_0[35:35], drlgt_0[35:35]);
  NOR2 I259 (df_0[36:36], dt_0[36:36], drlgt_0[36:36]);
  NOR2 I260 (df_0[37:37], dt_0[37:37], drlgt_0[37:37]);
  NOR2 I261 (df_0[38:38], dt_0[38:38], drlgt_0[38:38]);
  NOR2 I262 (df_0[39:39], dt_0[39:39], drlgt_0[39:39]);
  NOR2 I263 (df_0[40:40], dt_0[40:40], drlgt_0[40:40]);
  NOR2 I264 (df_0[41:41], dt_0[41:41], drlgt_0[41:41]);
  NOR2 I265 (df_0[42:42], dt_0[42:42], drlgt_0[42:42]);
  NOR2 I266 (df_0[43:43], dt_0[43:43], drlgt_0[43:43]);
  NOR2 I267 (df_0[44:44], dt_0[44:44], drlgt_0[44:44]);
  NOR2 I268 (df_0[45:45], dt_0[45:45], drlgt_0[45:45]);
  NOR2 I269 (df_0[46:46], dt_0[46:46], drlgt_0[46:46]);
  NOR2 I270 (df_0[47:47], dt_0[47:47], drlgt_0[47:47]);
  NOR2 I271 (df_0[48:48], dt_0[48:48], drlgt_0[48:48]);
  NOR2 I272 (df_0[49:49], dt_0[49:49], drlgt_0[49:49]);
  NOR2 I273 (df_0[50:50], dt_0[50:50], drlgt_0[50:50]);
  NOR2 I274 (df_0[51:51], dt_0[51:51], drlgt_0[51:51]);
  NOR2 I275 (df_0[52:52], dt_0[52:52], drlgt_0[52:52]);
  NOR2 I276 (df_0[53:53], dt_0[53:53], drlgt_0[53:53]);
  NOR2 I277 (df_0[54:54], dt_0[54:54], drlgt_0[54:54]);
  NOR2 I278 (df_0[55:55], dt_0[55:55], drlgt_0[55:55]);
  NOR2 I279 (df_0[56:56], dt_0[56:56], drlgt_0[56:56]);
  NOR2 I280 (df_0[57:57], dt_0[57:57], drlgt_0[57:57]);
  NOR2 I281 (df_0[58:58], dt_0[58:58], drlgt_0[58:58]);
  NOR2 I282 (df_0[59:59], dt_0[59:59], drlgt_0[59:59]);
  NOR2 I283 (df_0[60:60], dt_0[60:60], drlgt_0[60:60]);
  NOR2 I284 (df_0[61:61], dt_0[61:61], drlgt_0[61:61]);
  NOR2 I285 (df_0[62:62], dt_0[62:62], drlgt_0[62:62]);
  NOR2 I286 (df_0[63:63], dt_0[63:63], drlgt_0[63:63]);
  NOR2 I287 (df_0[64:64], dt_0[64:64], drlgt_0[64:64]);
  NOR2 I288 (df_0[65:65], dt_0[65:65], drlgt_0[65:65]);
  NOR2 I289 (df_0[66:66], dt_0[66:66], drlgt_0[66:66]);
  NOR2 I290 (df_0[67:67], dt_0[67:67], drlgt_0[67:67]);
  NOR2 I291 (df_0[68:68], dt_0[68:68], drlgt_0[68:68]);
  NOR2 I292 (df_0[69:69], dt_0[69:69], drlgt_0[69:69]);
  NOR2 I293 (df_0[70:70], dt_0[70:70], drlgt_0[70:70]);
  NOR2 I294 (df_0[71:71], dt_0[71:71], drlgt_0[71:71]);
  NOR2 I295 (df_0[72:72], dt_0[72:72], drlgt_0[72:72]);
  NOR2 I296 (df_0[73:73], dt_0[73:73], drlgt_0[73:73]);
  NOR3 I297 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I298 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I299 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I300 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I301 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I302 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I303 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I304 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I305 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I306 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I307 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I308 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I309 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I310 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I311 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I312 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I313 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I314 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I315 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I316 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I317 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I318 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I319 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I320 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I321 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I322 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I323 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I324 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I325 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I326 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I327 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I328 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  NOR3 I329 (dt_0[32:32], df_0[32:32], drlgf_0[32:32], reset);
  NOR3 I330 (dt_0[33:33], df_0[33:33], drlgf_0[33:33], reset);
  NOR3 I331 (dt_0[34:34], df_0[34:34], drlgf_0[34:34], reset);
  NOR3 I332 (dt_0[35:35], df_0[35:35], drlgf_0[35:35], reset);
  NOR3 I333 (dt_0[36:36], df_0[36:36], drlgf_0[36:36], reset);
  NOR3 I334 (dt_0[37:37], df_0[37:37], drlgf_0[37:37], reset);
  NOR3 I335 (dt_0[38:38], df_0[38:38], drlgf_0[38:38], reset);
  NOR3 I336 (dt_0[39:39], df_0[39:39], drlgf_0[39:39], reset);
  NOR3 I337 (dt_0[40:40], df_0[40:40], drlgf_0[40:40], reset);
  NOR3 I338 (dt_0[41:41], df_0[41:41], drlgf_0[41:41], reset);
  NOR3 I339 (dt_0[42:42], df_0[42:42], drlgf_0[42:42], reset);
  NOR3 I340 (dt_0[43:43], df_0[43:43], drlgf_0[43:43], reset);
  NOR3 I341 (dt_0[44:44], df_0[44:44], drlgf_0[44:44], reset);
  NOR3 I342 (dt_0[45:45], df_0[45:45], drlgf_0[45:45], reset);
  NOR3 I343 (dt_0[46:46], df_0[46:46], drlgf_0[46:46], reset);
  NOR3 I344 (dt_0[47:47], df_0[47:47], drlgf_0[47:47], reset);
  NOR3 I345 (dt_0[48:48], df_0[48:48], drlgf_0[48:48], reset);
  NOR3 I346 (dt_0[49:49], df_0[49:49], drlgf_0[49:49], reset);
  NOR3 I347 (dt_0[50:50], df_0[50:50], drlgf_0[50:50], reset);
  NOR3 I348 (dt_0[51:51], df_0[51:51], drlgf_0[51:51], reset);
  NOR3 I349 (dt_0[52:52], df_0[52:52], drlgf_0[52:52], reset);
  NOR3 I350 (dt_0[53:53], df_0[53:53], drlgf_0[53:53], reset);
  NOR3 I351 (dt_0[54:54], df_0[54:54], drlgf_0[54:54], reset);
  NOR3 I352 (dt_0[55:55], df_0[55:55], drlgf_0[55:55], reset);
  NOR3 I353 (dt_0[56:56], df_0[56:56], drlgf_0[56:56], reset);
  NOR3 I354 (dt_0[57:57], df_0[57:57], drlgf_0[57:57], reset);
  NOR3 I355 (dt_0[58:58], df_0[58:58], drlgf_0[58:58], reset);
  NOR3 I356 (dt_0[59:59], df_0[59:59], drlgf_0[59:59], reset);
  NOR3 I357 (dt_0[60:60], df_0[60:60], drlgf_0[60:60], reset);
  NOR3 I358 (dt_0[61:61], df_0[61:61], drlgf_0[61:61], reset);
  NOR3 I359 (dt_0[62:62], df_0[62:62], drlgf_0[62:62], reset);
  NOR3 I360 (dt_0[63:63], df_0[63:63], drlgf_0[63:63], reset);
  NOR3 I361 (dt_0[64:64], df_0[64:64], drlgf_0[64:64], reset);
  NOR3 I362 (dt_0[65:65], df_0[65:65], drlgf_0[65:65], reset);
  NOR3 I363 (dt_0[66:66], df_0[66:66], drlgf_0[66:66], reset);
  NOR3 I364 (dt_0[67:67], df_0[67:67], drlgf_0[67:67], reset);
  NOR3 I365 (dt_0[68:68], df_0[68:68], drlgf_0[68:68], reset);
  NOR3 I366 (dt_0[69:69], df_0[69:69], drlgf_0[69:69], reset);
  NOR3 I367 (dt_0[70:70], df_0[70:70], drlgf_0[70:70], reset);
  NOR3 I368 (dt_0[71:71], df_0[71:71], drlgf_0[71:71], reset);
  NOR3 I369 (dt_0[72:72], df_0[72:72], drlgf_0[72:72], reset);
  NOR3 I370 (dt_0[73:73], df_0[73:73], drlgf_0[73:73], reset);
  AO22 I371 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I372 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I373 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I374 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I375 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I376 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I377 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I378 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I379 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I380 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I381 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I382 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I383 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I384 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I385 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I386 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I387 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I388 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I389 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I390 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I391 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I392 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I393 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I394 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I395 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I396 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I397 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I398 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I399 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I400 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I401 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I402 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  AO22 I403 (wacks_0[32:32], drlgf_0[32:32], df_0[32:32], drlgt_0[32:32], dt_0[32:32]);
  AO22 I404 (wacks_0[33:33], drlgf_0[33:33], df_0[33:33], drlgt_0[33:33], dt_0[33:33]);
  AO22 I405 (wacks_0[34:34], drlgf_0[34:34], df_0[34:34], drlgt_0[34:34], dt_0[34:34]);
  AO22 I406 (wacks_0[35:35], drlgf_0[35:35], df_0[35:35], drlgt_0[35:35], dt_0[35:35]);
  AO22 I407 (wacks_0[36:36], drlgf_0[36:36], df_0[36:36], drlgt_0[36:36], dt_0[36:36]);
  AO22 I408 (wacks_0[37:37], drlgf_0[37:37], df_0[37:37], drlgt_0[37:37], dt_0[37:37]);
  AO22 I409 (wacks_0[38:38], drlgf_0[38:38], df_0[38:38], drlgt_0[38:38], dt_0[38:38]);
  AO22 I410 (wacks_0[39:39], drlgf_0[39:39], df_0[39:39], drlgt_0[39:39], dt_0[39:39]);
  AO22 I411 (wacks_0[40:40], drlgf_0[40:40], df_0[40:40], drlgt_0[40:40], dt_0[40:40]);
  AO22 I412 (wacks_0[41:41], drlgf_0[41:41], df_0[41:41], drlgt_0[41:41], dt_0[41:41]);
  AO22 I413 (wacks_0[42:42], drlgf_0[42:42], df_0[42:42], drlgt_0[42:42], dt_0[42:42]);
  AO22 I414 (wacks_0[43:43], drlgf_0[43:43], df_0[43:43], drlgt_0[43:43], dt_0[43:43]);
  AO22 I415 (wacks_0[44:44], drlgf_0[44:44], df_0[44:44], drlgt_0[44:44], dt_0[44:44]);
  AO22 I416 (wacks_0[45:45], drlgf_0[45:45], df_0[45:45], drlgt_0[45:45], dt_0[45:45]);
  AO22 I417 (wacks_0[46:46], drlgf_0[46:46], df_0[46:46], drlgt_0[46:46], dt_0[46:46]);
  AO22 I418 (wacks_0[47:47], drlgf_0[47:47], df_0[47:47], drlgt_0[47:47], dt_0[47:47]);
  AO22 I419 (wacks_0[48:48], drlgf_0[48:48], df_0[48:48], drlgt_0[48:48], dt_0[48:48]);
  AO22 I420 (wacks_0[49:49], drlgf_0[49:49], df_0[49:49], drlgt_0[49:49], dt_0[49:49]);
  AO22 I421 (wacks_0[50:50], drlgf_0[50:50], df_0[50:50], drlgt_0[50:50], dt_0[50:50]);
  AO22 I422 (wacks_0[51:51], drlgf_0[51:51], df_0[51:51], drlgt_0[51:51], dt_0[51:51]);
  AO22 I423 (wacks_0[52:52], drlgf_0[52:52], df_0[52:52], drlgt_0[52:52], dt_0[52:52]);
  AO22 I424 (wacks_0[53:53], drlgf_0[53:53], df_0[53:53], drlgt_0[53:53], dt_0[53:53]);
  AO22 I425 (wacks_0[54:54], drlgf_0[54:54], df_0[54:54], drlgt_0[54:54], dt_0[54:54]);
  AO22 I426 (wacks_0[55:55], drlgf_0[55:55], df_0[55:55], drlgt_0[55:55], dt_0[55:55]);
  AO22 I427 (wacks_0[56:56], drlgf_0[56:56], df_0[56:56], drlgt_0[56:56], dt_0[56:56]);
  AO22 I428 (wacks_0[57:57], drlgf_0[57:57], df_0[57:57], drlgt_0[57:57], dt_0[57:57]);
  AO22 I429 (wacks_0[58:58], drlgf_0[58:58], df_0[58:58], drlgt_0[58:58], dt_0[58:58]);
  AO22 I430 (wacks_0[59:59], drlgf_0[59:59], df_0[59:59], drlgt_0[59:59], dt_0[59:59]);
  AO22 I431 (wacks_0[60:60], drlgf_0[60:60], df_0[60:60], drlgt_0[60:60], dt_0[60:60]);
  AO22 I432 (wacks_0[61:61], drlgf_0[61:61], df_0[61:61], drlgt_0[61:61], dt_0[61:61]);
  AO22 I433 (wacks_0[62:62], drlgf_0[62:62], df_0[62:62], drlgt_0[62:62], dt_0[62:62]);
  AO22 I434 (wacks_0[63:63], drlgf_0[63:63], df_0[63:63], drlgt_0[63:63], dt_0[63:63]);
  AO22 I435 (wacks_0[64:64], drlgf_0[64:64], df_0[64:64], drlgt_0[64:64], dt_0[64:64]);
  AO22 I436 (wacks_0[65:65], drlgf_0[65:65], df_0[65:65], drlgt_0[65:65], dt_0[65:65]);
  AO22 I437 (wacks_0[66:66], drlgf_0[66:66], df_0[66:66], drlgt_0[66:66], dt_0[66:66]);
  AO22 I438 (wacks_0[67:67], drlgf_0[67:67], df_0[67:67], drlgt_0[67:67], dt_0[67:67]);
  AO22 I439 (wacks_0[68:68], drlgf_0[68:68], df_0[68:68], drlgt_0[68:68], dt_0[68:68]);
  AO22 I440 (wacks_0[69:69], drlgf_0[69:69], df_0[69:69], drlgt_0[69:69], dt_0[69:69]);
  AO22 I441 (wacks_0[70:70], drlgf_0[70:70], df_0[70:70], drlgt_0[70:70], dt_0[70:70]);
  AO22 I442 (wacks_0[71:71], drlgf_0[71:71], df_0[71:71], drlgt_0[71:71], dt_0[71:71]);
  AO22 I443 (wacks_0[72:72], drlgf_0[72:72], df_0[72:72], drlgt_0[72:72], dt_0[72:72]);
  AO22 I444 (wacks_0[73:73], drlgf_0[73:73], df_0[73:73], drlgt_0[73:73], dt_0[73:73]);
  OR2 I445 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I446 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I447 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I448 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I449 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I450 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I451 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I452 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I453 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I454 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I455 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I456 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I457 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I458 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I459 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I460 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I461 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I462 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I463 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I464 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I465 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I466 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I467 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I468 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I469 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I470 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I471 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I472 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I473 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I474 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I475 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I476 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  OR2 I477 (comp0_0[32:32], wg_0r0[32:32], wg_0r1[32:32]);
  OR2 I478 (comp0_0[33:33], wg_0r0[33:33], wg_0r1[33:33]);
  OR2 I479 (comp0_0[34:34], wg_0r0[34:34], wg_0r1[34:34]);
  OR2 I480 (comp0_0[35:35], wg_0r0[35:35], wg_0r1[35:35]);
  OR2 I481 (comp0_0[36:36], wg_0r0[36:36], wg_0r1[36:36]);
  OR2 I482 (comp0_0[37:37], wg_0r0[37:37], wg_0r1[37:37]);
  OR2 I483 (comp0_0[38:38], wg_0r0[38:38], wg_0r1[38:38]);
  OR2 I484 (comp0_0[39:39], wg_0r0[39:39], wg_0r1[39:39]);
  OR2 I485 (comp0_0[40:40], wg_0r0[40:40], wg_0r1[40:40]);
  OR2 I486 (comp0_0[41:41], wg_0r0[41:41], wg_0r1[41:41]);
  OR2 I487 (comp0_0[42:42], wg_0r0[42:42], wg_0r1[42:42]);
  OR2 I488 (comp0_0[43:43], wg_0r0[43:43], wg_0r1[43:43]);
  OR2 I489 (comp0_0[44:44], wg_0r0[44:44], wg_0r1[44:44]);
  OR2 I490 (comp0_0[45:45], wg_0r0[45:45], wg_0r1[45:45]);
  OR2 I491 (comp0_0[46:46], wg_0r0[46:46], wg_0r1[46:46]);
  OR2 I492 (comp0_0[47:47], wg_0r0[47:47], wg_0r1[47:47]);
  OR2 I493 (comp0_0[48:48], wg_0r0[48:48], wg_0r1[48:48]);
  OR2 I494 (comp0_0[49:49], wg_0r0[49:49], wg_0r1[49:49]);
  OR2 I495 (comp0_0[50:50], wg_0r0[50:50], wg_0r1[50:50]);
  OR2 I496 (comp0_0[51:51], wg_0r0[51:51], wg_0r1[51:51]);
  OR2 I497 (comp0_0[52:52], wg_0r0[52:52], wg_0r1[52:52]);
  OR2 I498 (comp0_0[53:53], wg_0r0[53:53], wg_0r1[53:53]);
  OR2 I499 (comp0_0[54:54], wg_0r0[54:54], wg_0r1[54:54]);
  OR2 I500 (comp0_0[55:55], wg_0r0[55:55], wg_0r1[55:55]);
  OR2 I501 (comp0_0[56:56], wg_0r0[56:56], wg_0r1[56:56]);
  OR2 I502 (comp0_0[57:57], wg_0r0[57:57], wg_0r1[57:57]);
  OR2 I503 (comp0_0[58:58], wg_0r0[58:58], wg_0r1[58:58]);
  OR2 I504 (comp0_0[59:59], wg_0r0[59:59], wg_0r1[59:59]);
  OR2 I505 (comp0_0[60:60], wg_0r0[60:60], wg_0r1[60:60]);
  OR2 I506 (comp0_0[61:61], wg_0r0[61:61], wg_0r1[61:61]);
  OR2 I507 (comp0_0[62:62], wg_0r0[62:62], wg_0r1[62:62]);
  OR2 I508 (comp0_0[63:63], wg_0r0[63:63], wg_0r1[63:63]);
  OR2 I509 (comp0_0[64:64], wg_0r0[64:64], wg_0r1[64:64]);
  OR2 I510 (comp0_0[65:65], wg_0r0[65:65], wg_0r1[65:65]);
  OR2 I511 (comp0_0[66:66], wg_0r0[66:66], wg_0r1[66:66]);
  OR2 I512 (comp0_0[67:67], wg_0r0[67:67], wg_0r1[67:67]);
  OR2 I513 (comp0_0[68:68], wg_0r0[68:68], wg_0r1[68:68]);
  OR2 I514 (comp0_0[69:69], wg_0r0[69:69], wg_0r1[69:69]);
  OR2 I515 (comp0_0[70:70], wg_0r0[70:70], wg_0r1[70:70]);
  OR2 I516 (comp0_0[71:71], wg_0r0[71:71], wg_0r1[71:71]);
  OR2 I517 (comp0_0[72:72], wg_0r0[72:72], wg_0r1[72:72]);
  OR2 I518 (comp0_0[73:73], wg_0r0[73:73], wg_0r1[73:73]);
  C3 I519 (simp5321_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I520 (simp5321_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I521 (simp5321_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I522 (simp5321_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I523 (simp5321_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I524 (simp5321_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I525 (simp5321_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I526 (simp5321_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I527 (simp5321_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I528 (simp5321_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C3 I529 (simp5321_0[10:10], comp0_0[30:30], comp0_0[31:31], comp0_0[32:32]);
  C3 I530 (simp5321_0[11:11], comp0_0[33:33], comp0_0[34:34], comp0_0[35:35]);
  C3 I531 (simp5321_0[12:12], comp0_0[36:36], comp0_0[37:37], comp0_0[38:38]);
  C3 I532 (simp5321_0[13:13], comp0_0[39:39], comp0_0[40:40], comp0_0[41:41]);
  C3 I533 (simp5321_0[14:14], comp0_0[42:42], comp0_0[43:43], comp0_0[44:44]);
  C3 I534 (simp5321_0[15:15], comp0_0[45:45], comp0_0[46:46], comp0_0[47:47]);
  C3 I535 (simp5321_0[16:16], comp0_0[48:48], comp0_0[49:49], comp0_0[50:50]);
  C3 I536 (simp5321_0[17:17], comp0_0[51:51], comp0_0[52:52], comp0_0[53:53]);
  C3 I537 (simp5321_0[18:18], comp0_0[54:54], comp0_0[55:55], comp0_0[56:56]);
  C3 I538 (simp5321_0[19:19], comp0_0[57:57], comp0_0[58:58], comp0_0[59:59]);
  C3 I539 (simp5321_0[20:20], comp0_0[60:60], comp0_0[61:61], comp0_0[62:62]);
  C3 I540 (simp5321_0[21:21], comp0_0[63:63], comp0_0[64:64], comp0_0[65:65]);
  C3 I541 (simp5321_0[22:22], comp0_0[66:66], comp0_0[67:67], comp0_0[68:68]);
  C3 I542 (simp5321_0[23:23], comp0_0[69:69], comp0_0[70:70], comp0_0[71:71]);
  C2 I543 (simp5321_0[24:24], comp0_0[72:72], comp0_0[73:73]);
  C3 I544 (simp5322_0[0:0], simp5321_0[0:0], simp5321_0[1:1], simp5321_0[2:2]);
  C3 I545 (simp5322_0[1:1], simp5321_0[3:3], simp5321_0[4:4], simp5321_0[5:5]);
  C3 I546 (simp5322_0[2:2], simp5321_0[6:6], simp5321_0[7:7], simp5321_0[8:8]);
  C3 I547 (simp5322_0[3:3], simp5321_0[9:9], simp5321_0[10:10], simp5321_0[11:11]);
  C3 I548 (simp5322_0[4:4], simp5321_0[12:12], simp5321_0[13:13], simp5321_0[14:14]);
  C3 I549 (simp5322_0[5:5], simp5321_0[15:15], simp5321_0[16:16], simp5321_0[17:17]);
  C3 I550 (simp5322_0[6:6], simp5321_0[18:18], simp5321_0[19:19], simp5321_0[20:20]);
  C3 I551 (simp5322_0[7:7], simp5321_0[21:21], simp5321_0[22:22], simp5321_0[23:23]);
  BUFF I552 (simp5322_0[8:8], simp5321_0[24:24]);
  C3 I553 (simp5323_0[0:0], simp5322_0[0:0], simp5322_0[1:1], simp5322_0[2:2]);
  C3 I554 (simp5323_0[1:1], simp5322_0[3:3], simp5322_0[4:4], simp5322_0[5:5]);
  C3 I555 (simp5323_0[2:2], simp5322_0[6:6], simp5322_0[7:7], simp5322_0[8:8]);
  C3 I556 (wc_0, simp5323_0[0:0], simp5323_0[1:1], simp5323_0[2:2]);
  AND2 I557 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I558 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I559 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I560 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I561 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I562 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I563 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I564 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I565 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I566 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I567 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I568 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I569 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I570 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I571 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I572 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I573 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I574 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I575 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I576 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I577 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I578 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I579 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I580 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I581 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I582 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I583 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I584 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I585 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I586 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I587 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I588 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I589 (conwgif_0[32:32], wg_0r0[32:32], conwig_0);
  AND2 I590 (conwgif_0[33:33], wg_0r0[33:33], conwig_0);
  AND2 I591 (conwgif_0[34:34], wg_0r0[34:34], conwig_0);
  AND2 I592 (conwgif_0[35:35], wg_0r0[35:35], conwig_0);
  AND2 I593 (conwgif_0[36:36], wg_0r0[36:36], conwig_0);
  AND2 I594 (conwgif_0[37:37], wg_0r0[37:37], conwig_0);
  AND2 I595 (conwgif_0[38:38], wg_0r0[38:38], conwig_0);
  AND2 I596 (conwgif_0[39:39], wg_0r0[39:39], conwig_0);
  AND2 I597 (conwgif_0[40:40], wg_0r0[40:40], conwig_0);
  AND2 I598 (conwgif_0[41:41], wg_0r0[41:41], conwig_0);
  AND2 I599 (conwgif_0[42:42], wg_0r0[42:42], conwig_0);
  AND2 I600 (conwgif_0[43:43], wg_0r0[43:43], conwig_0);
  AND2 I601 (conwgif_0[44:44], wg_0r0[44:44], conwig_0);
  AND2 I602 (conwgif_0[45:45], wg_0r0[45:45], conwig_0);
  AND2 I603 (conwgif_0[46:46], wg_0r0[46:46], conwig_0);
  AND2 I604 (conwgif_0[47:47], wg_0r0[47:47], conwig_0);
  AND2 I605 (conwgif_0[48:48], wg_0r0[48:48], conwig_0);
  AND2 I606 (conwgif_0[49:49], wg_0r0[49:49], conwig_0);
  AND2 I607 (conwgif_0[50:50], wg_0r0[50:50], conwig_0);
  AND2 I608 (conwgif_0[51:51], wg_0r0[51:51], conwig_0);
  AND2 I609 (conwgif_0[52:52], wg_0r0[52:52], conwig_0);
  AND2 I610 (conwgif_0[53:53], wg_0r0[53:53], conwig_0);
  AND2 I611 (conwgif_0[54:54], wg_0r0[54:54], conwig_0);
  AND2 I612 (conwgif_0[55:55], wg_0r0[55:55], conwig_0);
  AND2 I613 (conwgif_0[56:56], wg_0r0[56:56], conwig_0);
  AND2 I614 (conwgif_0[57:57], wg_0r0[57:57], conwig_0);
  AND2 I615 (conwgif_0[58:58], wg_0r0[58:58], conwig_0);
  AND2 I616 (conwgif_0[59:59], wg_0r0[59:59], conwig_0);
  AND2 I617 (conwgif_0[60:60], wg_0r0[60:60], conwig_0);
  AND2 I618 (conwgif_0[61:61], wg_0r0[61:61], conwig_0);
  AND2 I619 (conwgif_0[62:62], wg_0r0[62:62], conwig_0);
  AND2 I620 (conwgif_0[63:63], wg_0r0[63:63], conwig_0);
  AND2 I621 (conwgif_0[64:64], wg_0r0[64:64], conwig_0);
  AND2 I622 (conwgif_0[65:65], wg_0r0[65:65], conwig_0);
  AND2 I623 (conwgif_0[66:66], wg_0r0[66:66], conwig_0);
  AND2 I624 (conwgif_0[67:67], wg_0r0[67:67], conwig_0);
  AND2 I625 (conwgif_0[68:68], wg_0r0[68:68], conwig_0);
  AND2 I626 (conwgif_0[69:69], wg_0r0[69:69], conwig_0);
  AND2 I627 (conwgif_0[70:70], wg_0r0[70:70], conwig_0);
  AND2 I628 (conwgif_0[71:71], wg_0r0[71:71], conwig_0);
  AND2 I629 (conwgif_0[72:72], wg_0r0[72:72], conwig_0);
  AND2 I630 (conwgif_0[73:73], wg_0r0[73:73], conwig_0);
  AND2 I631 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I632 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I633 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I634 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I635 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I636 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I637 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I638 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I639 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I640 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I641 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I642 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I643 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I644 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I645 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I646 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I647 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I648 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I649 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I650 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I651 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I652 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I653 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I654 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I655 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I656 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I657 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I658 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I659 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I660 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I661 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I662 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  AND2 I663 (conwgit_0[32:32], wg_0r1[32:32], conwig_0);
  AND2 I664 (conwgit_0[33:33], wg_0r1[33:33], conwig_0);
  AND2 I665 (conwgit_0[34:34], wg_0r1[34:34], conwig_0);
  AND2 I666 (conwgit_0[35:35], wg_0r1[35:35], conwig_0);
  AND2 I667 (conwgit_0[36:36], wg_0r1[36:36], conwig_0);
  AND2 I668 (conwgit_0[37:37], wg_0r1[37:37], conwig_0);
  AND2 I669 (conwgit_0[38:38], wg_0r1[38:38], conwig_0);
  AND2 I670 (conwgit_0[39:39], wg_0r1[39:39], conwig_0);
  AND2 I671 (conwgit_0[40:40], wg_0r1[40:40], conwig_0);
  AND2 I672 (conwgit_0[41:41], wg_0r1[41:41], conwig_0);
  AND2 I673 (conwgit_0[42:42], wg_0r1[42:42], conwig_0);
  AND2 I674 (conwgit_0[43:43], wg_0r1[43:43], conwig_0);
  AND2 I675 (conwgit_0[44:44], wg_0r1[44:44], conwig_0);
  AND2 I676 (conwgit_0[45:45], wg_0r1[45:45], conwig_0);
  AND2 I677 (conwgit_0[46:46], wg_0r1[46:46], conwig_0);
  AND2 I678 (conwgit_0[47:47], wg_0r1[47:47], conwig_0);
  AND2 I679 (conwgit_0[48:48], wg_0r1[48:48], conwig_0);
  AND2 I680 (conwgit_0[49:49], wg_0r1[49:49], conwig_0);
  AND2 I681 (conwgit_0[50:50], wg_0r1[50:50], conwig_0);
  AND2 I682 (conwgit_0[51:51], wg_0r1[51:51], conwig_0);
  AND2 I683 (conwgit_0[52:52], wg_0r1[52:52], conwig_0);
  AND2 I684 (conwgit_0[53:53], wg_0r1[53:53], conwig_0);
  AND2 I685 (conwgit_0[54:54], wg_0r1[54:54], conwig_0);
  AND2 I686 (conwgit_0[55:55], wg_0r1[55:55], conwig_0);
  AND2 I687 (conwgit_0[56:56], wg_0r1[56:56], conwig_0);
  AND2 I688 (conwgit_0[57:57], wg_0r1[57:57], conwig_0);
  AND2 I689 (conwgit_0[58:58], wg_0r1[58:58], conwig_0);
  AND2 I690 (conwgit_0[59:59], wg_0r1[59:59], conwig_0);
  AND2 I691 (conwgit_0[60:60], wg_0r1[60:60], conwig_0);
  AND2 I692 (conwgit_0[61:61], wg_0r1[61:61], conwig_0);
  AND2 I693 (conwgit_0[62:62], wg_0r1[62:62], conwig_0);
  AND2 I694 (conwgit_0[63:63], wg_0r1[63:63], conwig_0);
  AND2 I695 (conwgit_0[64:64], wg_0r1[64:64], conwig_0);
  AND2 I696 (conwgit_0[65:65], wg_0r1[65:65], conwig_0);
  AND2 I697 (conwgit_0[66:66], wg_0r1[66:66], conwig_0);
  AND2 I698 (conwgit_0[67:67], wg_0r1[67:67], conwig_0);
  AND2 I699 (conwgit_0[68:68], wg_0r1[68:68], conwig_0);
  AND2 I700 (conwgit_0[69:69], wg_0r1[69:69], conwig_0);
  AND2 I701 (conwgit_0[70:70], wg_0r1[70:70], conwig_0);
  AND2 I702 (conwgit_0[71:71], wg_0r1[71:71], conwig_0);
  AND2 I703 (conwgit_0[72:72], wg_0r1[72:72], conwig_0);
  AND2 I704 (conwgit_0[73:73], wg_0r1[73:73], conwig_0);
  BUFF I705 (conwigc_0, wc_0);
  AO22 I706 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I707 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I708 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I709 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I710 (wenr_0[0:0], wc_0);
  BUFF I711 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I712 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I713 (wenr_0[1:1], wc_0);
  BUFF I714 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I715 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I716 (wenr_0[2:2], wc_0);
  BUFF I717 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I718 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I719 (wenr_0[3:3], wc_0);
  BUFF I720 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I721 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I722 (wenr_0[4:4], wc_0);
  BUFF I723 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I724 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I725 (wenr_0[5:5], wc_0);
  BUFF I726 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I727 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I728 (wenr_0[6:6], wc_0);
  BUFF I729 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I730 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I731 (wenr_0[7:7], wc_0);
  BUFF I732 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I733 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I734 (wenr_0[8:8], wc_0);
  BUFF I735 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I736 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I737 (wenr_0[9:9], wc_0);
  BUFF I738 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I739 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I740 (wenr_0[10:10], wc_0);
  BUFF I741 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I742 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I743 (wenr_0[11:11], wc_0);
  BUFF I744 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I745 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I746 (wenr_0[12:12], wc_0);
  BUFF I747 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I748 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I749 (wenr_0[13:13], wc_0);
  BUFF I750 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I751 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I752 (wenr_0[14:14], wc_0);
  BUFF I753 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I754 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I755 (wenr_0[15:15], wc_0);
  BUFF I756 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I757 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I758 (wenr_0[16:16], wc_0);
  BUFF I759 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I760 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I761 (wenr_0[17:17], wc_0);
  BUFF I762 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I763 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I764 (wenr_0[18:18], wc_0);
  BUFF I765 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I766 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I767 (wenr_0[19:19], wc_0);
  BUFF I768 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I769 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I770 (wenr_0[20:20], wc_0);
  BUFF I771 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I772 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I773 (wenr_0[21:21], wc_0);
  BUFF I774 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I775 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I776 (wenr_0[22:22], wc_0);
  BUFF I777 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I778 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I779 (wenr_0[23:23], wc_0);
  BUFF I780 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I781 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I782 (wenr_0[24:24], wc_0);
  BUFF I783 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I784 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I785 (wenr_0[25:25], wc_0);
  BUFF I786 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I787 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I788 (wenr_0[26:26], wc_0);
  BUFF I789 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I790 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I791 (wenr_0[27:27], wc_0);
  BUFF I792 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I793 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I794 (wenr_0[28:28], wc_0);
  BUFF I795 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I796 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I797 (wenr_0[29:29], wc_0);
  BUFF I798 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I799 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I800 (wenr_0[30:30], wc_0);
  BUFF I801 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I802 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I803 (wenr_0[31:31], wc_0);
  BUFF I804 (wf_0[32:32], conwgif_0[32:32]);
  BUFF I805 (wt_0[32:32], conwgit_0[32:32]);
  BUFF I806 (wenr_0[32:32], wc_0);
  BUFF I807 (wf_0[33:33], conwgif_0[33:33]);
  BUFF I808 (wt_0[33:33], conwgit_0[33:33]);
  BUFF I809 (wenr_0[33:33], wc_0);
  BUFF I810 (wf_0[34:34], conwgif_0[34:34]);
  BUFF I811 (wt_0[34:34], conwgit_0[34:34]);
  BUFF I812 (wenr_0[34:34], wc_0);
  BUFF I813 (wf_0[35:35], conwgif_0[35:35]);
  BUFF I814 (wt_0[35:35], conwgit_0[35:35]);
  BUFF I815 (wenr_0[35:35], wc_0);
  BUFF I816 (wf_0[36:36], conwgif_0[36:36]);
  BUFF I817 (wt_0[36:36], conwgit_0[36:36]);
  BUFF I818 (wenr_0[36:36], wc_0);
  BUFF I819 (wf_0[37:37], conwgif_0[37:37]);
  BUFF I820 (wt_0[37:37], conwgit_0[37:37]);
  BUFF I821 (wenr_0[37:37], wc_0);
  BUFF I822 (wf_0[38:38], conwgif_0[38:38]);
  BUFF I823 (wt_0[38:38], conwgit_0[38:38]);
  BUFF I824 (wenr_0[38:38], wc_0);
  BUFF I825 (wf_0[39:39], conwgif_0[39:39]);
  BUFF I826 (wt_0[39:39], conwgit_0[39:39]);
  BUFF I827 (wenr_0[39:39], wc_0);
  BUFF I828 (wf_0[40:40], conwgif_0[40:40]);
  BUFF I829 (wt_0[40:40], conwgit_0[40:40]);
  BUFF I830 (wenr_0[40:40], wc_0);
  BUFF I831 (wf_0[41:41], conwgif_0[41:41]);
  BUFF I832 (wt_0[41:41], conwgit_0[41:41]);
  BUFF I833 (wenr_0[41:41], wc_0);
  BUFF I834 (wf_0[42:42], conwgif_0[42:42]);
  BUFF I835 (wt_0[42:42], conwgit_0[42:42]);
  BUFF I836 (wenr_0[42:42], wc_0);
  BUFF I837 (wf_0[43:43], conwgif_0[43:43]);
  BUFF I838 (wt_0[43:43], conwgit_0[43:43]);
  BUFF I839 (wenr_0[43:43], wc_0);
  BUFF I840 (wf_0[44:44], conwgif_0[44:44]);
  BUFF I841 (wt_0[44:44], conwgit_0[44:44]);
  BUFF I842 (wenr_0[44:44], wc_0);
  BUFF I843 (wf_0[45:45], conwgif_0[45:45]);
  BUFF I844 (wt_0[45:45], conwgit_0[45:45]);
  BUFF I845 (wenr_0[45:45], wc_0);
  BUFF I846 (wf_0[46:46], conwgif_0[46:46]);
  BUFF I847 (wt_0[46:46], conwgit_0[46:46]);
  BUFF I848 (wenr_0[46:46], wc_0);
  BUFF I849 (wf_0[47:47], conwgif_0[47:47]);
  BUFF I850 (wt_0[47:47], conwgit_0[47:47]);
  BUFF I851 (wenr_0[47:47], wc_0);
  BUFF I852 (wf_0[48:48], conwgif_0[48:48]);
  BUFF I853 (wt_0[48:48], conwgit_0[48:48]);
  BUFF I854 (wenr_0[48:48], wc_0);
  BUFF I855 (wf_0[49:49], conwgif_0[49:49]);
  BUFF I856 (wt_0[49:49], conwgit_0[49:49]);
  BUFF I857 (wenr_0[49:49], wc_0);
  BUFF I858 (wf_0[50:50], conwgif_0[50:50]);
  BUFF I859 (wt_0[50:50], conwgit_0[50:50]);
  BUFF I860 (wenr_0[50:50], wc_0);
  BUFF I861 (wf_0[51:51], conwgif_0[51:51]);
  BUFF I862 (wt_0[51:51], conwgit_0[51:51]);
  BUFF I863 (wenr_0[51:51], wc_0);
  BUFF I864 (wf_0[52:52], conwgif_0[52:52]);
  BUFF I865 (wt_0[52:52], conwgit_0[52:52]);
  BUFF I866 (wenr_0[52:52], wc_0);
  BUFF I867 (wf_0[53:53], conwgif_0[53:53]);
  BUFF I868 (wt_0[53:53], conwgit_0[53:53]);
  BUFF I869 (wenr_0[53:53], wc_0);
  BUFF I870 (wf_0[54:54], conwgif_0[54:54]);
  BUFF I871 (wt_0[54:54], conwgit_0[54:54]);
  BUFF I872 (wenr_0[54:54], wc_0);
  BUFF I873 (wf_0[55:55], conwgif_0[55:55]);
  BUFF I874 (wt_0[55:55], conwgit_0[55:55]);
  BUFF I875 (wenr_0[55:55], wc_0);
  BUFF I876 (wf_0[56:56], conwgif_0[56:56]);
  BUFF I877 (wt_0[56:56], conwgit_0[56:56]);
  BUFF I878 (wenr_0[56:56], wc_0);
  BUFF I879 (wf_0[57:57], conwgif_0[57:57]);
  BUFF I880 (wt_0[57:57], conwgit_0[57:57]);
  BUFF I881 (wenr_0[57:57], wc_0);
  BUFF I882 (wf_0[58:58], conwgif_0[58:58]);
  BUFF I883 (wt_0[58:58], conwgit_0[58:58]);
  BUFF I884 (wenr_0[58:58], wc_0);
  BUFF I885 (wf_0[59:59], conwgif_0[59:59]);
  BUFF I886 (wt_0[59:59], conwgit_0[59:59]);
  BUFF I887 (wenr_0[59:59], wc_0);
  BUFF I888 (wf_0[60:60], conwgif_0[60:60]);
  BUFF I889 (wt_0[60:60], conwgit_0[60:60]);
  BUFF I890 (wenr_0[60:60], wc_0);
  BUFF I891 (wf_0[61:61], conwgif_0[61:61]);
  BUFF I892 (wt_0[61:61], conwgit_0[61:61]);
  BUFF I893 (wenr_0[61:61], wc_0);
  BUFF I894 (wf_0[62:62], conwgif_0[62:62]);
  BUFF I895 (wt_0[62:62], conwgit_0[62:62]);
  BUFF I896 (wenr_0[62:62], wc_0);
  BUFF I897 (wf_0[63:63], conwgif_0[63:63]);
  BUFF I898 (wt_0[63:63], conwgit_0[63:63]);
  BUFF I899 (wenr_0[63:63], wc_0);
  BUFF I900 (wf_0[64:64], conwgif_0[64:64]);
  BUFF I901 (wt_0[64:64], conwgit_0[64:64]);
  BUFF I902 (wenr_0[64:64], wc_0);
  BUFF I903 (wf_0[65:65], conwgif_0[65:65]);
  BUFF I904 (wt_0[65:65], conwgit_0[65:65]);
  BUFF I905 (wenr_0[65:65], wc_0);
  BUFF I906 (wf_0[66:66], conwgif_0[66:66]);
  BUFF I907 (wt_0[66:66], conwgit_0[66:66]);
  BUFF I908 (wenr_0[66:66], wc_0);
  BUFF I909 (wf_0[67:67], conwgif_0[67:67]);
  BUFF I910 (wt_0[67:67], conwgit_0[67:67]);
  BUFF I911 (wenr_0[67:67], wc_0);
  BUFF I912 (wf_0[68:68], conwgif_0[68:68]);
  BUFF I913 (wt_0[68:68], conwgit_0[68:68]);
  BUFF I914 (wenr_0[68:68], wc_0);
  BUFF I915 (wf_0[69:69], conwgif_0[69:69]);
  BUFF I916 (wt_0[69:69], conwgit_0[69:69]);
  BUFF I917 (wenr_0[69:69], wc_0);
  BUFF I918 (wf_0[70:70], conwgif_0[70:70]);
  BUFF I919 (wt_0[70:70], conwgit_0[70:70]);
  BUFF I920 (wenr_0[70:70], wc_0);
  BUFF I921 (wf_0[71:71], conwgif_0[71:71]);
  BUFF I922 (wt_0[71:71], conwgit_0[71:71]);
  BUFF I923 (wenr_0[71:71], wc_0);
  BUFF I924 (wf_0[72:72], conwgif_0[72:72]);
  BUFF I925 (wt_0[72:72], conwgit_0[72:72]);
  BUFF I926 (wenr_0[72:72], wc_0);
  BUFF I927 (wf_0[73:73], conwgif_0[73:73]);
  BUFF I928 (wt_0[73:73], conwgit_0[73:73]);
  BUFF I929 (wenr_0[73:73], wc_0);
  C3 I930 (simp9111_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I931 (simp9111_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I932 (simp9111_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I933 (simp9111_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I934 (simp9111_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I935 (simp9111_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I936 (simp9111_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I937 (simp9111_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I938 (simp9111_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I939 (simp9111_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I940 (simp9111_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I941 (simp9111_0[11:11], wacks_0[32:32], wacks_0[33:33], wacks_0[34:34]);
  C3 I942 (simp9111_0[12:12], wacks_0[35:35], wacks_0[36:36], wacks_0[37:37]);
  C3 I943 (simp9111_0[13:13], wacks_0[38:38], wacks_0[39:39], wacks_0[40:40]);
  C3 I944 (simp9111_0[14:14], wacks_0[41:41], wacks_0[42:42], wacks_0[43:43]);
  C3 I945 (simp9111_0[15:15], wacks_0[44:44], wacks_0[45:45], wacks_0[46:46]);
  C3 I946 (simp9111_0[16:16], wacks_0[47:47], wacks_0[48:48], wacks_0[49:49]);
  C3 I947 (simp9111_0[17:17], wacks_0[50:50], wacks_0[51:51], wacks_0[52:52]);
  C3 I948 (simp9111_0[18:18], wacks_0[53:53], wacks_0[54:54], wacks_0[55:55]);
  C3 I949 (simp9111_0[19:19], wacks_0[56:56], wacks_0[57:57], wacks_0[58:58]);
  C3 I950 (simp9111_0[20:20], wacks_0[59:59], wacks_0[60:60], wacks_0[61:61]);
  C3 I951 (simp9111_0[21:21], wacks_0[62:62], wacks_0[63:63], wacks_0[64:64]);
  C3 I952 (simp9111_0[22:22], wacks_0[65:65], wacks_0[66:66], wacks_0[67:67]);
  C3 I953 (simp9111_0[23:23], wacks_0[68:68], wacks_0[69:69], wacks_0[70:70]);
  C3 I954 (simp9111_0[24:24], wacks_0[71:71], wacks_0[72:72], wacks_0[73:73]);
  C3 I955 (simp9112_0[0:0], simp9111_0[0:0], simp9111_0[1:1], simp9111_0[2:2]);
  C3 I956 (simp9112_0[1:1], simp9111_0[3:3], simp9111_0[4:4], simp9111_0[5:5]);
  C3 I957 (simp9112_0[2:2], simp9111_0[6:6], simp9111_0[7:7], simp9111_0[8:8]);
  C3 I958 (simp9112_0[3:3], simp9111_0[9:9], simp9111_0[10:10], simp9111_0[11:11]);
  C3 I959 (simp9112_0[4:4], simp9111_0[12:12], simp9111_0[13:13], simp9111_0[14:14]);
  C3 I960 (simp9112_0[5:5], simp9111_0[15:15], simp9111_0[16:16], simp9111_0[17:17]);
  C3 I961 (simp9112_0[6:6], simp9111_0[18:18], simp9111_0[19:19], simp9111_0[20:20]);
  C3 I962 (simp9112_0[7:7], simp9111_0[21:21], simp9111_0[22:22], simp9111_0[23:23]);
  BUFF I963 (simp9112_0[8:8], simp9111_0[24:24]);
  C3 I964 (simp9113_0[0:0], simp9112_0[0:0], simp9112_0[1:1], simp9112_0[2:2]);
  C3 I965 (simp9113_0[1:1], simp9112_0[3:3], simp9112_0[4:4], simp9112_0[5:5]);
  C3 I966 (simp9113_0[2:2], simp9112_0[6:6], simp9112_0[7:7], simp9112_0[8:8]);
  C3 I967 (wd_0r, simp9113_0[0:0], simp9113_0[1:1], simp9113_0[2:2]);
  AND2 I968 (rd_0r0[0:0], df_0[26:26], rg_0r);
  AND2 I969 (rd_0r0[1:1], df_0[27:27], rg_0r);
  AND2 I970 (rd_0r0[2:2], df_0[28:28], rg_0r);
  AND2 I971 (rd_0r0[3:3], df_0[29:29], rg_0r);
  AND2 I972 (rd_0r0[4:4], df_0[30:30], rg_0r);
  AND2 I973 (rd_1r0, df_0[25:25], rg_1r);
  AND2 I974 (rd_2r0, df_0[25:25], rg_2r);
  AND2 I975 (rd_3r0[0:0], df_0[20:20], rg_3r);
  AND2 I976 (rd_3r0[1:1], df_0[21:21], rg_3r);
  AND2 I977 (rd_3r0[2:2], df_0[22:22], rg_3r);
  AND2 I978 (rd_3r0[3:3], df_0[23:23], rg_3r);
  AND2 I979 (rd_3r0[4:4], df_0[24:24], rg_3r);
  AND2 I980 (rd_4r0, df_0[9:9], rg_4r);
  AND2 I981 (rd_5r0[0:0], df_0[15:15], rg_5r);
  AND2 I982 (rd_5r0[1:1], df_0[16:16], rg_5r);
  AND2 I983 (rd_5r0[2:2], df_0[17:17], rg_5r);
  AND2 I984 (rd_5r0[3:3], df_0[18:18], rg_5r);
  AND2 I985 (rd_5r0[4:4], df_0[19:19], rg_5r);
  AND2 I986 (rd_6r0, df_0[8:8], rg_6r);
  AND2 I987 (rd_7r0[0:0], df_0[10:10], rg_7r);
  AND2 I988 (rd_7r0[1:1], df_0[11:11], rg_7r);
  AND2 I989 (rd_7r0[2:2], df_0[12:12], rg_7r);
  AND2 I990 (rd_7r0[3:3], df_0[13:13], rg_7r);
  AND2 I991 (rd_7r0[4:4], df_0[14:14], rg_7r);
  AND2 I992 (rd_8r0, df_0[7:7], rg_8r);
  AND2 I993 (rd_9r0[0:0], df_0[7:7], rg_9r);
  AND2 I994 (rd_9r0[1:1], df_0[8:8], rg_9r);
  AND2 I995 (rd_9r0[2:2], df_0[9:9], rg_9r);
  AND2 I996 (rd_10r0[0:0], df_0[38:38], rg_10r);
  AND2 I997 (rd_10r0[1:1], df_0[39:39], rg_10r);
  AND2 I998 (rd_10r0[2:2], df_0[40:40], rg_10r);
  AND2 I999 (rd_10r0[3:3], df_0[41:41], rg_10r);
  AND2 I1000 (rd_10r0[4:4], df_0[42:42], rg_10r);
  AND2 I1001 (rd_10r0[5:5], df_0[43:43], rg_10r);
  AND2 I1002 (rd_10r0[6:6], df_0[44:44], rg_10r);
  AND2 I1003 (rd_10r0[7:7], df_0[45:45], rg_10r);
  AND2 I1004 (rd_10r0[8:8], df_0[46:46], rg_10r);
  AND2 I1005 (rd_10r0[9:9], df_0[47:47], rg_10r);
  AND2 I1006 (rd_10r0[10:10], df_0[48:48], rg_10r);
  AND2 I1007 (rd_10r0[11:11], df_0[49:49], rg_10r);
  AND2 I1008 (rd_10r0[12:12], df_0[50:50], rg_10r);
  AND2 I1009 (rd_10r0[13:13], df_0[51:51], rg_10r);
  AND2 I1010 (rd_10r0[14:14], df_0[52:52], rg_10r);
  AND2 I1011 (rd_10r0[15:15], df_0[53:53], rg_10r);
  AND2 I1012 (rd_10r0[16:16], df_0[54:54], rg_10r);
  AND2 I1013 (rd_10r0[17:17], df_0[55:55], rg_10r);
  AND2 I1014 (rd_10r0[18:18], df_0[56:56], rg_10r);
  AND2 I1015 (rd_10r0[19:19], df_0[57:57], rg_10r);
  AND2 I1016 (rd_10r0[20:20], df_0[58:58], rg_10r);
  AND2 I1017 (rd_10r0[21:21], df_0[59:59], rg_10r);
  AND2 I1018 (rd_10r0[22:22], df_0[60:60], rg_10r);
  AND2 I1019 (rd_10r0[23:23], df_0[61:61], rg_10r);
  AND2 I1020 (rd_10r0[24:24], df_0[62:62], rg_10r);
  AND2 I1021 (rd_10r0[25:25], df_0[63:63], rg_10r);
  AND2 I1022 (rd_10r0[26:26], df_0[64:64], rg_10r);
  AND2 I1023 (rd_10r0[27:27], df_0[65:65], rg_10r);
  AND2 I1024 (rd_10r0[28:28], df_0[66:66], rg_10r);
  AND2 I1025 (rd_10r0[29:29], df_0[67:67], rg_10r);
  AND2 I1026 (rd_10r0[30:30], df_0[68:68], rg_10r);
  AND2 I1027 (rd_10r0[31:31], df_0[69:69], rg_10r);
  AND2 I1028 (rd_11r0, df_0[37:37], rg_11r);
  AND2 I1029 (rd_12r0[0:0], df_0[71:71], rg_12r);
  AND2 I1030 (rd_12r0[1:1], df_0[72:72], rg_12r);
  AND2 I1031 (rd_13r0[0:0], df_0[71:71], rg_13r);
  AND2 I1032 (rd_13r0[1:1], df_0[72:72], rg_13r);
  AND2 I1033 (rd_14r0, df_0[25:25], rg_14r);
  AND2 I1034 (rd_15r0[0:0], df_0[31:31], rg_15r);
  AND2 I1035 (rd_15r0[1:1], df_0[32:32], rg_15r);
  AND2 I1036 (rd_15r0[2:2], df_0[33:33], rg_15r);
  AND2 I1037 (rd_15r0[3:3], df_0[34:34], rg_15r);
  AND2 I1038 (rd_15r0[4:4], df_0[35:35], rg_15r);
  AND2 I1039 (rd_15r0[5:5], df_0[36:36], rg_15r);
  AND2 I1040 (rd_16r0[0:0], df_0[38:38], rg_16r);
  AND2 I1041 (rd_16r0[1:1], df_0[39:39], rg_16r);
  AND2 I1042 (rd_16r0[2:2], df_0[40:40], rg_16r);
  AND2 I1043 (rd_16r0[3:3], df_0[41:41], rg_16r);
  AND2 I1044 (rd_16r0[4:4], df_0[42:42], rg_16r);
  AND2 I1045 (rd_16r0[5:5], df_0[43:43], rg_16r);
  AND2 I1046 (rd_16r0[6:6], df_0[44:44], rg_16r);
  AND2 I1047 (rd_16r0[7:7], df_0[45:45], rg_16r);
  AND2 I1048 (rd_16r0[8:8], df_0[46:46], rg_16r);
  AND2 I1049 (rd_16r0[9:9], df_0[47:47], rg_16r);
  AND2 I1050 (rd_16r0[10:10], df_0[48:48], rg_16r);
  AND2 I1051 (rd_16r0[11:11], df_0[49:49], rg_16r);
  AND2 I1052 (rd_16r0[12:12], df_0[50:50], rg_16r);
  AND2 I1053 (rd_16r0[13:13], df_0[51:51], rg_16r);
  AND2 I1054 (rd_16r0[14:14], df_0[52:52], rg_16r);
  AND2 I1055 (rd_16r0[15:15], df_0[53:53], rg_16r);
  AND2 I1056 (rd_16r0[16:16], df_0[54:54], rg_16r);
  AND2 I1057 (rd_16r0[17:17], df_0[55:55], rg_16r);
  AND2 I1058 (rd_16r0[18:18], df_0[56:56], rg_16r);
  AND2 I1059 (rd_16r0[19:19], df_0[57:57], rg_16r);
  AND2 I1060 (rd_16r0[20:20], df_0[58:58], rg_16r);
  AND2 I1061 (rd_16r0[21:21], df_0[59:59], rg_16r);
  AND2 I1062 (rd_16r0[22:22], df_0[60:60], rg_16r);
  AND2 I1063 (rd_16r0[23:23], df_0[61:61], rg_16r);
  AND2 I1064 (rd_16r0[24:24], df_0[62:62], rg_16r);
  AND2 I1065 (rd_16r0[25:25], df_0[63:63], rg_16r);
  AND2 I1066 (rd_16r0[26:26], df_0[64:64], rg_16r);
  AND2 I1067 (rd_16r0[27:27], df_0[65:65], rg_16r);
  AND2 I1068 (rd_16r0[28:28], df_0[66:66], rg_16r);
  AND2 I1069 (rd_16r0[29:29], df_0[67:67], rg_16r);
  AND2 I1070 (rd_16r0[30:30], df_0[68:68], rg_16r);
  AND2 I1071 (rd_16r0[31:31], df_0[69:69], rg_16r);
  AND2 I1072 (rd_17r0, df_0[6:6], rg_17r);
  AND2 I1073 (rd_18r0[0:0], df_0[3:3], rg_18r);
  AND2 I1074 (rd_18r0[1:1], df_0[4:4], rg_18r);
  AND2 I1075 (rd_18r0[2:2], df_0[5:5], rg_18r);
  AND2 I1076 (rd_18r0[3:3], df_0[6:6], rg_18r);
  AND2 I1077 (rd_19r0[0:0], df_0[0:0], rg_19r);
  AND2 I1078 (rd_19r0[1:1], df_0[1:1], rg_19r);
  AND2 I1079 (rd_19r0[2:2], df_0[2:2], rg_19r);
  AND2 I1080 (rd_0r1[0:0], dt_0[26:26], rg_0r);
  AND2 I1081 (rd_0r1[1:1], dt_0[27:27], rg_0r);
  AND2 I1082 (rd_0r1[2:2], dt_0[28:28], rg_0r);
  AND2 I1083 (rd_0r1[3:3], dt_0[29:29], rg_0r);
  AND2 I1084 (rd_0r1[4:4], dt_0[30:30], rg_0r);
  AND2 I1085 (rd_1r1, dt_0[25:25], rg_1r);
  AND2 I1086 (rd_2r1, dt_0[25:25], rg_2r);
  AND2 I1087 (rd_3r1[0:0], dt_0[20:20], rg_3r);
  AND2 I1088 (rd_3r1[1:1], dt_0[21:21], rg_3r);
  AND2 I1089 (rd_3r1[2:2], dt_0[22:22], rg_3r);
  AND2 I1090 (rd_3r1[3:3], dt_0[23:23], rg_3r);
  AND2 I1091 (rd_3r1[4:4], dt_0[24:24], rg_3r);
  AND2 I1092 (rd_4r1, dt_0[9:9], rg_4r);
  AND2 I1093 (rd_5r1[0:0], dt_0[15:15], rg_5r);
  AND2 I1094 (rd_5r1[1:1], dt_0[16:16], rg_5r);
  AND2 I1095 (rd_5r1[2:2], dt_0[17:17], rg_5r);
  AND2 I1096 (rd_5r1[3:3], dt_0[18:18], rg_5r);
  AND2 I1097 (rd_5r1[4:4], dt_0[19:19], rg_5r);
  AND2 I1098 (rd_6r1, dt_0[8:8], rg_6r);
  AND2 I1099 (rd_7r1[0:0], dt_0[10:10], rg_7r);
  AND2 I1100 (rd_7r1[1:1], dt_0[11:11], rg_7r);
  AND2 I1101 (rd_7r1[2:2], dt_0[12:12], rg_7r);
  AND2 I1102 (rd_7r1[3:3], dt_0[13:13], rg_7r);
  AND2 I1103 (rd_7r1[4:4], dt_0[14:14], rg_7r);
  AND2 I1104 (rd_8r1, dt_0[7:7], rg_8r);
  AND2 I1105 (rd_9r1[0:0], dt_0[7:7], rg_9r);
  AND2 I1106 (rd_9r1[1:1], dt_0[8:8], rg_9r);
  AND2 I1107 (rd_9r1[2:2], dt_0[9:9], rg_9r);
  AND2 I1108 (rd_10r1[0:0], dt_0[38:38], rg_10r);
  AND2 I1109 (rd_10r1[1:1], dt_0[39:39], rg_10r);
  AND2 I1110 (rd_10r1[2:2], dt_0[40:40], rg_10r);
  AND2 I1111 (rd_10r1[3:3], dt_0[41:41], rg_10r);
  AND2 I1112 (rd_10r1[4:4], dt_0[42:42], rg_10r);
  AND2 I1113 (rd_10r1[5:5], dt_0[43:43], rg_10r);
  AND2 I1114 (rd_10r1[6:6], dt_0[44:44], rg_10r);
  AND2 I1115 (rd_10r1[7:7], dt_0[45:45], rg_10r);
  AND2 I1116 (rd_10r1[8:8], dt_0[46:46], rg_10r);
  AND2 I1117 (rd_10r1[9:9], dt_0[47:47], rg_10r);
  AND2 I1118 (rd_10r1[10:10], dt_0[48:48], rg_10r);
  AND2 I1119 (rd_10r1[11:11], dt_0[49:49], rg_10r);
  AND2 I1120 (rd_10r1[12:12], dt_0[50:50], rg_10r);
  AND2 I1121 (rd_10r1[13:13], dt_0[51:51], rg_10r);
  AND2 I1122 (rd_10r1[14:14], dt_0[52:52], rg_10r);
  AND2 I1123 (rd_10r1[15:15], dt_0[53:53], rg_10r);
  AND2 I1124 (rd_10r1[16:16], dt_0[54:54], rg_10r);
  AND2 I1125 (rd_10r1[17:17], dt_0[55:55], rg_10r);
  AND2 I1126 (rd_10r1[18:18], dt_0[56:56], rg_10r);
  AND2 I1127 (rd_10r1[19:19], dt_0[57:57], rg_10r);
  AND2 I1128 (rd_10r1[20:20], dt_0[58:58], rg_10r);
  AND2 I1129 (rd_10r1[21:21], dt_0[59:59], rg_10r);
  AND2 I1130 (rd_10r1[22:22], dt_0[60:60], rg_10r);
  AND2 I1131 (rd_10r1[23:23], dt_0[61:61], rg_10r);
  AND2 I1132 (rd_10r1[24:24], dt_0[62:62], rg_10r);
  AND2 I1133 (rd_10r1[25:25], dt_0[63:63], rg_10r);
  AND2 I1134 (rd_10r1[26:26], dt_0[64:64], rg_10r);
  AND2 I1135 (rd_10r1[27:27], dt_0[65:65], rg_10r);
  AND2 I1136 (rd_10r1[28:28], dt_0[66:66], rg_10r);
  AND2 I1137 (rd_10r1[29:29], dt_0[67:67], rg_10r);
  AND2 I1138 (rd_10r1[30:30], dt_0[68:68], rg_10r);
  AND2 I1139 (rd_10r1[31:31], dt_0[69:69], rg_10r);
  AND2 I1140 (rd_11r1, dt_0[37:37], rg_11r);
  AND2 I1141 (rd_12r1[0:0], dt_0[71:71], rg_12r);
  AND2 I1142 (rd_12r1[1:1], dt_0[72:72], rg_12r);
  AND2 I1143 (rd_13r1[0:0], dt_0[71:71], rg_13r);
  AND2 I1144 (rd_13r1[1:1], dt_0[72:72], rg_13r);
  AND2 I1145 (rd_14r1, dt_0[25:25], rg_14r);
  AND2 I1146 (rd_15r1[0:0], dt_0[31:31], rg_15r);
  AND2 I1147 (rd_15r1[1:1], dt_0[32:32], rg_15r);
  AND2 I1148 (rd_15r1[2:2], dt_0[33:33], rg_15r);
  AND2 I1149 (rd_15r1[3:3], dt_0[34:34], rg_15r);
  AND2 I1150 (rd_15r1[4:4], dt_0[35:35], rg_15r);
  AND2 I1151 (rd_15r1[5:5], dt_0[36:36], rg_15r);
  AND2 I1152 (rd_16r1[0:0], dt_0[38:38], rg_16r);
  AND2 I1153 (rd_16r1[1:1], dt_0[39:39], rg_16r);
  AND2 I1154 (rd_16r1[2:2], dt_0[40:40], rg_16r);
  AND2 I1155 (rd_16r1[3:3], dt_0[41:41], rg_16r);
  AND2 I1156 (rd_16r1[4:4], dt_0[42:42], rg_16r);
  AND2 I1157 (rd_16r1[5:5], dt_0[43:43], rg_16r);
  AND2 I1158 (rd_16r1[6:6], dt_0[44:44], rg_16r);
  AND2 I1159 (rd_16r1[7:7], dt_0[45:45], rg_16r);
  AND2 I1160 (rd_16r1[8:8], dt_0[46:46], rg_16r);
  AND2 I1161 (rd_16r1[9:9], dt_0[47:47], rg_16r);
  AND2 I1162 (rd_16r1[10:10], dt_0[48:48], rg_16r);
  AND2 I1163 (rd_16r1[11:11], dt_0[49:49], rg_16r);
  AND2 I1164 (rd_16r1[12:12], dt_0[50:50], rg_16r);
  AND2 I1165 (rd_16r1[13:13], dt_0[51:51], rg_16r);
  AND2 I1166 (rd_16r1[14:14], dt_0[52:52], rg_16r);
  AND2 I1167 (rd_16r1[15:15], dt_0[53:53], rg_16r);
  AND2 I1168 (rd_16r1[16:16], dt_0[54:54], rg_16r);
  AND2 I1169 (rd_16r1[17:17], dt_0[55:55], rg_16r);
  AND2 I1170 (rd_16r1[18:18], dt_0[56:56], rg_16r);
  AND2 I1171 (rd_16r1[19:19], dt_0[57:57], rg_16r);
  AND2 I1172 (rd_16r1[20:20], dt_0[58:58], rg_16r);
  AND2 I1173 (rd_16r1[21:21], dt_0[59:59], rg_16r);
  AND2 I1174 (rd_16r1[22:22], dt_0[60:60], rg_16r);
  AND2 I1175 (rd_16r1[23:23], dt_0[61:61], rg_16r);
  AND2 I1176 (rd_16r1[24:24], dt_0[62:62], rg_16r);
  AND2 I1177 (rd_16r1[25:25], dt_0[63:63], rg_16r);
  AND2 I1178 (rd_16r1[26:26], dt_0[64:64], rg_16r);
  AND2 I1179 (rd_16r1[27:27], dt_0[65:65], rg_16r);
  AND2 I1180 (rd_16r1[28:28], dt_0[66:66], rg_16r);
  AND2 I1181 (rd_16r1[29:29], dt_0[67:67], rg_16r);
  AND2 I1182 (rd_16r1[30:30], dt_0[68:68], rg_16r);
  AND2 I1183 (rd_16r1[31:31], dt_0[69:69], rg_16r);
  AND2 I1184 (rd_17r1, dt_0[6:6], rg_17r);
  AND2 I1185 (rd_18r1[0:0], dt_0[3:3], rg_18r);
  AND2 I1186 (rd_18r1[1:1], dt_0[4:4], rg_18r);
  AND2 I1187 (rd_18r1[2:2], dt_0[5:5], rg_18r);
  AND2 I1188 (rd_18r1[3:3], dt_0[6:6], rg_18r);
  AND2 I1189 (rd_19r1[0:0], dt_0[0:0], rg_19r);
  AND2 I1190 (rd_19r1[1:1], dt_0[1:1], rg_19r);
  AND2 I1191 (rd_19r1[2:2], dt_0[2:2], rg_19r);
  NOR3 I1192 (simp11361_0[0:0], rg_0r, rg_1r, rg_2r);
  NOR3 I1193 (simp11361_0[1:1], rg_3r, rg_4r, rg_5r);
  NOR3 I1194 (simp11361_0[2:2], rg_6r, rg_7r, rg_8r);
  NOR3 I1195 (simp11361_0[3:3], rg_9r, rg_10r, rg_11r);
  NOR3 I1196 (simp11361_0[4:4], rg_12r, rg_13r, rg_14r);
  NOR3 I1197 (simp11361_0[5:5], rg_15r, rg_16r, rg_17r);
  NOR3 I1198 (simp11361_0[6:6], rg_18r, rg_19r, rg_0a);
  NOR3 I1199 (simp11361_0[7:7], rg_1a, rg_2a, rg_3a);
  NOR3 I1200 (simp11361_0[8:8], rg_4a, rg_5a, rg_6a);
  NOR3 I1201 (simp11361_0[9:9], rg_7a, rg_8a, rg_9a);
  NOR3 I1202 (simp11361_0[10:10], rg_10a, rg_11a, rg_12a);
  NOR3 I1203 (simp11361_0[11:11], rg_13a, rg_14a, rg_15a);
  NOR3 I1204 (simp11361_0[12:12], rg_16a, rg_17a, rg_18a);
  INV I1205 (simp11361_0[13:13], rg_19a);
  NAND3 I1206 (simp11362_0[0:0], simp11361_0[0:0], simp11361_0[1:1], simp11361_0[2:2]);
  NAND3 I1207 (simp11362_0[1:1], simp11361_0[3:3], simp11361_0[4:4], simp11361_0[5:5]);
  NAND3 I1208 (simp11362_0[2:2], simp11361_0[6:6], simp11361_0[7:7], simp11361_0[8:8]);
  NAND3 I1209 (simp11362_0[3:3], simp11361_0[9:9], simp11361_0[10:10], simp11361_0[11:11]);
  NAND2 I1210 (simp11362_0[4:4], simp11361_0[12:12], simp11361_0[13:13]);
  NOR3 I1211 (simp11363_0[0:0], simp11362_0[0:0], simp11362_0[1:1], simp11362_0[2:2]);
  NOR2 I1212 (simp11363_0[1:1], simp11362_0[3:3], simp11362_0[4:4]);
  NAND2 I1213 (anyread_0, simp11363_0[0:0], simp11363_0[1:1]);
  BUFF I1214 (wg_0a, wd_0a);
  BUFF I1215 (rg_0a, rd_0a);
  BUFF I1216 (rg_1a, rd_1a);
  BUFF I1217 (rg_2a, rd_2a);
  BUFF I1218 (rg_3a, rd_3a);
  BUFF I1219 (rg_4a, rd_4a);
  BUFF I1220 (rg_5a, rd_5a);
  BUFF I1221 (rg_6a, rd_6a);
  BUFF I1222 (rg_7a, rd_7a);
  BUFF I1223 (rg_8a, rd_8a);
  BUFF I1224 (rg_9a, rd_9a);
  BUFF I1225 (rg_10a, rd_10a);
  BUFF I1226 (rg_11a, rd_11a);
  BUFF I1227 (rg_12a, rd_12a);
  BUFF I1228 (rg_13a, rd_13a);
  BUFF I1229 (rg_14a, rd_14a);
  BUFF I1230 (rg_15a, rd_15a);
  BUFF I1231 (rg_16a, rd_16a);
  BUFF I1232 (rg_17a, rd_17a);
  BUFF I1233 (rg_18a, rd_18a);
  BUFF I1234 (rg_19a, rd_19a);
endmodule

// tkj74m74_0 TeakJ [Many [74,0],One 74]
module tkj74m74_0 (i_0r0, i_0r1, i_0a, i_1r, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [73:0] i_0r0;
  input [73:0] i_0r1;
  output i_0a;
  input i_1r;
  output i_1a;
  output [73:0] o_0r0;
  output [73:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [73:0] joinf_0;
  wire [73:0] joint_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joinf_0[32:32], i_0r0[32:32]);
  BUFF I33 (joinf_0[33:33], i_0r0[33:33]);
  BUFF I34 (joinf_0[34:34], i_0r0[34:34]);
  BUFF I35 (joinf_0[35:35], i_0r0[35:35]);
  BUFF I36 (joinf_0[36:36], i_0r0[36:36]);
  BUFF I37 (joinf_0[37:37], i_0r0[37:37]);
  BUFF I38 (joinf_0[38:38], i_0r0[38:38]);
  BUFF I39 (joinf_0[39:39], i_0r0[39:39]);
  BUFF I40 (joinf_0[40:40], i_0r0[40:40]);
  BUFF I41 (joinf_0[41:41], i_0r0[41:41]);
  BUFF I42 (joinf_0[42:42], i_0r0[42:42]);
  BUFF I43 (joinf_0[43:43], i_0r0[43:43]);
  BUFF I44 (joinf_0[44:44], i_0r0[44:44]);
  BUFF I45 (joinf_0[45:45], i_0r0[45:45]);
  BUFF I46 (joinf_0[46:46], i_0r0[46:46]);
  BUFF I47 (joinf_0[47:47], i_0r0[47:47]);
  BUFF I48 (joinf_0[48:48], i_0r0[48:48]);
  BUFF I49 (joinf_0[49:49], i_0r0[49:49]);
  BUFF I50 (joinf_0[50:50], i_0r0[50:50]);
  BUFF I51 (joinf_0[51:51], i_0r0[51:51]);
  BUFF I52 (joinf_0[52:52], i_0r0[52:52]);
  BUFF I53 (joinf_0[53:53], i_0r0[53:53]);
  BUFF I54 (joinf_0[54:54], i_0r0[54:54]);
  BUFF I55 (joinf_0[55:55], i_0r0[55:55]);
  BUFF I56 (joinf_0[56:56], i_0r0[56:56]);
  BUFF I57 (joinf_0[57:57], i_0r0[57:57]);
  BUFF I58 (joinf_0[58:58], i_0r0[58:58]);
  BUFF I59 (joinf_0[59:59], i_0r0[59:59]);
  BUFF I60 (joinf_0[60:60], i_0r0[60:60]);
  BUFF I61 (joinf_0[61:61], i_0r0[61:61]);
  BUFF I62 (joinf_0[62:62], i_0r0[62:62]);
  BUFF I63 (joinf_0[63:63], i_0r0[63:63]);
  BUFF I64 (joinf_0[64:64], i_0r0[64:64]);
  BUFF I65 (joinf_0[65:65], i_0r0[65:65]);
  BUFF I66 (joinf_0[66:66], i_0r0[66:66]);
  BUFF I67 (joinf_0[67:67], i_0r0[67:67]);
  BUFF I68 (joinf_0[68:68], i_0r0[68:68]);
  BUFF I69 (joinf_0[69:69], i_0r0[69:69]);
  BUFF I70 (joinf_0[70:70], i_0r0[70:70]);
  BUFF I71 (joinf_0[71:71], i_0r0[71:71]);
  BUFF I72 (joinf_0[72:72], i_0r0[72:72]);
  BUFF I73 (joinf_0[73:73], i_0r0[73:73]);
  BUFF I74 (joint_0[0:0], i_0r1[0:0]);
  BUFF I75 (joint_0[1:1], i_0r1[1:1]);
  BUFF I76 (joint_0[2:2], i_0r1[2:2]);
  BUFF I77 (joint_0[3:3], i_0r1[3:3]);
  BUFF I78 (joint_0[4:4], i_0r1[4:4]);
  BUFF I79 (joint_0[5:5], i_0r1[5:5]);
  BUFF I80 (joint_0[6:6], i_0r1[6:6]);
  BUFF I81 (joint_0[7:7], i_0r1[7:7]);
  BUFF I82 (joint_0[8:8], i_0r1[8:8]);
  BUFF I83 (joint_0[9:9], i_0r1[9:9]);
  BUFF I84 (joint_0[10:10], i_0r1[10:10]);
  BUFF I85 (joint_0[11:11], i_0r1[11:11]);
  BUFF I86 (joint_0[12:12], i_0r1[12:12]);
  BUFF I87 (joint_0[13:13], i_0r1[13:13]);
  BUFF I88 (joint_0[14:14], i_0r1[14:14]);
  BUFF I89 (joint_0[15:15], i_0r1[15:15]);
  BUFF I90 (joint_0[16:16], i_0r1[16:16]);
  BUFF I91 (joint_0[17:17], i_0r1[17:17]);
  BUFF I92 (joint_0[18:18], i_0r1[18:18]);
  BUFF I93 (joint_0[19:19], i_0r1[19:19]);
  BUFF I94 (joint_0[20:20], i_0r1[20:20]);
  BUFF I95 (joint_0[21:21], i_0r1[21:21]);
  BUFF I96 (joint_0[22:22], i_0r1[22:22]);
  BUFF I97 (joint_0[23:23], i_0r1[23:23]);
  BUFF I98 (joint_0[24:24], i_0r1[24:24]);
  BUFF I99 (joint_0[25:25], i_0r1[25:25]);
  BUFF I100 (joint_0[26:26], i_0r1[26:26]);
  BUFF I101 (joint_0[27:27], i_0r1[27:27]);
  BUFF I102 (joint_0[28:28], i_0r1[28:28]);
  BUFF I103 (joint_0[29:29], i_0r1[29:29]);
  BUFF I104 (joint_0[30:30], i_0r1[30:30]);
  BUFF I105 (joint_0[31:31], i_0r1[31:31]);
  BUFF I106 (joint_0[32:32], i_0r1[32:32]);
  BUFF I107 (joint_0[33:33], i_0r1[33:33]);
  BUFF I108 (joint_0[34:34], i_0r1[34:34]);
  BUFF I109 (joint_0[35:35], i_0r1[35:35]);
  BUFF I110 (joint_0[36:36], i_0r1[36:36]);
  BUFF I111 (joint_0[37:37], i_0r1[37:37]);
  BUFF I112 (joint_0[38:38], i_0r1[38:38]);
  BUFF I113 (joint_0[39:39], i_0r1[39:39]);
  BUFF I114 (joint_0[40:40], i_0r1[40:40]);
  BUFF I115 (joint_0[41:41], i_0r1[41:41]);
  BUFF I116 (joint_0[42:42], i_0r1[42:42]);
  BUFF I117 (joint_0[43:43], i_0r1[43:43]);
  BUFF I118 (joint_0[44:44], i_0r1[44:44]);
  BUFF I119 (joint_0[45:45], i_0r1[45:45]);
  BUFF I120 (joint_0[46:46], i_0r1[46:46]);
  BUFF I121 (joint_0[47:47], i_0r1[47:47]);
  BUFF I122 (joint_0[48:48], i_0r1[48:48]);
  BUFF I123 (joint_0[49:49], i_0r1[49:49]);
  BUFF I124 (joint_0[50:50], i_0r1[50:50]);
  BUFF I125 (joint_0[51:51], i_0r1[51:51]);
  BUFF I126 (joint_0[52:52], i_0r1[52:52]);
  BUFF I127 (joint_0[53:53], i_0r1[53:53]);
  BUFF I128 (joint_0[54:54], i_0r1[54:54]);
  BUFF I129 (joint_0[55:55], i_0r1[55:55]);
  BUFF I130 (joint_0[56:56], i_0r1[56:56]);
  BUFF I131 (joint_0[57:57], i_0r1[57:57]);
  BUFF I132 (joint_0[58:58], i_0r1[58:58]);
  BUFF I133 (joint_0[59:59], i_0r1[59:59]);
  BUFF I134 (joint_0[60:60], i_0r1[60:60]);
  BUFF I135 (joint_0[61:61], i_0r1[61:61]);
  BUFF I136 (joint_0[62:62], i_0r1[62:62]);
  BUFF I137 (joint_0[63:63], i_0r1[63:63]);
  BUFF I138 (joint_0[64:64], i_0r1[64:64]);
  BUFF I139 (joint_0[65:65], i_0r1[65:65]);
  BUFF I140 (joint_0[66:66], i_0r1[66:66]);
  BUFF I141 (joint_0[67:67], i_0r1[67:67]);
  BUFF I142 (joint_0[68:68], i_0r1[68:68]);
  BUFF I143 (joint_0[69:69], i_0r1[69:69]);
  BUFF I144 (joint_0[70:70], i_0r1[70:70]);
  BUFF I145 (joint_0[71:71], i_0r1[71:71]);
  BUFF I146 (joint_0[72:72], i_0r1[72:72]);
  BUFF I147 (joint_0[73:73], i_0r1[73:73]);
  BUFF I148 (icomplete_0, i_1r);
  C2 I149 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I150 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I151 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I152 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I153 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I154 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I155 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I156 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I157 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I158 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I159 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I160 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I161 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I162 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I163 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I164 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I165 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I166 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I167 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I168 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I169 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I170 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I171 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I172 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I173 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I174 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I175 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I176 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I177 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I178 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I179 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I180 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I181 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I182 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I183 (o_0r0[33:33], joinf_0[33:33]);
  BUFF I184 (o_0r0[34:34], joinf_0[34:34]);
  BUFF I185 (o_0r0[35:35], joinf_0[35:35]);
  BUFF I186 (o_0r0[36:36], joinf_0[36:36]);
  BUFF I187 (o_0r0[37:37], joinf_0[37:37]);
  BUFF I188 (o_0r0[38:38], joinf_0[38:38]);
  BUFF I189 (o_0r0[39:39], joinf_0[39:39]);
  BUFF I190 (o_0r0[40:40], joinf_0[40:40]);
  BUFF I191 (o_0r0[41:41], joinf_0[41:41]);
  BUFF I192 (o_0r0[42:42], joinf_0[42:42]);
  BUFF I193 (o_0r0[43:43], joinf_0[43:43]);
  BUFF I194 (o_0r0[44:44], joinf_0[44:44]);
  BUFF I195 (o_0r0[45:45], joinf_0[45:45]);
  BUFF I196 (o_0r0[46:46], joinf_0[46:46]);
  BUFF I197 (o_0r0[47:47], joinf_0[47:47]);
  BUFF I198 (o_0r0[48:48], joinf_0[48:48]);
  BUFF I199 (o_0r0[49:49], joinf_0[49:49]);
  BUFF I200 (o_0r0[50:50], joinf_0[50:50]);
  BUFF I201 (o_0r0[51:51], joinf_0[51:51]);
  BUFF I202 (o_0r0[52:52], joinf_0[52:52]);
  BUFF I203 (o_0r0[53:53], joinf_0[53:53]);
  BUFF I204 (o_0r0[54:54], joinf_0[54:54]);
  BUFF I205 (o_0r0[55:55], joinf_0[55:55]);
  BUFF I206 (o_0r0[56:56], joinf_0[56:56]);
  BUFF I207 (o_0r0[57:57], joinf_0[57:57]);
  BUFF I208 (o_0r0[58:58], joinf_0[58:58]);
  BUFF I209 (o_0r0[59:59], joinf_0[59:59]);
  BUFF I210 (o_0r0[60:60], joinf_0[60:60]);
  BUFF I211 (o_0r0[61:61], joinf_0[61:61]);
  BUFF I212 (o_0r0[62:62], joinf_0[62:62]);
  BUFF I213 (o_0r0[63:63], joinf_0[63:63]);
  BUFF I214 (o_0r0[64:64], joinf_0[64:64]);
  BUFF I215 (o_0r0[65:65], joinf_0[65:65]);
  BUFF I216 (o_0r0[66:66], joinf_0[66:66]);
  BUFF I217 (o_0r0[67:67], joinf_0[67:67]);
  BUFF I218 (o_0r0[68:68], joinf_0[68:68]);
  BUFF I219 (o_0r0[69:69], joinf_0[69:69]);
  BUFF I220 (o_0r0[70:70], joinf_0[70:70]);
  BUFF I221 (o_0r0[71:71], joinf_0[71:71]);
  BUFF I222 (o_0r0[72:72], joinf_0[72:72]);
  BUFF I223 (o_0r0[73:73], joinf_0[73:73]);
  BUFF I224 (o_0r1[1:1], joint_0[1:1]);
  BUFF I225 (o_0r1[2:2], joint_0[2:2]);
  BUFF I226 (o_0r1[3:3], joint_0[3:3]);
  BUFF I227 (o_0r1[4:4], joint_0[4:4]);
  BUFF I228 (o_0r1[5:5], joint_0[5:5]);
  BUFF I229 (o_0r1[6:6], joint_0[6:6]);
  BUFF I230 (o_0r1[7:7], joint_0[7:7]);
  BUFF I231 (o_0r1[8:8], joint_0[8:8]);
  BUFF I232 (o_0r1[9:9], joint_0[9:9]);
  BUFF I233 (o_0r1[10:10], joint_0[10:10]);
  BUFF I234 (o_0r1[11:11], joint_0[11:11]);
  BUFF I235 (o_0r1[12:12], joint_0[12:12]);
  BUFF I236 (o_0r1[13:13], joint_0[13:13]);
  BUFF I237 (o_0r1[14:14], joint_0[14:14]);
  BUFF I238 (o_0r1[15:15], joint_0[15:15]);
  BUFF I239 (o_0r1[16:16], joint_0[16:16]);
  BUFF I240 (o_0r1[17:17], joint_0[17:17]);
  BUFF I241 (o_0r1[18:18], joint_0[18:18]);
  BUFF I242 (o_0r1[19:19], joint_0[19:19]);
  BUFF I243 (o_0r1[20:20], joint_0[20:20]);
  BUFF I244 (o_0r1[21:21], joint_0[21:21]);
  BUFF I245 (o_0r1[22:22], joint_0[22:22]);
  BUFF I246 (o_0r1[23:23], joint_0[23:23]);
  BUFF I247 (o_0r1[24:24], joint_0[24:24]);
  BUFF I248 (o_0r1[25:25], joint_0[25:25]);
  BUFF I249 (o_0r1[26:26], joint_0[26:26]);
  BUFF I250 (o_0r1[27:27], joint_0[27:27]);
  BUFF I251 (o_0r1[28:28], joint_0[28:28]);
  BUFF I252 (o_0r1[29:29], joint_0[29:29]);
  BUFF I253 (o_0r1[30:30], joint_0[30:30]);
  BUFF I254 (o_0r1[31:31], joint_0[31:31]);
  BUFF I255 (o_0r1[32:32], joint_0[32:32]);
  BUFF I256 (o_0r1[33:33], joint_0[33:33]);
  BUFF I257 (o_0r1[34:34], joint_0[34:34]);
  BUFF I258 (o_0r1[35:35], joint_0[35:35]);
  BUFF I259 (o_0r1[36:36], joint_0[36:36]);
  BUFF I260 (o_0r1[37:37], joint_0[37:37]);
  BUFF I261 (o_0r1[38:38], joint_0[38:38]);
  BUFF I262 (o_0r1[39:39], joint_0[39:39]);
  BUFF I263 (o_0r1[40:40], joint_0[40:40]);
  BUFF I264 (o_0r1[41:41], joint_0[41:41]);
  BUFF I265 (o_0r1[42:42], joint_0[42:42]);
  BUFF I266 (o_0r1[43:43], joint_0[43:43]);
  BUFF I267 (o_0r1[44:44], joint_0[44:44]);
  BUFF I268 (o_0r1[45:45], joint_0[45:45]);
  BUFF I269 (o_0r1[46:46], joint_0[46:46]);
  BUFF I270 (o_0r1[47:47], joint_0[47:47]);
  BUFF I271 (o_0r1[48:48], joint_0[48:48]);
  BUFF I272 (o_0r1[49:49], joint_0[49:49]);
  BUFF I273 (o_0r1[50:50], joint_0[50:50]);
  BUFF I274 (o_0r1[51:51], joint_0[51:51]);
  BUFF I275 (o_0r1[52:52], joint_0[52:52]);
  BUFF I276 (o_0r1[53:53], joint_0[53:53]);
  BUFF I277 (o_0r1[54:54], joint_0[54:54]);
  BUFF I278 (o_0r1[55:55], joint_0[55:55]);
  BUFF I279 (o_0r1[56:56], joint_0[56:56]);
  BUFF I280 (o_0r1[57:57], joint_0[57:57]);
  BUFF I281 (o_0r1[58:58], joint_0[58:58]);
  BUFF I282 (o_0r1[59:59], joint_0[59:59]);
  BUFF I283 (o_0r1[60:60], joint_0[60:60]);
  BUFF I284 (o_0r1[61:61], joint_0[61:61]);
  BUFF I285 (o_0r1[62:62], joint_0[62:62]);
  BUFF I286 (o_0r1[63:63], joint_0[63:63]);
  BUFF I287 (o_0r1[64:64], joint_0[64:64]);
  BUFF I288 (o_0r1[65:65], joint_0[65:65]);
  BUFF I289 (o_0r1[66:66], joint_0[66:66]);
  BUFF I290 (o_0r1[67:67], joint_0[67:67]);
  BUFF I291 (o_0r1[68:68], joint_0[68:68]);
  BUFF I292 (o_0r1[69:69], joint_0[69:69]);
  BUFF I293 (o_0r1[70:70], joint_0[70:70]);
  BUFF I294 (o_0r1[71:71], joint_0[71:71]);
  BUFF I295 (o_0r1[72:72], joint_0[72:72]);
  BUFF I296 (o_0r1[73:73], joint_0[73:73]);
  BUFF I297 (i_0a, o_0a);
  BUFF I298 (i_1a, o_0a);
endmodule

// tkf7mo0w0_o0w7 TeakF [0,0] [One 7,Many [0,7]]
module tkf7mo0w0_o0w7 (i_0r0, i_0r1, i_0a, o_0r, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [6:0] i_0r0;
  input [6:0] i_0r1;
  output i_0a;
  output o_0r;
  input o_0a;
  output [6:0] o_1r0;
  output [6:0] o_1r1;
  input o_1a;
  input reset;
  wire acomplete_0;
  wire icomplete_0;
  OR2 I0 (icomplete_0, i_0r0[0:0], i_0r1[0:0]);
  BUFF I1 (acomplete_0, icomplete_0);
  BUFF I2 (o_1r0[0:0], i_0r0[0:0]);
  BUFF I3 (o_1r0[1:1], i_0r0[1:1]);
  BUFF I4 (o_1r0[2:2], i_0r0[2:2]);
  BUFF I5 (o_1r0[3:3], i_0r0[3:3]);
  BUFF I6 (o_1r0[4:4], i_0r0[4:4]);
  BUFF I7 (o_1r0[5:5], i_0r0[5:5]);
  BUFF I8 (o_1r0[6:6], i_0r0[6:6]);
  BUFF I9 (o_1r1[0:0], i_0r1[0:0]);
  BUFF I10 (o_1r1[1:1], i_0r1[1:1]);
  BUFF I11 (o_1r1[2:2], i_0r1[2:2]);
  BUFF I12 (o_1r1[3:3], i_0r1[3:3]);
  BUFF I13 (o_1r1[4:4], i_0r1[4:4]);
  BUFF I14 (o_1r1[5:5], i_0r1[5:5]);
  BUFF I15 (o_1r1[6:6], i_0r1[6:6]);
  BUFF I16 (o_0r, icomplete_0);
  C3 I17 (i_0a, acomplete_0, o_0a, o_1a);
endmodule

// tkm3x7b TeakM [Many [7,7,7],One 7]
module tkm3x7b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, i_2r0, i_2r1, i_2a, o_0r0, o_0r1, o_0a, reset);
  input [6:0] i_0r0;
  input [6:0] i_0r1;
  output i_0a;
  input [6:0] i_1r0;
  input [6:0] i_1r1;
  output i_1a;
  input [6:0] i_2r0;
  input [6:0] i_2r1;
  output i_2a;
  output [6:0] o_0r0;
  output [6:0] o_0r1;
  input o_0a;
  input reset;
  wire [6:0] gfint_0;
  wire [6:0] gfint_1;
  wire [6:0] gfint_2;
  wire [6:0] gtint_0;
  wire [6:0] gtint_1;
  wire [6:0] gtint_2;
  wire choice_0;
  wire choice_1;
  wire choice_2;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire icomp_2;
  wire nchosen_0;
  wire [6:0] comp0_0;
  wire [2:0] simp781_0;
  wire [6:0] comp1_0;
  wire [2:0] simp871_0;
  wire [6:0] comp2_0;
  wire [2:0] simp961_0;
  OR3 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0], gfint_2[0:0]);
  OR3 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1], gfint_2[1:1]);
  OR3 I2 (o_0r0[2:2], gfint_0[2:2], gfint_1[2:2], gfint_2[2:2]);
  OR3 I3 (o_0r0[3:3], gfint_0[3:3], gfint_1[3:3], gfint_2[3:3]);
  OR3 I4 (o_0r0[4:4], gfint_0[4:4], gfint_1[4:4], gfint_2[4:4]);
  OR3 I5 (o_0r0[5:5], gfint_0[5:5], gfint_1[5:5], gfint_2[5:5]);
  OR3 I6 (o_0r0[6:6], gfint_0[6:6], gfint_1[6:6], gfint_2[6:6]);
  OR3 I7 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0], gtint_2[0:0]);
  OR3 I8 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1], gtint_2[1:1]);
  OR3 I9 (o_0r1[2:2], gtint_0[2:2], gtint_1[2:2], gtint_2[2:2]);
  OR3 I10 (o_0r1[3:3], gtint_0[3:3], gtint_1[3:3], gtint_2[3:3]);
  OR3 I11 (o_0r1[4:4], gtint_0[4:4], gtint_1[4:4], gtint_2[4:4]);
  OR3 I12 (o_0r1[5:5], gtint_0[5:5], gtint_1[5:5], gtint_2[5:5]);
  OR3 I13 (o_0r1[6:6], gtint_0[6:6], gtint_1[6:6], gtint_2[6:6]);
  AND2 I14 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I15 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I16 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I17 (gtint_0[3:3], choice_0, i_0r1[3:3]);
  AND2 I18 (gtint_0[4:4], choice_0, i_0r1[4:4]);
  AND2 I19 (gtint_0[5:5], choice_0, i_0r1[5:5]);
  AND2 I20 (gtint_0[6:6], choice_0, i_0r1[6:6]);
  AND2 I21 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I22 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I23 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I24 (gtint_1[3:3], choice_1, i_1r1[3:3]);
  AND2 I25 (gtint_1[4:4], choice_1, i_1r1[4:4]);
  AND2 I26 (gtint_1[5:5], choice_1, i_1r1[5:5]);
  AND2 I27 (gtint_1[6:6], choice_1, i_1r1[6:6]);
  AND2 I28 (gtint_2[0:0], choice_2, i_2r1[0:0]);
  AND2 I29 (gtint_2[1:1], choice_2, i_2r1[1:1]);
  AND2 I30 (gtint_2[2:2], choice_2, i_2r1[2:2]);
  AND2 I31 (gtint_2[3:3], choice_2, i_2r1[3:3]);
  AND2 I32 (gtint_2[4:4], choice_2, i_2r1[4:4]);
  AND2 I33 (gtint_2[5:5], choice_2, i_2r1[5:5]);
  AND2 I34 (gtint_2[6:6], choice_2, i_2r1[6:6]);
  AND2 I35 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I36 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I37 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I38 (gfint_0[3:3], choice_0, i_0r0[3:3]);
  AND2 I39 (gfint_0[4:4], choice_0, i_0r0[4:4]);
  AND2 I40 (gfint_0[5:5], choice_0, i_0r0[5:5]);
  AND2 I41 (gfint_0[6:6], choice_0, i_0r0[6:6]);
  AND2 I42 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I43 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I44 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  AND2 I45 (gfint_1[3:3], choice_1, i_1r0[3:3]);
  AND2 I46 (gfint_1[4:4], choice_1, i_1r0[4:4]);
  AND2 I47 (gfint_1[5:5], choice_1, i_1r0[5:5]);
  AND2 I48 (gfint_1[6:6], choice_1, i_1r0[6:6]);
  AND2 I49 (gfint_2[0:0], choice_2, i_2r0[0:0]);
  AND2 I50 (gfint_2[1:1], choice_2, i_2r0[1:1]);
  AND2 I51 (gfint_2[2:2], choice_2, i_2r0[2:2]);
  AND2 I52 (gfint_2[3:3], choice_2, i_2r0[3:3]);
  AND2 I53 (gfint_2[4:4], choice_2, i_2r0[4:4]);
  AND2 I54 (gfint_2[5:5], choice_2, i_2r0[5:5]);
  AND2 I55 (gfint_2[6:6], choice_2, i_2r0[6:6]);
  OR2 I56 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I57 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I58 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I59 (comp0_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I60 (comp0_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I61 (comp0_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I62 (comp0_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  C3 I63 (simp781_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I64 (simp781_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  BUFF I65 (simp781_0[2:2], comp0_0[6:6]);
  C3 I66 (icomp_0, simp781_0[0:0], simp781_0[1:1], simp781_0[2:2]);
  OR2 I67 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I68 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I69 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  OR2 I70 (comp1_0[3:3], i_1r0[3:3], i_1r1[3:3]);
  OR2 I71 (comp1_0[4:4], i_1r0[4:4], i_1r1[4:4]);
  OR2 I72 (comp1_0[5:5], i_1r0[5:5], i_1r1[5:5]);
  OR2 I73 (comp1_0[6:6], i_1r0[6:6], i_1r1[6:6]);
  C3 I74 (simp871_0[0:0], comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C3 I75 (simp871_0[1:1], comp1_0[3:3], comp1_0[4:4], comp1_0[5:5]);
  BUFF I76 (simp871_0[2:2], comp1_0[6:6]);
  C3 I77 (icomp_1, simp871_0[0:0], simp871_0[1:1], simp871_0[2:2]);
  OR2 I78 (comp2_0[0:0], i_2r0[0:0], i_2r1[0:0]);
  OR2 I79 (comp2_0[1:1], i_2r0[1:1], i_2r1[1:1]);
  OR2 I80 (comp2_0[2:2], i_2r0[2:2], i_2r1[2:2]);
  OR2 I81 (comp2_0[3:3], i_2r0[3:3], i_2r1[3:3]);
  OR2 I82 (comp2_0[4:4], i_2r0[4:4], i_2r1[4:4]);
  OR2 I83 (comp2_0[5:5], i_2r0[5:5], i_2r1[5:5]);
  OR2 I84 (comp2_0[6:6], i_2r0[6:6], i_2r1[6:6]);
  C3 I85 (simp961_0[0:0], comp2_0[0:0], comp2_0[1:1], comp2_0[2:2]);
  C3 I86 (simp961_0[1:1], comp2_0[3:3], comp2_0[4:4], comp2_0[5:5]);
  BUFF I87 (simp961_0[2:2], comp2_0[6:6]);
  C3 I88 (icomp_2, simp961_0[0:0], simp961_0[1:1], simp961_0[2:2]);
  C2R I89 (choice_0, icomp_0, nchosen_0, reset);
  C2R I90 (choice_1, icomp_1, nchosen_0, reset);
  C2R I91 (choice_2, icomp_2, nchosen_0, reset);
  OR3 I92 (anychoice_0, choice_0, choice_1, choice_2);
  NOR2 I93 (nchosen_0, anychoice_0, o_0a);
  C2R I94 (i_0a, choice_0, o_0a, reset);
  C2R I95 (i_1a, choice_1, o_0a, reset);
  C2R I96 (i_2a, choice_2, o_0a, reset);
endmodule

// tks35_o32w3_1o0w32_2o0w32_4o0w32 TeakS (32+:3) [([Imp 1 0],0),([Imp 2 0],0),([Imp 4 0],0)] [One 35,M
//   any [32,32,32]]
module tks35_o32w3_1o0w32_2o0w32_4o0w32 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r0, o_1r1, o_1a, o_2r0, o_2r1, o_2a, reset);
  input [34:0] i_0r0;
  input [34:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  output [31:0] o_1r0;
  output [31:0] o_1r1;
  input o_1a;
  output [31:0] o_2r0;
  output [31:0] o_2r1;
  input o_2a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire match2_0;
  wire [34:0] comp_0;
  wire [11:0] simp561_0;
  wire [3:0] simp562_0;
  wire [1:0] simp563_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (match0_0, i_0r1[32:32], i_0r0[33:33], i_0r0[34:34]);
  BUFF I2 (sel_1, match1_0);
  C3 I3 (match1_0, i_0r0[32:32], i_0r1[33:33], i_0r0[34:34]);
  BUFF I4 (sel_2, match2_0);
  C3 I5 (match2_0, i_0r0[32:32], i_0r0[33:33], i_0r1[34:34]);
  C2 I6 (gsel_0, sel_0, icomplete_0);
  C2 I7 (gsel_1, sel_1, icomplete_0);
  C2 I8 (gsel_2, sel_2, icomplete_0);
  OR2 I9 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I10 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I11 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I12 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I13 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I14 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I15 (comp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I16 (comp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I17 (comp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I18 (comp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I19 (comp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I20 (comp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I21 (comp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I22 (comp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I23 (comp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I24 (comp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I25 (comp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I26 (comp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I27 (comp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I28 (comp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I29 (comp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I30 (comp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I31 (comp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I32 (comp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I33 (comp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I34 (comp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I35 (comp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I36 (comp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I37 (comp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I38 (comp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I39 (comp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I40 (comp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I41 (comp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  OR2 I42 (comp_0[33:33], i_0r0[33:33], i_0r1[33:33]);
  OR2 I43 (comp_0[34:34], i_0r0[34:34], i_0r1[34:34]);
  C3 I44 (simp561_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I45 (simp561_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C3 I46 (simp561_0[2:2], comp_0[6:6], comp_0[7:7], comp_0[8:8]);
  C3 I47 (simp561_0[3:3], comp_0[9:9], comp_0[10:10], comp_0[11:11]);
  C3 I48 (simp561_0[4:4], comp_0[12:12], comp_0[13:13], comp_0[14:14]);
  C3 I49 (simp561_0[5:5], comp_0[15:15], comp_0[16:16], comp_0[17:17]);
  C3 I50 (simp561_0[6:6], comp_0[18:18], comp_0[19:19], comp_0[20:20]);
  C3 I51 (simp561_0[7:7], comp_0[21:21], comp_0[22:22], comp_0[23:23]);
  C3 I52 (simp561_0[8:8], comp_0[24:24], comp_0[25:25], comp_0[26:26]);
  C3 I53 (simp561_0[9:9], comp_0[27:27], comp_0[28:28], comp_0[29:29]);
  C3 I54 (simp561_0[10:10], comp_0[30:30], comp_0[31:31], comp_0[32:32]);
  C2 I55 (simp561_0[11:11], comp_0[33:33], comp_0[34:34]);
  C3 I56 (simp562_0[0:0], simp561_0[0:0], simp561_0[1:1], simp561_0[2:2]);
  C3 I57 (simp562_0[1:1], simp561_0[3:3], simp561_0[4:4], simp561_0[5:5]);
  C3 I58 (simp562_0[2:2], simp561_0[6:6], simp561_0[7:7], simp561_0[8:8]);
  C3 I59 (simp562_0[3:3], simp561_0[9:9], simp561_0[10:10], simp561_0[11:11]);
  C3 I60 (simp563_0[0:0], simp562_0[0:0], simp562_0[1:1], simp562_0[2:2]);
  BUFF I61 (simp563_0[1:1], simp562_0[3:3]);
  C2 I62 (icomplete_0, simp563_0[0:0], simp563_0[1:1]);
  C2 I63 (o_0r0[0:0], i_0r0[0:0], gsel_0);
  C2 I64 (o_0r0[1:1], i_0r0[1:1], gsel_0);
  C2 I65 (o_0r0[2:2], i_0r0[2:2], gsel_0);
  C2 I66 (o_0r0[3:3], i_0r0[3:3], gsel_0);
  C2 I67 (o_0r0[4:4], i_0r0[4:4], gsel_0);
  C2 I68 (o_0r0[5:5], i_0r0[5:5], gsel_0);
  C2 I69 (o_0r0[6:6], i_0r0[6:6], gsel_0);
  C2 I70 (o_0r0[7:7], i_0r0[7:7], gsel_0);
  C2 I71 (o_0r0[8:8], i_0r0[8:8], gsel_0);
  C2 I72 (o_0r0[9:9], i_0r0[9:9], gsel_0);
  C2 I73 (o_0r0[10:10], i_0r0[10:10], gsel_0);
  C2 I74 (o_0r0[11:11], i_0r0[11:11], gsel_0);
  C2 I75 (o_0r0[12:12], i_0r0[12:12], gsel_0);
  C2 I76 (o_0r0[13:13], i_0r0[13:13], gsel_0);
  C2 I77 (o_0r0[14:14], i_0r0[14:14], gsel_0);
  C2 I78 (o_0r0[15:15], i_0r0[15:15], gsel_0);
  C2 I79 (o_0r0[16:16], i_0r0[16:16], gsel_0);
  C2 I80 (o_0r0[17:17], i_0r0[17:17], gsel_0);
  C2 I81 (o_0r0[18:18], i_0r0[18:18], gsel_0);
  C2 I82 (o_0r0[19:19], i_0r0[19:19], gsel_0);
  C2 I83 (o_0r0[20:20], i_0r0[20:20], gsel_0);
  C2 I84 (o_0r0[21:21], i_0r0[21:21], gsel_0);
  C2 I85 (o_0r0[22:22], i_0r0[22:22], gsel_0);
  C2 I86 (o_0r0[23:23], i_0r0[23:23], gsel_0);
  C2 I87 (o_0r0[24:24], i_0r0[24:24], gsel_0);
  C2 I88 (o_0r0[25:25], i_0r0[25:25], gsel_0);
  C2 I89 (o_0r0[26:26], i_0r0[26:26], gsel_0);
  C2 I90 (o_0r0[27:27], i_0r0[27:27], gsel_0);
  C2 I91 (o_0r0[28:28], i_0r0[28:28], gsel_0);
  C2 I92 (o_0r0[29:29], i_0r0[29:29], gsel_0);
  C2 I93 (o_0r0[30:30], i_0r0[30:30], gsel_0);
  C2 I94 (o_0r0[31:31], i_0r0[31:31], gsel_0);
  C2 I95 (o_1r0[0:0], i_0r0[0:0], gsel_1);
  C2 I96 (o_1r0[1:1], i_0r0[1:1], gsel_1);
  C2 I97 (o_1r0[2:2], i_0r0[2:2], gsel_1);
  C2 I98 (o_1r0[3:3], i_0r0[3:3], gsel_1);
  C2 I99 (o_1r0[4:4], i_0r0[4:4], gsel_1);
  C2 I100 (o_1r0[5:5], i_0r0[5:5], gsel_1);
  C2 I101 (o_1r0[6:6], i_0r0[6:6], gsel_1);
  C2 I102 (o_1r0[7:7], i_0r0[7:7], gsel_1);
  C2 I103 (o_1r0[8:8], i_0r0[8:8], gsel_1);
  C2 I104 (o_1r0[9:9], i_0r0[9:9], gsel_1);
  C2 I105 (o_1r0[10:10], i_0r0[10:10], gsel_1);
  C2 I106 (o_1r0[11:11], i_0r0[11:11], gsel_1);
  C2 I107 (o_1r0[12:12], i_0r0[12:12], gsel_1);
  C2 I108 (o_1r0[13:13], i_0r0[13:13], gsel_1);
  C2 I109 (o_1r0[14:14], i_0r0[14:14], gsel_1);
  C2 I110 (o_1r0[15:15], i_0r0[15:15], gsel_1);
  C2 I111 (o_1r0[16:16], i_0r0[16:16], gsel_1);
  C2 I112 (o_1r0[17:17], i_0r0[17:17], gsel_1);
  C2 I113 (o_1r0[18:18], i_0r0[18:18], gsel_1);
  C2 I114 (o_1r0[19:19], i_0r0[19:19], gsel_1);
  C2 I115 (o_1r0[20:20], i_0r0[20:20], gsel_1);
  C2 I116 (o_1r0[21:21], i_0r0[21:21], gsel_1);
  C2 I117 (o_1r0[22:22], i_0r0[22:22], gsel_1);
  C2 I118 (o_1r0[23:23], i_0r0[23:23], gsel_1);
  C2 I119 (o_1r0[24:24], i_0r0[24:24], gsel_1);
  C2 I120 (o_1r0[25:25], i_0r0[25:25], gsel_1);
  C2 I121 (o_1r0[26:26], i_0r0[26:26], gsel_1);
  C2 I122 (o_1r0[27:27], i_0r0[27:27], gsel_1);
  C2 I123 (o_1r0[28:28], i_0r0[28:28], gsel_1);
  C2 I124 (o_1r0[29:29], i_0r0[29:29], gsel_1);
  C2 I125 (o_1r0[30:30], i_0r0[30:30], gsel_1);
  C2 I126 (o_1r0[31:31], i_0r0[31:31], gsel_1);
  C2 I127 (o_2r0[0:0], i_0r0[0:0], gsel_2);
  C2 I128 (o_2r0[1:1], i_0r0[1:1], gsel_2);
  C2 I129 (o_2r0[2:2], i_0r0[2:2], gsel_2);
  C2 I130 (o_2r0[3:3], i_0r0[3:3], gsel_2);
  C2 I131 (o_2r0[4:4], i_0r0[4:4], gsel_2);
  C2 I132 (o_2r0[5:5], i_0r0[5:5], gsel_2);
  C2 I133 (o_2r0[6:6], i_0r0[6:6], gsel_2);
  C2 I134 (o_2r0[7:7], i_0r0[7:7], gsel_2);
  C2 I135 (o_2r0[8:8], i_0r0[8:8], gsel_2);
  C2 I136 (o_2r0[9:9], i_0r0[9:9], gsel_2);
  C2 I137 (o_2r0[10:10], i_0r0[10:10], gsel_2);
  C2 I138 (o_2r0[11:11], i_0r0[11:11], gsel_2);
  C2 I139 (o_2r0[12:12], i_0r0[12:12], gsel_2);
  C2 I140 (o_2r0[13:13], i_0r0[13:13], gsel_2);
  C2 I141 (o_2r0[14:14], i_0r0[14:14], gsel_2);
  C2 I142 (o_2r0[15:15], i_0r0[15:15], gsel_2);
  C2 I143 (o_2r0[16:16], i_0r0[16:16], gsel_2);
  C2 I144 (o_2r0[17:17], i_0r0[17:17], gsel_2);
  C2 I145 (o_2r0[18:18], i_0r0[18:18], gsel_2);
  C2 I146 (o_2r0[19:19], i_0r0[19:19], gsel_2);
  C2 I147 (o_2r0[20:20], i_0r0[20:20], gsel_2);
  C2 I148 (o_2r0[21:21], i_0r0[21:21], gsel_2);
  C2 I149 (o_2r0[22:22], i_0r0[22:22], gsel_2);
  C2 I150 (o_2r0[23:23], i_0r0[23:23], gsel_2);
  C2 I151 (o_2r0[24:24], i_0r0[24:24], gsel_2);
  C2 I152 (o_2r0[25:25], i_0r0[25:25], gsel_2);
  C2 I153 (o_2r0[26:26], i_0r0[26:26], gsel_2);
  C2 I154 (o_2r0[27:27], i_0r0[27:27], gsel_2);
  C2 I155 (o_2r0[28:28], i_0r0[28:28], gsel_2);
  C2 I156 (o_2r0[29:29], i_0r0[29:29], gsel_2);
  C2 I157 (o_2r0[30:30], i_0r0[30:30], gsel_2);
  C2 I158 (o_2r0[31:31], i_0r0[31:31], gsel_2);
  C2 I159 (o_0r1[0:0], i_0r1[0:0], gsel_0);
  C2 I160 (o_0r1[1:1], i_0r1[1:1], gsel_0);
  C2 I161 (o_0r1[2:2], i_0r1[2:2], gsel_0);
  C2 I162 (o_0r1[3:3], i_0r1[3:3], gsel_0);
  C2 I163 (o_0r1[4:4], i_0r1[4:4], gsel_0);
  C2 I164 (o_0r1[5:5], i_0r1[5:5], gsel_0);
  C2 I165 (o_0r1[6:6], i_0r1[6:6], gsel_0);
  C2 I166 (o_0r1[7:7], i_0r1[7:7], gsel_0);
  C2 I167 (o_0r1[8:8], i_0r1[8:8], gsel_0);
  C2 I168 (o_0r1[9:9], i_0r1[9:9], gsel_0);
  C2 I169 (o_0r1[10:10], i_0r1[10:10], gsel_0);
  C2 I170 (o_0r1[11:11], i_0r1[11:11], gsel_0);
  C2 I171 (o_0r1[12:12], i_0r1[12:12], gsel_0);
  C2 I172 (o_0r1[13:13], i_0r1[13:13], gsel_0);
  C2 I173 (o_0r1[14:14], i_0r1[14:14], gsel_0);
  C2 I174 (o_0r1[15:15], i_0r1[15:15], gsel_0);
  C2 I175 (o_0r1[16:16], i_0r1[16:16], gsel_0);
  C2 I176 (o_0r1[17:17], i_0r1[17:17], gsel_0);
  C2 I177 (o_0r1[18:18], i_0r1[18:18], gsel_0);
  C2 I178 (o_0r1[19:19], i_0r1[19:19], gsel_0);
  C2 I179 (o_0r1[20:20], i_0r1[20:20], gsel_0);
  C2 I180 (o_0r1[21:21], i_0r1[21:21], gsel_0);
  C2 I181 (o_0r1[22:22], i_0r1[22:22], gsel_0);
  C2 I182 (o_0r1[23:23], i_0r1[23:23], gsel_0);
  C2 I183 (o_0r1[24:24], i_0r1[24:24], gsel_0);
  C2 I184 (o_0r1[25:25], i_0r1[25:25], gsel_0);
  C2 I185 (o_0r1[26:26], i_0r1[26:26], gsel_0);
  C2 I186 (o_0r1[27:27], i_0r1[27:27], gsel_0);
  C2 I187 (o_0r1[28:28], i_0r1[28:28], gsel_0);
  C2 I188 (o_0r1[29:29], i_0r1[29:29], gsel_0);
  C2 I189 (o_0r1[30:30], i_0r1[30:30], gsel_0);
  C2 I190 (o_0r1[31:31], i_0r1[31:31], gsel_0);
  C2 I191 (o_1r1[0:0], i_0r1[0:0], gsel_1);
  C2 I192 (o_1r1[1:1], i_0r1[1:1], gsel_1);
  C2 I193 (o_1r1[2:2], i_0r1[2:2], gsel_1);
  C2 I194 (o_1r1[3:3], i_0r1[3:3], gsel_1);
  C2 I195 (o_1r1[4:4], i_0r1[4:4], gsel_1);
  C2 I196 (o_1r1[5:5], i_0r1[5:5], gsel_1);
  C2 I197 (o_1r1[6:6], i_0r1[6:6], gsel_1);
  C2 I198 (o_1r1[7:7], i_0r1[7:7], gsel_1);
  C2 I199 (o_1r1[8:8], i_0r1[8:8], gsel_1);
  C2 I200 (o_1r1[9:9], i_0r1[9:9], gsel_1);
  C2 I201 (o_1r1[10:10], i_0r1[10:10], gsel_1);
  C2 I202 (o_1r1[11:11], i_0r1[11:11], gsel_1);
  C2 I203 (o_1r1[12:12], i_0r1[12:12], gsel_1);
  C2 I204 (o_1r1[13:13], i_0r1[13:13], gsel_1);
  C2 I205 (o_1r1[14:14], i_0r1[14:14], gsel_1);
  C2 I206 (o_1r1[15:15], i_0r1[15:15], gsel_1);
  C2 I207 (o_1r1[16:16], i_0r1[16:16], gsel_1);
  C2 I208 (o_1r1[17:17], i_0r1[17:17], gsel_1);
  C2 I209 (o_1r1[18:18], i_0r1[18:18], gsel_1);
  C2 I210 (o_1r1[19:19], i_0r1[19:19], gsel_1);
  C2 I211 (o_1r1[20:20], i_0r1[20:20], gsel_1);
  C2 I212 (o_1r1[21:21], i_0r1[21:21], gsel_1);
  C2 I213 (o_1r1[22:22], i_0r1[22:22], gsel_1);
  C2 I214 (o_1r1[23:23], i_0r1[23:23], gsel_1);
  C2 I215 (o_1r1[24:24], i_0r1[24:24], gsel_1);
  C2 I216 (o_1r1[25:25], i_0r1[25:25], gsel_1);
  C2 I217 (o_1r1[26:26], i_0r1[26:26], gsel_1);
  C2 I218 (o_1r1[27:27], i_0r1[27:27], gsel_1);
  C2 I219 (o_1r1[28:28], i_0r1[28:28], gsel_1);
  C2 I220 (o_1r1[29:29], i_0r1[29:29], gsel_1);
  C2 I221 (o_1r1[30:30], i_0r1[30:30], gsel_1);
  C2 I222 (o_1r1[31:31], i_0r1[31:31], gsel_1);
  C2 I223 (o_2r1[0:0], i_0r1[0:0], gsel_2);
  C2 I224 (o_2r1[1:1], i_0r1[1:1], gsel_2);
  C2 I225 (o_2r1[2:2], i_0r1[2:2], gsel_2);
  C2 I226 (o_2r1[3:3], i_0r1[3:3], gsel_2);
  C2 I227 (o_2r1[4:4], i_0r1[4:4], gsel_2);
  C2 I228 (o_2r1[5:5], i_0r1[5:5], gsel_2);
  C2 I229 (o_2r1[6:6], i_0r1[6:6], gsel_2);
  C2 I230 (o_2r1[7:7], i_0r1[7:7], gsel_2);
  C2 I231 (o_2r1[8:8], i_0r1[8:8], gsel_2);
  C2 I232 (o_2r1[9:9], i_0r1[9:9], gsel_2);
  C2 I233 (o_2r1[10:10], i_0r1[10:10], gsel_2);
  C2 I234 (o_2r1[11:11], i_0r1[11:11], gsel_2);
  C2 I235 (o_2r1[12:12], i_0r1[12:12], gsel_2);
  C2 I236 (o_2r1[13:13], i_0r1[13:13], gsel_2);
  C2 I237 (o_2r1[14:14], i_0r1[14:14], gsel_2);
  C2 I238 (o_2r1[15:15], i_0r1[15:15], gsel_2);
  C2 I239 (o_2r1[16:16], i_0r1[16:16], gsel_2);
  C2 I240 (o_2r1[17:17], i_0r1[17:17], gsel_2);
  C2 I241 (o_2r1[18:18], i_0r1[18:18], gsel_2);
  C2 I242 (o_2r1[19:19], i_0r1[19:19], gsel_2);
  C2 I243 (o_2r1[20:20], i_0r1[20:20], gsel_2);
  C2 I244 (o_2r1[21:21], i_0r1[21:21], gsel_2);
  C2 I245 (o_2r1[22:22], i_0r1[22:22], gsel_2);
  C2 I246 (o_2r1[23:23], i_0r1[23:23], gsel_2);
  C2 I247 (o_2r1[24:24], i_0r1[24:24], gsel_2);
  C2 I248 (o_2r1[25:25], i_0r1[25:25], gsel_2);
  C2 I249 (o_2r1[26:26], i_0r1[26:26], gsel_2);
  C2 I250 (o_2r1[27:27], i_0r1[27:27], gsel_2);
  C2 I251 (o_2r1[28:28], i_0r1[28:28], gsel_2);
  C2 I252 (o_2r1[29:29], i_0r1[29:29], gsel_2);
  C2 I253 (o_2r1[30:30], i_0r1[30:30], gsel_2);
  C2 I254 (o_2r1[31:31], i_0r1[31:31], gsel_2);
  OR3 I255 (oack_0, o_0a, o_1a, o_2a);
  C2 I256 (i_0a, oack_0, icomplete_0);
endmodule

// tkj7m4_3 TeakJ [Many [4,3],One 7]
module tkj7m4_3 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [3:0] i_0r0;
  input [3:0] i_0r1;
  output i_0a;
  input [2:0] i_1r0;
  input [2:0] i_1r1;
  output i_1a;
  output [6:0] o_0r0;
  output [6:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [6:0] joinf_0;
  wire [6:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_1r0[0:0]);
  BUFF I5 (joinf_0[5:5], i_1r0[1:1]);
  BUFF I6 (joinf_0[6:6], i_1r0[2:2]);
  BUFF I7 (joint_0[0:0], i_0r1[0:0]);
  BUFF I8 (joint_0[1:1], i_0r1[1:1]);
  BUFF I9 (joint_0[2:2], i_0r1[2:2]);
  BUFF I10 (joint_0[3:3], i_0r1[3:3]);
  BUFF I11 (joint_0[4:4], i_1r1[0:0]);
  BUFF I12 (joint_0[5:5], i_1r1[1:1]);
  BUFF I13 (joint_0[6:6], i_1r1[2:2]);
  OR2 I14 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I15 (icomplete_0, dcomplete_0);
  C2 I16 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I17 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I18 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I19 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I20 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I21 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I22 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I23 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I24 (o_0r1[1:1], joint_0[1:1]);
  BUFF I25 (o_0r1[2:2], joint_0[2:2]);
  BUFF I26 (o_0r1[3:3], joint_0[3:3]);
  BUFF I27 (o_0r1[4:4], joint_0[4:4]);
  BUFF I28 (o_0r1[5:5], joint_0[5:5]);
  BUFF I29 (o_0r1[6:6], joint_0[6:6]);
  BUFF I30 (i_0a, o_0a);
  BUFF I31 (i_1a, o_0a);
endmodule

// tks7_o4w3_1o0w4_2o0w4_4o0w4 TeakS (4+:3) [([Imp 1 0],0),([Imp 2 0],0),([Imp 4 0],0)] [One 7,Many [4,
//   4,4]]
module tks7_o4w3_1o0w4_2o0w4_4o0w4 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r0, o_1r1, o_1a, o_2r0, o_2r1, o_2a, reset);
  input [6:0] i_0r0;
  input [6:0] i_0r1;
  output i_0a;
  output [3:0] o_0r0;
  output [3:0] o_0r1;
  input o_0a;
  output [3:0] o_1r0;
  output [3:0] o_1r1;
  input o_1a;
  output [3:0] o_2r0;
  output [3:0] o_2r1;
  input o_2a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire sel_2;
  wire gsel_0;
  wire gsel_1;
  wire gsel_2;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire match2_0;
  wire [6:0] comp_0;
  wire [2:0] simp281_0;
  BUFF I0 (sel_0, match0_0);
  C3 I1 (match0_0, i_0r1[4:4], i_0r0[5:5], i_0r0[6:6]);
  BUFF I2 (sel_1, match1_0);
  C3 I3 (match1_0, i_0r0[4:4], i_0r1[5:5], i_0r0[6:6]);
  BUFF I4 (sel_2, match2_0);
  C3 I5 (match2_0, i_0r0[4:4], i_0r0[5:5], i_0r1[6:6]);
  C2 I6 (gsel_0, sel_0, icomplete_0);
  C2 I7 (gsel_1, sel_1, icomplete_0);
  C2 I8 (gsel_2, sel_2, icomplete_0);
  OR2 I9 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I10 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I11 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I12 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I13 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I14 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I15 (comp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  C3 I16 (simp281_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I17 (simp281_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  BUFF I18 (simp281_0[2:2], comp_0[6:6]);
  C3 I19 (icomplete_0, simp281_0[0:0], simp281_0[1:1], simp281_0[2:2]);
  C2 I20 (o_0r0[0:0], i_0r0[0:0], gsel_0);
  C2 I21 (o_0r0[1:1], i_0r0[1:1], gsel_0);
  C2 I22 (o_0r0[2:2], i_0r0[2:2], gsel_0);
  C2 I23 (o_0r0[3:3], i_0r0[3:3], gsel_0);
  C2 I24 (o_1r0[0:0], i_0r0[0:0], gsel_1);
  C2 I25 (o_1r0[1:1], i_0r0[1:1], gsel_1);
  C2 I26 (o_1r0[2:2], i_0r0[2:2], gsel_1);
  C2 I27 (o_1r0[3:3], i_0r0[3:3], gsel_1);
  C2 I28 (o_2r0[0:0], i_0r0[0:0], gsel_2);
  C2 I29 (o_2r0[1:1], i_0r0[1:1], gsel_2);
  C2 I30 (o_2r0[2:2], i_0r0[2:2], gsel_2);
  C2 I31 (o_2r0[3:3], i_0r0[3:3], gsel_2);
  C2 I32 (o_0r1[0:0], i_0r1[0:0], gsel_0);
  C2 I33 (o_0r1[1:1], i_0r1[1:1], gsel_0);
  C2 I34 (o_0r1[2:2], i_0r1[2:2], gsel_0);
  C2 I35 (o_0r1[3:3], i_0r1[3:3], gsel_0);
  C2 I36 (o_1r1[0:0], i_0r1[0:0], gsel_1);
  C2 I37 (o_1r1[1:1], i_0r1[1:1], gsel_1);
  C2 I38 (o_1r1[2:2], i_0r1[2:2], gsel_1);
  C2 I39 (o_1r1[3:3], i_0r1[3:3], gsel_1);
  C2 I40 (o_2r1[0:0], i_0r1[0:0], gsel_2);
  C2 I41 (o_2r1[1:1], i_0r1[1:1], gsel_2);
  C2 I42 (o_2r1[2:2], i_0r1[2:2], gsel_2);
  C2 I43 (o_2r1[3:3], i_0r1[3:3], gsel_2);
  OR3 I44 (oack_0, o_0a, o_1a, o_2a);
  C2 I45 (i_0a, oack_0, icomplete_0);
endmodule

// tkm2x3b TeakM [Many [3,3],One 3]
module tkm2x3b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [2:0] i_0r0;
  input [2:0] i_0r1;
  output i_0a;
  input [2:0] i_1r0;
  input [2:0] i_1r1;
  output i_1a;
  output [2:0] o_0r0;
  output [2:0] o_0r1;
  input o_0a;
  input reset;
  wire [2:0] gfint_0;
  wire [2:0] gfint_1;
  wire [2:0] gtint_0;
  wire [2:0] gtint_1;
  wire choice_0;
  wire choice_1;
  wire anychoice_0;
  wire icomp_0;
  wire icomp_1;
  wire nchosen_0;
  wire [2:0] comp0_0;
  wire [2:0] comp1_0;
  OR2 I0 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0]);
  OR2 I1 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1]);
  OR2 I2 (o_0r0[2:2], gfint_0[2:2], gfint_1[2:2]);
  OR2 I3 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0]);
  OR2 I4 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1]);
  OR2 I5 (o_0r1[2:2], gtint_0[2:2], gtint_1[2:2]);
  AND2 I6 (gtint_0[0:0], choice_0, i_0r1[0:0]);
  AND2 I7 (gtint_0[1:1], choice_0, i_0r1[1:1]);
  AND2 I8 (gtint_0[2:2], choice_0, i_0r1[2:2]);
  AND2 I9 (gtint_1[0:0], choice_1, i_1r1[0:0]);
  AND2 I10 (gtint_1[1:1], choice_1, i_1r1[1:1]);
  AND2 I11 (gtint_1[2:2], choice_1, i_1r1[2:2]);
  AND2 I12 (gfint_0[0:0], choice_0, i_0r0[0:0]);
  AND2 I13 (gfint_0[1:1], choice_0, i_0r0[1:1]);
  AND2 I14 (gfint_0[2:2], choice_0, i_0r0[2:2]);
  AND2 I15 (gfint_1[0:0], choice_1, i_1r0[0:0]);
  AND2 I16 (gfint_1[1:1], choice_1, i_1r0[1:1]);
  AND2 I17 (gfint_1[2:2], choice_1, i_1r0[2:2]);
  OR2 I18 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I19 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I20 (comp0_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  C3 I21 (icomp_0, comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  OR2 I22 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I23 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  OR2 I24 (comp1_0[2:2], i_1r0[2:2], i_1r1[2:2]);
  C3 I25 (icomp_1, comp1_0[0:0], comp1_0[1:1], comp1_0[2:2]);
  C2R I26 (choice_0, icomp_0, nchosen_0, reset);
  C2R I27 (choice_1, icomp_1, nchosen_0, reset);
  OR2 I28 (anychoice_0, choice_0, choice_1);
  NOR2 I29 (nchosen_0, anychoice_0, o_0a);
  C2R I30 (i_0a, choice_0, o_0a, reset);
  C2R I31 (i_1a, choice_1, o_0a, reset);
endmodule

// tkvv32_wo0w32_ro0w32 TeakV "v" 32 [] [0] [0] [Many [32],Many [0],Many [0],Many [32]]
module tkvv32_wo0w32_ro0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I457 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I458 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I459 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I460 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I461 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I462 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I463 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I464 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I465 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I466 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I467 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I468 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I469 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I470 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I471 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I472 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I473 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I474 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I475 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I476 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I477 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I478 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I479 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I480 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I481 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I482 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I483 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I484 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I485 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I486 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I487 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  OR2 I488 (anyread_0, rg_0r, rg_0a);
  BUFF I489 (wg_0a, wd_0a);
  BUFF I490 (rg_0a, rd_0a);
endmodule

// tkvmread32_wo0w32_ro0w32 TeakV "mread" 32 [] [0] [0] [Many [32],Many [0],Many [0],Many [32]]
module tkvmread32_wo0w32_ro0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I457 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I458 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I459 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I460 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I461 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I462 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I463 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I464 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I465 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I466 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I467 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I468 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I469 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I470 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I471 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I472 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I473 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I474 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I475 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I476 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I477 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I478 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I479 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I480 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I481 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I482 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I483 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I484 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I485 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I486 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I487 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  OR2 I488 (anyread_0, rg_0r, rg_0a);
  BUFF I489 (wg_0a, wd_0a);
  BUFF I490 (rg_0a, rd_0a);
endmodule

// tkvfaddr32_wo0w32_ro0w32 TeakV "faddr" 32 [] [0] [0] [Many [32],Many [0],Many [0],Many [32]]
module tkvfaddr32_wo0w32_ro0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I457 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I458 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I459 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I460 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I461 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I462 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I463 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I464 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I465 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I466 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I467 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I468 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I469 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I470 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I471 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I472 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I473 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I474 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I475 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I476 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I477 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I478 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I479 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I480 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I481 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I482 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I483 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I484 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I485 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I486 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I487 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  OR2 I488 (anyread_0, rg_0r, rg_0a);
  BUFF I489 (wg_0a, wd_0a);
  BUFF I490 (rg_0a, rd_0a);
endmodule

// tkvdwrite32_wo0w32_ro0w32 TeakV "dwrite" 32 [] [0] [0] [Many [32],Many [0],Many [0],Many [32]]
module tkvdwrite32_wo0w32_ro0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I457 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I458 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I459 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I460 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I461 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I462 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I463 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I464 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I465 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I466 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I467 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I468 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I469 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I470 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I471 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I472 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I473 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I474 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I475 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I476 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I477 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I478 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I479 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I480 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I481 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I482 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I483 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I484 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I485 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I486 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I487 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  OR2 I488 (anyread_0, rg_0r, rg_0a);
  BUFF I489 (wg_0a, wd_0a);
  BUFF I490 (rg_0a, rd_0a);
endmodule

// tkvdaddr32_wo0w32_ro0w32 TeakV "daddr" 32 [] [0] [0] [Many [32],Many [0],Many [0],Many [32]]
module tkvdaddr32_wo0w32_ro0w32 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [31:0] wg_0r0;
  input [31:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [31:0] rd_0r0;
  output [31:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [31:0] wf_0;
  wire [31:0] wt_0;
  wire [31:0] df_0;
  wire [31:0] dt_0;
  wire wc_0;
  wire [31:0] wacks_0;
  wire [31:0] wenr_0;
  wire [31:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [31:0] drlgf_0;
  wire [31:0] drlgt_0;
  wire [31:0] comp0_0;
  wire [10:0] simp2381_0;
  wire [3:0] simp2382_0;
  wire [1:0] simp2383_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [31:0] conwgit_0;
  wire [31:0] conwgif_0;
  wire conwig_0;
  wire [10:0] simp4071_0;
  wire [3:0] simp4072_0;
  wire [1:0] simp4073_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I34 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I35 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I36 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I37 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I38 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I39 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I40 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I41 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I42 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I43 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I44 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I45 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I46 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I47 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I48 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I49 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I50 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I51 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I52 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I53 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I54 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I55 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I56 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I57 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I58 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I59 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I60 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I61 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I62 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I63 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I64 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I65 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I66 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I67 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I68 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I69 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I70 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I71 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I72 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I73 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I74 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I75 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I76 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I77 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I78 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I79 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I80 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I81 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I82 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I83 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I84 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I85 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I86 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I87 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I88 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I89 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I90 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I91 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I92 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I93 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I94 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I95 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I96 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  NOR2 I97 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I98 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I99 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I100 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I101 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I102 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I103 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I104 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I105 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I106 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I107 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I108 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I109 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I110 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I111 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I112 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I113 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I114 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I115 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I116 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I117 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I118 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I119 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I120 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I121 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I122 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I123 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I124 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I125 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I126 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I127 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I128 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR3 I129 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I130 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I131 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I132 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I133 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I134 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I135 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I136 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I137 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I138 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I139 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I140 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I141 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I142 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I143 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I144 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I145 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I146 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I147 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I148 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I149 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I150 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I151 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I152 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I153 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I154 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I155 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I156 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I157 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I158 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I159 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I160 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  AO22 I161 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I162 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I163 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I164 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I165 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I166 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I167 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I168 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I169 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I170 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I171 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I172 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I173 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I174 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I175 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I176 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I177 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I178 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I179 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I180 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I181 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I182 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I183 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I184 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I185 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I186 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I187 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I188 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I189 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I190 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I191 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I192 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  OR2 I193 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I194 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I195 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I196 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I197 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I198 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I199 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I200 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I201 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I202 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I203 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I204 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I205 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I206 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I207 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I208 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I209 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I210 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I211 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I212 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I213 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I214 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I215 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I216 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I217 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I218 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I219 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I220 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I221 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I222 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I223 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I224 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  C3 I225 (simp2381_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I226 (simp2381_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I227 (simp2381_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I228 (simp2381_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I229 (simp2381_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I230 (simp2381_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I231 (simp2381_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I232 (simp2381_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I233 (simp2381_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I234 (simp2381_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C2 I235 (simp2381_0[10:10], comp0_0[30:30], comp0_0[31:31]);
  C3 I236 (simp2382_0[0:0], simp2381_0[0:0], simp2381_0[1:1], simp2381_0[2:2]);
  C3 I237 (simp2382_0[1:1], simp2381_0[3:3], simp2381_0[4:4], simp2381_0[5:5]);
  C3 I238 (simp2382_0[2:2], simp2381_0[6:6], simp2381_0[7:7], simp2381_0[8:8]);
  C2 I239 (simp2382_0[3:3], simp2381_0[9:9], simp2381_0[10:10]);
  C3 I240 (simp2383_0[0:0], simp2382_0[0:0], simp2382_0[1:1], simp2382_0[2:2]);
  BUFF I241 (simp2383_0[1:1], simp2382_0[3:3]);
  C2 I242 (wc_0, simp2383_0[0:0], simp2383_0[1:1]);
  AND2 I243 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I244 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I245 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I246 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I247 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I248 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I249 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I250 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I251 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I252 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I253 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I254 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I255 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I256 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I257 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I258 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I259 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I260 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I261 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I262 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I263 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I264 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I265 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I266 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I267 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I268 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I269 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I270 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I271 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I272 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I273 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I274 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I275 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I276 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I277 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I278 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I279 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I280 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I281 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I282 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I283 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I284 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I285 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I286 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I287 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I288 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I289 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I290 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I291 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I292 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I293 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I294 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I295 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I296 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I297 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I298 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I299 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I300 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I301 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I302 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I303 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I304 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I305 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I306 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  BUFF I307 (conwigc_0, wc_0);
  AO22 I308 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I309 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I310 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I311 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I312 (wenr_0[0:0], wc_0);
  BUFF I313 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I314 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I315 (wenr_0[1:1], wc_0);
  BUFF I316 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I317 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I318 (wenr_0[2:2], wc_0);
  BUFF I319 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I320 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I321 (wenr_0[3:3], wc_0);
  BUFF I322 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I323 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I324 (wenr_0[4:4], wc_0);
  BUFF I325 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I326 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I327 (wenr_0[5:5], wc_0);
  BUFF I328 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I329 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I330 (wenr_0[6:6], wc_0);
  BUFF I331 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I332 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I333 (wenr_0[7:7], wc_0);
  BUFF I334 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I335 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I336 (wenr_0[8:8], wc_0);
  BUFF I337 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I338 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I339 (wenr_0[9:9], wc_0);
  BUFF I340 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I341 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I342 (wenr_0[10:10], wc_0);
  BUFF I343 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I344 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I345 (wenr_0[11:11], wc_0);
  BUFF I346 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I347 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I348 (wenr_0[12:12], wc_0);
  BUFF I349 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I350 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I351 (wenr_0[13:13], wc_0);
  BUFF I352 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I353 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I354 (wenr_0[14:14], wc_0);
  BUFF I355 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I356 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I357 (wenr_0[15:15], wc_0);
  BUFF I358 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I359 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I360 (wenr_0[16:16], wc_0);
  BUFF I361 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I362 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I363 (wenr_0[17:17], wc_0);
  BUFF I364 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I365 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I366 (wenr_0[18:18], wc_0);
  BUFF I367 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I368 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I369 (wenr_0[19:19], wc_0);
  BUFF I370 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I371 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I372 (wenr_0[20:20], wc_0);
  BUFF I373 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I374 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I375 (wenr_0[21:21], wc_0);
  BUFF I376 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I377 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I378 (wenr_0[22:22], wc_0);
  BUFF I379 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I380 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I381 (wenr_0[23:23], wc_0);
  BUFF I382 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I383 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I384 (wenr_0[24:24], wc_0);
  BUFF I385 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I386 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I387 (wenr_0[25:25], wc_0);
  BUFF I388 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I389 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I390 (wenr_0[26:26], wc_0);
  BUFF I391 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I392 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I393 (wenr_0[27:27], wc_0);
  BUFF I394 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I395 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I396 (wenr_0[28:28], wc_0);
  BUFF I397 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I398 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I399 (wenr_0[29:29], wc_0);
  BUFF I400 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I401 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I402 (wenr_0[30:30], wc_0);
  BUFF I403 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I404 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I405 (wenr_0[31:31], wc_0);
  C3 I406 (simp4071_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I407 (simp4071_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I408 (simp4071_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I409 (simp4071_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I410 (simp4071_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I411 (simp4071_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I412 (simp4071_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I413 (simp4071_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I414 (simp4071_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I415 (simp4071_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I416 (simp4071_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I417 (simp4072_0[0:0], simp4071_0[0:0], simp4071_0[1:1], simp4071_0[2:2]);
  C3 I418 (simp4072_0[1:1], simp4071_0[3:3], simp4071_0[4:4], simp4071_0[5:5]);
  C3 I419 (simp4072_0[2:2], simp4071_0[6:6], simp4071_0[7:7], simp4071_0[8:8]);
  C2 I420 (simp4072_0[3:3], simp4071_0[9:9], simp4071_0[10:10]);
  C3 I421 (simp4073_0[0:0], simp4072_0[0:0], simp4072_0[1:1], simp4072_0[2:2]);
  BUFF I422 (simp4073_0[1:1], simp4072_0[3:3]);
  C2 I423 (wd_0r, simp4073_0[0:0], simp4073_0[1:1]);
  AND2 I424 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I425 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I426 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I427 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I428 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I429 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I430 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I431 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I432 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I433 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I434 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I435 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I436 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I437 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I438 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I439 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I440 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I441 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I442 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I443 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I444 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I445 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I446 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I447 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I448 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I449 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I450 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I451 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I452 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I453 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I454 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I455 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I456 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I457 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I458 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I459 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I460 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I461 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I462 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I463 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I464 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I465 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I466 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I467 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I468 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I469 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I470 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I471 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I472 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I473 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I474 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I475 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I476 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I477 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I478 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I479 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I480 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I481 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I482 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I483 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I484 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I485 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I486 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I487 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  OR2 I488 (anyread_0, rg_0r, rg_0a);
  BUFF I489 (wg_0a, wd_0a);
  BUFF I490 (rg_0a, rd_0a);
endmodule

// tkvdaccess3_wo0w3_ro0w3o0w1 TeakV "daccess" 3 [] [0] [0,0] [Many [3],Many [0],Many [0,0],Many [3,1]]
module tkvdaccess3_wo0w3_ro0w3o0w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rg_1r, rg_1a, rd_0r0, rd_0r1, rd_0a, rd_1r0, rd_1r1, rd_1a, reset);
  input [2:0] wg_0r0;
  input [2:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  input rg_1r;
  output rg_1a;
  output [2:0] rd_0r0;
  output [2:0] rd_0r1;
  input rd_0a;
  output rd_1r0;
  output rd_1r1;
  input rd_1a;
  input reset;
  wire [2:0] wf_0;
  wire [2:0] wt_0;
  wire [2:0] df_0;
  wire [2:0] dt_0;
  wire wc_0;
  wire [2:0] wacks_0;
  wire [2:0] wenr_0;
  wire [2:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [2:0] drlgf_0;
  wire [2:0] drlgt_0;
  wire [2:0] comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [2:0] conwgit_0;
  wire [2:0] conwgif_0;
  wire conwig_0;
  wire [1:0] simp591_0;
  wire [1:0] simp681_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I5 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I6 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I7 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I8 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I9 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  NOR2 I10 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I11 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I12 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR3 I13 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I14 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I15 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  AO22 I16 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I17 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I18 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  OR2 I19 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I20 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I21 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  C3 I22 (wc_0, comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  AND2 I23 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I24 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I25 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I26 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I27 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I28 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  BUFF I29 (conwigc_0, wc_0);
  AO22 I30 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I31 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I32 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I33 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I34 (wenr_0[0:0], wc_0);
  BUFF I35 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I36 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I37 (wenr_0[1:1], wc_0);
  BUFF I38 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I39 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I40 (wenr_0[2:2], wc_0);
  C3 I41 (simp591_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  BUFF I42 (simp591_0[1:1], wacks_0[2:2]);
  C2 I43 (wd_0r, simp591_0[0:0], simp591_0[1:1]);
  AND2 I44 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I45 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I46 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I47 (rd_1r0, df_0[0:0], rg_1r);
  AND2 I48 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I49 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I50 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I51 (rd_1r1, dt_0[0:0], rg_1r);
  NOR3 I52 (simp681_0[0:0], rg_0r, rg_1r, rg_0a);
  INV I53 (simp681_0[1:1], rg_1a);
  NAND2 I54 (anyread_0, simp681_0[0:0], simp681_0[1:1]);
  BUFF I55 (wg_0a, wd_0a);
  BUFF I56 (rg_0a, rd_0a);
  BUFF I57 (rg_1a, rd_1a);
endmodule

// tka2x2b TeakA [Many [2,2],One 2]
module tka2x2b (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [1:0] i_0r0;
  input [1:0] i_0r1;
  output i_0a;
  input [1:0] i_1r0;
  input [1:0] i_1r1;
  output i_1a;
  output [1:0] o_0r0;
  output [1:0] o_0r1;
  input o_0a;
  input reset;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire nia_0;
  wire nia_1;
  wire selcomp_0;
  wire selcomp_1;
  wire [1:0] gfint_0;
  wire [1:0] gfint_1;
  wire [1:0] gtint_0;
  wire [1:0] gtint_1;
  wire [1:0] comp0_0;
  wire [1:0] comp1_0;
  OR2 I0 (comp0_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I1 (comp0_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  C2 I2 (selcomp_0, comp0_0[0:0], comp0_0[1:1]);
  OR2 I3 (comp1_0[0:0], i_1r0[0:0], i_1r1[0:0]);
  OR2 I4 (comp1_0[1:1], i_1r0[1:1], i_1r1[1:1]);
  C2 I5 (selcomp_1, comp1_0[0:0], comp1_0[1:1]);
  INV I6 (nia_0, i_0a);
  INV I7 (nia_1, i_1a);
  AND2 I8 (sel_0, nia_1, gsel_0);
  AND2 I9 (sel_1, nia_0, gsel_1);
  MUTEX I10 (selcomp_0, selcomp_1, gsel_0, gsel_1);
  OR2 I11 (o_0r0[0:0], gfint_0[0:0], gfint_1[0:0]);
  OR2 I12 (o_0r0[1:1], gfint_0[1:1], gfint_1[1:1]);
  OR2 I13 (o_0r1[0:0], gtint_0[0:0], gtint_1[0:0]);
  OR2 I14 (o_0r1[1:1], gtint_0[1:1], gtint_1[1:1]);
  AND2 I15 (gtint_0[0:0], sel_0, i_0r1[0:0]);
  AND2 I16 (gtint_0[1:1], sel_0, i_0r1[1:1]);
  AND2 I17 (gtint_1[0:0], sel_1, i_1r1[0:0]);
  AND2 I18 (gtint_1[1:1], sel_1, i_1r1[1:1]);
  AND2 I19 (gfint_0[0:0], sel_0, i_0r0[0:0]);
  AND2 I20 (gfint_0[1:1], sel_0, i_0r0[1:1]);
  AND2 I21 (gfint_1[0:0], sel_1, i_1r0[0:0]);
  AND2 I22 (gfint_1[1:1], sel_1, i_1r0[1:1]);
  C2R I23 (i_0a, sel_0, o_0a, reset);
  C2R I24 (i_1a, sel_1, o_0a, reset);
endmodule

// tkj34m32_2 TeakJ [Many [32,2],One 34]
module tkj34m32_2 (i_0r0, i_0r1, i_0a, i_1r0, i_1r1, i_1a, o_0r0, o_0r1, o_0a, reset);
  input [31:0] i_0r0;
  input [31:0] i_0r1;
  output i_0a;
  input [1:0] i_1r0;
  input [1:0] i_1r1;
  output i_1a;
  output [33:0] o_0r0;
  output [33:0] o_0r1;
  input o_0a;
  input reset;
  wire icomplete_0;
  wire [33:0] joinf_0;
  wire [33:0] joint_0;
  wire dcomplete_0;
  BUFF I0 (joinf_0[0:0], i_0r0[0:0]);
  BUFF I1 (joinf_0[1:1], i_0r0[1:1]);
  BUFF I2 (joinf_0[2:2], i_0r0[2:2]);
  BUFF I3 (joinf_0[3:3], i_0r0[3:3]);
  BUFF I4 (joinf_0[4:4], i_0r0[4:4]);
  BUFF I5 (joinf_0[5:5], i_0r0[5:5]);
  BUFF I6 (joinf_0[6:6], i_0r0[6:6]);
  BUFF I7 (joinf_0[7:7], i_0r0[7:7]);
  BUFF I8 (joinf_0[8:8], i_0r0[8:8]);
  BUFF I9 (joinf_0[9:9], i_0r0[9:9]);
  BUFF I10 (joinf_0[10:10], i_0r0[10:10]);
  BUFF I11 (joinf_0[11:11], i_0r0[11:11]);
  BUFF I12 (joinf_0[12:12], i_0r0[12:12]);
  BUFF I13 (joinf_0[13:13], i_0r0[13:13]);
  BUFF I14 (joinf_0[14:14], i_0r0[14:14]);
  BUFF I15 (joinf_0[15:15], i_0r0[15:15]);
  BUFF I16 (joinf_0[16:16], i_0r0[16:16]);
  BUFF I17 (joinf_0[17:17], i_0r0[17:17]);
  BUFF I18 (joinf_0[18:18], i_0r0[18:18]);
  BUFF I19 (joinf_0[19:19], i_0r0[19:19]);
  BUFF I20 (joinf_0[20:20], i_0r0[20:20]);
  BUFF I21 (joinf_0[21:21], i_0r0[21:21]);
  BUFF I22 (joinf_0[22:22], i_0r0[22:22]);
  BUFF I23 (joinf_0[23:23], i_0r0[23:23]);
  BUFF I24 (joinf_0[24:24], i_0r0[24:24]);
  BUFF I25 (joinf_0[25:25], i_0r0[25:25]);
  BUFF I26 (joinf_0[26:26], i_0r0[26:26]);
  BUFF I27 (joinf_0[27:27], i_0r0[27:27]);
  BUFF I28 (joinf_0[28:28], i_0r0[28:28]);
  BUFF I29 (joinf_0[29:29], i_0r0[29:29]);
  BUFF I30 (joinf_0[30:30], i_0r0[30:30]);
  BUFF I31 (joinf_0[31:31], i_0r0[31:31]);
  BUFF I32 (joinf_0[32:32], i_1r0[0:0]);
  BUFF I33 (joinf_0[33:33], i_1r0[1:1]);
  BUFF I34 (joint_0[0:0], i_0r1[0:0]);
  BUFF I35 (joint_0[1:1], i_0r1[1:1]);
  BUFF I36 (joint_0[2:2], i_0r1[2:2]);
  BUFF I37 (joint_0[3:3], i_0r1[3:3]);
  BUFF I38 (joint_0[4:4], i_0r1[4:4]);
  BUFF I39 (joint_0[5:5], i_0r1[5:5]);
  BUFF I40 (joint_0[6:6], i_0r1[6:6]);
  BUFF I41 (joint_0[7:7], i_0r1[7:7]);
  BUFF I42 (joint_0[8:8], i_0r1[8:8]);
  BUFF I43 (joint_0[9:9], i_0r1[9:9]);
  BUFF I44 (joint_0[10:10], i_0r1[10:10]);
  BUFF I45 (joint_0[11:11], i_0r1[11:11]);
  BUFF I46 (joint_0[12:12], i_0r1[12:12]);
  BUFF I47 (joint_0[13:13], i_0r1[13:13]);
  BUFF I48 (joint_0[14:14], i_0r1[14:14]);
  BUFF I49 (joint_0[15:15], i_0r1[15:15]);
  BUFF I50 (joint_0[16:16], i_0r1[16:16]);
  BUFF I51 (joint_0[17:17], i_0r1[17:17]);
  BUFF I52 (joint_0[18:18], i_0r1[18:18]);
  BUFF I53 (joint_0[19:19], i_0r1[19:19]);
  BUFF I54 (joint_0[20:20], i_0r1[20:20]);
  BUFF I55 (joint_0[21:21], i_0r1[21:21]);
  BUFF I56 (joint_0[22:22], i_0r1[22:22]);
  BUFF I57 (joint_0[23:23], i_0r1[23:23]);
  BUFF I58 (joint_0[24:24], i_0r1[24:24]);
  BUFF I59 (joint_0[25:25], i_0r1[25:25]);
  BUFF I60 (joint_0[26:26], i_0r1[26:26]);
  BUFF I61 (joint_0[27:27], i_0r1[27:27]);
  BUFF I62 (joint_0[28:28], i_0r1[28:28]);
  BUFF I63 (joint_0[29:29], i_0r1[29:29]);
  BUFF I64 (joint_0[30:30], i_0r1[30:30]);
  BUFF I65 (joint_0[31:31], i_0r1[31:31]);
  BUFF I66 (joint_0[32:32], i_1r1[0:0]);
  BUFF I67 (joint_0[33:33], i_1r1[1:1]);
  OR2 I68 (dcomplete_0, i_1r0[0:0], i_1r1[0:0]);
  BUFF I69 (icomplete_0, dcomplete_0);
  C2 I70 (o_0r0[0:0], joinf_0[0:0], icomplete_0);
  C2 I71 (o_0r1[0:0], joint_0[0:0], icomplete_0);
  BUFF I72 (o_0r0[1:1], joinf_0[1:1]);
  BUFF I73 (o_0r0[2:2], joinf_0[2:2]);
  BUFF I74 (o_0r0[3:3], joinf_0[3:3]);
  BUFF I75 (o_0r0[4:4], joinf_0[4:4]);
  BUFF I76 (o_0r0[5:5], joinf_0[5:5]);
  BUFF I77 (o_0r0[6:6], joinf_0[6:6]);
  BUFF I78 (o_0r0[7:7], joinf_0[7:7]);
  BUFF I79 (o_0r0[8:8], joinf_0[8:8]);
  BUFF I80 (o_0r0[9:9], joinf_0[9:9]);
  BUFF I81 (o_0r0[10:10], joinf_0[10:10]);
  BUFF I82 (o_0r0[11:11], joinf_0[11:11]);
  BUFF I83 (o_0r0[12:12], joinf_0[12:12]);
  BUFF I84 (o_0r0[13:13], joinf_0[13:13]);
  BUFF I85 (o_0r0[14:14], joinf_0[14:14]);
  BUFF I86 (o_0r0[15:15], joinf_0[15:15]);
  BUFF I87 (o_0r0[16:16], joinf_0[16:16]);
  BUFF I88 (o_0r0[17:17], joinf_0[17:17]);
  BUFF I89 (o_0r0[18:18], joinf_0[18:18]);
  BUFF I90 (o_0r0[19:19], joinf_0[19:19]);
  BUFF I91 (o_0r0[20:20], joinf_0[20:20]);
  BUFF I92 (o_0r0[21:21], joinf_0[21:21]);
  BUFF I93 (o_0r0[22:22], joinf_0[22:22]);
  BUFF I94 (o_0r0[23:23], joinf_0[23:23]);
  BUFF I95 (o_0r0[24:24], joinf_0[24:24]);
  BUFF I96 (o_0r0[25:25], joinf_0[25:25]);
  BUFF I97 (o_0r0[26:26], joinf_0[26:26]);
  BUFF I98 (o_0r0[27:27], joinf_0[27:27]);
  BUFF I99 (o_0r0[28:28], joinf_0[28:28]);
  BUFF I100 (o_0r0[29:29], joinf_0[29:29]);
  BUFF I101 (o_0r0[30:30], joinf_0[30:30]);
  BUFF I102 (o_0r0[31:31], joinf_0[31:31]);
  BUFF I103 (o_0r0[32:32], joinf_0[32:32]);
  BUFF I104 (o_0r0[33:33], joinf_0[33:33]);
  BUFF I105 (o_0r1[1:1], joint_0[1:1]);
  BUFF I106 (o_0r1[2:2], joint_0[2:2]);
  BUFF I107 (o_0r1[3:3], joint_0[3:3]);
  BUFF I108 (o_0r1[4:4], joint_0[4:4]);
  BUFF I109 (o_0r1[5:5], joint_0[5:5]);
  BUFF I110 (o_0r1[6:6], joint_0[6:6]);
  BUFF I111 (o_0r1[7:7], joint_0[7:7]);
  BUFF I112 (o_0r1[8:8], joint_0[8:8]);
  BUFF I113 (o_0r1[9:9], joint_0[9:9]);
  BUFF I114 (o_0r1[10:10], joint_0[10:10]);
  BUFF I115 (o_0r1[11:11], joint_0[11:11]);
  BUFF I116 (o_0r1[12:12], joint_0[12:12]);
  BUFF I117 (o_0r1[13:13], joint_0[13:13]);
  BUFF I118 (o_0r1[14:14], joint_0[14:14]);
  BUFF I119 (o_0r1[15:15], joint_0[15:15]);
  BUFF I120 (o_0r1[16:16], joint_0[16:16]);
  BUFF I121 (o_0r1[17:17], joint_0[17:17]);
  BUFF I122 (o_0r1[18:18], joint_0[18:18]);
  BUFF I123 (o_0r1[19:19], joint_0[19:19]);
  BUFF I124 (o_0r1[20:20], joint_0[20:20]);
  BUFF I125 (o_0r1[21:21], joint_0[21:21]);
  BUFF I126 (o_0r1[22:22], joint_0[22:22]);
  BUFF I127 (o_0r1[23:23], joint_0[23:23]);
  BUFF I128 (o_0r1[24:24], joint_0[24:24]);
  BUFF I129 (o_0r1[25:25], joint_0[25:25]);
  BUFF I130 (o_0r1[26:26], joint_0[26:26]);
  BUFF I131 (o_0r1[27:27], joint_0[27:27]);
  BUFF I132 (o_0r1[28:28], joint_0[28:28]);
  BUFF I133 (o_0r1[29:29], joint_0[29:29]);
  BUFF I134 (o_0r1[30:30], joint_0[30:30]);
  BUFF I135 (o_0r1[31:31], joint_0[31:31]);
  BUFF I136 (o_0r1[32:32], joint_0[32:32]);
  BUFF I137 (o_0r1[33:33], joint_0[33:33]);
  BUFF I138 (i_0a, o_0a);
  BUFF I139 (i_1a, o_0a);
endmodule

// tks34_o32w2_1o0w32_2o0w32 TeakS (32+:2) [([Imp 1 0],0),([Imp 2 0],0)] [One 34,Many [32,32]]
module tks34_o32w2_1o0w32_2o0w32 (i_0r0, i_0r1, i_0a, o_0r0, o_0r1, o_0a, o_1r0, o_1r1, o_1a, reset);
  input [33:0] i_0r0;
  input [33:0] i_0r1;
  output i_0a;
  output [31:0] o_0r0;
  output [31:0] o_0r1;
  input o_0a;
  output [31:0] o_1r0;
  output [31:0] o_1r1;
  input o_1a;
  input reset;
  wire icomplete_0;
  wire sel_0;
  wire sel_1;
  wire gsel_0;
  wire gsel_1;
  wire oack_0;
  wire match0_0;
  wire match1_0;
  wire [33:0] comp_0;
  wire [11:0] simp491_0;
  wire [3:0] simp492_0;
  wire [1:0] simp493_0;
  BUFF I0 (sel_0, match0_0);
  C2 I1 (match0_0, i_0r1[32:32], i_0r0[33:33]);
  BUFF I2 (sel_1, match1_0);
  C2 I3 (match1_0, i_0r0[32:32], i_0r1[33:33]);
  C2 I4 (gsel_0, sel_0, icomplete_0);
  C2 I5 (gsel_1, sel_1, icomplete_0);
  OR2 I6 (comp_0[0:0], i_0r0[0:0], i_0r1[0:0]);
  OR2 I7 (comp_0[1:1], i_0r0[1:1], i_0r1[1:1]);
  OR2 I8 (comp_0[2:2], i_0r0[2:2], i_0r1[2:2]);
  OR2 I9 (comp_0[3:3], i_0r0[3:3], i_0r1[3:3]);
  OR2 I10 (comp_0[4:4], i_0r0[4:4], i_0r1[4:4]);
  OR2 I11 (comp_0[5:5], i_0r0[5:5], i_0r1[5:5]);
  OR2 I12 (comp_0[6:6], i_0r0[6:6], i_0r1[6:6]);
  OR2 I13 (comp_0[7:7], i_0r0[7:7], i_0r1[7:7]);
  OR2 I14 (comp_0[8:8], i_0r0[8:8], i_0r1[8:8]);
  OR2 I15 (comp_0[9:9], i_0r0[9:9], i_0r1[9:9]);
  OR2 I16 (comp_0[10:10], i_0r0[10:10], i_0r1[10:10]);
  OR2 I17 (comp_0[11:11], i_0r0[11:11], i_0r1[11:11]);
  OR2 I18 (comp_0[12:12], i_0r0[12:12], i_0r1[12:12]);
  OR2 I19 (comp_0[13:13], i_0r0[13:13], i_0r1[13:13]);
  OR2 I20 (comp_0[14:14], i_0r0[14:14], i_0r1[14:14]);
  OR2 I21 (comp_0[15:15], i_0r0[15:15], i_0r1[15:15]);
  OR2 I22 (comp_0[16:16], i_0r0[16:16], i_0r1[16:16]);
  OR2 I23 (comp_0[17:17], i_0r0[17:17], i_0r1[17:17]);
  OR2 I24 (comp_0[18:18], i_0r0[18:18], i_0r1[18:18]);
  OR2 I25 (comp_0[19:19], i_0r0[19:19], i_0r1[19:19]);
  OR2 I26 (comp_0[20:20], i_0r0[20:20], i_0r1[20:20]);
  OR2 I27 (comp_0[21:21], i_0r0[21:21], i_0r1[21:21]);
  OR2 I28 (comp_0[22:22], i_0r0[22:22], i_0r1[22:22]);
  OR2 I29 (comp_0[23:23], i_0r0[23:23], i_0r1[23:23]);
  OR2 I30 (comp_0[24:24], i_0r0[24:24], i_0r1[24:24]);
  OR2 I31 (comp_0[25:25], i_0r0[25:25], i_0r1[25:25]);
  OR2 I32 (comp_0[26:26], i_0r0[26:26], i_0r1[26:26]);
  OR2 I33 (comp_0[27:27], i_0r0[27:27], i_0r1[27:27]);
  OR2 I34 (comp_0[28:28], i_0r0[28:28], i_0r1[28:28]);
  OR2 I35 (comp_0[29:29], i_0r0[29:29], i_0r1[29:29]);
  OR2 I36 (comp_0[30:30], i_0r0[30:30], i_0r1[30:30]);
  OR2 I37 (comp_0[31:31], i_0r0[31:31], i_0r1[31:31]);
  OR2 I38 (comp_0[32:32], i_0r0[32:32], i_0r1[32:32]);
  OR2 I39 (comp_0[33:33], i_0r0[33:33], i_0r1[33:33]);
  C3 I40 (simp491_0[0:0], comp_0[0:0], comp_0[1:1], comp_0[2:2]);
  C3 I41 (simp491_0[1:1], comp_0[3:3], comp_0[4:4], comp_0[5:5]);
  C3 I42 (simp491_0[2:2], comp_0[6:6], comp_0[7:7], comp_0[8:8]);
  C3 I43 (simp491_0[3:3], comp_0[9:9], comp_0[10:10], comp_0[11:11]);
  C3 I44 (simp491_0[4:4], comp_0[12:12], comp_0[13:13], comp_0[14:14]);
  C3 I45 (simp491_0[5:5], comp_0[15:15], comp_0[16:16], comp_0[17:17]);
  C3 I46 (simp491_0[6:6], comp_0[18:18], comp_0[19:19], comp_0[20:20]);
  C3 I47 (simp491_0[7:7], comp_0[21:21], comp_0[22:22], comp_0[23:23]);
  C3 I48 (simp491_0[8:8], comp_0[24:24], comp_0[25:25], comp_0[26:26]);
  C3 I49 (simp491_0[9:9], comp_0[27:27], comp_0[28:28], comp_0[29:29]);
  C3 I50 (simp491_0[10:10], comp_0[30:30], comp_0[31:31], comp_0[32:32]);
  BUFF I51 (simp491_0[11:11], comp_0[33:33]);
  C3 I52 (simp492_0[0:0], simp491_0[0:0], simp491_0[1:1], simp491_0[2:2]);
  C3 I53 (simp492_0[1:1], simp491_0[3:3], simp491_0[4:4], simp491_0[5:5]);
  C3 I54 (simp492_0[2:2], simp491_0[6:6], simp491_0[7:7], simp491_0[8:8]);
  C3 I55 (simp492_0[3:3], simp491_0[9:9], simp491_0[10:10], simp491_0[11:11]);
  C3 I56 (simp493_0[0:0], simp492_0[0:0], simp492_0[1:1], simp492_0[2:2]);
  BUFF I57 (simp493_0[1:1], simp492_0[3:3]);
  C2 I58 (icomplete_0, simp493_0[0:0], simp493_0[1:1]);
  C2 I59 (o_0r0[0:0], i_0r0[0:0], gsel_0);
  C2 I60 (o_0r0[1:1], i_0r0[1:1], gsel_0);
  C2 I61 (o_0r0[2:2], i_0r0[2:2], gsel_0);
  C2 I62 (o_0r0[3:3], i_0r0[3:3], gsel_0);
  C2 I63 (o_0r0[4:4], i_0r0[4:4], gsel_0);
  C2 I64 (o_0r0[5:5], i_0r0[5:5], gsel_0);
  C2 I65 (o_0r0[6:6], i_0r0[6:6], gsel_0);
  C2 I66 (o_0r0[7:7], i_0r0[7:7], gsel_0);
  C2 I67 (o_0r0[8:8], i_0r0[8:8], gsel_0);
  C2 I68 (o_0r0[9:9], i_0r0[9:9], gsel_0);
  C2 I69 (o_0r0[10:10], i_0r0[10:10], gsel_0);
  C2 I70 (o_0r0[11:11], i_0r0[11:11], gsel_0);
  C2 I71 (o_0r0[12:12], i_0r0[12:12], gsel_0);
  C2 I72 (o_0r0[13:13], i_0r0[13:13], gsel_0);
  C2 I73 (o_0r0[14:14], i_0r0[14:14], gsel_0);
  C2 I74 (o_0r0[15:15], i_0r0[15:15], gsel_0);
  C2 I75 (o_0r0[16:16], i_0r0[16:16], gsel_0);
  C2 I76 (o_0r0[17:17], i_0r0[17:17], gsel_0);
  C2 I77 (o_0r0[18:18], i_0r0[18:18], gsel_0);
  C2 I78 (o_0r0[19:19], i_0r0[19:19], gsel_0);
  C2 I79 (o_0r0[20:20], i_0r0[20:20], gsel_0);
  C2 I80 (o_0r0[21:21], i_0r0[21:21], gsel_0);
  C2 I81 (o_0r0[22:22], i_0r0[22:22], gsel_0);
  C2 I82 (o_0r0[23:23], i_0r0[23:23], gsel_0);
  C2 I83 (o_0r0[24:24], i_0r0[24:24], gsel_0);
  C2 I84 (o_0r0[25:25], i_0r0[25:25], gsel_0);
  C2 I85 (o_0r0[26:26], i_0r0[26:26], gsel_0);
  C2 I86 (o_0r0[27:27], i_0r0[27:27], gsel_0);
  C2 I87 (o_0r0[28:28], i_0r0[28:28], gsel_0);
  C2 I88 (o_0r0[29:29], i_0r0[29:29], gsel_0);
  C2 I89 (o_0r0[30:30], i_0r0[30:30], gsel_0);
  C2 I90 (o_0r0[31:31], i_0r0[31:31], gsel_0);
  C2 I91 (o_1r0[0:0], i_0r0[0:0], gsel_1);
  C2 I92 (o_1r0[1:1], i_0r0[1:1], gsel_1);
  C2 I93 (o_1r0[2:2], i_0r0[2:2], gsel_1);
  C2 I94 (o_1r0[3:3], i_0r0[3:3], gsel_1);
  C2 I95 (o_1r0[4:4], i_0r0[4:4], gsel_1);
  C2 I96 (o_1r0[5:5], i_0r0[5:5], gsel_1);
  C2 I97 (o_1r0[6:6], i_0r0[6:6], gsel_1);
  C2 I98 (o_1r0[7:7], i_0r0[7:7], gsel_1);
  C2 I99 (o_1r0[8:8], i_0r0[8:8], gsel_1);
  C2 I100 (o_1r0[9:9], i_0r0[9:9], gsel_1);
  C2 I101 (o_1r0[10:10], i_0r0[10:10], gsel_1);
  C2 I102 (o_1r0[11:11], i_0r0[11:11], gsel_1);
  C2 I103 (o_1r0[12:12], i_0r0[12:12], gsel_1);
  C2 I104 (o_1r0[13:13], i_0r0[13:13], gsel_1);
  C2 I105 (o_1r0[14:14], i_0r0[14:14], gsel_1);
  C2 I106 (o_1r0[15:15], i_0r0[15:15], gsel_1);
  C2 I107 (o_1r0[16:16], i_0r0[16:16], gsel_1);
  C2 I108 (o_1r0[17:17], i_0r0[17:17], gsel_1);
  C2 I109 (o_1r0[18:18], i_0r0[18:18], gsel_1);
  C2 I110 (o_1r0[19:19], i_0r0[19:19], gsel_1);
  C2 I111 (o_1r0[20:20], i_0r0[20:20], gsel_1);
  C2 I112 (o_1r0[21:21], i_0r0[21:21], gsel_1);
  C2 I113 (o_1r0[22:22], i_0r0[22:22], gsel_1);
  C2 I114 (o_1r0[23:23], i_0r0[23:23], gsel_1);
  C2 I115 (o_1r0[24:24], i_0r0[24:24], gsel_1);
  C2 I116 (o_1r0[25:25], i_0r0[25:25], gsel_1);
  C2 I117 (o_1r0[26:26], i_0r0[26:26], gsel_1);
  C2 I118 (o_1r0[27:27], i_0r0[27:27], gsel_1);
  C2 I119 (o_1r0[28:28], i_0r0[28:28], gsel_1);
  C2 I120 (o_1r0[29:29], i_0r0[29:29], gsel_1);
  C2 I121 (o_1r0[30:30], i_0r0[30:30], gsel_1);
  C2 I122 (o_1r0[31:31], i_0r0[31:31], gsel_1);
  C2 I123 (o_0r1[0:0], i_0r1[0:0], gsel_0);
  C2 I124 (o_0r1[1:1], i_0r1[1:1], gsel_0);
  C2 I125 (o_0r1[2:2], i_0r1[2:2], gsel_0);
  C2 I126 (o_0r1[3:3], i_0r1[3:3], gsel_0);
  C2 I127 (o_0r1[4:4], i_0r1[4:4], gsel_0);
  C2 I128 (o_0r1[5:5], i_0r1[5:5], gsel_0);
  C2 I129 (o_0r1[6:6], i_0r1[6:6], gsel_0);
  C2 I130 (o_0r1[7:7], i_0r1[7:7], gsel_0);
  C2 I131 (o_0r1[8:8], i_0r1[8:8], gsel_0);
  C2 I132 (o_0r1[9:9], i_0r1[9:9], gsel_0);
  C2 I133 (o_0r1[10:10], i_0r1[10:10], gsel_0);
  C2 I134 (o_0r1[11:11], i_0r1[11:11], gsel_0);
  C2 I135 (o_0r1[12:12], i_0r1[12:12], gsel_0);
  C2 I136 (o_0r1[13:13], i_0r1[13:13], gsel_0);
  C2 I137 (o_0r1[14:14], i_0r1[14:14], gsel_0);
  C2 I138 (o_0r1[15:15], i_0r1[15:15], gsel_0);
  C2 I139 (o_0r1[16:16], i_0r1[16:16], gsel_0);
  C2 I140 (o_0r1[17:17], i_0r1[17:17], gsel_0);
  C2 I141 (o_0r1[18:18], i_0r1[18:18], gsel_0);
  C2 I142 (o_0r1[19:19], i_0r1[19:19], gsel_0);
  C2 I143 (o_0r1[20:20], i_0r1[20:20], gsel_0);
  C2 I144 (o_0r1[21:21], i_0r1[21:21], gsel_0);
  C2 I145 (o_0r1[22:22], i_0r1[22:22], gsel_0);
  C2 I146 (o_0r1[23:23], i_0r1[23:23], gsel_0);
  C2 I147 (o_0r1[24:24], i_0r1[24:24], gsel_0);
  C2 I148 (o_0r1[25:25], i_0r1[25:25], gsel_0);
  C2 I149 (o_0r1[26:26], i_0r1[26:26], gsel_0);
  C2 I150 (o_0r1[27:27], i_0r1[27:27], gsel_0);
  C2 I151 (o_0r1[28:28], i_0r1[28:28], gsel_0);
  C2 I152 (o_0r1[29:29], i_0r1[29:29], gsel_0);
  C2 I153 (o_0r1[30:30], i_0r1[30:30], gsel_0);
  C2 I154 (o_0r1[31:31], i_0r1[31:31], gsel_0);
  C2 I155 (o_1r1[0:0], i_0r1[0:0], gsel_1);
  C2 I156 (o_1r1[1:1], i_0r1[1:1], gsel_1);
  C2 I157 (o_1r1[2:2], i_0r1[2:2], gsel_1);
  C2 I158 (o_1r1[3:3], i_0r1[3:3], gsel_1);
  C2 I159 (o_1r1[4:4], i_0r1[4:4], gsel_1);
  C2 I160 (o_1r1[5:5], i_0r1[5:5], gsel_1);
  C2 I161 (o_1r1[6:6], i_0r1[6:6], gsel_1);
  C2 I162 (o_1r1[7:7], i_0r1[7:7], gsel_1);
  C2 I163 (o_1r1[8:8], i_0r1[8:8], gsel_1);
  C2 I164 (o_1r1[9:9], i_0r1[9:9], gsel_1);
  C2 I165 (o_1r1[10:10], i_0r1[10:10], gsel_1);
  C2 I166 (o_1r1[11:11], i_0r1[11:11], gsel_1);
  C2 I167 (o_1r1[12:12], i_0r1[12:12], gsel_1);
  C2 I168 (o_1r1[13:13], i_0r1[13:13], gsel_1);
  C2 I169 (o_1r1[14:14], i_0r1[14:14], gsel_1);
  C2 I170 (o_1r1[15:15], i_0r1[15:15], gsel_1);
  C2 I171 (o_1r1[16:16], i_0r1[16:16], gsel_1);
  C2 I172 (o_1r1[17:17], i_0r1[17:17], gsel_1);
  C2 I173 (o_1r1[18:18], i_0r1[18:18], gsel_1);
  C2 I174 (o_1r1[19:19], i_0r1[19:19], gsel_1);
  C2 I175 (o_1r1[20:20], i_0r1[20:20], gsel_1);
  C2 I176 (o_1r1[21:21], i_0r1[21:21], gsel_1);
  C2 I177 (o_1r1[22:22], i_0r1[22:22], gsel_1);
  C2 I178 (o_1r1[23:23], i_0r1[23:23], gsel_1);
  C2 I179 (o_1r1[24:24], i_0r1[24:24], gsel_1);
  C2 I180 (o_1r1[25:25], i_0r1[25:25], gsel_1);
  C2 I181 (o_1r1[26:26], i_0r1[26:26], gsel_1);
  C2 I182 (o_1r1[27:27], i_0r1[27:27], gsel_1);
  C2 I183 (o_1r1[28:28], i_0r1[28:28], gsel_1);
  C2 I184 (o_1r1[29:29], i_0r1[29:29], gsel_1);
  C2 I185 (o_1r1[30:30], i_0r1[30:30], gsel_1);
  C2 I186 (o_1r1[31:31], i_0r1[31:31], gsel_1);
  OR2 I187 (oack_0, o_0a, o_1a);
  C2 I188 (i_0a, oack_0, icomplete_0);
endmodule

// tkvv65_wo0w65_ro0w65 TeakV "v" 65 [] [0] [0] [Many [65],Many [0],Many [0],Many [65]]
module tkvv65_wo0w65_ro0w65 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [64:0] wg_0r0;
  input [64:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [64:0] rd_0r0;
  output [64:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [64:0] wf_0;
  wire [64:0] wt_0;
  wire [64:0] df_0;
  wire [64:0] dt_0;
  wire wc_0;
  wire [64:0] wacks_0;
  wire [64:0] wenr_0;
  wire [64:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [64:0] drlgf_0;
  wire [64:0] drlgt_0;
  wire [64:0] comp0_0;
  wire [21:0] simp4691_0;
  wire [7:0] simp4692_0;
  wire [2:0] simp4693_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [64:0] conwgit_0;
  wire [64:0] conwgif_0;
  wire conwig_0;
  wire [21:0] simp8031_0;
  wire [7:0] simp8032_0;
  wire [2:0] simp8033_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (wen_0[32:32], wenr_0[32:32], nreset_0);
  AND2 I34 (wen_0[33:33], wenr_0[33:33], nreset_0);
  AND2 I35 (wen_0[34:34], wenr_0[34:34], nreset_0);
  AND2 I36 (wen_0[35:35], wenr_0[35:35], nreset_0);
  AND2 I37 (wen_0[36:36], wenr_0[36:36], nreset_0);
  AND2 I38 (wen_0[37:37], wenr_0[37:37], nreset_0);
  AND2 I39 (wen_0[38:38], wenr_0[38:38], nreset_0);
  AND2 I40 (wen_0[39:39], wenr_0[39:39], nreset_0);
  AND2 I41 (wen_0[40:40], wenr_0[40:40], nreset_0);
  AND2 I42 (wen_0[41:41], wenr_0[41:41], nreset_0);
  AND2 I43 (wen_0[42:42], wenr_0[42:42], nreset_0);
  AND2 I44 (wen_0[43:43], wenr_0[43:43], nreset_0);
  AND2 I45 (wen_0[44:44], wenr_0[44:44], nreset_0);
  AND2 I46 (wen_0[45:45], wenr_0[45:45], nreset_0);
  AND2 I47 (wen_0[46:46], wenr_0[46:46], nreset_0);
  AND2 I48 (wen_0[47:47], wenr_0[47:47], nreset_0);
  AND2 I49 (wen_0[48:48], wenr_0[48:48], nreset_0);
  AND2 I50 (wen_0[49:49], wenr_0[49:49], nreset_0);
  AND2 I51 (wen_0[50:50], wenr_0[50:50], nreset_0);
  AND2 I52 (wen_0[51:51], wenr_0[51:51], nreset_0);
  AND2 I53 (wen_0[52:52], wenr_0[52:52], nreset_0);
  AND2 I54 (wen_0[53:53], wenr_0[53:53], nreset_0);
  AND2 I55 (wen_0[54:54], wenr_0[54:54], nreset_0);
  AND2 I56 (wen_0[55:55], wenr_0[55:55], nreset_0);
  AND2 I57 (wen_0[56:56], wenr_0[56:56], nreset_0);
  AND2 I58 (wen_0[57:57], wenr_0[57:57], nreset_0);
  AND2 I59 (wen_0[58:58], wenr_0[58:58], nreset_0);
  AND2 I60 (wen_0[59:59], wenr_0[59:59], nreset_0);
  AND2 I61 (wen_0[60:60], wenr_0[60:60], nreset_0);
  AND2 I62 (wen_0[61:61], wenr_0[61:61], nreset_0);
  AND2 I63 (wen_0[62:62], wenr_0[62:62], nreset_0);
  AND2 I64 (wen_0[63:63], wenr_0[63:63], nreset_0);
  AND2 I65 (wen_0[64:64], wenr_0[64:64], nreset_0);
  AND2 I66 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I67 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I68 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I69 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I70 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I71 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I72 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I73 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I74 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I75 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I76 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I77 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I78 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I79 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I80 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I81 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I82 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I83 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I84 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I85 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I86 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I87 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I88 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I89 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I90 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I91 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I92 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I93 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I94 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I95 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I96 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I97 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I98 (drlgf_0[32:32], wf_0[32:32], wen_0[32:32]);
  AND2 I99 (drlgf_0[33:33], wf_0[33:33], wen_0[33:33]);
  AND2 I100 (drlgf_0[34:34], wf_0[34:34], wen_0[34:34]);
  AND2 I101 (drlgf_0[35:35], wf_0[35:35], wen_0[35:35]);
  AND2 I102 (drlgf_0[36:36], wf_0[36:36], wen_0[36:36]);
  AND2 I103 (drlgf_0[37:37], wf_0[37:37], wen_0[37:37]);
  AND2 I104 (drlgf_0[38:38], wf_0[38:38], wen_0[38:38]);
  AND2 I105 (drlgf_0[39:39], wf_0[39:39], wen_0[39:39]);
  AND2 I106 (drlgf_0[40:40], wf_0[40:40], wen_0[40:40]);
  AND2 I107 (drlgf_0[41:41], wf_0[41:41], wen_0[41:41]);
  AND2 I108 (drlgf_0[42:42], wf_0[42:42], wen_0[42:42]);
  AND2 I109 (drlgf_0[43:43], wf_0[43:43], wen_0[43:43]);
  AND2 I110 (drlgf_0[44:44], wf_0[44:44], wen_0[44:44]);
  AND2 I111 (drlgf_0[45:45], wf_0[45:45], wen_0[45:45]);
  AND2 I112 (drlgf_0[46:46], wf_0[46:46], wen_0[46:46]);
  AND2 I113 (drlgf_0[47:47], wf_0[47:47], wen_0[47:47]);
  AND2 I114 (drlgf_0[48:48], wf_0[48:48], wen_0[48:48]);
  AND2 I115 (drlgf_0[49:49], wf_0[49:49], wen_0[49:49]);
  AND2 I116 (drlgf_0[50:50], wf_0[50:50], wen_0[50:50]);
  AND2 I117 (drlgf_0[51:51], wf_0[51:51], wen_0[51:51]);
  AND2 I118 (drlgf_0[52:52], wf_0[52:52], wen_0[52:52]);
  AND2 I119 (drlgf_0[53:53], wf_0[53:53], wen_0[53:53]);
  AND2 I120 (drlgf_0[54:54], wf_0[54:54], wen_0[54:54]);
  AND2 I121 (drlgf_0[55:55], wf_0[55:55], wen_0[55:55]);
  AND2 I122 (drlgf_0[56:56], wf_0[56:56], wen_0[56:56]);
  AND2 I123 (drlgf_0[57:57], wf_0[57:57], wen_0[57:57]);
  AND2 I124 (drlgf_0[58:58], wf_0[58:58], wen_0[58:58]);
  AND2 I125 (drlgf_0[59:59], wf_0[59:59], wen_0[59:59]);
  AND2 I126 (drlgf_0[60:60], wf_0[60:60], wen_0[60:60]);
  AND2 I127 (drlgf_0[61:61], wf_0[61:61], wen_0[61:61]);
  AND2 I128 (drlgf_0[62:62], wf_0[62:62], wen_0[62:62]);
  AND2 I129 (drlgf_0[63:63], wf_0[63:63], wen_0[63:63]);
  AND2 I130 (drlgf_0[64:64], wf_0[64:64], wen_0[64:64]);
  AND2 I131 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I132 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I133 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I134 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I135 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I136 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I137 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I138 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I139 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I140 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I141 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I142 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I143 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I144 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I145 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I146 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I147 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I148 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I149 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I150 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I151 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I152 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I153 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I154 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I155 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I156 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I157 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I158 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I159 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I160 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I161 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I162 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  AND2 I163 (drlgt_0[32:32], wt_0[32:32], wen_0[32:32]);
  AND2 I164 (drlgt_0[33:33], wt_0[33:33], wen_0[33:33]);
  AND2 I165 (drlgt_0[34:34], wt_0[34:34], wen_0[34:34]);
  AND2 I166 (drlgt_0[35:35], wt_0[35:35], wen_0[35:35]);
  AND2 I167 (drlgt_0[36:36], wt_0[36:36], wen_0[36:36]);
  AND2 I168 (drlgt_0[37:37], wt_0[37:37], wen_0[37:37]);
  AND2 I169 (drlgt_0[38:38], wt_0[38:38], wen_0[38:38]);
  AND2 I170 (drlgt_0[39:39], wt_0[39:39], wen_0[39:39]);
  AND2 I171 (drlgt_0[40:40], wt_0[40:40], wen_0[40:40]);
  AND2 I172 (drlgt_0[41:41], wt_0[41:41], wen_0[41:41]);
  AND2 I173 (drlgt_0[42:42], wt_0[42:42], wen_0[42:42]);
  AND2 I174 (drlgt_0[43:43], wt_0[43:43], wen_0[43:43]);
  AND2 I175 (drlgt_0[44:44], wt_0[44:44], wen_0[44:44]);
  AND2 I176 (drlgt_0[45:45], wt_0[45:45], wen_0[45:45]);
  AND2 I177 (drlgt_0[46:46], wt_0[46:46], wen_0[46:46]);
  AND2 I178 (drlgt_0[47:47], wt_0[47:47], wen_0[47:47]);
  AND2 I179 (drlgt_0[48:48], wt_0[48:48], wen_0[48:48]);
  AND2 I180 (drlgt_0[49:49], wt_0[49:49], wen_0[49:49]);
  AND2 I181 (drlgt_0[50:50], wt_0[50:50], wen_0[50:50]);
  AND2 I182 (drlgt_0[51:51], wt_0[51:51], wen_0[51:51]);
  AND2 I183 (drlgt_0[52:52], wt_0[52:52], wen_0[52:52]);
  AND2 I184 (drlgt_0[53:53], wt_0[53:53], wen_0[53:53]);
  AND2 I185 (drlgt_0[54:54], wt_0[54:54], wen_0[54:54]);
  AND2 I186 (drlgt_0[55:55], wt_0[55:55], wen_0[55:55]);
  AND2 I187 (drlgt_0[56:56], wt_0[56:56], wen_0[56:56]);
  AND2 I188 (drlgt_0[57:57], wt_0[57:57], wen_0[57:57]);
  AND2 I189 (drlgt_0[58:58], wt_0[58:58], wen_0[58:58]);
  AND2 I190 (drlgt_0[59:59], wt_0[59:59], wen_0[59:59]);
  AND2 I191 (drlgt_0[60:60], wt_0[60:60], wen_0[60:60]);
  AND2 I192 (drlgt_0[61:61], wt_0[61:61], wen_0[61:61]);
  AND2 I193 (drlgt_0[62:62], wt_0[62:62], wen_0[62:62]);
  AND2 I194 (drlgt_0[63:63], wt_0[63:63], wen_0[63:63]);
  AND2 I195 (drlgt_0[64:64], wt_0[64:64], wen_0[64:64]);
  NOR2 I196 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I197 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I198 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I199 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I200 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I201 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I202 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I203 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I204 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I205 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I206 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I207 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I208 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I209 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I210 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I211 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I212 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I213 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I214 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I215 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I216 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I217 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I218 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I219 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I220 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I221 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I222 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I223 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I224 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I225 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I226 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I227 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR2 I228 (df_0[32:32], dt_0[32:32], drlgt_0[32:32]);
  NOR2 I229 (df_0[33:33], dt_0[33:33], drlgt_0[33:33]);
  NOR2 I230 (df_0[34:34], dt_0[34:34], drlgt_0[34:34]);
  NOR2 I231 (df_0[35:35], dt_0[35:35], drlgt_0[35:35]);
  NOR2 I232 (df_0[36:36], dt_0[36:36], drlgt_0[36:36]);
  NOR2 I233 (df_0[37:37], dt_0[37:37], drlgt_0[37:37]);
  NOR2 I234 (df_0[38:38], dt_0[38:38], drlgt_0[38:38]);
  NOR2 I235 (df_0[39:39], dt_0[39:39], drlgt_0[39:39]);
  NOR2 I236 (df_0[40:40], dt_0[40:40], drlgt_0[40:40]);
  NOR2 I237 (df_0[41:41], dt_0[41:41], drlgt_0[41:41]);
  NOR2 I238 (df_0[42:42], dt_0[42:42], drlgt_0[42:42]);
  NOR2 I239 (df_0[43:43], dt_0[43:43], drlgt_0[43:43]);
  NOR2 I240 (df_0[44:44], dt_0[44:44], drlgt_0[44:44]);
  NOR2 I241 (df_0[45:45], dt_0[45:45], drlgt_0[45:45]);
  NOR2 I242 (df_0[46:46], dt_0[46:46], drlgt_0[46:46]);
  NOR2 I243 (df_0[47:47], dt_0[47:47], drlgt_0[47:47]);
  NOR2 I244 (df_0[48:48], dt_0[48:48], drlgt_0[48:48]);
  NOR2 I245 (df_0[49:49], dt_0[49:49], drlgt_0[49:49]);
  NOR2 I246 (df_0[50:50], dt_0[50:50], drlgt_0[50:50]);
  NOR2 I247 (df_0[51:51], dt_0[51:51], drlgt_0[51:51]);
  NOR2 I248 (df_0[52:52], dt_0[52:52], drlgt_0[52:52]);
  NOR2 I249 (df_0[53:53], dt_0[53:53], drlgt_0[53:53]);
  NOR2 I250 (df_0[54:54], dt_0[54:54], drlgt_0[54:54]);
  NOR2 I251 (df_0[55:55], dt_0[55:55], drlgt_0[55:55]);
  NOR2 I252 (df_0[56:56], dt_0[56:56], drlgt_0[56:56]);
  NOR2 I253 (df_0[57:57], dt_0[57:57], drlgt_0[57:57]);
  NOR2 I254 (df_0[58:58], dt_0[58:58], drlgt_0[58:58]);
  NOR2 I255 (df_0[59:59], dt_0[59:59], drlgt_0[59:59]);
  NOR2 I256 (df_0[60:60], dt_0[60:60], drlgt_0[60:60]);
  NOR2 I257 (df_0[61:61], dt_0[61:61], drlgt_0[61:61]);
  NOR2 I258 (df_0[62:62], dt_0[62:62], drlgt_0[62:62]);
  NOR2 I259 (df_0[63:63], dt_0[63:63], drlgt_0[63:63]);
  NOR2 I260 (df_0[64:64], dt_0[64:64], drlgt_0[64:64]);
  NOR3 I261 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I262 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I263 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I264 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I265 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I266 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I267 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I268 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I269 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I270 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I271 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I272 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I273 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I274 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I275 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I276 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I277 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I278 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I279 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I280 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I281 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I282 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I283 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I284 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I285 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I286 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I287 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I288 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I289 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I290 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I291 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I292 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  NOR3 I293 (dt_0[32:32], df_0[32:32], drlgf_0[32:32], reset);
  NOR3 I294 (dt_0[33:33], df_0[33:33], drlgf_0[33:33], reset);
  NOR3 I295 (dt_0[34:34], df_0[34:34], drlgf_0[34:34], reset);
  NOR3 I296 (dt_0[35:35], df_0[35:35], drlgf_0[35:35], reset);
  NOR3 I297 (dt_0[36:36], df_0[36:36], drlgf_0[36:36], reset);
  NOR3 I298 (dt_0[37:37], df_0[37:37], drlgf_0[37:37], reset);
  NOR3 I299 (dt_0[38:38], df_0[38:38], drlgf_0[38:38], reset);
  NOR3 I300 (dt_0[39:39], df_0[39:39], drlgf_0[39:39], reset);
  NOR3 I301 (dt_0[40:40], df_0[40:40], drlgf_0[40:40], reset);
  NOR3 I302 (dt_0[41:41], df_0[41:41], drlgf_0[41:41], reset);
  NOR3 I303 (dt_0[42:42], df_0[42:42], drlgf_0[42:42], reset);
  NOR3 I304 (dt_0[43:43], df_0[43:43], drlgf_0[43:43], reset);
  NOR3 I305 (dt_0[44:44], df_0[44:44], drlgf_0[44:44], reset);
  NOR3 I306 (dt_0[45:45], df_0[45:45], drlgf_0[45:45], reset);
  NOR3 I307 (dt_0[46:46], df_0[46:46], drlgf_0[46:46], reset);
  NOR3 I308 (dt_0[47:47], df_0[47:47], drlgf_0[47:47], reset);
  NOR3 I309 (dt_0[48:48], df_0[48:48], drlgf_0[48:48], reset);
  NOR3 I310 (dt_0[49:49], df_0[49:49], drlgf_0[49:49], reset);
  NOR3 I311 (dt_0[50:50], df_0[50:50], drlgf_0[50:50], reset);
  NOR3 I312 (dt_0[51:51], df_0[51:51], drlgf_0[51:51], reset);
  NOR3 I313 (dt_0[52:52], df_0[52:52], drlgf_0[52:52], reset);
  NOR3 I314 (dt_0[53:53], df_0[53:53], drlgf_0[53:53], reset);
  NOR3 I315 (dt_0[54:54], df_0[54:54], drlgf_0[54:54], reset);
  NOR3 I316 (dt_0[55:55], df_0[55:55], drlgf_0[55:55], reset);
  NOR3 I317 (dt_0[56:56], df_0[56:56], drlgf_0[56:56], reset);
  NOR3 I318 (dt_0[57:57], df_0[57:57], drlgf_0[57:57], reset);
  NOR3 I319 (dt_0[58:58], df_0[58:58], drlgf_0[58:58], reset);
  NOR3 I320 (dt_0[59:59], df_0[59:59], drlgf_0[59:59], reset);
  NOR3 I321 (dt_0[60:60], df_0[60:60], drlgf_0[60:60], reset);
  NOR3 I322 (dt_0[61:61], df_0[61:61], drlgf_0[61:61], reset);
  NOR3 I323 (dt_0[62:62], df_0[62:62], drlgf_0[62:62], reset);
  NOR3 I324 (dt_0[63:63], df_0[63:63], drlgf_0[63:63], reset);
  NOR3 I325 (dt_0[64:64], df_0[64:64], drlgf_0[64:64], reset);
  AO22 I326 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I327 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I328 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I329 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I330 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I331 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I332 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I333 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I334 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I335 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I336 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I337 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I338 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I339 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I340 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I341 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I342 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I343 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I344 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I345 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I346 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I347 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I348 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I349 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I350 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I351 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I352 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I353 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I354 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I355 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I356 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I357 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  AO22 I358 (wacks_0[32:32], drlgf_0[32:32], df_0[32:32], drlgt_0[32:32], dt_0[32:32]);
  AO22 I359 (wacks_0[33:33], drlgf_0[33:33], df_0[33:33], drlgt_0[33:33], dt_0[33:33]);
  AO22 I360 (wacks_0[34:34], drlgf_0[34:34], df_0[34:34], drlgt_0[34:34], dt_0[34:34]);
  AO22 I361 (wacks_0[35:35], drlgf_0[35:35], df_0[35:35], drlgt_0[35:35], dt_0[35:35]);
  AO22 I362 (wacks_0[36:36], drlgf_0[36:36], df_0[36:36], drlgt_0[36:36], dt_0[36:36]);
  AO22 I363 (wacks_0[37:37], drlgf_0[37:37], df_0[37:37], drlgt_0[37:37], dt_0[37:37]);
  AO22 I364 (wacks_0[38:38], drlgf_0[38:38], df_0[38:38], drlgt_0[38:38], dt_0[38:38]);
  AO22 I365 (wacks_0[39:39], drlgf_0[39:39], df_0[39:39], drlgt_0[39:39], dt_0[39:39]);
  AO22 I366 (wacks_0[40:40], drlgf_0[40:40], df_0[40:40], drlgt_0[40:40], dt_0[40:40]);
  AO22 I367 (wacks_0[41:41], drlgf_0[41:41], df_0[41:41], drlgt_0[41:41], dt_0[41:41]);
  AO22 I368 (wacks_0[42:42], drlgf_0[42:42], df_0[42:42], drlgt_0[42:42], dt_0[42:42]);
  AO22 I369 (wacks_0[43:43], drlgf_0[43:43], df_0[43:43], drlgt_0[43:43], dt_0[43:43]);
  AO22 I370 (wacks_0[44:44], drlgf_0[44:44], df_0[44:44], drlgt_0[44:44], dt_0[44:44]);
  AO22 I371 (wacks_0[45:45], drlgf_0[45:45], df_0[45:45], drlgt_0[45:45], dt_0[45:45]);
  AO22 I372 (wacks_0[46:46], drlgf_0[46:46], df_0[46:46], drlgt_0[46:46], dt_0[46:46]);
  AO22 I373 (wacks_0[47:47], drlgf_0[47:47], df_0[47:47], drlgt_0[47:47], dt_0[47:47]);
  AO22 I374 (wacks_0[48:48], drlgf_0[48:48], df_0[48:48], drlgt_0[48:48], dt_0[48:48]);
  AO22 I375 (wacks_0[49:49], drlgf_0[49:49], df_0[49:49], drlgt_0[49:49], dt_0[49:49]);
  AO22 I376 (wacks_0[50:50], drlgf_0[50:50], df_0[50:50], drlgt_0[50:50], dt_0[50:50]);
  AO22 I377 (wacks_0[51:51], drlgf_0[51:51], df_0[51:51], drlgt_0[51:51], dt_0[51:51]);
  AO22 I378 (wacks_0[52:52], drlgf_0[52:52], df_0[52:52], drlgt_0[52:52], dt_0[52:52]);
  AO22 I379 (wacks_0[53:53], drlgf_0[53:53], df_0[53:53], drlgt_0[53:53], dt_0[53:53]);
  AO22 I380 (wacks_0[54:54], drlgf_0[54:54], df_0[54:54], drlgt_0[54:54], dt_0[54:54]);
  AO22 I381 (wacks_0[55:55], drlgf_0[55:55], df_0[55:55], drlgt_0[55:55], dt_0[55:55]);
  AO22 I382 (wacks_0[56:56], drlgf_0[56:56], df_0[56:56], drlgt_0[56:56], dt_0[56:56]);
  AO22 I383 (wacks_0[57:57], drlgf_0[57:57], df_0[57:57], drlgt_0[57:57], dt_0[57:57]);
  AO22 I384 (wacks_0[58:58], drlgf_0[58:58], df_0[58:58], drlgt_0[58:58], dt_0[58:58]);
  AO22 I385 (wacks_0[59:59], drlgf_0[59:59], df_0[59:59], drlgt_0[59:59], dt_0[59:59]);
  AO22 I386 (wacks_0[60:60], drlgf_0[60:60], df_0[60:60], drlgt_0[60:60], dt_0[60:60]);
  AO22 I387 (wacks_0[61:61], drlgf_0[61:61], df_0[61:61], drlgt_0[61:61], dt_0[61:61]);
  AO22 I388 (wacks_0[62:62], drlgf_0[62:62], df_0[62:62], drlgt_0[62:62], dt_0[62:62]);
  AO22 I389 (wacks_0[63:63], drlgf_0[63:63], df_0[63:63], drlgt_0[63:63], dt_0[63:63]);
  AO22 I390 (wacks_0[64:64], drlgf_0[64:64], df_0[64:64], drlgt_0[64:64], dt_0[64:64]);
  OR2 I391 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I392 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I393 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I394 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I395 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I396 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I397 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I398 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I399 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I400 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I401 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I402 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I403 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I404 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I405 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I406 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I407 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I408 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I409 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I410 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I411 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I412 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I413 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I414 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I415 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I416 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I417 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I418 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I419 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I420 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I421 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I422 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  OR2 I423 (comp0_0[32:32], wg_0r0[32:32], wg_0r1[32:32]);
  OR2 I424 (comp0_0[33:33], wg_0r0[33:33], wg_0r1[33:33]);
  OR2 I425 (comp0_0[34:34], wg_0r0[34:34], wg_0r1[34:34]);
  OR2 I426 (comp0_0[35:35], wg_0r0[35:35], wg_0r1[35:35]);
  OR2 I427 (comp0_0[36:36], wg_0r0[36:36], wg_0r1[36:36]);
  OR2 I428 (comp0_0[37:37], wg_0r0[37:37], wg_0r1[37:37]);
  OR2 I429 (comp0_0[38:38], wg_0r0[38:38], wg_0r1[38:38]);
  OR2 I430 (comp0_0[39:39], wg_0r0[39:39], wg_0r1[39:39]);
  OR2 I431 (comp0_0[40:40], wg_0r0[40:40], wg_0r1[40:40]);
  OR2 I432 (comp0_0[41:41], wg_0r0[41:41], wg_0r1[41:41]);
  OR2 I433 (comp0_0[42:42], wg_0r0[42:42], wg_0r1[42:42]);
  OR2 I434 (comp0_0[43:43], wg_0r0[43:43], wg_0r1[43:43]);
  OR2 I435 (comp0_0[44:44], wg_0r0[44:44], wg_0r1[44:44]);
  OR2 I436 (comp0_0[45:45], wg_0r0[45:45], wg_0r1[45:45]);
  OR2 I437 (comp0_0[46:46], wg_0r0[46:46], wg_0r1[46:46]);
  OR2 I438 (comp0_0[47:47], wg_0r0[47:47], wg_0r1[47:47]);
  OR2 I439 (comp0_0[48:48], wg_0r0[48:48], wg_0r1[48:48]);
  OR2 I440 (comp0_0[49:49], wg_0r0[49:49], wg_0r1[49:49]);
  OR2 I441 (comp0_0[50:50], wg_0r0[50:50], wg_0r1[50:50]);
  OR2 I442 (comp0_0[51:51], wg_0r0[51:51], wg_0r1[51:51]);
  OR2 I443 (comp0_0[52:52], wg_0r0[52:52], wg_0r1[52:52]);
  OR2 I444 (comp0_0[53:53], wg_0r0[53:53], wg_0r1[53:53]);
  OR2 I445 (comp0_0[54:54], wg_0r0[54:54], wg_0r1[54:54]);
  OR2 I446 (comp0_0[55:55], wg_0r0[55:55], wg_0r1[55:55]);
  OR2 I447 (comp0_0[56:56], wg_0r0[56:56], wg_0r1[56:56]);
  OR2 I448 (comp0_0[57:57], wg_0r0[57:57], wg_0r1[57:57]);
  OR2 I449 (comp0_0[58:58], wg_0r0[58:58], wg_0r1[58:58]);
  OR2 I450 (comp0_0[59:59], wg_0r0[59:59], wg_0r1[59:59]);
  OR2 I451 (comp0_0[60:60], wg_0r0[60:60], wg_0r1[60:60]);
  OR2 I452 (comp0_0[61:61], wg_0r0[61:61], wg_0r1[61:61]);
  OR2 I453 (comp0_0[62:62], wg_0r0[62:62], wg_0r1[62:62]);
  OR2 I454 (comp0_0[63:63], wg_0r0[63:63], wg_0r1[63:63]);
  OR2 I455 (comp0_0[64:64], wg_0r0[64:64], wg_0r1[64:64]);
  C3 I456 (simp4691_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I457 (simp4691_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I458 (simp4691_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I459 (simp4691_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I460 (simp4691_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I461 (simp4691_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I462 (simp4691_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I463 (simp4691_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I464 (simp4691_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I465 (simp4691_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C3 I466 (simp4691_0[10:10], comp0_0[30:30], comp0_0[31:31], comp0_0[32:32]);
  C3 I467 (simp4691_0[11:11], comp0_0[33:33], comp0_0[34:34], comp0_0[35:35]);
  C3 I468 (simp4691_0[12:12], comp0_0[36:36], comp0_0[37:37], comp0_0[38:38]);
  C3 I469 (simp4691_0[13:13], comp0_0[39:39], comp0_0[40:40], comp0_0[41:41]);
  C3 I470 (simp4691_0[14:14], comp0_0[42:42], comp0_0[43:43], comp0_0[44:44]);
  C3 I471 (simp4691_0[15:15], comp0_0[45:45], comp0_0[46:46], comp0_0[47:47]);
  C3 I472 (simp4691_0[16:16], comp0_0[48:48], comp0_0[49:49], comp0_0[50:50]);
  C3 I473 (simp4691_0[17:17], comp0_0[51:51], comp0_0[52:52], comp0_0[53:53]);
  C3 I474 (simp4691_0[18:18], comp0_0[54:54], comp0_0[55:55], comp0_0[56:56]);
  C3 I475 (simp4691_0[19:19], comp0_0[57:57], comp0_0[58:58], comp0_0[59:59]);
  C3 I476 (simp4691_0[20:20], comp0_0[60:60], comp0_0[61:61], comp0_0[62:62]);
  C2 I477 (simp4691_0[21:21], comp0_0[63:63], comp0_0[64:64]);
  C3 I478 (simp4692_0[0:0], simp4691_0[0:0], simp4691_0[1:1], simp4691_0[2:2]);
  C3 I479 (simp4692_0[1:1], simp4691_0[3:3], simp4691_0[4:4], simp4691_0[5:5]);
  C3 I480 (simp4692_0[2:2], simp4691_0[6:6], simp4691_0[7:7], simp4691_0[8:8]);
  C3 I481 (simp4692_0[3:3], simp4691_0[9:9], simp4691_0[10:10], simp4691_0[11:11]);
  C3 I482 (simp4692_0[4:4], simp4691_0[12:12], simp4691_0[13:13], simp4691_0[14:14]);
  C3 I483 (simp4692_0[5:5], simp4691_0[15:15], simp4691_0[16:16], simp4691_0[17:17]);
  C3 I484 (simp4692_0[6:6], simp4691_0[18:18], simp4691_0[19:19], simp4691_0[20:20]);
  BUFF I485 (simp4692_0[7:7], simp4691_0[21:21]);
  C3 I486 (simp4693_0[0:0], simp4692_0[0:0], simp4692_0[1:1], simp4692_0[2:2]);
  C3 I487 (simp4693_0[1:1], simp4692_0[3:3], simp4692_0[4:4], simp4692_0[5:5]);
  C2 I488 (simp4693_0[2:2], simp4692_0[6:6], simp4692_0[7:7]);
  C3 I489 (wc_0, simp4693_0[0:0], simp4693_0[1:1], simp4693_0[2:2]);
  AND2 I490 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I491 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I492 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I493 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I494 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I495 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I496 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I497 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I498 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I499 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I500 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I501 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I502 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I503 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I504 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I505 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I506 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I507 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I508 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I509 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I510 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I511 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I512 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I513 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I514 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I515 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I516 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I517 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I518 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I519 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I520 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I521 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I522 (conwgif_0[32:32], wg_0r0[32:32], conwig_0);
  AND2 I523 (conwgif_0[33:33], wg_0r0[33:33], conwig_0);
  AND2 I524 (conwgif_0[34:34], wg_0r0[34:34], conwig_0);
  AND2 I525 (conwgif_0[35:35], wg_0r0[35:35], conwig_0);
  AND2 I526 (conwgif_0[36:36], wg_0r0[36:36], conwig_0);
  AND2 I527 (conwgif_0[37:37], wg_0r0[37:37], conwig_0);
  AND2 I528 (conwgif_0[38:38], wg_0r0[38:38], conwig_0);
  AND2 I529 (conwgif_0[39:39], wg_0r0[39:39], conwig_0);
  AND2 I530 (conwgif_0[40:40], wg_0r0[40:40], conwig_0);
  AND2 I531 (conwgif_0[41:41], wg_0r0[41:41], conwig_0);
  AND2 I532 (conwgif_0[42:42], wg_0r0[42:42], conwig_0);
  AND2 I533 (conwgif_0[43:43], wg_0r0[43:43], conwig_0);
  AND2 I534 (conwgif_0[44:44], wg_0r0[44:44], conwig_0);
  AND2 I535 (conwgif_0[45:45], wg_0r0[45:45], conwig_0);
  AND2 I536 (conwgif_0[46:46], wg_0r0[46:46], conwig_0);
  AND2 I537 (conwgif_0[47:47], wg_0r0[47:47], conwig_0);
  AND2 I538 (conwgif_0[48:48], wg_0r0[48:48], conwig_0);
  AND2 I539 (conwgif_0[49:49], wg_0r0[49:49], conwig_0);
  AND2 I540 (conwgif_0[50:50], wg_0r0[50:50], conwig_0);
  AND2 I541 (conwgif_0[51:51], wg_0r0[51:51], conwig_0);
  AND2 I542 (conwgif_0[52:52], wg_0r0[52:52], conwig_0);
  AND2 I543 (conwgif_0[53:53], wg_0r0[53:53], conwig_0);
  AND2 I544 (conwgif_0[54:54], wg_0r0[54:54], conwig_0);
  AND2 I545 (conwgif_0[55:55], wg_0r0[55:55], conwig_0);
  AND2 I546 (conwgif_0[56:56], wg_0r0[56:56], conwig_0);
  AND2 I547 (conwgif_0[57:57], wg_0r0[57:57], conwig_0);
  AND2 I548 (conwgif_0[58:58], wg_0r0[58:58], conwig_0);
  AND2 I549 (conwgif_0[59:59], wg_0r0[59:59], conwig_0);
  AND2 I550 (conwgif_0[60:60], wg_0r0[60:60], conwig_0);
  AND2 I551 (conwgif_0[61:61], wg_0r0[61:61], conwig_0);
  AND2 I552 (conwgif_0[62:62], wg_0r0[62:62], conwig_0);
  AND2 I553 (conwgif_0[63:63], wg_0r0[63:63], conwig_0);
  AND2 I554 (conwgif_0[64:64], wg_0r0[64:64], conwig_0);
  AND2 I555 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I556 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I557 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I558 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I559 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I560 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I561 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I562 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I563 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I564 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I565 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I566 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I567 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I568 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I569 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I570 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I571 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I572 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I573 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I574 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I575 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I576 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I577 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I578 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I579 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I580 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I581 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I582 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I583 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I584 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I585 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I586 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  AND2 I587 (conwgit_0[32:32], wg_0r1[32:32], conwig_0);
  AND2 I588 (conwgit_0[33:33], wg_0r1[33:33], conwig_0);
  AND2 I589 (conwgit_0[34:34], wg_0r1[34:34], conwig_0);
  AND2 I590 (conwgit_0[35:35], wg_0r1[35:35], conwig_0);
  AND2 I591 (conwgit_0[36:36], wg_0r1[36:36], conwig_0);
  AND2 I592 (conwgit_0[37:37], wg_0r1[37:37], conwig_0);
  AND2 I593 (conwgit_0[38:38], wg_0r1[38:38], conwig_0);
  AND2 I594 (conwgit_0[39:39], wg_0r1[39:39], conwig_0);
  AND2 I595 (conwgit_0[40:40], wg_0r1[40:40], conwig_0);
  AND2 I596 (conwgit_0[41:41], wg_0r1[41:41], conwig_0);
  AND2 I597 (conwgit_0[42:42], wg_0r1[42:42], conwig_0);
  AND2 I598 (conwgit_0[43:43], wg_0r1[43:43], conwig_0);
  AND2 I599 (conwgit_0[44:44], wg_0r1[44:44], conwig_0);
  AND2 I600 (conwgit_0[45:45], wg_0r1[45:45], conwig_0);
  AND2 I601 (conwgit_0[46:46], wg_0r1[46:46], conwig_0);
  AND2 I602 (conwgit_0[47:47], wg_0r1[47:47], conwig_0);
  AND2 I603 (conwgit_0[48:48], wg_0r1[48:48], conwig_0);
  AND2 I604 (conwgit_0[49:49], wg_0r1[49:49], conwig_0);
  AND2 I605 (conwgit_0[50:50], wg_0r1[50:50], conwig_0);
  AND2 I606 (conwgit_0[51:51], wg_0r1[51:51], conwig_0);
  AND2 I607 (conwgit_0[52:52], wg_0r1[52:52], conwig_0);
  AND2 I608 (conwgit_0[53:53], wg_0r1[53:53], conwig_0);
  AND2 I609 (conwgit_0[54:54], wg_0r1[54:54], conwig_0);
  AND2 I610 (conwgit_0[55:55], wg_0r1[55:55], conwig_0);
  AND2 I611 (conwgit_0[56:56], wg_0r1[56:56], conwig_0);
  AND2 I612 (conwgit_0[57:57], wg_0r1[57:57], conwig_0);
  AND2 I613 (conwgit_0[58:58], wg_0r1[58:58], conwig_0);
  AND2 I614 (conwgit_0[59:59], wg_0r1[59:59], conwig_0);
  AND2 I615 (conwgit_0[60:60], wg_0r1[60:60], conwig_0);
  AND2 I616 (conwgit_0[61:61], wg_0r1[61:61], conwig_0);
  AND2 I617 (conwgit_0[62:62], wg_0r1[62:62], conwig_0);
  AND2 I618 (conwgit_0[63:63], wg_0r1[63:63], conwig_0);
  AND2 I619 (conwgit_0[64:64], wg_0r1[64:64], conwig_0);
  BUFF I620 (conwigc_0, wc_0);
  AO22 I621 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I622 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I623 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I624 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I625 (wenr_0[0:0], wc_0);
  BUFF I626 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I627 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I628 (wenr_0[1:1], wc_0);
  BUFF I629 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I630 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I631 (wenr_0[2:2], wc_0);
  BUFF I632 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I633 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I634 (wenr_0[3:3], wc_0);
  BUFF I635 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I636 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I637 (wenr_0[4:4], wc_0);
  BUFF I638 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I639 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I640 (wenr_0[5:5], wc_0);
  BUFF I641 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I642 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I643 (wenr_0[6:6], wc_0);
  BUFF I644 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I645 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I646 (wenr_0[7:7], wc_0);
  BUFF I647 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I648 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I649 (wenr_0[8:8], wc_0);
  BUFF I650 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I651 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I652 (wenr_0[9:9], wc_0);
  BUFF I653 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I654 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I655 (wenr_0[10:10], wc_0);
  BUFF I656 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I657 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I658 (wenr_0[11:11], wc_0);
  BUFF I659 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I660 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I661 (wenr_0[12:12], wc_0);
  BUFF I662 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I663 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I664 (wenr_0[13:13], wc_0);
  BUFF I665 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I666 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I667 (wenr_0[14:14], wc_0);
  BUFF I668 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I669 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I670 (wenr_0[15:15], wc_0);
  BUFF I671 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I672 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I673 (wenr_0[16:16], wc_0);
  BUFF I674 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I675 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I676 (wenr_0[17:17], wc_0);
  BUFF I677 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I678 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I679 (wenr_0[18:18], wc_0);
  BUFF I680 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I681 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I682 (wenr_0[19:19], wc_0);
  BUFF I683 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I684 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I685 (wenr_0[20:20], wc_0);
  BUFF I686 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I687 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I688 (wenr_0[21:21], wc_0);
  BUFF I689 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I690 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I691 (wenr_0[22:22], wc_0);
  BUFF I692 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I693 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I694 (wenr_0[23:23], wc_0);
  BUFF I695 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I696 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I697 (wenr_0[24:24], wc_0);
  BUFF I698 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I699 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I700 (wenr_0[25:25], wc_0);
  BUFF I701 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I702 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I703 (wenr_0[26:26], wc_0);
  BUFF I704 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I705 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I706 (wenr_0[27:27], wc_0);
  BUFF I707 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I708 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I709 (wenr_0[28:28], wc_0);
  BUFF I710 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I711 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I712 (wenr_0[29:29], wc_0);
  BUFF I713 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I714 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I715 (wenr_0[30:30], wc_0);
  BUFF I716 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I717 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I718 (wenr_0[31:31], wc_0);
  BUFF I719 (wf_0[32:32], conwgif_0[32:32]);
  BUFF I720 (wt_0[32:32], conwgit_0[32:32]);
  BUFF I721 (wenr_0[32:32], wc_0);
  BUFF I722 (wf_0[33:33], conwgif_0[33:33]);
  BUFF I723 (wt_0[33:33], conwgit_0[33:33]);
  BUFF I724 (wenr_0[33:33], wc_0);
  BUFF I725 (wf_0[34:34], conwgif_0[34:34]);
  BUFF I726 (wt_0[34:34], conwgit_0[34:34]);
  BUFF I727 (wenr_0[34:34], wc_0);
  BUFF I728 (wf_0[35:35], conwgif_0[35:35]);
  BUFF I729 (wt_0[35:35], conwgit_0[35:35]);
  BUFF I730 (wenr_0[35:35], wc_0);
  BUFF I731 (wf_0[36:36], conwgif_0[36:36]);
  BUFF I732 (wt_0[36:36], conwgit_0[36:36]);
  BUFF I733 (wenr_0[36:36], wc_0);
  BUFF I734 (wf_0[37:37], conwgif_0[37:37]);
  BUFF I735 (wt_0[37:37], conwgit_0[37:37]);
  BUFF I736 (wenr_0[37:37], wc_0);
  BUFF I737 (wf_0[38:38], conwgif_0[38:38]);
  BUFF I738 (wt_0[38:38], conwgit_0[38:38]);
  BUFF I739 (wenr_0[38:38], wc_0);
  BUFF I740 (wf_0[39:39], conwgif_0[39:39]);
  BUFF I741 (wt_0[39:39], conwgit_0[39:39]);
  BUFF I742 (wenr_0[39:39], wc_0);
  BUFF I743 (wf_0[40:40], conwgif_0[40:40]);
  BUFF I744 (wt_0[40:40], conwgit_0[40:40]);
  BUFF I745 (wenr_0[40:40], wc_0);
  BUFF I746 (wf_0[41:41], conwgif_0[41:41]);
  BUFF I747 (wt_0[41:41], conwgit_0[41:41]);
  BUFF I748 (wenr_0[41:41], wc_0);
  BUFF I749 (wf_0[42:42], conwgif_0[42:42]);
  BUFF I750 (wt_0[42:42], conwgit_0[42:42]);
  BUFF I751 (wenr_0[42:42], wc_0);
  BUFF I752 (wf_0[43:43], conwgif_0[43:43]);
  BUFF I753 (wt_0[43:43], conwgit_0[43:43]);
  BUFF I754 (wenr_0[43:43], wc_0);
  BUFF I755 (wf_0[44:44], conwgif_0[44:44]);
  BUFF I756 (wt_0[44:44], conwgit_0[44:44]);
  BUFF I757 (wenr_0[44:44], wc_0);
  BUFF I758 (wf_0[45:45], conwgif_0[45:45]);
  BUFF I759 (wt_0[45:45], conwgit_0[45:45]);
  BUFF I760 (wenr_0[45:45], wc_0);
  BUFF I761 (wf_0[46:46], conwgif_0[46:46]);
  BUFF I762 (wt_0[46:46], conwgit_0[46:46]);
  BUFF I763 (wenr_0[46:46], wc_0);
  BUFF I764 (wf_0[47:47], conwgif_0[47:47]);
  BUFF I765 (wt_0[47:47], conwgit_0[47:47]);
  BUFF I766 (wenr_0[47:47], wc_0);
  BUFF I767 (wf_0[48:48], conwgif_0[48:48]);
  BUFF I768 (wt_0[48:48], conwgit_0[48:48]);
  BUFF I769 (wenr_0[48:48], wc_0);
  BUFF I770 (wf_0[49:49], conwgif_0[49:49]);
  BUFF I771 (wt_0[49:49], conwgit_0[49:49]);
  BUFF I772 (wenr_0[49:49], wc_0);
  BUFF I773 (wf_0[50:50], conwgif_0[50:50]);
  BUFF I774 (wt_0[50:50], conwgit_0[50:50]);
  BUFF I775 (wenr_0[50:50], wc_0);
  BUFF I776 (wf_0[51:51], conwgif_0[51:51]);
  BUFF I777 (wt_0[51:51], conwgit_0[51:51]);
  BUFF I778 (wenr_0[51:51], wc_0);
  BUFF I779 (wf_0[52:52], conwgif_0[52:52]);
  BUFF I780 (wt_0[52:52], conwgit_0[52:52]);
  BUFF I781 (wenr_0[52:52], wc_0);
  BUFF I782 (wf_0[53:53], conwgif_0[53:53]);
  BUFF I783 (wt_0[53:53], conwgit_0[53:53]);
  BUFF I784 (wenr_0[53:53], wc_0);
  BUFF I785 (wf_0[54:54], conwgif_0[54:54]);
  BUFF I786 (wt_0[54:54], conwgit_0[54:54]);
  BUFF I787 (wenr_0[54:54], wc_0);
  BUFF I788 (wf_0[55:55], conwgif_0[55:55]);
  BUFF I789 (wt_0[55:55], conwgit_0[55:55]);
  BUFF I790 (wenr_0[55:55], wc_0);
  BUFF I791 (wf_0[56:56], conwgif_0[56:56]);
  BUFF I792 (wt_0[56:56], conwgit_0[56:56]);
  BUFF I793 (wenr_0[56:56], wc_0);
  BUFF I794 (wf_0[57:57], conwgif_0[57:57]);
  BUFF I795 (wt_0[57:57], conwgit_0[57:57]);
  BUFF I796 (wenr_0[57:57], wc_0);
  BUFF I797 (wf_0[58:58], conwgif_0[58:58]);
  BUFF I798 (wt_0[58:58], conwgit_0[58:58]);
  BUFF I799 (wenr_0[58:58], wc_0);
  BUFF I800 (wf_0[59:59], conwgif_0[59:59]);
  BUFF I801 (wt_0[59:59], conwgit_0[59:59]);
  BUFF I802 (wenr_0[59:59], wc_0);
  BUFF I803 (wf_0[60:60], conwgif_0[60:60]);
  BUFF I804 (wt_0[60:60], conwgit_0[60:60]);
  BUFF I805 (wenr_0[60:60], wc_0);
  BUFF I806 (wf_0[61:61], conwgif_0[61:61]);
  BUFF I807 (wt_0[61:61], conwgit_0[61:61]);
  BUFF I808 (wenr_0[61:61], wc_0);
  BUFF I809 (wf_0[62:62], conwgif_0[62:62]);
  BUFF I810 (wt_0[62:62], conwgit_0[62:62]);
  BUFF I811 (wenr_0[62:62], wc_0);
  BUFF I812 (wf_0[63:63], conwgif_0[63:63]);
  BUFF I813 (wt_0[63:63], conwgit_0[63:63]);
  BUFF I814 (wenr_0[63:63], wc_0);
  BUFF I815 (wf_0[64:64], conwgif_0[64:64]);
  BUFF I816 (wt_0[64:64], conwgit_0[64:64]);
  BUFF I817 (wenr_0[64:64], wc_0);
  C3 I818 (simp8031_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I819 (simp8031_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I820 (simp8031_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I821 (simp8031_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I822 (simp8031_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I823 (simp8031_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I824 (simp8031_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I825 (simp8031_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I826 (simp8031_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I827 (simp8031_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I828 (simp8031_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I829 (simp8031_0[11:11], wacks_0[32:32], wacks_0[33:33], wacks_0[34:34]);
  C3 I830 (simp8031_0[12:12], wacks_0[35:35], wacks_0[36:36], wacks_0[37:37]);
  C3 I831 (simp8031_0[13:13], wacks_0[38:38], wacks_0[39:39], wacks_0[40:40]);
  C3 I832 (simp8031_0[14:14], wacks_0[41:41], wacks_0[42:42], wacks_0[43:43]);
  C3 I833 (simp8031_0[15:15], wacks_0[44:44], wacks_0[45:45], wacks_0[46:46]);
  C3 I834 (simp8031_0[16:16], wacks_0[47:47], wacks_0[48:48], wacks_0[49:49]);
  C3 I835 (simp8031_0[17:17], wacks_0[50:50], wacks_0[51:51], wacks_0[52:52]);
  C3 I836 (simp8031_0[18:18], wacks_0[53:53], wacks_0[54:54], wacks_0[55:55]);
  C3 I837 (simp8031_0[19:19], wacks_0[56:56], wacks_0[57:57], wacks_0[58:58]);
  C3 I838 (simp8031_0[20:20], wacks_0[59:59], wacks_0[60:60], wacks_0[61:61]);
  C3 I839 (simp8031_0[21:21], wacks_0[62:62], wacks_0[63:63], wacks_0[64:64]);
  C3 I840 (simp8032_0[0:0], simp8031_0[0:0], simp8031_0[1:1], simp8031_0[2:2]);
  C3 I841 (simp8032_0[1:1], simp8031_0[3:3], simp8031_0[4:4], simp8031_0[5:5]);
  C3 I842 (simp8032_0[2:2], simp8031_0[6:6], simp8031_0[7:7], simp8031_0[8:8]);
  C3 I843 (simp8032_0[3:3], simp8031_0[9:9], simp8031_0[10:10], simp8031_0[11:11]);
  C3 I844 (simp8032_0[4:4], simp8031_0[12:12], simp8031_0[13:13], simp8031_0[14:14]);
  C3 I845 (simp8032_0[5:5], simp8031_0[15:15], simp8031_0[16:16], simp8031_0[17:17]);
  C3 I846 (simp8032_0[6:6], simp8031_0[18:18], simp8031_0[19:19], simp8031_0[20:20]);
  BUFF I847 (simp8032_0[7:7], simp8031_0[21:21]);
  C3 I848 (simp8033_0[0:0], simp8032_0[0:0], simp8032_0[1:1], simp8032_0[2:2]);
  C3 I849 (simp8033_0[1:1], simp8032_0[3:3], simp8032_0[4:4], simp8032_0[5:5]);
  C2 I850 (simp8033_0[2:2], simp8032_0[6:6], simp8032_0[7:7]);
  C3 I851 (wd_0r, simp8033_0[0:0], simp8033_0[1:1], simp8033_0[2:2]);
  AND2 I852 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I853 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I854 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I855 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I856 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I857 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I858 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I859 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I860 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I861 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I862 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I863 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I864 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I865 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I866 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I867 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I868 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I869 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I870 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I871 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I872 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I873 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I874 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I875 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I876 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I877 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I878 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I879 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I880 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I881 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I882 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I883 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I884 (rd_0r0[32:32], df_0[32:32], rg_0r);
  AND2 I885 (rd_0r0[33:33], df_0[33:33], rg_0r);
  AND2 I886 (rd_0r0[34:34], df_0[34:34], rg_0r);
  AND2 I887 (rd_0r0[35:35], df_0[35:35], rg_0r);
  AND2 I888 (rd_0r0[36:36], df_0[36:36], rg_0r);
  AND2 I889 (rd_0r0[37:37], df_0[37:37], rg_0r);
  AND2 I890 (rd_0r0[38:38], df_0[38:38], rg_0r);
  AND2 I891 (rd_0r0[39:39], df_0[39:39], rg_0r);
  AND2 I892 (rd_0r0[40:40], df_0[40:40], rg_0r);
  AND2 I893 (rd_0r0[41:41], df_0[41:41], rg_0r);
  AND2 I894 (rd_0r0[42:42], df_0[42:42], rg_0r);
  AND2 I895 (rd_0r0[43:43], df_0[43:43], rg_0r);
  AND2 I896 (rd_0r0[44:44], df_0[44:44], rg_0r);
  AND2 I897 (rd_0r0[45:45], df_0[45:45], rg_0r);
  AND2 I898 (rd_0r0[46:46], df_0[46:46], rg_0r);
  AND2 I899 (rd_0r0[47:47], df_0[47:47], rg_0r);
  AND2 I900 (rd_0r0[48:48], df_0[48:48], rg_0r);
  AND2 I901 (rd_0r0[49:49], df_0[49:49], rg_0r);
  AND2 I902 (rd_0r0[50:50], df_0[50:50], rg_0r);
  AND2 I903 (rd_0r0[51:51], df_0[51:51], rg_0r);
  AND2 I904 (rd_0r0[52:52], df_0[52:52], rg_0r);
  AND2 I905 (rd_0r0[53:53], df_0[53:53], rg_0r);
  AND2 I906 (rd_0r0[54:54], df_0[54:54], rg_0r);
  AND2 I907 (rd_0r0[55:55], df_0[55:55], rg_0r);
  AND2 I908 (rd_0r0[56:56], df_0[56:56], rg_0r);
  AND2 I909 (rd_0r0[57:57], df_0[57:57], rg_0r);
  AND2 I910 (rd_0r0[58:58], df_0[58:58], rg_0r);
  AND2 I911 (rd_0r0[59:59], df_0[59:59], rg_0r);
  AND2 I912 (rd_0r0[60:60], df_0[60:60], rg_0r);
  AND2 I913 (rd_0r0[61:61], df_0[61:61], rg_0r);
  AND2 I914 (rd_0r0[62:62], df_0[62:62], rg_0r);
  AND2 I915 (rd_0r0[63:63], df_0[63:63], rg_0r);
  AND2 I916 (rd_0r0[64:64], df_0[64:64], rg_0r);
  AND2 I917 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I918 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I919 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I920 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I921 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I922 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I923 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I924 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I925 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I926 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I927 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I928 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I929 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I930 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I931 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I932 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I933 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I934 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I935 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I936 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I937 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I938 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I939 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I940 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I941 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I942 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I943 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I944 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I945 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I946 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I947 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I948 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I949 (rd_0r1[32:32], dt_0[32:32], rg_0r);
  AND2 I950 (rd_0r1[33:33], dt_0[33:33], rg_0r);
  AND2 I951 (rd_0r1[34:34], dt_0[34:34], rg_0r);
  AND2 I952 (rd_0r1[35:35], dt_0[35:35], rg_0r);
  AND2 I953 (rd_0r1[36:36], dt_0[36:36], rg_0r);
  AND2 I954 (rd_0r1[37:37], dt_0[37:37], rg_0r);
  AND2 I955 (rd_0r1[38:38], dt_0[38:38], rg_0r);
  AND2 I956 (rd_0r1[39:39], dt_0[39:39], rg_0r);
  AND2 I957 (rd_0r1[40:40], dt_0[40:40], rg_0r);
  AND2 I958 (rd_0r1[41:41], dt_0[41:41], rg_0r);
  AND2 I959 (rd_0r1[42:42], dt_0[42:42], rg_0r);
  AND2 I960 (rd_0r1[43:43], dt_0[43:43], rg_0r);
  AND2 I961 (rd_0r1[44:44], dt_0[44:44], rg_0r);
  AND2 I962 (rd_0r1[45:45], dt_0[45:45], rg_0r);
  AND2 I963 (rd_0r1[46:46], dt_0[46:46], rg_0r);
  AND2 I964 (rd_0r1[47:47], dt_0[47:47], rg_0r);
  AND2 I965 (rd_0r1[48:48], dt_0[48:48], rg_0r);
  AND2 I966 (rd_0r1[49:49], dt_0[49:49], rg_0r);
  AND2 I967 (rd_0r1[50:50], dt_0[50:50], rg_0r);
  AND2 I968 (rd_0r1[51:51], dt_0[51:51], rg_0r);
  AND2 I969 (rd_0r1[52:52], dt_0[52:52], rg_0r);
  AND2 I970 (rd_0r1[53:53], dt_0[53:53], rg_0r);
  AND2 I971 (rd_0r1[54:54], dt_0[54:54], rg_0r);
  AND2 I972 (rd_0r1[55:55], dt_0[55:55], rg_0r);
  AND2 I973 (rd_0r1[56:56], dt_0[56:56], rg_0r);
  AND2 I974 (rd_0r1[57:57], dt_0[57:57], rg_0r);
  AND2 I975 (rd_0r1[58:58], dt_0[58:58], rg_0r);
  AND2 I976 (rd_0r1[59:59], dt_0[59:59], rg_0r);
  AND2 I977 (rd_0r1[60:60], dt_0[60:60], rg_0r);
  AND2 I978 (rd_0r1[61:61], dt_0[61:61], rg_0r);
  AND2 I979 (rd_0r1[62:62], dt_0[62:62], rg_0r);
  AND2 I980 (rd_0r1[63:63], dt_0[63:63], rg_0r);
  AND2 I981 (rd_0r1[64:64], dt_0[64:64], rg_0r);
  OR2 I982 (anyread_0, rg_0r, rg_0a);
  BUFF I983 (wg_0a, wd_0a);
  BUFF I984 (rg_0a, rd_0a);
endmodule

// tkvv74_wo0w74_ro0w74 TeakV "v" 74 [] [0] [0] [Many [74],Many [0],Many [0],Many [74]]
module tkvv74_wo0w74_ro0w74 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [73:0] wg_0r0;
  input [73:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [73:0] rd_0r0;
  output [73:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [73:0] wf_0;
  wire [73:0] wt_0;
  wire [73:0] df_0;
  wire [73:0] dt_0;
  wire wc_0;
  wire [73:0] wacks_0;
  wire [73:0] wenr_0;
  wire [73:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [73:0] drlgf_0;
  wire [73:0] drlgt_0;
  wire [73:0] comp0_0;
  wire [24:0] simp5321_0;
  wire [8:0] simp5322_0;
  wire [2:0] simp5323_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [73:0] conwgit_0;
  wire [73:0] conwgif_0;
  wire conwig_0;
  wire [24:0] simp9111_0;
  wire [8:0] simp9112_0;
  wire [2:0] simp9113_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (wen_0[32:32], wenr_0[32:32], nreset_0);
  AND2 I34 (wen_0[33:33], wenr_0[33:33], nreset_0);
  AND2 I35 (wen_0[34:34], wenr_0[34:34], nreset_0);
  AND2 I36 (wen_0[35:35], wenr_0[35:35], nreset_0);
  AND2 I37 (wen_0[36:36], wenr_0[36:36], nreset_0);
  AND2 I38 (wen_0[37:37], wenr_0[37:37], nreset_0);
  AND2 I39 (wen_0[38:38], wenr_0[38:38], nreset_0);
  AND2 I40 (wen_0[39:39], wenr_0[39:39], nreset_0);
  AND2 I41 (wen_0[40:40], wenr_0[40:40], nreset_0);
  AND2 I42 (wen_0[41:41], wenr_0[41:41], nreset_0);
  AND2 I43 (wen_0[42:42], wenr_0[42:42], nreset_0);
  AND2 I44 (wen_0[43:43], wenr_0[43:43], nreset_0);
  AND2 I45 (wen_0[44:44], wenr_0[44:44], nreset_0);
  AND2 I46 (wen_0[45:45], wenr_0[45:45], nreset_0);
  AND2 I47 (wen_0[46:46], wenr_0[46:46], nreset_0);
  AND2 I48 (wen_0[47:47], wenr_0[47:47], nreset_0);
  AND2 I49 (wen_0[48:48], wenr_0[48:48], nreset_0);
  AND2 I50 (wen_0[49:49], wenr_0[49:49], nreset_0);
  AND2 I51 (wen_0[50:50], wenr_0[50:50], nreset_0);
  AND2 I52 (wen_0[51:51], wenr_0[51:51], nreset_0);
  AND2 I53 (wen_0[52:52], wenr_0[52:52], nreset_0);
  AND2 I54 (wen_0[53:53], wenr_0[53:53], nreset_0);
  AND2 I55 (wen_0[54:54], wenr_0[54:54], nreset_0);
  AND2 I56 (wen_0[55:55], wenr_0[55:55], nreset_0);
  AND2 I57 (wen_0[56:56], wenr_0[56:56], nreset_0);
  AND2 I58 (wen_0[57:57], wenr_0[57:57], nreset_0);
  AND2 I59 (wen_0[58:58], wenr_0[58:58], nreset_0);
  AND2 I60 (wen_0[59:59], wenr_0[59:59], nreset_0);
  AND2 I61 (wen_0[60:60], wenr_0[60:60], nreset_0);
  AND2 I62 (wen_0[61:61], wenr_0[61:61], nreset_0);
  AND2 I63 (wen_0[62:62], wenr_0[62:62], nreset_0);
  AND2 I64 (wen_0[63:63], wenr_0[63:63], nreset_0);
  AND2 I65 (wen_0[64:64], wenr_0[64:64], nreset_0);
  AND2 I66 (wen_0[65:65], wenr_0[65:65], nreset_0);
  AND2 I67 (wen_0[66:66], wenr_0[66:66], nreset_0);
  AND2 I68 (wen_0[67:67], wenr_0[67:67], nreset_0);
  AND2 I69 (wen_0[68:68], wenr_0[68:68], nreset_0);
  AND2 I70 (wen_0[69:69], wenr_0[69:69], nreset_0);
  AND2 I71 (wen_0[70:70], wenr_0[70:70], nreset_0);
  AND2 I72 (wen_0[71:71], wenr_0[71:71], nreset_0);
  AND2 I73 (wen_0[72:72], wenr_0[72:72], nreset_0);
  AND2 I74 (wen_0[73:73], wenr_0[73:73], nreset_0);
  AND2 I75 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I76 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I77 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I78 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I79 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I80 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I81 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I82 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I83 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I84 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I85 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I86 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I87 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I88 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I89 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I90 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I91 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I92 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I93 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I94 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I95 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I96 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I97 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I98 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I99 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I100 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I101 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I102 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I103 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I104 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I105 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I106 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I107 (drlgf_0[32:32], wf_0[32:32], wen_0[32:32]);
  AND2 I108 (drlgf_0[33:33], wf_0[33:33], wen_0[33:33]);
  AND2 I109 (drlgf_0[34:34], wf_0[34:34], wen_0[34:34]);
  AND2 I110 (drlgf_0[35:35], wf_0[35:35], wen_0[35:35]);
  AND2 I111 (drlgf_0[36:36], wf_0[36:36], wen_0[36:36]);
  AND2 I112 (drlgf_0[37:37], wf_0[37:37], wen_0[37:37]);
  AND2 I113 (drlgf_0[38:38], wf_0[38:38], wen_0[38:38]);
  AND2 I114 (drlgf_0[39:39], wf_0[39:39], wen_0[39:39]);
  AND2 I115 (drlgf_0[40:40], wf_0[40:40], wen_0[40:40]);
  AND2 I116 (drlgf_0[41:41], wf_0[41:41], wen_0[41:41]);
  AND2 I117 (drlgf_0[42:42], wf_0[42:42], wen_0[42:42]);
  AND2 I118 (drlgf_0[43:43], wf_0[43:43], wen_0[43:43]);
  AND2 I119 (drlgf_0[44:44], wf_0[44:44], wen_0[44:44]);
  AND2 I120 (drlgf_0[45:45], wf_0[45:45], wen_0[45:45]);
  AND2 I121 (drlgf_0[46:46], wf_0[46:46], wen_0[46:46]);
  AND2 I122 (drlgf_0[47:47], wf_0[47:47], wen_0[47:47]);
  AND2 I123 (drlgf_0[48:48], wf_0[48:48], wen_0[48:48]);
  AND2 I124 (drlgf_0[49:49], wf_0[49:49], wen_0[49:49]);
  AND2 I125 (drlgf_0[50:50], wf_0[50:50], wen_0[50:50]);
  AND2 I126 (drlgf_0[51:51], wf_0[51:51], wen_0[51:51]);
  AND2 I127 (drlgf_0[52:52], wf_0[52:52], wen_0[52:52]);
  AND2 I128 (drlgf_0[53:53], wf_0[53:53], wen_0[53:53]);
  AND2 I129 (drlgf_0[54:54], wf_0[54:54], wen_0[54:54]);
  AND2 I130 (drlgf_0[55:55], wf_0[55:55], wen_0[55:55]);
  AND2 I131 (drlgf_0[56:56], wf_0[56:56], wen_0[56:56]);
  AND2 I132 (drlgf_0[57:57], wf_0[57:57], wen_0[57:57]);
  AND2 I133 (drlgf_0[58:58], wf_0[58:58], wen_0[58:58]);
  AND2 I134 (drlgf_0[59:59], wf_0[59:59], wen_0[59:59]);
  AND2 I135 (drlgf_0[60:60], wf_0[60:60], wen_0[60:60]);
  AND2 I136 (drlgf_0[61:61], wf_0[61:61], wen_0[61:61]);
  AND2 I137 (drlgf_0[62:62], wf_0[62:62], wen_0[62:62]);
  AND2 I138 (drlgf_0[63:63], wf_0[63:63], wen_0[63:63]);
  AND2 I139 (drlgf_0[64:64], wf_0[64:64], wen_0[64:64]);
  AND2 I140 (drlgf_0[65:65], wf_0[65:65], wen_0[65:65]);
  AND2 I141 (drlgf_0[66:66], wf_0[66:66], wen_0[66:66]);
  AND2 I142 (drlgf_0[67:67], wf_0[67:67], wen_0[67:67]);
  AND2 I143 (drlgf_0[68:68], wf_0[68:68], wen_0[68:68]);
  AND2 I144 (drlgf_0[69:69], wf_0[69:69], wen_0[69:69]);
  AND2 I145 (drlgf_0[70:70], wf_0[70:70], wen_0[70:70]);
  AND2 I146 (drlgf_0[71:71], wf_0[71:71], wen_0[71:71]);
  AND2 I147 (drlgf_0[72:72], wf_0[72:72], wen_0[72:72]);
  AND2 I148 (drlgf_0[73:73], wf_0[73:73], wen_0[73:73]);
  AND2 I149 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I150 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I151 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I152 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I153 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I154 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I155 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I156 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I157 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I158 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I159 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I160 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I161 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I162 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I163 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I164 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I165 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I166 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I167 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I168 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I169 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I170 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I171 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I172 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I173 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I174 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I175 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I176 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I177 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I178 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I179 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I180 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  AND2 I181 (drlgt_0[32:32], wt_0[32:32], wen_0[32:32]);
  AND2 I182 (drlgt_0[33:33], wt_0[33:33], wen_0[33:33]);
  AND2 I183 (drlgt_0[34:34], wt_0[34:34], wen_0[34:34]);
  AND2 I184 (drlgt_0[35:35], wt_0[35:35], wen_0[35:35]);
  AND2 I185 (drlgt_0[36:36], wt_0[36:36], wen_0[36:36]);
  AND2 I186 (drlgt_0[37:37], wt_0[37:37], wen_0[37:37]);
  AND2 I187 (drlgt_0[38:38], wt_0[38:38], wen_0[38:38]);
  AND2 I188 (drlgt_0[39:39], wt_0[39:39], wen_0[39:39]);
  AND2 I189 (drlgt_0[40:40], wt_0[40:40], wen_0[40:40]);
  AND2 I190 (drlgt_0[41:41], wt_0[41:41], wen_0[41:41]);
  AND2 I191 (drlgt_0[42:42], wt_0[42:42], wen_0[42:42]);
  AND2 I192 (drlgt_0[43:43], wt_0[43:43], wen_0[43:43]);
  AND2 I193 (drlgt_0[44:44], wt_0[44:44], wen_0[44:44]);
  AND2 I194 (drlgt_0[45:45], wt_0[45:45], wen_0[45:45]);
  AND2 I195 (drlgt_0[46:46], wt_0[46:46], wen_0[46:46]);
  AND2 I196 (drlgt_0[47:47], wt_0[47:47], wen_0[47:47]);
  AND2 I197 (drlgt_0[48:48], wt_0[48:48], wen_0[48:48]);
  AND2 I198 (drlgt_0[49:49], wt_0[49:49], wen_0[49:49]);
  AND2 I199 (drlgt_0[50:50], wt_0[50:50], wen_0[50:50]);
  AND2 I200 (drlgt_0[51:51], wt_0[51:51], wen_0[51:51]);
  AND2 I201 (drlgt_0[52:52], wt_0[52:52], wen_0[52:52]);
  AND2 I202 (drlgt_0[53:53], wt_0[53:53], wen_0[53:53]);
  AND2 I203 (drlgt_0[54:54], wt_0[54:54], wen_0[54:54]);
  AND2 I204 (drlgt_0[55:55], wt_0[55:55], wen_0[55:55]);
  AND2 I205 (drlgt_0[56:56], wt_0[56:56], wen_0[56:56]);
  AND2 I206 (drlgt_0[57:57], wt_0[57:57], wen_0[57:57]);
  AND2 I207 (drlgt_0[58:58], wt_0[58:58], wen_0[58:58]);
  AND2 I208 (drlgt_0[59:59], wt_0[59:59], wen_0[59:59]);
  AND2 I209 (drlgt_0[60:60], wt_0[60:60], wen_0[60:60]);
  AND2 I210 (drlgt_0[61:61], wt_0[61:61], wen_0[61:61]);
  AND2 I211 (drlgt_0[62:62], wt_0[62:62], wen_0[62:62]);
  AND2 I212 (drlgt_0[63:63], wt_0[63:63], wen_0[63:63]);
  AND2 I213 (drlgt_0[64:64], wt_0[64:64], wen_0[64:64]);
  AND2 I214 (drlgt_0[65:65], wt_0[65:65], wen_0[65:65]);
  AND2 I215 (drlgt_0[66:66], wt_0[66:66], wen_0[66:66]);
  AND2 I216 (drlgt_0[67:67], wt_0[67:67], wen_0[67:67]);
  AND2 I217 (drlgt_0[68:68], wt_0[68:68], wen_0[68:68]);
  AND2 I218 (drlgt_0[69:69], wt_0[69:69], wen_0[69:69]);
  AND2 I219 (drlgt_0[70:70], wt_0[70:70], wen_0[70:70]);
  AND2 I220 (drlgt_0[71:71], wt_0[71:71], wen_0[71:71]);
  AND2 I221 (drlgt_0[72:72], wt_0[72:72], wen_0[72:72]);
  AND2 I222 (drlgt_0[73:73], wt_0[73:73], wen_0[73:73]);
  NOR2 I223 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I224 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I225 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I226 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I227 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I228 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I229 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I230 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I231 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I232 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I233 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I234 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I235 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I236 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I237 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I238 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I239 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I240 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I241 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I242 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I243 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I244 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I245 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I246 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I247 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I248 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I249 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I250 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I251 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I252 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I253 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I254 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR2 I255 (df_0[32:32], dt_0[32:32], drlgt_0[32:32]);
  NOR2 I256 (df_0[33:33], dt_0[33:33], drlgt_0[33:33]);
  NOR2 I257 (df_0[34:34], dt_0[34:34], drlgt_0[34:34]);
  NOR2 I258 (df_0[35:35], dt_0[35:35], drlgt_0[35:35]);
  NOR2 I259 (df_0[36:36], dt_0[36:36], drlgt_0[36:36]);
  NOR2 I260 (df_0[37:37], dt_0[37:37], drlgt_0[37:37]);
  NOR2 I261 (df_0[38:38], dt_0[38:38], drlgt_0[38:38]);
  NOR2 I262 (df_0[39:39], dt_0[39:39], drlgt_0[39:39]);
  NOR2 I263 (df_0[40:40], dt_0[40:40], drlgt_0[40:40]);
  NOR2 I264 (df_0[41:41], dt_0[41:41], drlgt_0[41:41]);
  NOR2 I265 (df_0[42:42], dt_0[42:42], drlgt_0[42:42]);
  NOR2 I266 (df_0[43:43], dt_0[43:43], drlgt_0[43:43]);
  NOR2 I267 (df_0[44:44], dt_0[44:44], drlgt_0[44:44]);
  NOR2 I268 (df_0[45:45], dt_0[45:45], drlgt_0[45:45]);
  NOR2 I269 (df_0[46:46], dt_0[46:46], drlgt_0[46:46]);
  NOR2 I270 (df_0[47:47], dt_0[47:47], drlgt_0[47:47]);
  NOR2 I271 (df_0[48:48], dt_0[48:48], drlgt_0[48:48]);
  NOR2 I272 (df_0[49:49], dt_0[49:49], drlgt_0[49:49]);
  NOR2 I273 (df_0[50:50], dt_0[50:50], drlgt_0[50:50]);
  NOR2 I274 (df_0[51:51], dt_0[51:51], drlgt_0[51:51]);
  NOR2 I275 (df_0[52:52], dt_0[52:52], drlgt_0[52:52]);
  NOR2 I276 (df_0[53:53], dt_0[53:53], drlgt_0[53:53]);
  NOR2 I277 (df_0[54:54], dt_0[54:54], drlgt_0[54:54]);
  NOR2 I278 (df_0[55:55], dt_0[55:55], drlgt_0[55:55]);
  NOR2 I279 (df_0[56:56], dt_0[56:56], drlgt_0[56:56]);
  NOR2 I280 (df_0[57:57], dt_0[57:57], drlgt_0[57:57]);
  NOR2 I281 (df_0[58:58], dt_0[58:58], drlgt_0[58:58]);
  NOR2 I282 (df_0[59:59], dt_0[59:59], drlgt_0[59:59]);
  NOR2 I283 (df_0[60:60], dt_0[60:60], drlgt_0[60:60]);
  NOR2 I284 (df_0[61:61], dt_0[61:61], drlgt_0[61:61]);
  NOR2 I285 (df_0[62:62], dt_0[62:62], drlgt_0[62:62]);
  NOR2 I286 (df_0[63:63], dt_0[63:63], drlgt_0[63:63]);
  NOR2 I287 (df_0[64:64], dt_0[64:64], drlgt_0[64:64]);
  NOR2 I288 (df_0[65:65], dt_0[65:65], drlgt_0[65:65]);
  NOR2 I289 (df_0[66:66], dt_0[66:66], drlgt_0[66:66]);
  NOR2 I290 (df_0[67:67], dt_0[67:67], drlgt_0[67:67]);
  NOR2 I291 (df_0[68:68], dt_0[68:68], drlgt_0[68:68]);
  NOR2 I292 (df_0[69:69], dt_0[69:69], drlgt_0[69:69]);
  NOR2 I293 (df_0[70:70], dt_0[70:70], drlgt_0[70:70]);
  NOR2 I294 (df_0[71:71], dt_0[71:71], drlgt_0[71:71]);
  NOR2 I295 (df_0[72:72], dt_0[72:72], drlgt_0[72:72]);
  NOR2 I296 (df_0[73:73], dt_0[73:73], drlgt_0[73:73]);
  NOR3 I297 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I298 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I299 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I300 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I301 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I302 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I303 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I304 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I305 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I306 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I307 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I308 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I309 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I310 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I311 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I312 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I313 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I314 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I315 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I316 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I317 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I318 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I319 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I320 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I321 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I322 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I323 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I324 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I325 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I326 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I327 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I328 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  NOR3 I329 (dt_0[32:32], df_0[32:32], drlgf_0[32:32], reset);
  NOR3 I330 (dt_0[33:33], df_0[33:33], drlgf_0[33:33], reset);
  NOR3 I331 (dt_0[34:34], df_0[34:34], drlgf_0[34:34], reset);
  NOR3 I332 (dt_0[35:35], df_0[35:35], drlgf_0[35:35], reset);
  NOR3 I333 (dt_0[36:36], df_0[36:36], drlgf_0[36:36], reset);
  NOR3 I334 (dt_0[37:37], df_0[37:37], drlgf_0[37:37], reset);
  NOR3 I335 (dt_0[38:38], df_0[38:38], drlgf_0[38:38], reset);
  NOR3 I336 (dt_0[39:39], df_0[39:39], drlgf_0[39:39], reset);
  NOR3 I337 (dt_0[40:40], df_0[40:40], drlgf_0[40:40], reset);
  NOR3 I338 (dt_0[41:41], df_0[41:41], drlgf_0[41:41], reset);
  NOR3 I339 (dt_0[42:42], df_0[42:42], drlgf_0[42:42], reset);
  NOR3 I340 (dt_0[43:43], df_0[43:43], drlgf_0[43:43], reset);
  NOR3 I341 (dt_0[44:44], df_0[44:44], drlgf_0[44:44], reset);
  NOR3 I342 (dt_0[45:45], df_0[45:45], drlgf_0[45:45], reset);
  NOR3 I343 (dt_0[46:46], df_0[46:46], drlgf_0[46:46], reset);
  NOR3 I344 (dt_0[47:47], df_0[47:47], drlgf_0[47:47], reset);
  NOR3 I345 (dt_0[48:48], df_0[48:48], drlgf_0[48:48], reset);
  NOR3 I346 (dt_0[49:49], df_0[49:49], drlgf_0[49:49], reset);
  NOR3 I347 (dt_0[50:50], df_0[50:50], drlgf_0[50:50], reset);
  NOR3 I348 (dt_0[51:51], df_0[51:51], drlgf_0[51:51], reset);
  NOR3 I349 (dt_0[52:52], df_0[52:52], drlgf_0[52:52], reset);
  NOR3 I350 (dt_0[53:53], df_0[53:53], drlgf_0[53:53], reset);
  NOR3 I351 (dt_0[54:54], df_0[54:54], drlgf_0[54:54], reset);
  NOR3 I352 (dt_0[55:55], df_0[55:55], drlgf_0[55:55], reset);
  NOR3 I353 (dt_0[56:56], df_0[56:56], drlgf_0[56:56], reset);
  NOR3 I354 (dt_0[57:57], df_0[57:57], drlgf_0[57:57], reset);
  NOR3 I355 (dt_0[58:58], df_0[58:58], drlgf_0[58:58], reset);
  NOR3 I356 (dt_0[59:59], df_0[59:59], drlgf_0[59:59], reset);
  NOR3 I357 (dt_0[60:60], df_0[60:60], drlgf_0[60:60], reset);
  NOR3 I358 (dt_0[61:61], df_0[61:61], drlgf_0[61:61], reset);
  NOR3 I359 (dt_0[62:62], df_0[62:62], drlgf_0[62:62], reset);
  NOR3 I360 (dt_0[63:63], df_0[63:63], drlgf_0[63:63], reset);
  NOR3 I361 (dt_0[64:64], df_0[64:64], drlgf_0[64:64], reset);
  NOR3 I362 (dt_0[65:65], df_0[65:65], drlgf_0[65:65], reset);
  NOR3 I363 (dt_0[66:66], df_0[66:66], drlgf_0[66:66], reset);
  NOR3 I364 (dt_0[67:67], df_0[67:67], drlgf_0[67:67], reset);
  NOR3 I365 (dt_0[68:68], df_0[68:68], drlgf_0[68:68], reset);
  NOR3 I366 (dt_0[69:69], df_0[69:69], drlgf_0[69:69], reset);
  NOR3 I367 (dt_0[70:70], df_0[70:70], drlgf_0[70:70], reset);
  NOR3 I368 (dt_0[71:71], df_0[71:71], drlgf_0[71:71], reset);
  NOR3 I369 (dt_0[72:72], df_0[72:72], drlgf_0[72:72], reset);
  NOR3 I370 (dt_0[73:73], df_0[73:73], drlgf_0[73:73], reset);
  AO22 I371 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I372 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I373 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I374 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I375 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I376 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I377 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I378 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I379 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I380 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I381 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I382 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I383 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I384 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I385 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I386 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I387 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I388 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I389 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I390 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I391 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I392 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I393 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I394 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I395 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I396 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I397 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I398 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I399 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I400 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I401 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I402 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  AO22 I403 (wacks_0[32:32], drlgf_0[32:32], df_0[32:32], drlgt_0[32:32], dt_0[32:32]);
  AO22 I404 (wacks_0[33:33], drlgf_0[33:33], df_0[33:33], drlgt_0[33:33], dt_0[33:33]);
  AO22 I405 (wacks_0[34:34], drlgf_0[34:34], df_0[34:34], drlgt_0[34:34], dt_0[34:34]);
  AO22 I406 (wacks_0[35:35], drlgf_0[35:35], df_0[35:35], drlgt_0[35:35], dt_0[35:35]);
  AO22 I407 (wacks_0[36:36], drlgf_0[36:36], df_0[36:36], drlgt_0[36:36], dt_0[36:36]);
  AO22 I408 (wacks_0[37:37], drlgf_0[37:37], df_0[37:37], drlgt_0[37:37], dt_0[37:37]);
  AO22 I409 (wacks_0[38:38], drlgf_0[38:38], df_0[38:38], drlgt_0[38:38], dt_0[38:38]);
  AO22 I410 (wacks_0[39:39], drlgf_0[39:39], df_0[39:39], drlgt_0[39:39], dt_0[39:39]);
  AO22 I411 (wacks_0[40:40], drlgf_0[40:40], df_0[40:40], drlgt_0[40:40], dt_0[40:40]);
  AO22 I412 (wacks_0[41:41], drlgf_0[41:41], df_0[41:41], drlgt_0[41:41], dt_0[41:41]);
  AO22 I413 (wacks_0[42:42], drlgf_0[42:42], df_0[42:42], drlgt_0[42:42], dt_0[42:42]);
  AO22 I414 (wacks_0[43:43], drlgf_0[43:43], df_0[43:43], drlgt_0[43:43], dt_0[43:43]);
  AO22 I415 (wacks_0[44:44], drlgf_0[44:44], df_0[44:44], drlgt_0[44:44], dt_0[44:44]);
  AO22 I416 (wacks_0[45:45], drlgf_0[45:45], df_0[45:45], drlgt_0[45:45], dt_0[45:45]);
  AO22 I417 (wacks_0[46:46], drlgf_0[46:46], df_0[46:46], drlgt_0[46:46], dt_0[46:46]);
  AO22 I418 (wacks_0[47:47], drlgf_0[47:47], df_0[47:47], drlgt_0[47:47], dt_0[47:47]);
  AO22 I419 (wacks_0[48:48], drlgf_0[48:48], df_0[48:48], drlgt_0[48:48], dt_0[48:48]);
  AO22 I420 (wacks_0[49:49], drlgf_0[49:49], df_0[49:49], drlgt_0[49:49], dt_0[49:49]);
  AO22 I421 (wacks_0[50:50], drlgf_0[50:50], df_0[50:50], drlgt_0[50:50], dt_0[50:50]);
  AO22 I422 (wacks_0[51:51], drlgf_0[51:51], df_0[51:51], drlgt_0[51:51], dt_0[51:51]);
  AO22 I423 (wacks_0[52:52], drlgf_0[52:52], df_0[52:52], drlgt_0[52:52], dt_0[52:52]);
  AO22 I424 (wacks_0[53:53], drlgf_0[53:53], df_0[53:53], drlgt_0[53:53], dt_0[53:53]);
  AO22 I425 (wacks_0[54:54], drlgf_0[54:54], df_0[54:54], drlgt_0[54:54], dt_0[54:54]);
  AO22 I426 (wacks_0[55:55], drlgf_0[55:55], df_0[55:55], drlgt_0[55:55], dt_0[55:55]);
  AO22 I427 (wacks_0[56:56], drlgf_0[56:56], df_0[56:56], drlgt_0[56:56], dt_0[56:56]);
  AO22 I428 (wacks_0[57:57], drlgf_0[57:57], df_0[57:57], drlgt_0[57:57], dt_0[57:57]);
  AO22 I429 (wacks_0[58:58], drlgf_0[58:58], df_0[58:58], drlgt_0[58:58], dt_0[58:58]);
  AO22 I430 (wacks_0[59:59], drlgf_0[59:59], df_0[59:59], drlgt_0[59:59], dt_0[59:59]);
  AO22 I431 (wacks_0[60:60], drlgf_0[60:60], df_0[60:60], drlgt_0[60:60], dt_0[60:60]);
  AO22 I432 (wacks_0[61:61], drlgf_0[61:61], df_0[61:61], drlgt_0[61:61], dt_0[61:61]);
  AO22 I433 (wacks_0[62:62], drlgf_0[62:62], df_0[62:62], drlgt_0[62:62], dt_0[62:62]);
  AO22 I434 (wacks_0[63:63], drlgf_0[63:63], df_0[63:63], drlgt_0[63:63], dt_0[63:63]);
  AO22 I435 (wacks_0[64:64], drlgf_0[64:64], df_0[64:64], drlgt_0[64:64], dt_0[64:64]);
  AO22 I436 (wacks_0[65:65], drlgf_0[65:65], df_0[65:65], drlgt_0[65:65], dt_0[65:65]);
  AO22 I437 (wacks_0[66:66], drlgf_0[66:66], df_0[66:66], drlgt_0[66:66], dt_0[66:66]);
  AO22 I438 (wacks_0[67:67], drlgf_0[67:67], df_0[67:67], drlgt_0[67:67], dt_0[67:67]);
  AO22 I439 (wacks_0[68:68], drlgf_0[68:68], df_0[68:68], drlgt_0[68:68], dt_0[68:68]);
  AO22 I440 (wacks_0[69:69], drlgf_0[69:69], df_0[69:69], drlgt_0[69:69], dt_0[69:69]);
  AO22 I441 (wacks_0[70:70], drlgf_0[70:70], df_0[70:70], drlgt_0[70:70], dt_0[70:70]);
  AO22 I442 (wacks_0[71:71], drlgf_0[71:71], df_0[71:71], drlgt_0[71:71], dt_0[71:71]);
  AO22 I443 (wacks_0[72:72], drlgf_0[72:72], df_0[72:72], drlgt_0[72:72], dt_0[72:72]);
  AO22 I444 (wacks_0[73:73], drlgf_0[73:73], df_0[73:73], drlgt_0[73:73], dt_0[73:73]);
  OR2 I445 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I446 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I447 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I448 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I449 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I450 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I451 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I452 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I453 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I454 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I455 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I456 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I457 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I458 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I459 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I460 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I461 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I462 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I463 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I464 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I465 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I466 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I467 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I468 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I469 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I470 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I471 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I472 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I473 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I474 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I475 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I476 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  OR2 I477 (comp0_0[32:32], wg_0r0[32:32], wg_0r1[32:32]);
  OR2 I478 (comp0_0[33:33], wg_0r0[33:33], wg_0r1[33:33]);
  OR2 I479 (comp0_0[34:34], wg_0r0[34:34], wg_0r1[34:34]);
  OR2 I480 (comp0_0[35:35], wg_0r0[35:35], wg_0r1[35:35]);
  OR2 I481 (comp0_0[36:36], wg_0r0[36:36], wg_0r1[36:36]);
  OR2 I482 (comp0_0[37:37], wg_0r0[37:37], wg_0r1[37:37]);
  OR2 I483 (comp0_0[38:38], wg_0r0[38:38], wg_0r1[38:38]);
  OR2 I484 (comp0_0[39:39], wg_0r0[39:39], wg_0r1[39:39]);
  OR2 I485 (comp0_0[40:40], wg_0r0[40:40], wg_0r1[40:40]);
  OR2 I486 (comp0_0[41:41], wg_0r0[41:41], wg_0r1[41:41]);
  OR2 I487 (comp0_0[42:42], wg_0r0[42:42], wg_0r1[42:42]);
  OR2 I488 (comp0_0[43:43], wg_0r0[43:43], wg_0r1[43:43]);
  OR2 I489 (comp0_0[44:44], wg_0r0[44:44], wg_0r1[44:44]);
  OR2 I490 (comp0_0[45:45], wg_0r0[45:45], wg_0r1[45:45]);
  OR2 I491 (comp0_0[46:46], wg_0r0[46:46], wg_0r1[46:46]);
  OR2 I492 (comp0_0[47:47], wg_0r0[47:47], wg_0r1[47:47]);
  OR2 I493 (comp0_0[48:48], wg_0r0[48:48], wg_0r1[48:48]);
  OR2 I494 (comp0_0[49:49], wg_0r0[49:49], wg_0r1[49:49]);
  OR2 I495 (comp0_0[50:50], wg_0r0[50:50], wg_0r1[50:50]);
  OR2 I496 (comp0_0[51:51], wg_0r0[51:51], wg_0r1[51:51]);
  OR2 I497 (comp0_0[52:52], wg_0r0[52:52], wg_0r1[52:52]);
  OR2 I498 (comp0_0[53:53], wg_0r0[53:53], wg_0r1[53:53]);
  OR2 I499 (comp0_0[54:54], wg_0r0[54:54], wg_0r1[54:54]);
  OR2 I500 (comp0_0[55:55], wg_0r0[55:55], wg_0r1[55:55]);
  OR2 I501 (comp0_0[56:56], wg_0r0[56:56], wg_0r1[56:56]);
  OR2 I502 (comp0_0[57:57], wg_0r0[57:57], wg_0r1[57:57]);
  OR2 I503 (comp0_0[58:58], wg_0r0[58:58], wg_0r1[58:58]);
  OR2 I504 (comp0_0[59:59], wg_0r0[59:59], wg_0r1[59:59]);
  OR2 I505 (comp0_0[60:60], wg_0r0[60:60], wg_0r1[60:60]);
  OR2 I506 (comp0_0[61:61], wg_0r0[61:61], wg_0r1[61:61]);
  OR2 I507 (comp0_0[62:62], wg_0r0[62:62], wg_0r1[62:62]);
  OR2 I508 (comp0_0[63:63], wg_0r0[63:63], wg_0r1[63:63]);
  OR2 I509 (comp0_0[64:64], wg_0r0[64:64], wg_0r1[64:64]);
  OR2 I510 (comp0_0[65:65], wg_0r0[65:65], wg_0r1[65:65]);
  OR2 I511 (comp0_0[66:66], wg_0r0[66:66], wg_0r1[66:66]);
  OR2 I512 (comp0_0[67:67], wg_0r0[67:67], wg_0r1[67:67]);
  OR2 I513 (comp0_0[68:68], wg_0r0[68:68], wg_0r1[68:68]);
  OR2 I514 (comp0_0[69:69], wg_0r0[69:69], wg_0r1[69:69]);
  OR2 I515 (comp0_0[70:70], wg_0r0[70:70], wg_0r1[70:70]);
  OR2 I516 (comp0_0[71:71], wg_0r0[71:71], wg_0r1[71:71]);
  OR2 I517 (comp0_0[72:72], wg_0r0[72:72], wg_0r1[72:72]);
  OR2 I518 (comp0_0[73:73], wg_0r0[73:73], wg_0r1[73:73]);
  C3 I519 (simp5321_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I520 (simp5321_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I521 (simp5321_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I522 (simp5321_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I523 (simp5321_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I524 (simp5321_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I525 (simp5321_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I526 (simp5321_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I527 (simp5321_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I528 (simp5321_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C3 I529 (simp5321_0[10:10], comp0_0[30:30], comp0_0[31:31], comp0_0[32:32]);
  C3 I530 (simp5321_0[11:11], comp0_0[33:33], comp0_0[34:34], comp0_0[35:35]);
  C3 I531 (simp5321_0[12:12], comp0_0[36:36], comp0_0[37:37], comp0_0[38:38]);
  C3 I532 (simp5321_0[13:13], comp0_0[39:39], comp0_0[40:40], comp0_0[41:41]);
  C3 I533 (simp5321_0[14:14], comp0_0[42:42], comp0_0[43:43], comp0_0[44:44]);
  C3 I534 (simp5321_0[15:15], comp0_0[45:45], comp0_0[46:46], comp0_0[47:47]);
  C3 I535 (simp5321_0[16:16], comp0_0[48:48], comp0_0[49:49], comp0_0[50:50]);
  C3 I536 (simp5321_0[17:17], comp0_0[51:51], comp0_0[52:52], comp0_0[53:53]);
  C3 I537 (simp5321_0[18:18], comp0_0[54:54], comp0_0[55:55], comp0_0[56:56]);
  C3 I538 (simp5321_0[19:19], comp0_0[57:57], comp0_0[58:58], comp0_0[59:59]);
  C3 I539 (simp5321_0[20:20], comp0_0[60:60], comp0_0[61:61], comp0_0[62:62]);
  C3 I540 (simp5321_0[21:21], comp0_0[63:63], comp0_0[64:64], comp0_0[65:65]);
  C3 I541 (simp5321_0[22:22], comp0_0[66:66], comp0_0[67:67], comp0_0[68:68]);
  C3 I542 (simp5321_0[23:23], comp0_0[69:69], comp0_0[70:70], comp0_0[71:71]);
  C2 I543 (simp5321_0[24:24], comp0_0[72:72], comp0_0[73:73]);
  C3 I544 (simp5322_0[0:0], simp5321_0[0:0], simp5321_0[1:1], simp5321_0[2:2]);
  C3 I545 (simp5322_0[1:1], simp5321_0[3:3], simp5321_0[4:4], simp5321_0[5:5]);
  C3 I546 (simp5322_0[2:2], simp5321_0[6:6], simp5321_0[7:7], simp5321_0[8:8]);
  C3 I547 (simp5322_0[3:3], simp5321_0[9:9], simp5321_0[10:10], simp5321_0[11:11]);
  C3 I548 (simp5322_0[4:4], simp5321_0[12:12], simp5321_0[13:13], simp5321_0[14:14]);
  C3 I549 (simp5322_0[5:5], simp5321_0[15:15], simp5321_0[16:16], simp5321_0[17:17]);
  C3 I550 (simp5322_0[6:6], simp5321_0[18:18], simp5321_0[19:19], simp5321_0[20:20]);
  C3 I551 (simp5322_0[7:7], simp5321_0[21:21], simp5321_0[22:22], simp5321_0[23:23]);
  BUFF I552 (simp5322_0[8:8], simp5321_0[24:24]);
  C3 I553 (simp5323_0[0:0], simp5322_0[0:0], simp5322_0[1:1], simp5322_0[2:2]);
  C3 I554 (simp5323_0[1:1], simp5322_0[3:3], simp5322_0[4:4], simp5322_0[5:5]);
  C3 I555 (simp5323_0[2:2], simp5322_0[6:6], simp5322_0[7:7], simp5322_0[8:8]);
  C3 I556 (wc_0, simp5323_0[0:0], simp5323_0[1:1], simp5323_0[2:2]);
  AND2 I557 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I558 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I559 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I560 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I561 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I562 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I563 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I564 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I565 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I566 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I567 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I568 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I569 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I570 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I571 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I572 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I573 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I574 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I575 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I576 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I577 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I578 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I579 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I580 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I581 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I582 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I583 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I584 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I585 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I586 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I587 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I588 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I589 (conwgif_0[32:32], wg_0r0[32:32], conwig_0);
  AND2 I590 (conwgif_0[33:33], wg_0r0[33:33], conwig_0);
  AND2 I591 (conwgif_0[34:34], wg_0r0[34:34], conwig_0);
  AND2 I592 (conwgif_0[35:35], wg_0r0[35:35], conwig_0);
  AND2 I593 (conwgif_0[36:36], wg_0r0[36:36], conwig_0);
  AND2 I594 (conwgif_0[37:37], wg_0r0[37:37], conwig_0);
  AND2 I595 (conwgif_0[38:38], wg_0r0[38:38], conwig_0);
  AND2 I596 (conwgif_0[39:39], wg_0r0[39:39], conwig_0);
  AND2 I597 (conwgif_0[40:40], wg_0r0[40:40], conwig_0);
  AND2 I598 (conwgif_0[41:41], wg_0r0[41:41], conwig_0);
  AND2 I599 (conwgif_0[42:42], wg_0r0[42:42], conwig_0);
  AND2 I600 (conwgif_0[43:43], wg_0r0[43:43], conwig_0);
  AND2 I601 (conwgif_0[44:44], wg_0r0[44:44], conwig_0);
  AND2 I602 (conwgif_0[45:45], wg_0r0[45:45], conwig_0);
  AND2 I603 (conwgif_0[46:46], wg_0r0[46:46], conwig_0);
  AND2 I604 (conwgif_0[47:47], wg_0r0[47:47], conwig_0);
  AND2 I605 (conwgif_0[48:48], wg_0r0[48:48], conwig_0);
  AND2 I606 (conwgif_0[49:49], wg_0r0[49:49], conwig_0);
  AND2 I607 (conwgif_0[50:50], wg_0r0[50:50], conwig_0);
  AND2 I608 (conwgif_0[51:51], wg_0r0[51:51], conwig_0);
  AND2 I609 (conwgif_0[52:52], wg_0r0[52:52], conwig_0);
  AND2 I610 (conwgif_0[53:53], wg_0r0[53:53], conwig_0);
  AND2 I611 (conwgif_0[54:54], wg_0r0[54:54], conwig_0);
  AND2 I612 (conwgif_0[55:55], wg_0r0[55:55], conwig_0);
  AND2 I613 (conwgif_0[56:56], wg_0r0[56:56], conwig_0);
  AND2 I614 (conwgif_0[57:57], wg_0r0[57:57], conwig_0);
  AND2 I615 (conwgif_0[58:58], wg_0r0[58:58], conwig_0);
  AND2 I616 (conwgif_0[59:59], wg_0r0[59:59], conwig_0);
  AND2 I617 (conwgif_0[60:60], wg_0r0[60:60], conwig_0);
  AND2 I618 (conwgif_0[61:61], wg_0r0[61:61], conwig_0);
  AND2 I619 (conwgif_0[62:62], wg_0r0[62:62], conwig_0);
  AND2 I620 (conwgif_0[63:63], wg_0r0[63:63], conwig_0);
  AND2 I621 (conwgif_0[64:64], wg_0r0[64:64], conwig_0);
  AND2 I622 (conwgif_0[65:65], wg_0r0[65:65], conwig_0);
  AND2 I623 (conwgif_0[66:66], wg_0r0[66:66], conwig_0);
  AND2 I624 (conwgif_0[67:67], wg_0r0[67:67], conwig_0);
  AND2 I625 (conwgif_0[68:68], wg_0r0[68:68], conwig_0);
  AND2 I626 (conwgif_0[69:69], wg_0r0[69:69], conwig_0);
  AND2 I627 (conwgif_0[70:70], wg_0r0[70:70], conwig_0);
  AND2 I628 (conwgif_0[71:71], wg_0r0[71:71], conwig_0);
  AND2 I629 (conwgif_0[72:72], wg_0r0[72:72], conwig_0);
  AND2 I630 (conwgif_0[73:73], wg_0r0[73:73], conwig_0);
  AND2 I631 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I632 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I633 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I634 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I635 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I636 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I637 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I638 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I639 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I640 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I641 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I642 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I643 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I644 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I645 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I646 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I647 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I648 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I649 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I650 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I651 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I652 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I653 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I654 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I655 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I656 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I657 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I658 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I659 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I660 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I661 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I662 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  AND2 I663 (conwgit_0[32:32], wg_0r1[32:32], conwig_0);
  AND2 I664 (conwgit_0[33:33], wg_0r1[33:33], conwig_0);
  AND2 I665 (conwgit_0[34:34], wg_0r1[34:34], conwig_0);
  AND2 I666 (conwgit_0[35:35], wg_0r1[35:35], conwig_0);
  AND2 I667 (conwgit_0[36:36], wg_0r1[36:36], conwig_0);
  AND2 I668 (conwgit_0[37:37], wg_0r1[37:37], conwig_0);
  AND2 I669 (conwgit_0[38:38], wg_0r1[38:38], conwig_0);
  AND2 I670 (conwgit_0[39:39], wg_0r1[39:39], conwig_0);
  AND2 I671 (conwgit_0[40:40], wg_0r1[40:40], conwig_0);
  AND2 I672 (conwgit_0[41:41], wg_0r1[41:41], conwig_0);
  AND2 I673 (conwgit_0[42:42], wg_0r1[42:42], conwig_0);
  AND2 I674 (conwgit_0[43:43], wg_0r1[43:43], conwig_0);
  AND2 I675 (conwgit_0[44:44], wg_0r1[44:44], conwig_0);
  AND2 I676 (conwgit_0[45:45], wg_0r1[45:45], conwig_0);
  AND2 I677 (conwgit_0[46:46], wg_0r1[46:46], conwig_0);
  AND2 I678 (conwgit_0[47:47], wg_0r1[47:47], conwig_0);
  AND2 I679 (conwgit_0[48:48], wg_0r1[48:48], conwig_0);
  AND2 I680 (conwgit_0[49:49], wg_0r1[49:49], conwig_0);
  AND2 I681 (conwgit_0[50:50], wg_0r1[50:50], conwig_0);
  AND2 I682 (conwgit_0[51:51], wg_0r1[51:51], conwig_0);
  AND2 I683 (conwgit_0[52:52], wg_0r1[52:52], conwig_0);
  AND2 I684 (conwgit_0[53:53], wg_0r1[53:53], conwig_0);
  AND2 I685 (conwgit_0[54:54], wg_0r1[54:54], conwig_0);
  AND2 I686 (conwgit_0[55:55], wg_0r1[55:55], conwig_0);
  AND2 I687 (conwgit_0[56:56], wg_0r1[56:56], conwig_0);
  AND2 I688 (conwgit_0[57:57], wg_0r1[57:57], conwig_0);
  AND2 I689 (conwgit_0[58:58], wg_0r1[58:58], conwig_0);
  AND2 I690 (conwgit_0[59:59], wg_0r1[59:59], conwig_0);
  AND2 I691 (conwgit_0[60:60], wg_0r1[60:60], conwig_0);
  AND2 I692 (conwgit_0[61:61], wg_0r1[61:61], conwig_0);
  AND2 I693 (conwgit_0[62:62], wg_0r1[62:62], conwig_0);
  AND2 I694 (conwgit_0[63:63], wg_0r1[63:63], conwig_0);
  AND2 I695 (conwgit_0[64:64], wg_0r1[64:64], conwig_0);
  AND2 I696 (conwgit_0[65:65], wg_0r1[65:65], conwig_0);
  AND2 I697 (conwgit_0[66:66], wg_0r1[66:66], conwig_0);
  AND2 I698 (conwgit_0[67:67], wg_0r1[67:67], conwig_0);
  AND2 I699 (conwgit_0[68:68], wg_0r1[68:68], conwig_0);
  AND2 I700 (conwgit_0[69:69], wg_0r1[69:69], conwig_0);
  AND2 I701 (conwgit_0[70:70], wg_0r1[70:70], conwig_0);
  AND2 I702 (conwgit_0[71:71], wg_0r1[71:71], conwig_0);
  AND2 I703 (conwgit_0[72:72], wg_0r1[72:72], conwig_0);
  AND2 I704 (conwgit_0[73:73], wg_0r1[73:73], conwig_0);
  BUFF I705 (conwigc_0, wc_0);
  AO22 I706 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I707 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I708 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I709 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I710 (wenr_0[0:0], wc_0);
  BUFF I711 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I712 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I713 (wenr_0[1:1], wc_0);
  BUFF I714 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I715 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I716 (wenr_0[2:2], wc_0);
  BUFF I717 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I718 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I719 (wenr_0[3:3], wc_0);
  BUFF I720 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I721 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I722 (wenr_0[4:4], wc_0);
  BUFF I723 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I724 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I725 (wenr_0[5:5], wc_0);
  BUFF I726 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I727 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I728 (wenr_0[6:6], wc_0);
  BUFF I729 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I730 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I731 (wenr_0[7:7], wc_0);
  BUFF I732 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I733 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I734 (wenr_0[8:8], wc_0);
  BUFF I735 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I736 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I737 (wenr_0[9:9], wc_0);
  BUFF I738 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I739 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I740 (wenr_0[10:10], wc_0);
  BUFF I741 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I742 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I743 (wenr_0[11:11], wc_0);
  BUFF I744 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I745 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I746 (wenr_0[12:12], wc_0);
  BUFF I747 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I748 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I749 (wenr_0[13:13], wc_0);
  BUFF I750 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I751 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I752 (wenr_0[14:14], wc_0);
  BUFF I753 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I754 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I755 (wenr_0[15:15], wc_0);
  BUFF I756 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I757 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I758 (wenr_0[16:16], wc_0);
  BUFF I759 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I760 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I761 (wenr_0[17:17], wc_0);
  BUFF I762 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I763 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I764 (wenr_0[18:18], wc_0);
  BUFF I765 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I766 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I767 (wenr_0[19:19], wc_0);
  BUFF I768 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I769 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I770 (wenr_0[20:20], wc_0);
  BUFF I771 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I772 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I773 (wenr_0[21:21], wc_0);
  BUFF I774 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I775 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I776 (wenr_0[22:22], wc_0);
  BUFF I777 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I778 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I779 (wenr_0[23:23], wc_0);
  BUFF I780 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I781 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I782 (wenr_0[24:24], wc_0);
  BUFF I783 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I784 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I785 (wenr_0[25:25], wc_0);
  BUFF I786 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I787 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I788 (wenr_0[26:26], wc_0);
  BUFF I789 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I790 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I791 (wenr_0[27:27], wc_0);
  BUFF I792 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I793 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I794 (wenr_0[28:28], wc_0);
  BUFF I795 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I796 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I797 (wenr_0[29:29], wc_0);
  BUFF I798 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I799 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I800 (wenr_0[30:30], wc_0);
  BUFF I801 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I802 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I803 (wenr_0[31:31], wc_0);
  BUFF I804 (wf_0[32:32], conwgif_0[32:32]);
  BUFF I805 (wt_0[32:32], conwgit_0[32:32]);
  BUFF I806 (wenr_0[32:32], wc_0);
  BUFF I807 (wf_0[33:33], conwgif_0[33:33]);
  BUFF I808 (wt_0[33:33], conwgit_0[33:33]);
  BUFF I809 (wenr_0[33:33], wc_0);
  BUFF I810 (wf_0[34:34], conwgif_0[34:34]);
  BUFF I811 (wt_0[34:34], conwgit_0[34:34]);
  BUFF I812 (wenr_0[34:34], wc_0);
  BUFF I813 (wf_0[35:35], conwgif_0[35:35]);
  BUFF I814 (wt_0[35:35], conwgit_0[35:35]);
  BUFF I815 (wenr_0[35:35], wc_0);
  BUFF I816 (wf_0[36:36], conwgif_0[36:36]);
  BUFF I817 (wt_0[36:36], conwgit_0[36:36]);
  BUFF I818 (wenr_0[36:36], wc_0);
  BUFF I819 (wf_0[37:37], conwgif_0[37:37]);
  BUFF I820 (wt_0[37:37], conwgit_0[37:37]);
  BUFF I821 (wenr_0[37:37], wc_0);
  BUFF I822 (wf_0[38:38], conwgif_0[38:38]);
  BUFF I823 (wt_0[38:38], conwgit_0[38:38]);
  BUFF I824 (wenr_0[38:38], wc_0);
  BUFF I825 (wf_0[39:39], conwgif_0[39:39]);
  BUFF I826 (wt_0[39:39], conwgit_0[39:39]);
  BUFF I827 (wenr_0[39:39], wc_0);
  BUFF I828 (wf_0[40:40], conwgif_0[40:40]);
  BUFF I829 (wt_0[40:40], conwgit_0[40:40]);
  BUFF I830 (wenr_0[40:40], wc_0);
  BUFF I831 (wf_0[41:41], conwgif_0[41:41]);
  BUFF I832 (wt_0[41:41], conwgit_0[41:41]);
  BUFF I833 (wenr_0[41:41], wc_0);
  BUFF I834 (wf_0[42:42], conwgif_0[42:42]);
  BUFF I835 (wt_0[42:42], conwgit_0[42:42]);
  BUFF I836 (wenr_0[42:42], wc_0);
  BUFF I837 (wf_0[43:43], conwgif_0[43:43]);
  BUFF I838 (wt_0[43:43], conwgit_0[43:43]);
  BUFF I839 (wenr_0[43:43], wc_0);
  BUFF I840 (wf_0[44:44], conwgif_0[44:44]);
  BUFF I841 (wt_0[44:44], conwgit_0[44:44]);
  BUFF I842 (wenr_0[44:44], wc_0);
  BUFF I843 (wf_0[45:45], conwgif_0[45:45]);
  BUFF I844 (wt_0[45:45], conwgit_0[45:45]);
  BUFF I845 (wenr_0[45:45], wc_0);
  BUFF I846 (wf_0[46:46], conwgif_0[46:46]);
  BUFF I847 (wt_0[46:46], conwgit_0[46:46]);
  BUFF I848 (wenr_0[46:46], wc_0);
  BUFF I849 (wf_0[47:47], conwgif_0[47:47]);
  BUFF I850 (wt_0[47:47], conwgit_0[47:47]);
  BUFF I851 (wenr_0[47:47], wc_0);
  BUFF I852 (wf_0[48:48], conwgif_0[48:48]);
  BUFF I853 (wt_0[48:48], conwgit_0[48:48]);
  BUFF I854 (wenr_0[48:48], wc_0);
  BUFF I855 (wf_0[49:49], conwgif_0[49:49]);
  BUFF I856 (wt_0[49:49], conwgit_0[49:49]);
  BUFF I857 (wenr_0[49:49], wc_0);
  BUFF I858 (wf_0[50:50], conwgif_0[50:50]);
  BUFF I859 (wt_0[50:50], conwgit_0[50:50]);
  BUFF I860 (wenr_0[50:50], wc_0);
  BUFF I861 (wf_0[51:51], conwgif_0[51:51]);
  BUFF I862 (wt_0[51:51], conwgit_0[51:51]);
  BUFF I863 (wenr_0[51:51], wc_0);
  BUFF I864 (wf_0[52:52], conwgif_0[52:52]);
  BUFF I865 (wt_0[52:52], conwgit_0[52:52]);
  BUFF I866 (wenr_0[52:52], wc_0);
  BUFF I867 (wf_0[53:53], conwgif_0[53:53]);
  BUFF I868 (wt_0[53:53], conwgit_0[53:53]);
  BUFF I869 (wenr_0[53:53], wc_0);
  BUFF I870 (wf_0[54:54], conwgif_0[54:54]);
  BUFF I871 (wt_0[54:54], conwgit_0[54:54]);
  BUFF I872 (wenr_0[54:54], wc_0);
  BUFF I873 (wf_0[55:55], conwgif_0[55:55]);
  BUFF I874 (wt_0[55:55], conwgit_0[55:55]);
  BUFF I875 (wenr_0[55:55], wc_0);
  BUFF I876 (wf_0[56:56], conwgif_0[56:56]);
  BUFF I877 (wt_0[56:56], conwgit_0[56:56]);
  BUFF I878 (wenr_0[56:56], wc_0);
  BUFF I879 (wf_0[57:57], conwgif_0[57:57]);
  BUFF I880 (wt_0[57:57], conwgit_0[57:57]);
  BUFF I881 (wenr_0[57:57], wc_0);
  BUFF I882 (wf_0[58:58], conwgif_0[58:58]);
  BUFF I883 (wt_0[58:58], conwgit_0[58:58]);
  BUFF I884 (wenr_0[58:58], wc_0);
  BUFF I885 (wf_0[59:59], conwgif_0[59:59]);
  BUFF I886 (wt_0[59:59], conwgit_0[59:59]);
  BUFF I887 (wenr_0[59:59], wc_0);
  BUFF I888 (wf_0[60:60], conwgif_0[60:60]);
  BUFF I889 (wt_0[60:60], conwgit_0[60:60]);
  BUFF I890 (wenr_0[60:60], wc_0);
  BUFF I891 (wf_0[61:61], conwgif_0[61:61]);
  BUFF I892 (wt_0[61:61], conwgit_0[61:61]);
  BUFF I893 (wenr_0[61:61], wc_0);
  BUFF I894 (wf_0[62:62], conwgif_0[62:62]);
  BUFF I895 (wt_0[62:62], conwgit_0[62:62]);
  BUFF I896 (wenr_0[62:62], wc_0);
  BUFF I897 (wf_0[63:63], conwgif_0[63:63]);
  BUFF I898 (wt_0[63:63], conwgit_0[63:63]);
  BUFF I899 (wenr_0[63:63], wc_0);
  BUFF I900 (wf_0[64:64], conwgif_0[64:64]);
  BUFF I901 (wt_0[64:64], conwgit_0[64:64]);
  BUFF I902 (wenr_0[64:64], wc_0);
  BUFF I903 (wf_0[65:65], conwgif_0[65:65]);
  BUFF I904 (wt_0[65:65], conwgit_0[65:65]);
  BUFF I905 (wenr_0[65:65], wc_0);
  BUFF I906 (wf_0[66:66], conwgif_0[66:66]);
  BUFF I907 (wt_0[66:66], conwgit_0[66:66]);
  BUFF I908 (wenr_0[66:66], wc_0);
  BUFF I909 (wf_0[67:67], conwgif_0[67:67]);
  BUFF I910 (wt_0[67:67], conwgit_0[67:67]);
  BUFF I911 (wenr_0[67:67], wc_0);
  BUFF I912 (wf_0[68:68], conwgif_0[68:68]);
  BUFF I913 (wt_0[68:68], conwgit_0[68:68]);
  BUFF I914 (wenr_0[68:68], wc_0);
  BUFF I915 (wf_0[69:69], conwgif_0[69:69]);
  BUFF I916 (wt_0[69:69], conwgit_0[69:69]);
  BUFF I917 (wenr_0[69:69], wc_0);
  BUFF I918 (wf_0[70:70], conwgif_0[70:70]);
  BUFF I919 (wt_0[70:70], conwgit_0[70:70]);
  BUFF I920 (wenr_0[70:70], wc_0);
  BUFF I921 (wf_0[71:71], conwgif_0[71:71]);
  BUFF I922 (wt_0[71:71], conwgit_0[71:71]);
  BUFF I923 (wenr_0[71:71], wc_0);
  BUFF I924 (wf_0[72:72], conwgif_0[72:72]);
  BUFF I925 (wt_0[72:72], conwgit_0[72:72]);
  BUFF I926 (wenr_0[72:72], wc_0);
  BUFF I927 (wf_0[73:73], conwgif_0[73:73]);
  BUFF I928 (wt_0[73:73], conwgit_0[73:73]);
  BUFF I929 (wenr_0[73:73], wc_0);
  C3 I930 (simp9111_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I931 (simp9111_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I932 (simp9111_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I933 (simp9111_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I934 (simp9111_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I935 (simp9111_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I936 (simp9111_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I937 (simp9111_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I938 (simp9111_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I939 (simp9111_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I940 (simp9111_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  C3 I941 (simp9111_0[11:11], wacks_0[32:32], wacks_0[33:33], wacks_0[34:34]);
  C3 I942 (simp9111_0[12:12], wacks_0[35:35], wacks_0[36:36], wacks_0[37:37]);
  C3 I943 (simp9111_0[13:13], wacks_0[38:38], wacks_0[39:39], wacks_0[40:40]);
  C3 I944 (simp9111_0[14:14], wacks_0[41:41], wacks_0[42:42], wacks_0[43:43]);
  C3 I945 (simp9111_0[15:15], wacks_0[44:44], wacks_0[45:45], wacks_0[46:46]);
  C3 I946 (simp9111_0[16:16], wacks_0[47:47], wacks_0[48:48], wacks_0[49:49]);
  C3 I947 (simp9111_0[17:17], wacks_0[50:50], wacks_0[51:51], wacks_0[52:52]);
  C3 I948 (simp9111_0[18:18], wacks_0[53:53], wacks_0[54:54], wacks_0[55:55]);
  C3 I949 (simp9111_0[19:19], wacks_0[56:56], wacks_0[57:57], wacks_0[58:58]);
  C3 I950 (simp9111_0[20:20], wacks_0[59:59], wacks_0[60:60], wacks_0[61:61]);
  C3 I951 (simp9111_0[21:21], wacks_0[62:62], wacks_0[63:63], wacks_0[64:64]);
  C3 I952 (simp9111_0[22:22], wacks_0[65:65], wacks_0[66:66], wacks_0[67:67]);
  C3 I953 (simp9111_0[23:23], wacks_0[68:68], wacks_0[69:69], wacks_0[70:70]);
  C3 I954 (simp9111_0[24:24], wacks_0[71:71], wacks_0[72:72], wacks_0[73:73]);
  C3 I955 (simp9112_0[0:0], simp9111_0[0:0], simp9111_0[1:1], simp9111_0[2:2]);
  C3 I956 (simp9112_0[1:1], simp9111_0[3:3], simp9111_0[4:4], simp9111_0[5:5]);
  C3 I957 (simp9112_0[2:2], simp9111_0[6:6], simp9111_0[7:7], simp9111_0[8:8]);
  C3 I958 (simp9112_0[3:3], simp9111_0[9:9], simp9111_0[10:10], simp9111_0[11:11]);
  C3 I959 (simp9112_0[4:4], simp9111_0[12:12], simp9111_0[13:13], simp9111_0[14:14]);
  C3 I960 (simp9112_0[5:5], simp9111_0[15:15], simp9111_0[16:16], simp9111_0[17:17]);
  C3 I961 (simp9112_0[6:6], simp9111_0[18:18], simp9111_0[19:19], simp9111_0[20:20]);
  C3 I962 (simp9112_0[7:7], simp9111_0[21:21], simp9111_0[22:22], simp9111_0[23:23]);
  BUFF I963 (simp9112_0[8:8], simp9111_0[24:24]);
  C3 I964 (simp9113_0[0:0], simp9112_0[0:0], simp9112_0[1:1], simp9112_0[2:2]);
  C3 I965 (simp9113_0[1:1], simp9112_0[3:3], simp9112_0[4:4], simp9112_0[5:5]);
  C3 I966 (simp9113_0[2:2], simp9112_0[6:6], simp9112_0[7:7], simp9112_0[8:8]);
  C3 I967 (wd_0r, simp9113_0[0:0], simp9113_0[1:1], simp9113_0[2:2]);
  AND2 I968 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I969 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I970 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I971 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I972 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I973 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I974 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I975 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I976 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I977 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I978 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I979 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I980 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I981 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I982 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I983 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I984 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I985 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I986 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I987 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I988 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I989 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I990 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I991 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I992 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I993 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I994 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I995 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I996 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I997 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I998 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I999 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I1000 (rd_0r0[32:32], df_0[32:32], rg_0r);
  AND2 I1001 (rd_0r0[33:33], df_0[33:33], rg_0r);
  AND2 I1002 (rd_0r0[34:34], df_0[34:34], rg_0r);
  AND2 I1003 (rd_0r0[35:35], df_0[35:35], rg_0r);
  AND2 I1004 (rd_0r0[36:36], df_0[36:36], rg_0r);
  AND2 I1005 (rd_0r0[37:37], df_0[37:37], rg_0r);
  AND2 I1006 (rd_0r0[38:38], df_0[38:38], rg_0r);
  AND2 I1007 (rd_0r0[39:39], df_0[39:39], rg_0r);
  AND2 I1008 (rd_0r0[40:40], df_0[40:40], rg_0r);
  AND2 I1009 (rd_0r0[41:41], df_0[41:41], rg_0r);
  AND2 I1010 (rd_0r0[42:42], df_0[42:42], rg_0r);
  AND2 I1011 (rd_0r0[43:43], df_0[43:43], rg_0r);
  AND2 I1012 (rd_0r0[44:44], df_0[44:44], rg_0r);
  AND2 I1013 (rd_0r0[45:45], df_0[45:45], rg_0r);
  AND2 I1014 (rd_0r0[46:46], df_0[46:46], rg_0r);
  AND2 I1015 (rd_0r0[47:47], df_0[47:47], rg_0r);
  AND2 I1016 (rd_0r0[48:48], df_0[48:48], rg_0r);
  AND2 I1017 (rd_0r0[49:49], df_0[49:49], rg_0r);
  AND2 I1018 (rd_0r0[50:50], df_0[50:50], rg_0r);
  AND2 I1019 (rd_0r0[51:51], df_0[51:51], rg_0r);
  AND2 I1020 (rd_0r0[52:52], df_0[52:52], rg_0r);
  AND2 I1021 (rd_0r0[53:53], df_0[53:53], rg_0r);
  AND2 I1022 (rd_0r0[54:54], df_0[54:54], rg_0r);
  AND2 I1023 (rd_0r0[55:55], df_0[55:55], rg_0r);
  AND2 I1024 (rd_0r0[56:56], df_0[56:56], rg_0r);
  AND2 I1025 (rd_0r0[57:57], df_0[57:57], rg_0r);
  AND2 I1026 (rd_0r0[58:58], df_0[58:58], rg_0r);
  AND2 I1027 (rd_0r0[59:59], df_0[59:59], rg_0r);
  AND2 I1028 (rd_0r0[60:60], df_0[60:60], rg_0r);
  AND2 I1029 (rd_0r0[61:61], df_0[61:61], rg_0r);
  AND2 I1030 (rd_0r0[62:62], df_0[62:62], rg_0r);
  AND2 I1031 (rd_0r0[63:63], df_0[63:63], rg_0r);
  AND2 I1032 (rd_0r0[64:64], df_0[64:64], rg_0r);
  AND2 I1033 (rd_0r0[65:65], df_0[65:65], rg_0r);
  AND2 I1034 (rd_0r0[66:66], df_0[66:66], rg_0r);
  AND2 I1035 (rd_0r0[67:67], df_0[67:67], rg_0r);
  AND2 I1036 (rd_0r0[68:68], df_0[68:68], rg_0r);
  AND2 I1037 (rd_0r0[69:69], df_0[69:69], rg_0r);
  AND2 I1038 (rd_0r0[70:70], df_0[70:70], rg_0r);
  AND2 I1039 (rd_0r0[71:71], df_0[71:71], rg_0r);
  AND2 I1040 (rd_0r0[72:72], df_0[72:72], rg_0r);
  AND2 I1041 (rd_0r0[73:73], df_0[73:73], rg_0r);
  AND2 I1042 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I1043 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I1044 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I1045 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I1046 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I1047 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I1048 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I1049 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I1050 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I1051 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I1052 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I1053 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I1054 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I1055 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I1056 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I1057 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I1058 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I1059 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I1060 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I1061 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I1062 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I1063 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I1064 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I1065 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I1066 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I1067 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I1068 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I1069 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I1070 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I1071 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I1072 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I1073 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I1074 (rd_0r1[32:32], dt_0[32:32], rg_0r);
  AND2 I1075 (rd_0r1[33:33], dt_0[33:33], rg_0r);
  AND2 I1076 (rd_0r1[34:34], dt_0[34:34], rg_0r);
  AND2 I1077 (rd_0r1[35:35], dt_0[35:35], rg_0r);
  AND2 I1078 (rd_0r1[36:36], dt_0[36:36], rg_0r);
  AND2 I1079 (rd_0r1[37:37], dt_0[37:37], rg_0r);
  AND2 I1080 (rd_0r1[38:38], dt_0[38:38], rg_0r);
  AND2 I1081 (rd_0r1[39:39], dt_0[39:39], rg_0r);
  AND2 I1082 (rd_0r1[40:40], dt_0[40:40], rg_0r);
  AND2 I1083 (rd_0r1[41:41], dt_0[41:41], rg_0r);
  AND2 I1084 (rd_0r1[42:42], dt_0[42:42], rg_0r);
  AND2 I1085 (rd_0r1[43:43], dt_0[43:43], rg_0r);
  AND2 I1086 (rd_0r1[44:44], dt_0[44:44], rg_0r);
  AND2 I1087 (rd_0r1[45:45], dt_0[45:45], rg_0r);
  AND2 I1088 (rd_0r1[46:46], dt_0[46:46], rg_0r);
  AND2 I1089 (rd_0r1[47:47], dt_0[47:47], rg_0r);
  AND2 I1090 (rd_0r1[48:48], dt_0[48:48], rg_0r);
  AND2 I1091 (rd_0r1[49:49], dt_0[49:49], rg_0r);
  AND2 I1092 (rd_0r1[50:50], dt_0[50:50], rg_0r);
  AND2 I1093 (rd_0r1[51:51], dt_0[51:51], rg_0r);
  AND2 I1094 (rd_0r1[52:52], dt_0[52:52], rg_0r);
  AND2 I1095 (rd_0r1[53:53], dt_0[53:53], rg_0r);
  AND2 I1096 (rd_0r1[54:54], dt_0[54:54], rg_0r);
  AND2 I1097 (rd_0r1[55:55], dt_0[55:55], rg_0r);
  AND2 I1098 (rd_0r1[56:56], dt_0[56:56], rg_0r);
  AND2 I1099 (rd_0r1[57:57], dt_0[57:57], rg_0r);
  AND2 I1100 (rd_0r1[58:58], dt_0[58:58], rg_0r);
  AND2 I1101 (rd_0r1[59:59], dt_0[59:59], rg_0r);
  AND2 I1102 (rd_0r1[60:60], dt_0[60:60], rg_0r);
  AND2 I1103 (rd_0r1[61:61], dt_0[61:61], rg_0r);
  AND2 I1104 (rd_0r1[62:62], dt_0[62:62], rg_0r);
  AND2 I1105 (rd_0r1[63:63], dt_0[63:63], rg_0r);
  AND2 I1106 (rd_0r1[64:64], dt_0[64:64], rg_0r);
  AND2 I1107 (rd_0r1[65:65], dt_0[65:65], rg_0r);
  AND2 I1108 (rd_0r1[66:66], dt_0[66:66], rg_0r);
  AND2 I1109 (rd_0r1[67:67], dt_0[67:67], rg_0r);
  AND2 I1110 (rd_0r1[68:68], dt_0[68:68], rg_0r);
  AND2 I1111 (rd_0r1[69:69], dt_0[69:69], rg_0r);
  AND2 I1112 (rd_0r1[70:70], dt_0[70:70], rg_0r);
  AND2 I1113 (rd_0r1[71:71], dt_0[71:71], rg_0r);
  AND2 I1114 (rd_0r1[72:72], dt_0[72:72], rg_0r);
  AND2 I1115 (rd_0r1[73:73], dt_0[73:73], rg_0r);
  OR2 I1116 (anyread_0, rg_0r, rg_0a);
  BUFF I1117 (wg_0a, wd_0a);
  BUFF I1118 (rg_0a, rd_0a);
endmodule

// tkvv33_wo0w33_ro0w33 TeakV "v" 33 [] [0] [0] [Many [33],Many [0],Many [0],Many [33]]
module tkvv33_wo0w33_ro0w33 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input [32:0] wg_0r0;
  input [32:0] wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output [32:0] rd_0r0;
  output [32:0] rd_0r1;
  input rd_0a;
  input reset;
  wire [32:0] wf_0;
  wire [32:0] wt_0;
  wire [32:0] df_0;
  wire [32:0] dt_0;
  wire wc_0;
  wire [32:0] wacks_0;
  wire [32:0] wenr_0;
  wire [32:0] wen_0;
  wire anyread_0;
  wire nreset_0;
  wire [32:0] drlgf_0;
  wire [32:0] drlgt_0;
  wire [32:0] comp0_0;
  wire [10:0] simp2451_0;
  wire [3:0] simp2452_0;
  wire [1:0] simp2453_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire [32:0] conwgit_0;
  wire [32:0] conwgif_0;
  wire conwig_0;
  wire [11:0] simp4191_0;
  wire [3:0] simp4192_0;
  wire [1:0] simp4193_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0[0:0], wenr_0[0:0], nreset_0);
  AND2 I2 (wen_0[1:1], wenr_0[1:1], nreset_0);
  AND2 I3 (wen_0[2:2], wenr_0[2:2], nreset_0);
  AND2 I4 (wen_0[3:3], wenr_0[3:3], nreset_0);
  AND2 I5 (wen_0[4:4], wenr_0[4:4], nreset_0);
  AND2 I6 (wen_0[5:5], wenr_0[5:5], nreset_0);
  AND2 I7 (wen_0[6:6], wenr_0[6:6], nreset_0);
  AND2 I8 (wen_0[7:7], wenr_0[7:7], nreset_0);
  AND2 I9 (wen_0[8:8], wenr_0[8:8], nreset_0);
  AND2 I10 (wen_0[9:9], wenr_0[9:9], nreset_0);
  AND2 I11 (wen_0[10:10], wenr_0[10:10], nreset_0);
  AND2 I12 (wen_0[11:11], wenr_0[11:11], nreset_0);
  AND2 I13 (wen_0[12:12], wenr_0[12:12], nreset_0);
  AND2 I14 (wen_0[13:13], wenr_0[13:13], nreset_0);
  AND2 I15 (wen_0[14:14], wenr_0[14:14], nreset_0);
  AND2 I16 (wen_0[15:15], wenr_0[15:15], nreset_0);
  AND2 I17 (wen_0[16:16], wenr_0[16:16], nreset_0);
  AND2 I18 (wen_0[17:17], wenr_0[17:17], nreset_0);
  AND2 I19 (wen_0[18:18], wenr_0[18:18], nreset_0);
  AND2 I20 (wen_0[19:19], wenr_0[19:19], nreset_0);
  AND2 I21 (wen_0[20:20], wenr_0[20:20], nreset_0);
  AND2 I22 (wen_0[21:21], wenr_0[21:21], nreset_0);
  AND2 I23 (wen_0[22:22], wenr_0[22:22], nreset_0);
  AND2 I24 (wen_0[23:23], wenr_0[23:23], nreset_0);
  AND2 I25 (wen_0[24:24], wenr_0[24:24], nreset_0);
  AND2 I26 (wen_0[25:25], wenr_0[25:25], nreset_0);
  AND2 I27 (wen_0[26:26], wenr_0[26:26], nreset_0);
  AND2 I28 (wen_0[27:27], wenr_0[27:27], nreset_0);
  AND2 I29 (wen_0[28:28], wenr_0[28:28], nreset_0);
  AND2 I30 (wen_0[29:29], wenr_0[29:29], nreset_0);
  AND2 I31 (wen_0[30:30], wenr_0[30:30], nreset_0);
  AND2 I32 (wen_0[31:31], wenr_0[31:31], nreset_0);
  AND2 I33 (wen_0[32:32], wenr_0[32:32], nreset_0);
  AND2 I34 (drlgf_0[0:0], wf_0[0:0], wen_0[0:0]);
  AND2 I35 (drlgf_0[1:1], wf_0[1:1], wen_0[1:1]);
  AND2 I36 (drlgf_0[2:2], wf_0[2:2], wen_0[2:2]);
  AND2 I37 (drlgf_0[3:3], wf_0[3:3], wen_0[3:3]);
  AND2 I38 (drlgf_0[4:4], wf_0[4:4], wen_0[4:4]);
  AND2 I39 (drlgf_0[5:5], wf_0[5:5], wen_0[5:5]);
  AND2 I40 (drlgf_0[6:6], wf_0[6:6], wen_0[6:6]);
  AND2 I41 (drlgf_0[7:7], wf_0[7:7], wen_0[7:7]);
  AND2 I42 (drlgf_0[8:8], wf_0[8:8], wen_0[8:8]);
  AND2 I43 (drlgf_0[9:9], wf_0[9:9], wen_0[9:9]);
  AND2 I44 (drlgf_0[10:10], wf_0[10:10], wen_0[10:10]);
  AND2 I45 (drlgf_0[11:11], wf_0[11:11], wen_0[11:11]);
  AND2 I46 (drlgf_0[12:12], wf_0[12:12], wen_0[12:12]);
  AND2 I47 (drlgf_0[13:13], wf_0[13:13], wen_0[13:13]);
  AND2 I48 (drlgf_0[14:14], wf_0[14:14], wen_0[14:14]);
  AND2 I49 (drlgf_0[15:15], wf_0[15:15], wen_0[15:15]);
  AND2 I50 (drlgf_0[16:16], wf_0[16:16], wen_0[16:16]);
  AND2 I51 (drlgf_0[17:17], wf_0[17:17], wen_0[17:17]);
  AND2 I52 (drlgf_0[18:18], wf_0[18:18], wen_0[18:18]);
  AND2 I53 (drlgf_0[19:19], wf_0[19:19], wen_0[19:19]);
  AND2 I54 (drlgf_0[20:20], wf_0[20:20], wen_0[20:20]);
  AND2 I55 (drlgf_0[21:21], wf_0[21:21], wen_0[21:21]);
  AND2 I56 (drlgf_0[22:22], wf_0[22:22], wen_0[22:22]);
  AND2 I57 (drlgf_0[23:23], wf_0[23:23], wen_0[23:23]);
  AND2 I58 (drlgf_0[24:24], wf_0[24:24], wen_0[24:24]);
  AND2 I59 (drlgf_0[25:25], wf_0[25:25], wen_0[25:25]);
  AND2 I60 (drlgf_0[26:26], wf_0[26:26], wen_0[26:26]);
  AND2 I61 (drlgf_0[27:27], wf_0[27:27], wen_0[27:27]);
  AND2 I62 (drlgf_0[28:28], wf_0[28:28], wen_0[28:28]);
  AND2 I63 (drlgf_0[29:29], wf_0[29:29], wen_0[29:29]);
  AND2 I64 (drlgf_0[30:30], wf_0[30:30], wen_0[30:30]);
  AND2 I65 (drlgf_0[31:31], wf_0[31:31], wen_0[31:31]);
  AND2 I66 (drlgf_0[32:32], wf_0[32:32], wen_0[32:32]);
  AND2 I67 (drlgt_0[0:0], wt_0[0:0], wen_0[0:0]);
  AND2 I68 (drlgt_0[1:1], wt_0[1:1], wen_0[1:1]);
  AND2 I69 (drlgt_0[2:2], wt_0[2:2], wen_0[2:2]);
  AND2 I70 (drlgt_0[3:3], wt_0[3:3], wen_0[3:3]);
  AND2 I71 (drlgt_0[4:4], wt_0[4:4], wen_0[4:4]);
  AND2 I72 (drlgt_0[5:5], wt_0[5:5], wen_0[5:5]);
  AND2 I73 (drlgt_0[6:6], wt_0[6:6], wen_0[6:6]);
  AND2 I74 (drlgt_0[7:7], wt_0[7:7], wen_0[7:7]);
  AND2 I75 (drlgt_0[8:8], wt_0[8:8], wen_0[8:8]);
  AND2 I76 (drlgt_0[9:9], wt_0[9:9], wen_0[9:9]);
  AND2 I77 (drlgt_0[10:10], wt_0[10:10], wen_0[10:10]);
  AND2 I78 (drlgt_0[11:11], wt_0[11:11], wen_0[11:11]);
  AND2 I79 (drlgt_0[12:12], wt_0[12:12], wen_0[12:12]);
  AND2 I80 (drlgt_0[13:13], wt_0[13:13], wen_0[13:13]);
  AND2 I81 (drlgt_0[14:14], wt_0[14:14], wen_0[14:14]);
  AND2 I82 (drlgt_0[15:15], wt_0[15:15], wen_0[15:15]);
  AND2 I83 (drlgt_0[16:16], wt_0[16:16], wen_0[16:16]);
  AND2 I84 (drlgt_0[17:17], wt_0[17:17], wen_0[17:17]);
  AND2 I85 (drlgt_0[18:18], wt_0[18:18], wen_0[18:18]);
  AND2 I86 (drlgt_0[19:19], wt_0[19:19], wen_0[19:19]);
  AND2 I87 (drlgt_0[20:20], wt_0[20:20], wen_0[20:20]);
  AND2 I88 (drlgt_0[21:21], wt_0[21:21], wen_0[21:21]);
  AND2 I89 (drlgt_0[22:22], wt_0[22:22], wen_0[22:22]);
  AND2 I90 (drlgt_0[23:23], wt_0[23:23], wen_0[23:23]);
  AND2 I91 (drlgt_0[24:24], wt_0[24:24], wen_0[24:24]);
  AND2 I92 (drlgt_0[25:25], wt_0[25:25], wen_0[25:25]);
  AND2 I93 (drlgt_0[26:26], wt_0[26:26], wen_0[26:26]);
  AND2 I94 (drlgt_0[27:27], wt_0[27:27], wen_0[27:27]);
  AND2 I95 (drlgt_0[28:28], wt_0[28:28], wen_0[28:28]);
  AND2 I96 (drlgt_0[29:29], wt_0[29:29], wen_0[29:29]);
  AND2 I97 (drlgt_0[30:30], wt_0[30:30], wen_0[30:30]);
  AND2 I98 (drlgt_0[31:31], wt_0[31:31], wen_0[31:31]);
  AND2 I99 (drlgt_0[32:32], wt_0[32:32], wen_0[32:32]);
  NOR2 I100 (df_0[0:0], dt_0[0:0], drlgt_0[0:0]);
  NOR2 I101 (df_0[1:1], dt_0[1:1], drlgt_0[1:1]);
  NOR2 I102 (df_0[2:2], dt_0[2:2], drlgt_0[2:2]);
  NOR2 I103 (df_0[3:3], dt_0[3:3], drlgt_0[3:3]);
  NOR2 I104 (df_0[4:4], dt_0[4:4], drlgt_0[4:4]);
  NOR2 I105 (df_0[5:5], dt_0[5:5], drlgt_0[5:5]);
  NOR2 I106 (df_0[6:6], dt_0[6:6], drlgt_0[6:6]);
  NOR2 I107 (df_0[7:7], dt_0[7:7], drlgt_0[7:7]);
  NOR2 I108 (df_0[8:8], dt_0[8:8], drlgt_0[8:8]);
  NOR2 I109 (df_0[9:9], dt_0[9:9], drlgt_0[9:9]);
  NOR2 I110 (df_0[10:10], dt_0[10:10], drlgt_0[10:10]);
  NOR2 I111 (df_0[11:11], dt_0[11:11], drlgt_0[11:11]);
  NOR2 I112 (df_0[12:12], dt_0[12:12], drlgt_0[12:12]);
  NOR2 I113 (df_0[13:13], dt_0[13:13], drlgt_0[13:13]);
  NOR2 I114 (df_0[14:14], dt_0[14:14], drlgt_0[14:14]);
  NOR2 I115 (df_0[15:15], dt_0[15:15], drlgt_0[15:15]);
  NOR2 I116 (df_0[16:16], dt_0[16:16], drlgt_0[16:16]);
  NOR2 I117 (df_0[17:17], dt_0[17:17], drlgt_0[17:17]);
  NOR2 I118 (df_0[18:18], dt_0[18:18], drlgt_0[18:18]);
  NOR2 I119 (df_0[19:19], dt_0[19:19], drlgt_0[19:19]);
  NOR2 I120 (df_0[20:20], dt_0[20:20], drlgt_0[20:20]);
  NOR2 I121 (df_0[21:21], dt_0[21:21], drlgt_0[21:21]);
  NOR2 I122 (df_0[22:22], dt_0[22:22], drlgt_0[22:22]);
  NOR2 I123 (df_0[23:23], dt_0[23:23], drlgt_0[23:23]);
  NOR2 I124 (df_0[24:24], dt_0[24:24], drlgt_0[24:24]);
  NOR2 I125 (df_0[25:25], dt_0[25:25], drlgt_0[25:25]);
  NOR2 I126 (df_0[26:26], dt_0[26:26], drlgt_0[26:26]);
  NOR2 I127 (df_0[27:27], dt_0[27:27], drlgt_0[27:27]);
  NOR2 I128 (df_0[28:28], dt_0[28:28], drlgt_0[28:28]);
  NOR2 I129 (df_0[29:29], dt_0[29:29], drlgt_0[29:29]);
  NOR2 I130 (df_0[30:30], dt_0[30:30], drlgt_0[30:30]);
  NOR2 I131 (df_0[31:31], dt_0[31:31], drlgt_0[31:31]);
  NOR2 I132 (df_0[32:32], dt_0[32:32], drlgt_0[32:32]);
  NOR3 I133 (dt_0[0:0], df_0[0:0], drlgf_0[0:0], reset);
  NOR3 I134 (dt_0[1:1], df_0[1:1], drlgf_0[1:1], reset);
  NOR3 I135 (dt_0[2:2], df_0[2:2], drlgf_0[2:2], reset);
  NOR3 I136 (dt_0[3:3], df_0[3:3], drlgf_0[3:3], reset);
  NOR3 I137 (dt_0[4:4], df_0[4:4], drlgf_0[4:4], reset);
  NOR3 I138 (dt_0[5:5], df_0[5:5], drlgf_0[5:5], reset);
  NOR3 I139 (dt_0[6:6], df_0[6:6], drlgf_0[6:6], reset);
  NOR3 I140 (dt_0[7:7], df_0[7:7], drlgf_0[7:7], reset);
  NOR3 I141 (dt_0[8:8], df_0[8:8], drlgf_0[8:8], reset);
  NOR3 I142 (dt_0[9:9], df_0[9:9], drlgf_0[9:9], reset);
  NOR3 I143 (dt_0[10:10], df_0[10:10], drlgf_0[10:10], reset);
  NOR3 I144 (dt_0[11:11], df_0[11:11], drlgf_0[11:11], reset);
  NOR3 I145 (dt_0[12:12], df_0[12:12], drlgf_0[12:12], reset);
  NOR3 I146 (dt_0[13:13], df_0[13:13], drlgf_0[13:13], reset);
  NOR3 I147 (dt_0[14:14], df_0[14:14], drlgf_0[14:14], reset);
  NOR3 I148 (dt_0[15:15], df_0[15:15], drlgf_0[15:15], reset);
  NOR3 I149 (dt_0[16:16], df_0[16:16], drlgf_0[16:16], reset);
  NOR3 I150 (dt_0[17:17], df_0[17:17], drlgf_0[17:17], reset);
  NOR3 I151 (dt_0[18:18], df_0[18:18], drlgf_0[18:18], reset);
  NOR3 I152 (dt_0[19:19], df_0[19:19], drlgf_0[19:19], reset);
  NOR3 I153 (dt_0[20:20], df_0[20:20], drlgf_0[20:20], reset);
  NOR3 I154 (dt_0[21:21], df_0[21:21], drlgf_0[21:21], reset);
  NOR3 I155 (dt_0[22:22], df_0[22:22], drlgf_0[22:22], reset);
  NOR3 I156 (dt_0[23:23], df_0[23:23], drlgf_0[23:23], reset);
  NOR3 I157 (dt_0[24:24], df_0[24:24], drlgf_0[24:24], reset);
  NOR3 I158 (dt_0[25:25], df_0[25:25], drlgf_0[25:25], reset);
  NOR3 I159 (dt_0[26:26], df_0[26:26], drlgf_0[26:26], reset);
  NOR3 I160 (dt_0[27:27], df_0[27:27], drlgf_0[27:27], reset);
  NOR3 I161 (dt_0[28:28], df_0[28:28], drlgf_0[28:28], reset);
  NOR3 I162 (dt_0[29:29], df_0[29:29], drlgf_0[29:29], reset);
  NOR3 I163 (dt_0[30:30], df_0[30:30], drlgf_0[30:30], reset);
  NOR3 I164 (dt_0[31:31], df_0[31:31], drlgf_0[31:31], reset);
  NOR3 I165 (dt_0[32:32], df_0[32:32], drlgf_0[32:32], reset);
  AO22 I166 (wacks_0[0:0], drlgf_0[0:0], df_0[0:0], drlgt_0[0:0], dt_0[0:0]);
  AO22 I167 (wacks_0[1:1], drlgf_0[1:1], df_0[1:1], drlgt_0[1:1], dt_0[1:1]);
  AO22 I168 (wacks_0[2:2], drlgf_0[2:2], df_0[2:2], drlgt_0[2:2], dt_0[2:2]);
  AO22 I169 (wacks_0[3:3], drlgf_0[3:3], df_0[3:3], drlgt_0[3:3], dt_0[3:3]);
  AO22 I170 (wacks_0[4:4], drlgf_0[4:4], df_0[4:4], drlgt_0[4:4], dt_0[4:4]);
  AO22 I171 (wacks_0[5:5], drlgf_0[5:5], df_0[5:5], drlgt_0[5:5], dt_0[5:5]);
  AO22 I172 (wacks_0[6:6], drlgf_0[6:6], df_0[6:6], drlgt_0[6:6], dt_0[6:6]);
  AO22 I173 (wacks_0[7:7], drlgf_0[7:7], df_0[7:7], drlgt_0[7:7], dt_0[7:7]);
  AO22 I174 (wacks_0[8:8], drlgf_0[8:8], df_0[8:8], drlgt_0[8:8], dt_0[8:8]);
  AO22 I175 (wacks_0[9:9], drlgf_0[9:9], df_0[9:9], drlgt_0[9:9], dt_0[9:9]);
  AO22 I176 (wacks_0[10:10], drlgf_0[10:10], df_0[10:10], drlgt_0[10:10], dt_0[10:10]);
  AO22 I177 (wacks_0[11:11], drlgf_0[11:11], df_0[11:11], drlgt_0[11:11], dt_0[11:11]);
  AO22 I178 (wacks_0[12:12], drlgf_0[12:12], df_0[12:12], drlgt_0[12:12], dt_0[12:12]);
  AO22 I179 (wacks_0[13:13], drlgf_0[13:13], df_0[13:13], drlgt_0[13:13], dt_0[13:13]);
  AO22 I180 (wacks_0[14:14], drlgf_0[14:14], df_0[14:14], drlgt_0[14:14], dt_0[14:14]);
  AO22 I181 (wacks_0[15:15], drlgf_0[15:15], df_0[15:15], drlgt_0[15:15], dt_0[15:15]);
  AO22 I182 (wacks_0[16:16], drlgf_0[16:16], df_0[16:16], drlgt_0[16:16], dt_0[16:16]);
  AO22 I183 (wacks_0[17:17], drlgf_0[17:17], df_0[17:17], drlgt_0[17:17], dt_0[17:17]);
  AO22 I184 (wacks_0[18:18], drlgf_0[18:18], df_0[18:18], drlgt_0[18:18], dt_0[18:18]);
  AO22 I185 (wacks_0[19:19], drlgf_0[19:19], df_0[19:19], drlgt_0[19:19], dt_0[19:19]);
  AO22 I186 (wacks_0[20:20], drlgf_0[20:20], df_0[20:20], drlgt_0[20:20], dt_0[20:20]);
  AO22 I187 (wacks_0[21:21], drlgf_0[21:21], df_0[21:21], drlgt_0[21:21], dt_0[21:21]);
  AO22 I188 (wacks_0[22:22], drlgf_0[22:22], df_0[22:22], drlgt_0[22:22], dt_0[22:22]);
  AO22 I189 (wacks_0[23:23], drlgf_0[23:23], df_0[23:23], drlgt_0[23:23], dt_0[23:23]);
  AO22 I190 (wacks_0[24:24], drlgf_0[24:24], df_0[24:24], drlgt_0[24:24], dt_0[24:24]);
  AO22 I191 (wacks_0[25:25], drlgf_0[25:25], df_0[25:25], drlgt_0[25:25], dt_0[25:25]);
  AO22 I192 (wacks_0[26:26], drlgf_0[26:26], df_0[26:26], drlgt_0[26:26], dt_0[26:26]);
  AO22 I193 (wacks_0[27:27], drlgf_0[27:27], df_0[27:27], drlgt_0[27:27], dt_0[27:27]);
  AO22 I194 (wacks_0[28:28], drlgf_0[28:28], df_0[28:28], drlgt_0[28:28], dt_0[28:28]);
  AO22 I195 (wacks_0[29:29], drlgf_0[29:29], df_0[29:29], drlgt_0[29:29], dt_0[29:29]);
  AO22 I196 (wacks_0[30:30], drlgf_0[30:30], df_0[30:30], drlgt_0[30:30], dt_0[30:30]);
  AO22 I197 (wacks_0[31:31], drlgf_0[31:31], df_0[31:31], drlgt_0[31:31], dt_0[31:31]);
  AO22 I198 (wacks_0[32:32], drlgf_0[32:32], df_0[32:32], drlgt_0[32:32], dt_0[32:32]);
  OR2 I199 (comp0_0[0:0], wg_0r0[0:0], wg_0r1[0:0]);
  OR2 I200 (comp0_0[1:1], wg_0r0[1:1], wg_0r1[1:1]);
  OR2 I201 (comp0_0[2:2], wg_0r0[2:2], wg_0r1[2:2]);
  OR2 I202 (comp0_0[3:3], wg_0r0[3:3], wg_0r1[3:3]);
  OR2 I203 (comp0_0[4:4], wg_0r0[4:4], wg_0r1[4:4]);
  OR2 I204 (comp0_0[5:5], wg_0r0[5:5], wg_0r1[5:5]);
  OR2 I205 (comp0_0[6:6], wg_0r0[6:6], wg_0r1[6:6]);
  OR2 I206 (comp0_0[7:7], wg_0r0[7:7], wg_0r1[7:7]);
  OR2 I207 (comp0_0[8:8], wg_0r0[8:8], wg_0r1[8:8]);
  OR2 I208 (comp0_0[9:9], wg_0r0[9:9], wg_0r1[9:9]);
  OR2 I209 (comp0_0[10:10], wg_0r0[10:10], wg_0r1[10:10]);
  OR2 I210 (comp0_0[11:11], wg_0r0[11:11], wg_0r1[11:11]);
  OR2 I211 (comp0_0[12:12], wg_0r0[12:12], wg_0r1[12:12]);
  OR2 I212 (comp0_0[13:13], wg_0r0[13:13], wg_0r1[13:13]);
  OR2 I213 (comp0_0[14:14], wg_0r0[14:14], wg_0r1[14:14]);
  OR2 I214 (comp0_0[15:15], wg_0r0[15:15], wg_0r1[15:15]);
  OR2 I215 (comp0_0[16:16], wg_0r0[16:16], wg_0r1[16:16]);
  OR2 I216 (comp0_0[17:17], wg_0r0[17:17], wg_0r1[17:17]);
  OR2 I217 (comp0_0[18:18], wg_0r0[18:18], wg_0r1[18:18]);
  OR2 I218 (comp0_0[19:19], wg_0r0[19:19], wg_0r1[19:19]);
  OR2 I219 (comp0_0[20:20], wg_0r0[20:20], wg_0r1[20:20]);
  OR2 I220 (comp0_0[21:21], wg_0r0[21:21], wg_0r1[21:21]);
  OR2 I221 (comp0_0[22:22], wg_0r0[22:22], wg_0r1[22:22]);
  OR2 I222 (comp0_0[23:23], wg_0r0[23:23], wg_0r1[23:23]);
  OR2 I223 (comp0_0[24:24], wg_0r0[24:24], wg_0r1[24:24]);
  OR2 I224 (comp0_0[25:25], wg_0r0[25:25], wg_0r1[25:25]);
  OR2 I225 (comp0_0[26:26], wg_0r0[26:26], wg_0r1[26:26]);
  OR2 I226 (comp0_0[27:27], wg_0r0[27:27], wg_0r1[27:27]);
  OR2 I227 (comp0_0[28:28], wg_0r0[28:28], wg_0r1[28:28]);
  OR2 I228 (comp0_0[29:29], wg_0r0[29:29], wg_0r1[29:29]);
  OR2 I229 (comp0_0[30:30], wg_0r0[30:30], wg_0r1[30:30]);
  OR2 I230 (comp0_0[31:31], wg_0r0[31:31], wg_0r1[31:31]);
  OR2 I231 (comp0_0[32:32], wg_0r0[32:32], wg_0r1[32:32]);
  C3 I232 (simp2451_0[0:0], comp0_0[0:0], comp0_0[1:1], comp0_0[2:2]);
  C3 I233 (simp2451_0[1:1], comp0_0[3:3], comp0_0[4:4], comp0_0[5:5]);
  C3 I234 (simp2451_0[2:2], comp0_0[6:6], comp0_0[7:7], comp0_0[8:8]);
  C3 I235 (simp2451_0[3:3], comp0_0[9:9], comp0_0[10:10], comp0_0[11:11]);
  C3 I236 (simp2451_0[4:4], comp0_0[12:12], comp0_0[13:13], comp0_0[14:14]);
  C3 I237 (simp2451_0[5:5], comp0_0[15:15], comp0_0[16:16], comp0_0[17:17]);
  C3 I238 (simp2451_0[6:6], comp0_0[18:18], comp0_0[19:19], comp0_0[20:20]);
  C3 I239 (simp2451_0[7:7], comp0_0[21:21], comp0_0[22:22], comp0_0[23:23]);
  C3 I240 (simp2451_0[8:8], comp0_0[24:24], comp0_0[25:25], comp0_0[26:26]);
  C3 I241 (simp2451_0[9:9], comp0_0[27:27], comp0_0[28:28], comp0_0[29:29]);
  C3 I242 (simp2451_0[10:10], comp0_0[30:30], comp0_0[31:31], comp0_0[32:32]);
  C3 I243 (simp2452_0[0:0], simp2451_0[0:0], simp2451_0[1:1], simp2451_0[2:2]);
  C3 I244 (simp2452_0[1:1], simp2451_0[3:3], simp2451_0[4:4], simp2451_0[5:5]);
  C3 I245 (simp2452_0[2:2], simp2451_0[6:6], simp2451_0[7:7], simp2451_0[8:8]);
  C2 I246 (simp2452_0[3:3], simp2451_0[9:9], simp2451_0[10:10]);
  C3 I247 (simp2453_0[0:0], simp2452_0[0:0], simp2452_0[1:1], simp2452_0[2:2]);
  BUFF I248 (simp2453_0[1:1], simp2452_0[3:3]);
  C2 I249 (wc_0, simp2453_0[0:0], simp2453_0[1:1]);
  AND2 I250 (conwgif_0[0:0], wg_0r0[0:0], conwig_0);
  AND2 I251 (conwgif_0[1:1], wg_0r0[1:1], conwig_0);
  AND2 I252 (conwgif_0[2:2], wg_0r0[2:2], conwig_0);
  AND2 I253 (conwgif_0[3:3], wg_0r0[3:3], conwig_0);
  AND2 I254 (conwgif_0[4:4], wg_0r0[4:4], conwig_0);
  AND2 I255 (conwgif_0[5:5], wg_0r0[5:5], conwig_0);
  AND2 I256 (conwgif_0[6:6], wg_0r0[6:6], conwig_0);
  AND2 I257 (conwgif_0[7:7], wg_0r0[7:7], conwig_0);
  AND2 I258 (conwgif_0[8:8], wg_0r0[8:8], conwig_0);
  AND2 I259 (conwgif_0[9:9], wg_0r0[9:9], conwig_0);
  AND2 I260 (conwgif_0[10:10], wg_0r0[10:10], conwig_0);
  AND2 I261 (conwgif_0[11:11], wg_0r0[11:11], conwig_0);
  AND2 I262 (conwgif_0[12:12], wg_0r0[12:12], conwig_0);
  AND2 I263 (conwgif_0[13:13], wg_0r0[13:13], conwig_0);
  AND2 I264 (conwgif_0[14:14], wg_0r0[14:14], conwig_0);
  AND2 I265 (conwgif_0[15:15], wg_0r0[15:15], conwig_0);
  AND2 I266 (conwgif_0[16:16], wg_0r0[16:16], conwig_0);
  AND2 I267 (conwgif_0[17:17], wg_0r0[17:17], conwig_0);
  AND2 I268 (conwgif_0[18:18], wg_0r0[18:18], conwig_0);
  AND2 I269 (conwgif_0[19:19], wg_0r0[19:19], conwig_0);
  AND2 I270 (conwgif_0[20:20], wg_0r0[20:20], conwig_0);
  AND2 I271 (conwgif_0[21:21], wg_0r0[21:21], conwig_0);
  AND2 I272 (conwgif_0[22:22], wg_0r0[22:22], conwig_0);
  AND2 I273 (conwgif_0[23:23], wg_0r0[23:23], conwig_0);
  AND2 I274 (conwgif_0[24:24], wg_0r0[24:24], conwig_0);
  AND2 I275 (conwgif_0[25:25], wg_0r0[25:25], conwig_0);
  AND2 I276 (conwgif_0[26:26], wg_0r0[26:26], conwig_0);
  AND2 I277 (conwgif_0[27:27], wg_0r0[27:27], conwig_0);
  AND2 I278 (conwgif_0[28:28], wg_0r0[28:28], conwig_0);
  AND2 I279 (conwgif_0[29:29], wg_0r0[29:29], conwig_0);
  AND2 I280 (conwgif_0[30:30], wg_0r0[30:30], conwig_0);
  AND2 I281 (conwgif_0[31:31], wg_0r0[31:31], conwig_0);
  AND2 I282 (conwgif_0[32:32], wg_0r0[32:32], conwig_0);
  AND2 I283 (conwgit_0[0:0], wg_0r1[0:0], conwig_0);
  AND2 I284 (conwgit_0[1:1], wg_0r1[1:1], conwig_0);
  AND2 I285 (conwgit_0[2:2], wg_0r1[2:2], conwig_0);
  AND2 I286 (conwgit_0[3:3], wg_0r1[3:3], conwig_0);
  AND2 I287 (conwgit_0[4:4], wg_0r1[4:4], conwig_0);
  AND2 I288 (conwgit_0[5:5], wg_0r1[5:5], conwig_0);
  AND2 I289 (conwgit_0[6:6], wg_0r1[6:6], conwig_0);
  AND2 I290 (conwgit_0[7:7], wg_0r1[7:7], conwig_0);
  AND2 I291 (conwgit_0[8:8], wg_0r1[8:8], conwig_0);
  AND2 I292 (conwgit_0[9:9], wg_0r1[9:9], conwig_0);
  AND2 I293 (conwgit_0[10:10], wg_0r1[10:10], conwig_0);
  AND2 I294 (conwgit_0[11:11], wg_0r1[11:11], conwig_0);
  AND2 I295 (conwgit_0[12:12], wg_0r1[12:12], conwig_0);
  AND2 I296 (conwgit_0[13:13], wg_0r1[13:13], conwig_0);
  AND2 I297 (conwgit_0[14:14], wg_0r1[14:14], conwig_0);
  AND2 I298 (conwgit_0[15:15], wg_0r1[15:15], conwig_0);
  AND2 I299 (conwgit_0[16:16], wg_0r1[16:16], conwig_0);
  AND2 I300 (conwgit_0[17:17], wg_0r1[17:17], conwig_0);
  AND2 I301 (conwgit_0[18:18], wg_0r1[18:18], conwig_0);
  AND2 I302 (conwgit_0[19:19], wg_0r1[19:19], conwig_0);
  AND2 I303 (conwgit_0[20:20], wg_0r1[20:20], conwig_0);
  AND2 I304 (conwgit_0[21:21], wg_0r1[21:21], conwig_0);
  AND2 I305 (conwgit_0[22:22], wg_0r1[22:22], conwig_0);
  AND2 I306 (conwgit_0[23:23], wg_0r1[23:23], conwig_0);
  AND2 I307 (conwgit_0[24:24], wg_0r1[24:24], conwig_0);
  AND2 I308 (conwgit_0[25:25], wg_0r1[25:25], conwig_0);
  AND2 I309 (conwgit_0[26:26], wg_0r1[26:26], conwig_0);
  AND2 I310 (conwgit_0[27:27], wg_0r1[27:27], conwig_0);
  AND2 I311 (conwgit_0[28:28], wg_0r1[28:28], conwig_0);
  AND2 I312 (conwgit_0[29:29], wg_0r1[29:29], conwig_0);
  AND2 I313 (conwgit_0[30:30], wg_0r1[30:30], conwig_0);
  AND2 I314 (conwgit_0[31:31], wg_0r1[31:31], conwig_0);
  AND2 I315 (conwgit_0[32:32], wg_0r1[32:32], conwig_0);
  BUFF I316 (conwigc_0, wc_0);
  AO22 I317 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I318 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I319 (wf_0[0:0], conwgif_0[0:0]);
  BUFF I320 (wt_0[0:0], conwgit_0[0:0]);
  BUFF I321 (wenr_0[0:0], wc_0);
  BUFF I322 (wf_0[1:1], conwgif_0[1:1]);
  BUFF I323 (wt_0[1:1], conwgit_0[1:1]);
  BUFF I324 (wenr_0[1:1], wc_0);
  BUFF I325 (wf_0[2:2], conwgif_0[2:2]);
  BUFF I326 (wt_0[2:2], conwgit_0[2:2]);
  BUFF I327 (wenr_0[2:2], wc_0);
  BUFF I328 (wf_0[3:3], conwgif_0[3:3]);
  BUFF I329 (wt_0[3:3], conwgit_0[3:3]);
  BUFF I330 (wenr_0[3:3], wc_0);
  BUFF I331 (wf_0[4:4], conwgif_0[4:4]);
  BUFF I332 (wt_0[4:4], conwgit_0[4:4]);
  BUFF I333 (wenr_0[4:4], wc_0);
  BUFF I334 (wf_0[5:5], conwgif_0[5:5]);
  BUFF I335 (wt_0[5:5], conwgit_0[5:5]);
  BUFF I336 (wenr_0[5:5], wc_0);
  BUFF I337 (wf_0[6:6], conwgif_0[6:6]);
  BUFF I338 (wt_0[6:6], conwgit_0[6:6]);
  BUFF I339 (wenr_0[6:6], wc_0);
  BUFF I340 (wf_0[7:7], conwgif_0[7:7]);
  BUFF I341 (wt_0[7:7], conwgit_0[7:7]);
  BUFF I342 (wenr_0[7:7], wc_0);
  BUFF I343 (wf_0[8:8], conwgif_0[8:8]);
  BUFF I344 (wt_0[8:8], conwgit_0[8:8]);
  BUFF I345 (wenr_0[8:8], wc_0);
  BUFF I346 (wf_0[9:9], conwgif_0[9:9]);
  BUFF I347 (wt_0[9:9], conwgit_0[9:9]);
  BUFF I348 (wenr_0[9:9], wc_0);
  BUFF I349 (wf_0[10:10], conwgif_0[10:10]);
  BUFF I350 (wt_0[10:10], conwgit_0[10:10]);
  BUFF I351 (wenr_0[10:10], wc_0);
  BUFF I352 (wf_0[11:11], conwgif_0[11:11]);
  BUFF I353 (wt_0[11:11], conwgit_0[11:11]);
  BUFF I354 (wenr_0[11:11], wc_0);
  BUFF I355 (wf_0[12:12], conwgif_0[12:12]);
  BUFF I356 (wt_0[12:12], conwgit_0[12:12]);
  BUFF I357 (wenr_0[12:12], wc_0);
  BUFF I358 (wf_0[13:13], conwgif_0[13:13]);
  BUFF I359 (wt_0[13:13], conwgit_0[13:13]);
  BUFF I360 (wenr_0[13:13], wc_0);
  BUFF I361 (wf_0[14:14], conwgif_0[14:14]);
  BUFF I362 (wt_0[14:14], conwgit_0[14:14]);
  BUFF I363 (wenr_0[14:14], wc_0);
  BUFF I364 (wf_0[15:15], conwgif_0[15:15]);
  BUFF I365 (wt_0[15:15], conwgit_0[15:15]);
  BUFF I366 (wenr_0[15:15], wc_0);
  BUFF I367 (wf_0[16:16], conwgif_0[16:16]);
  BUFF I368 (wt_0[16:16], conwgit_0[16:16]);
  BUFF I369 (wenr_0[16:16], wc_0);
  BUFF I370 (wf_0[17:17], conwgif_0[17:17]);
  BUFF I371 (wt_0[17:17], conwgit_0[17:17]);
  BUFF I372 (wenr_0[17:17], wc_0);
  BUFF I373 (wf_0[18:18], conwgif_0[18:18]);
  BUFF I374 (wt_0[18:18], conwgit_0[18:18]);
  BUFF I375 (wenr_0[18:18], wc_0);
  BUFF I376 (wf_0[19:19], conwgif_0[19:19]);
  BUFF I377 (wt_0[19:19], conwgit_0[19:19]);
  BUFF I378 (wenr_0[19:19], wc_0);
  BUFF I379 (wf_0[20:20], conwgif_0[20:20]);
  BUFF I380 (wt_0[20:20], conwgit_0[20:20]);
  BUFF I381 (wenr_0[20:20], wc_0);
  BUFF I382 (wf_0[21:21], conwgif_0[21:21]);
  BUFF I383 (wt_0[21:21], conwgit_0[21:21]);
  BUFF I384 (wenr_0[21:21], wc_0);
  BUFF I385 (wf_0[22:22], conwgif_0[22:22]);
  BUFF I386 (wt_0[22:22], conwgit_0[22:22]);
  BUFF I387 (wenr_0[22:22], wc_0);
  BUFF I388 (wf_0[23:23], conwgif_0[23:23]);
  BUFF I389 (wt_0[23:23], conwgit_0[23:23]);
  BUFF I390 (wenr_0[23:23], wc_0);
  BUFF I391 (wf_0[24:24], conwgif_0[24:24]);
  BUFF I392 (wt_0[24:24], conwgit_0[24:24]);
  BUFF I393 (wenr_0[24:24], wc_0);
  BUFF I394 (wf_0[25:25], conwgif_0[25:25]);
  BUFF I395 (wt_0[25:25], conwgit_0[25:25]);
  BUFF I396 (wenr_0[25:25], wc_0);
  BUFF I397 (wf_0[26:26], conwgif_0[26:26]);
  BUFF I398 (wt_0[26:26], conwgit_0[26:26]);
  BUFF I399 (wenr_0[26:26], wc_0);
  BUFF I400 (wf_0[27:27], conwgif_0[27:27]);
  BUFF I401 (wt_0[27:27], conwgit_0[27:27]);
  BUFF I402 (wenr_0[27:27], wc_0);
  BUFF I403 (wf_0[28:28], conwgif_0[28:28]);
  BUFF I404 (wt_0[28:28], conwgit_0[28:28]);
  BUFF I405 (wenr_0[28:28], wc_0);
  BUFF I406 (wf_0[29:29], conwgif_0[29:29]);
  BUFF I407 (wt_0[29:29], conwgit_0[29:29]);
  BUFF I408 (wenr_0[29:29], wc_0);
  BUFF I409 (wf_0[30:30], conwgif_0[30:30]);
  BUFF I410 (wt_0[30:30], conwgit_0[30:30]);
  BUFF I411 (wenr_0[30:30], wc_0);
  BUFF I412 (wf_0[31:31], conwgif_0[31:31]);
  BUFF I413 (wt_0[31:31], conwgit_0[31:31]);
  BUFF I414 (wenr_0[31:31], wc_0);
  BUFF I415 (wf_0[32:32], conwgif_0[32:32]);
  BUFF I416 (wt_0[32:32], conwgit_0[32:32]);
  BUFF I417 (wenr_0[32:32], wc_0);
  C3 I418 (simp4191_0[0:0], conwig_0, wacks_0[0:0], wacks_0[1:1]);
  C3 I419 (simp4191_0[1:1], wacks_0[2:2], wacks_0[3:3], wacks_0[4:4]);
  C3 I420 (simp4191_0[2:2], wacks_0[5:5], wacks_0[6:6], wacks_0[7:7]);
  C3 I421 (simp4191_0[3:3], wacks_0[8:8], wacks_0[9:9], wacks_0[10:10]);
  C3 I422 (simp4191_0[4:4], wacks_0[11:11], wacks_0[12:12], wacks_0[13:13]);
  C3 I423 (simp4191_0[5:5], wacks_0[14:14], wacks_0[15:15], wacks_0[16:16]);
  C3 I424 (simp4191_0[6:6], wacks_0[17:17], wacks_0[18:18], wacks_0[19:19]);
  C3 I425 (simp4191_0[7:7], wacks_0[20:20], wacks_0[21:21], wacks_0[22:22]);
  C3 I426 (simp4191_0[8:8], wacks_0[23:23], wacks_0[24:24], wacks_0[25:25]);
  C3 I427 (simp4191_0[9:9], wacks_0[26:26], wacks_0[27:27], wacks_0[28:28]);
  C3 I428 (simp4191_0[10:10], wacks_0[29:29], wacks_0[30:30], wacks_0[31:31]);
  BUFF I429 (simp4191_0[11:11], wacks_0[32:32]);
  C3 I430 (simp4192_0[0:0], simp4191_0[0:0], simp4191_0[1:1], simp4191_0[2:2]);
  C3 I431 (simp4192_0[1:1], simp4191_0[3:3], simp4191_0[4:4], simp4191_0[5:5]);
  C3 I432 (simp4192_0[2:2], simp4191_0[6:6], simp4191_0[7:7], simp4191_0[8:8]);
  C3 I433 (simp4192_0[3:3], simp4191_0[9:9], simp4191_0[10:10], simp4191_0[11:11]);
  C3 I434 (simp4193_0[0:0], simp4192_0[0:0], simp4192_0[1:1], simp4192_0[2:2]);
  BUFF I435 (simp4193_0[1:1], simp4192_0[3:3]);
  C2 I436 (wd_0r, simp4193_0[0:0], simp4193_0[1:1]);
  AND2 I437 (rd_0r0[0:0], df_0[0:0], rg_0r);
  AND2 I438 (rd_0r0[1:1], df_0[1:1], rg_0r);
  AND2 I439 (rd_0r0[2:2], df_0[2:2], rg_0r);
  AND2 I440 (rd_0r0[3:3], df_0[3:3], rg_0r);
  AND2 I441 (rd_0r0[4:4], df_0[4:4], rg_0r);
  AND2 I442 (rd_0r0[5:5], df_0[5:5], rg_0r);
  AND2 I443 (rd_0r0[6:6], df_0[6:6], rg_0r);
  AND2 I444 (rd_0r0[7:7], df_0[7:7], rg_0r);
  AND2 I445 (rd_0r0[8:8], df_0[8:8], rg_0r);
  AND2 I446 (rd_0r0[9:9], df_0[9:9], rg_0r);
  AND2 I447 (rd_0r0[10:10], df_0[10:10], rg_0r);
  AND2 I448 (rd_0r0[11:11], df_0[11:11], rg_0r);
  AND2 I449 (rd_0r0[12:12], df_0[12:12], rg_0r);
  AND2 I450 (rd_0r0[13:13], df_0[13:13], rg_0r);
  AND2 I451 (rd_0r0[14:14], df_0[14:14], rg_0r);
  AND2 I452 (rd_0r0[15:15], df_0[15:15], rg_0r);
  AND2 I453 (rd_0r0[16:16], df_0[16:16], rg_0r);
  AND2 I454 (rd_0r0[17:17], df_0[17:17], rg_0r);
  AND2 I455 (rd_0r0[18:18], df_0[18:18], rg_0r);
  AND2 I456 (rd_0r0[19:19], df_0[19:19], rg_0r);
  AND2 I457 (rd_0r0[20:20], df_0[20:20], rg_0r);
  AND2 I458 (rd_0r0[21:21], df_0[21:21], rg_0r);
  AND2 I459 (rd_0r0[22:22], df_0[22:22], rg_0r);
  AND2 I460 (rd_0r0[23:23], df_0[23:23], rg_0r);
  AND2 I461 (rd_0r0[24:24], df_0[24:24], rg_0r);
  AND2 I462 (rd_0r0[25:25], df_0[25:25], rg_0r);
  AND2 I463 (rd_0r0[26:26], df_0[26:26], rg_0r);
  AND2 I464 (rd_0r0[27:27], df_0[27:27], rg_0r);
  AND2 I465 (rd_0r0[28:28], df_0[28:28], rg_0r);
  AND2 I466 (rd_0r0[29:29], df_0[29:29], rg_0r);
  AND2 I467 (rd_0r0[30:30], df_0[30:30], rg_0r);
  AND2 I468 (rd_0r0[31:31], df_0[31:31], rg_0r);
  AND2 I469 (rd_0r0[32:32], df_0[32:32], rg_0r);
  AND2 I470 (rd_0r1[0:0], dt_0[0:0], rg_0r);
  AND2 I471 (rd_0r1[1:1], dt_0[1:1], rg_0r);
  AND2 I472 (rd_0r1[2:2], dt_0[2:2], rg_0r);
  AND2 I473 (rd_0r1[3:3], dt_0[3:3], rg_0r);
  AND2 I474 (rd_0r1[4:4], dt_0[4:4], rg_0r);
  AND2 I475 (rd_0r1[5:5], dt_0[5:5], rg_0r);
  AND2 I476 (rd_0r1[6:6], dt_0[6:6], rg_0r);
  AND2 I477 (rd_0r1[7:7], dt_0[7:7], rg_0r);
  AND2 I478 (rd_0r1[8:8], dt_0[8:8], rg_0r);
  AND2 I479 (rd_0r1[9:9], dt_0[9:9], rg_0r);
  AND2 I480 (rd_0r1[10:10], dt_0[10:10], rg_0r);
  AND2 I481 (rd_0r1[11:11], dt_0[11:11], rg_0r);
  AND2 I482 (rd_0r1[12:12], dt_0[12:12], rg_0r);
  AND2 I483 (rd_0r1[13:13], dt_0[13:13], rg_0r);
  AND2 I484 (rd_0r1[14:14], dt_0[14:14], rg_0r);
  AND2 I485 (rd_0r1[15:15], dt_0[15:15], rg_0r);
  AND2 I486 (rd_0r1[16:16], dt_0[16:16], rg_0r);
  AND2 I487 (rd_0r1[17:17], dt_0[17:17], rg_0r);
  AND2 I488 (rd_0r1[18:18], dt_0[18:18], rg_0r);
  AND2 I489 (rd_0r1[19:19], dt_0[19:19], rg_0r);
  AND2 I490 (rd_0r1[20:20], dt_0[20:20], rg_0r);
  AND2 I491 (rd_0r1[21:21], dt_0[21:21], rg_0r);
  AND2 I492 (rd_0r1[22:22], dt_0[22:22], rg_0r);
  AND2 I493 (rd_0r1[23:23], dt_0[23:23], rg_0r);
  AND2 I494 (rd_0r1[24:24], dt_0[24:24], rg_0r);
  AND2 I495 (rd_0r1[25:25], dt_0[25:25], rg_0r);
  AND2 I496 (rd_0r1[26:26], dt_0[26:26], rg_0r);
  AND2 I497 (rd_0r1[27:27], dt_0[27:27], rg_0r);
  AND2 I498 (rd_0r1[28:28], dt_0[28:28], rg_0r);
  AND2 I499 (rd_0r1[29:29], dt_0[29:29], rg_0r);
  AND2 I500 (rd_0r1[30:30], dt_0[30:30], rg_0r);
  AND2 I501 (rd_0r1[31:31], dt_0[31:31], rg_0r);
  AND2 I502 (rd_0r1[32:32], dt_0[32:32], rg_0r);
  OR2 I503 (anyread_0, rg_0r, rg_0a);
  BUFF I504 (wg_0a, wd_0a);
  BUFF I505 (rg_0a, rd_0a);
endmodule

// tkvv1_wo0w1_ro0w1 TeakV "v" 1 [] [0] [0] [Many [1],Many [0],Many [0],Many [1]]
module tkvv1_wo0w1_ro0w1 (wg_0r0, wg_0r1, wg_0a, wd_0r, wd_0a, rg_0r, rg_0a, rd_0r0, rd_0r1, rd_0a, reset);
  input wg_0r0;
  input wg_0r1;
  output wg_0a;
  output wd_0r;
  input wd_0a;
  input rg_0r;
  output rg_0a;
  output rd_0r0;
  output rd_0r1;
  input rd_0a;
  input reset;
  wire wf_0;
  wire wt_0;
  wire df_0;
  wire dt_0;
  wire wc_0;
  wire wacks_0;
  wire wenr_0;
  wire wen_0;
  wire anyread_0;
  wire nreset_0;
  wire drlgf_0;
  wire drlgt_0;
  wire comp0_0;
  wire conwigc_0;
  wire conwigcanw_0;
  wire conwgit_0;
  wire conwgif_0;
  wire conwig_0;
  INV I0 (nreset_0, reset);
  AND2 I1 (wen_0, wenr_0, nreset_0);
  AND2 I2 (drlgf_0, wf_0, wen_0);
  AND2 I3 (drlgt_0, wt_0, wen_0);
  NOR2 I4 (df_0, dt_0, drlgt_0);
  NOR3 I5 (dt_0, df_0, drlgf_0, reset);
  AO22 I6 (wacks_0, drlgf_0, df_0, drlgt_0, dt_0);
  OR2 I7 (comp0_0, wg_0r0, wg_0r1);
  BUFF I8 (wc_0, comp0_0);
  AND2 I9 (conwgif_0, wg_0r0, conwig_0);
  AND2 I10 (conwgit_0, wg_0r1, conwig_0);
  BUFF I11 (conwigc_0, wc_0);
  AO22 I12 (conwig_0, conwigc_0, conwigcanw_0, conwigc_0, conwig_0);
  NOR2 I13 (conwigcanw_0, anyread_0, conwig_0);
  BUFF I14 (wf_0, conwgif_0);
  BUFF I15 (wt_0, conwgit_0);
  BUFF I16 (wenr_0, wc_0);
  C2 I17 (wd_0r, conwig_0, wacks_0);
  AND2 I18 (rd_0r0, df_0, rg_0r);
  AND2 I19 (rd_0r1, dt_0, rg_0r);
  OR2 I20 (anyread_0, rg_0r, rg_0a);
  BUFF I21 (wg_0a, wd_0a);
  BUFF I22 (rg_0a, rd_0a);
endmodule

module teak_FetchInitial (doFetchI_0r0, doFetchI_0r1, doFetchI_0a, doFetchO_0r0, doFetchO_0r1, doFetchO_0a, reset);
  input doFetchI_0r0;
  input doFetchI_0r1;
  output doFetchI_0a;
  output doFetchO_0r0;
  output doFetchO_0r1;
  input doFetchO_0a;
  input reset;
  wire L3_0r;
  wire L3_0a;
  wire L5_0r0;
  wire L5_0r1;
  wire L5_0a;
  wire L7_0r;
  wire L7_0a;
  wire L9_0r0;
  wire L9_0r1;
  wire L9_0a;
  wire L11_0r;
  wire L11_0a;
  wire L13_0r0;
  wire L13_0r1;
  wire L13_0a;
  wire L14_0r;
  wire L14_0a;
  wire L15_0r0;
  wire L15_0r1;
  wire L15_0a;
  wire L17_0r;
  wire L17_0a;
  wire L18_0r;
  wire L18_0a;
  wire L20_0r;
  wire L20_0a;
  wire L21_0r0;
  wire L21_0r1;
  wire L21_0a;
  wire L22_0r;
  wire L22_0a;
  wire L23_0r0;
  wire L23_0r1;
  wire L23_0a;
  wire L24_0r;
  wire L24_0a;
  wire L25_0r0;
  wire L25_0r1;
  wire L25_0a;
  wire L26_0r0;
  wire L26_0r1;
  wire L26_0a;
  wire L27_0r;
  wire L27_0a;
  wire [2:0] L29_0r0;
  wire [2:0] L29_0r1;
  wire L29_0a;
  wire [2:0] L30_0r0;
  wire [2:0] L30_0r1;
  wire L30_0a;
  wire [2:0] L31_0r0;
  wire [2:0] L31_0r1;
  wire L31_0a;
  wire [2:0] L32_0r0;
  wire [2:0] L32_0r1;
  wire L32_0a;
  wire [2:0] L33_0r0;
  wire [2:0] L33_0r1;
  wire L33_0a;
  tko0m1_1nm1b0 I0 (L3_0r, L3_0a, L5_0r0, L5_0r1, L5_0a, reset);
  tko0m1_1nm1b0 I1 (L7_0r, L7_0a, L9_0r0, L9_0r1, L9_0a, reset);
  tkvdoFetchI1_wo0w1_ro0w1 I2 (L15_0r0, L15_0r1, L15_0a, L11_0r, L11_0a, L11_0r, L11_0a, L13_0r0, L13_0r1, L13_0a, reset);
  tkm2x0b I3 (L18_0r, L18_0a, L14_0r, L14_0a, L17_0r, L17_0a, reset);
  tkj1m1_0 I4 (doFetchI_0r0, doFetchI_0r1, doFetchI_0a, L17_0r, L17_0a, L15_0r0, L15_0r1, L15_0a, reset);
  tkf1mo0w0_o0w1 I5 (L5_0r0, L5_0r1, L5_0a, L20_0r, L20_0a, L21_0r0, L21_0r1, L21_0a, reset);
  tkf1mo0w0_o0w1 I6 (L9_0r0, L9_0r1, L9_0a, L22_0r, L22_0a, L23_0r0, L23_0r1, L23_0a, reset);
  tkf1mo0w0_o0w1 I7 (L13_0r0, L13_0r1, L13_0a, L24_0r, L24_0a, L25_0r0, L25_0r1, L25_0a, reset);
  tkm3x1b I8 (L21_0r0, L21_0r1, L21_0a, L23_0r0, L23_0r1, L23_0a, L25_0r0, L25_0r1, L25_0a, L26_0r0, L26_0r1, L26_0a, reset);
  tkf1mo0w0_o0w1 I9 (L26_0r0, L26_0r1, L26_0a, L27_0r, L27_0a, doFetchO_0r0, doFetchO_0r1, doFetchO_0a, reset);
  tko0m3_1nm3b1 I10 (L20_0r, L20_0a, L29_0r0[2:0], L29_0r1[2:0], L29_0a, reset);
  tko0m3_1nm3b2 I11 (L22_0r, L22_0a, L30_0r0[2:0], L30_0r1[2:0], L30_0a, reset);
  tko0m3_1nm3b4 I12 (L24_0r, L24_0a, L31_0r0[2:0], L31_0r1[2:0], L31_0a, reset);
  tkm3x3b I13 (L29_0r0[2:0], L29_0r1[2:0], L29_0a, L30_0r0[2:0], L30_0r1[2:0], L30_0a, L31_0r0[2:0], L31_0r1[2:0], L31_0a, L32_0r0[2:0], L32_0r1[2:0], L32_0a, reset);
  tkj3m0_3 I14 (L27_0r, L27_0a, L32_0r0[2:0], L32_0r1[2:0], L32_0a, L33_0r0[2:0], L33_0r1[2:0], L33_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_4o0w0 I15 (L33_0r0[2:0], L33_0r1[2:0], L33_0a, L7_0r, L7_0a, L18_0r, L18_0a, L14_0r, L14_0a, reset);
  tkr I16 (L3_0r, L3_0a, reset);
endmodule

module teak_Fetch (doFetch_0r0, doFetch_0r1, doFetch_0a, newPc_0r0, newPc_0r1, newPc_0a, inst_0r0, inst_0r1, inst_0a, faddr_0r0, faddr_0r1, faddr_0a, finst_0r0, finst_0r1, finst_0a, reset);
  input doFetch_0r0;
  input doFetch_0r1;
  output doFetch_0a;
  input [31:0] newPc_0r0;
  input [31:0] newPc_0r1;
  output newPc_0a;
  output [64:0] inst_0r0;
  output [64:0] inst_0r1;
  input inst_0a;
  output [31:0] faddr_0r0;
  output [31:0] faddr_0r1;
  input faddr_0a;
  input [31:0] finst_0r0;
  input [31:0] finst_0r1;
  output finst_0a;
  input reset;
  wire L2_0r;
  wire L2_0a;
  wire [31:0] L4_0r0;
  wire [31:0] L4_0r1;
  wire L4_0a;
  wire L5_0r;
  wire L5_0a;
  wire L6_0r;
  wire L6_0a;
  wire L8_0r0;
  wire L8_0r1;
  wire L8_0a;
  wire L9_0r;
  wire L9_0a;
  wire L12_0r;
  wire L12_0a;
  wire L13_0r0;
  wire L13_0r1;
  wire L13_0a;
  wire L14_0r;
  wire L14_0a;
  wire L15_0r;
  wire L15_0a;
  wire L17_0r;
  wire L17_0a;
  wire [31:0] L19_0r0;
  wire [31:0] L19_0r1;
  wire L19_0a;
  wire L20_0r;
  wire L20_0a;
  wire L21_0r;
  wire L21_0a;
  wire L22_0r;
  wire L22_0a;
  wire L23_0r;
  wire L23_0a;
  wire [31:0] L24_0r0;
  wire [31:0] L24_0r1;
  wire L24_0a;
  wire L26_0r;
  wire L26_0a;
  wire L27_0r;
  wire L27_0a;
  wire L29_0r0;
  wire L29_0r1;
  wire L29_0a;
  wire L30_0r;
  wire L30_0a;
  wire L31_0r;
  wire L31_0a;
  wire L33_0r;
  wire L33_0a;
  wire L34_0r;
  wire L34_0a;
  wire L35_0r;
  wire L35_0a;
  wire L36_0r0;
  wire L36_0r1;
  wire L36_0a;
  wire L38_0r;
  wire L38_0a;
  wire L39_0r;
  wire L39_0a;
  wire L41_0r;
  wire L41_0a;
  wire [31:0] L43_0r0;
  wire [31:0] L43_0r1;
  wire L43_0a;
  wire L44_0r;
  wire L44_0a;
  wire L45_0r;
  wire L45_0a;
  wire [31:0] L46_0r0;
  wire [31:0] L46_0r1;
  wire L46_0a;
  wire L47_0r;
  wire L47_0a;
  wire [31:0] L48_0r0;
  wire [31:0] L48_0r1;
  wire L48_0a;
  wire L49_0r;
  wire L49_0a;
  wire L50_0r0;
  wire L50_0r1;
  wire L50_0a;
  wire [32:0] L51_0r0;
  wire [32:0] L51_0r1;
  wire L51_0a;
  wire L53_0r;
  wire L53_0a;
  wire [64:0] L54_0r0;
  wire [64:0] L54_0r1;
  wire L54_0a;
  wire L55_0r;
  wire L55_0a;
  wire L56_0r;
  wire L56_0a;
  wire L57_0r;
  wire L57_0a;
  wire L58_0r;
  wire L58_0a;
  wire [31:0] L59_0r0;
  wire [31:0] L59_0r1;
  wire L59_0a;
  wire L61_0r;
  wire L61_0a;
  wire L63_0r;
  wire L63_0a;
  wire [31:0] L64_0r0;
  wire [31:0] L64_0r1;
  wire L64_0a;
  wire L65_0r;
  wire L65_0a;
  wire [2:0] L66_0r0;
  wire [2:0] L66_0r1;
  wire L66_0a;
  wire [34:0] L67_0r0;
  wire [34:0] L67_0r1;
  wire L67_0a;
  wire [32:0] L68_0r0;
  wire [32:0] L68_0r1;
  wire L68_0a;
  wire L69_0r;
  wire L69_0a;
  wire [31:0] L70_0r0;
  wire [31:0] L70_0r1;
  wire L70_0a;
  wire L71_0r;
  wire L71_0a;
  wire L72_0r;
  wire L72_0a;
  wire L74_0r;
  wire L74_0a;
  wire [31:0] L76_0r0;
  wire [31:0] L76_0r1;
  wire L76_0a;
  wire L77_0r;
  wire L77_0a;
  wire L78_0r;
  wire L78_0a;
  wire L80_0r0;
  wire L80_0r1;
  wire L80_0a;
  wire L81_0r;
  wire L81_0a;
  wire L82_0r;
  wire L82_0a;
  wire L83_0r;
  wire L83_0a;
  wire L84_0r;
  wire L84_0a;
  wire L85_0r;
  wire L85_0a;
  wire L86_0r;
  wire L86_0a;
  wire L87_0r;
  wire L87_0a;
  wire [1:0] L88_0r0;
  wire [1:0] L88_0r1;
  wire L88_0a;
  wire [1:0] L89_0r0;
  wire [1:0] L89_0r1;
  wire L89_0a;
  wire [1:0] L90_0r0;
  wire [1:0] L90_0r1;
  wire L90_0a;
  wire [1:0] L91_0r0;
  wire [1:0] L91_0r1;
  wire L91_0a;
  wire L92_0r0;
  wire L92_0r1;
  wire L92_0a;
  wire L93_0r;
  wire L93_0a;
  wire L94_0r;
  wire L94_0a;
  wire L95_0r0;
  wire L95_0r1;
  wire L95_0a;
  wire L96_0r;
  wire L96_0a;
  wire L97_0r0;
  wire L97_0r1;
  wire L97_0a;
  wire L98_0r;
  wire L98_0a;
  wire L99_0r0;
  wire L99_0r1;
  wire L99_0a;
  wire [2:0] L100_0r0;
  wire [2:0] L100_0r1;
  wire L100_0a;
  wire [2:0] L101_0r0;
  wire [2:0] L101_0r1;
  wire L101_0a;
  wire [2:0] L102_0r0;
  wire [2:0] L102_0r1;
  wire L102_0a;
  wire [2:0] L103_0r0;
  wire [2:0] L103_0r1;
  wire L103_0a;
  wire [2:0] L104_0r0;
  wire [2:0] L104_0r1;
  wire L104_0a;
  wire [31:0] L105_0r0;
  wire [31:0] L105_0r1;
  wire L105_0a;
  wire L106_0r;
  wire L106_0a;
  wire L107_0r;
  wire L107_0a;
  wire [31:0] L108_0r0;
  wire [31:0] L108_0r1;
  wire L108_0a;
  wire L109_0r;
  wire L109_0a;
  wire [31:0] L110_0r0;
  wire [31:0] L110_0r1;
  wire L110_0a;
  wire L111_0r;
  wire L111_0a;
  wire [31:0] L112_0r0;
  wire [31:0] L112_0r1;
  wire L112_0a;
  wire [2:0] L113_0r0;
  wire [2:0] L113_0r1;
  wire L113_0a;
  wire [2:0] L114_0r0;
  wire [2:0] L114_0r1;
  wire L114_0a;
  wire [2:0] L115_0r0;
  wire [2:0] L115_0r1;
  wire L115_0a;
  wire [2:0] L116_0r0;
  wire [2:0] L116_0r1;
  wire L116_0a;
  wire [2:0] L117_0r0;
  wire [2:0] L117_0r1;
  wire L117_0a;
  tko0m32_1nm32b0 I0 (L2_0r, L2_0a, L4_0r0[31:0], L4_0r1[31:0], L4_0a, reset);
  tko0m1_1nm1b1 I1 (L6_0r, L6_0a, L8_0r0, L8_0r1, L8_0a, reset);
  tkj0m0_0 I2 (L5_0r, L5_0a, L9_0r, L9_0a, L39_0r, L39_0a, reset);
  tkf0mo0w0_o0w0 I3 (L22_0r, L22_0a, L17_0r, L17_0a, L21_0r, L21_0a, reset);
  tkj0m0_0 I4 (L20_0r, L20_0a, L21_0r, L21_0a, L23_0r, L23_0a, reset);
  tkvnewPc32_wo0w32_ro0w32 I5 (L24_0r0[31:0], L24_0r1[31:0], L24_0a, L22_0r, L22_0a, L17_0r, L17_0a, L19_0r0[31:0], L19_0r1[31:0], L19_0a, reset);
  tko0m1_1nm1b1 I6 (L27_0r, L27_0a, L29_0r0, L29_0r1, L29_0a, reset);
  tkf0mo0w0_o0w0 I7 (L31_0r, L31_0a, L26_0r, L26_0a, L27_0r, L27_0a, reset);
  tkj0m0_0 I8 (L23_0r, L23_0a, L30_0r, L30_0a, L33_0r, L33_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I9 (L13_0r0, L13_0r1, L13_0a, L14_0r, L14_0a, L31_0r, L31_0a, reset);
  tkm2x0b I10 (L15_0r, L15_0a, L34_0r, L34_0a, L35_0r, L35_0a, reset);
  tkvdoFetch1_wo0w1_ro0w1 I11 (L36_0r0, L36_0r1, L36_0a, L12_0r, L12_0a, L12_0r, L12_0a, L13_0r0, L13_0r1, L13_0a, reset);
  tkm2x0b I12 (L39_0r, L39_0a, L35_0r, L35_0a, L38_0r, L38_0a, reset);
  tkj33m32_1 I13 (L48_0r0[31:0], L48_0r1[31:0], L48_0a, L50_0r0, L50_0r1, L50_0a, L51_0r0[32:0], L51_0r1[32:0], L51_0a, reset);
  tkj65m32_33 I14 (L46_0r0[31:0], L46_0r1[31:0], L46_0a, L51_0r0[32:0], L51_0r1[32:0], L51_0a, L54_0r0[64:0], L54_0r1[64:0], L54_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I15 (L53_0r, L53_0a, L45_0r, L45_0a, L47_0r, L47_0a, L49_0r, L49_0a, reset);
  tkf0mo0w0_o0w0 I16 (L57_0r, L57_0a, L53_0r, L53_0a, L56_0r, L56_0a, reset);
  tkj0m0_0 I17 (L55_0r, L55_0a, L56_0r, L56_0a, L58_0r, L58_0a, reset);
  tkvfinst32_wo0w32_ro0w32 I18 (L59_0r0[31:0], L59_0r1[31:0], L59_0a, L57_0r, L57_0a, L45_0r, L45_0a, L46_0r0[31:0], L46_0r1[31:0], L46_0a, reset);
  tko0m3_1nm3b4 I19 (L65_0r, L65_0a, L66_0r0[2:0], L66_0r1[2:0], L66_0a, reset);
  tkj35m32_3 I20 (L64_0r0[31:0], L64_0r1[31:0], L64_0a, L66_0r0[2:0], L66_0r1[2:0], L66_0a, L67_0r0[34:0], L67_0r1[34:0], L67_0a, reset);
  tko35m33_1api0w32b_2api32w3b_3nm1b0_4apt1o0w32bt3o0w1b_5nm30b0_6apt2o0w3bt5o0w30b_7addt4o0w33bt6o0w33b I21 (L67_0r0[34:0], L67_0r1[34:0], L67_0a, L68_0r0[32:0], L68_0r1[32:0], L68_0a, reset);
  tkf33mo0w32 I22 (L68_0r0[32:0], L68_0r1[32:0], L68_0a, L70_0r0[31:0], L70_0r1[31:0], L70_0a, reset);
  tkf0mo0w0_o0w0 I23 (L69_0r, L69_0a, L63_0r, L63_0a, L65_0r, L65_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I24 (L72_0r, L72_0a, L41_0r, L41_0a, L61_0r, L61_0a, L69_0r, L69_0a, reset);
  tkj0m0_0_0 I25 (L44_0r, L44_0a, L58_0r, L58_0a, L71_0r, L71_0a, L82_0r, L82_0a, reset);
  tko0m1_1nm1b0 I26 (L78_0r, L78_0a, L80_0r0, L80_0r1, L80_0a, reset);
  tkf0mo0w0_o0w0 I27 (L82_0r, L82_0a, L74_0r, L74_0a, L78_0r, L78_0a, reset);
  tkj0m0_0 I28 (L77_0r, L77_0a, L81_0r, L81_0a, L83_0r, L83_0a, reset);
  tkf0mo0w0_o0w0 I29 (L14_0r, L14_0a, L84_0r, L84_0a, L85_0r, L85_0a, reset);
  tkf0mo0w0_o0w0 I30 (L33_0r, L33_0a, L86_0r, L86_0a, L87_0r, L87_0a, reset);
  tkm2x0b I31 (L84_0r, L84_0a, L86_0r, L86_0a, L72_0r, L72_0a, reset);
  tko0m2_1nm2b1 I32 (L85_0r, L85_0a, L88_0r0[1:0], L88_0r1[1:0], L88_0a, reset);
  tko0m2_1nm2b2 I33 (L87_0r, L87_0a, L89_0r0[1:0], L89_0r1[1:0], L89_0a, reset);
  tkm2x2b I34 (L88_0r0[1:0], L88_0r1[1:0], L88_0a, L89_0r0[1:0], L89_0r1[1:0], L89_0a, L90_0r0[1:0], L90_0r1[1:0], L90_0a, reset);
  tkj2m0_2 I35 (L83_0r, L83_0a, L90_0r0[1:0], L90_0r1[1:0], L90_0a, L91_0r0[1:0], L91_0r1[1:0], L91_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I36 (L91_0r0[1:0], L91_0r1[1:0], L91_0a, L15_0r, L15_0a, L34_0r, L34_0a, reset);
  tkf1mo0w0_o0w1 I37 (L80_0r0, L80_0r1, L80_0a, L94_0r, L94_0a, L95_0r0, L95_0r1, L95_0a, reset);
  tkf1mo0w0_o0w1 I38 (L29_0r0, L29_0r1, L29_0a, L96_0r, L96_0a, L97_0r0, L97_0r1, L97_0a, reset);
  tkf1mo0w0_o0w1 I39 (L8_0r0, L8_0r1, L8_0a, L98_0r, L98_0a, L99_0r0, L99_0r1, L99_0a, reset);
  tkm3x1b I40 (L95_0r0, L95_0r1, L95_0a, L97_0r0, L97_0r1, L97_0a, L99_0r0, L99_0r1, L99_0a, L92_0r0, L92_0r1, L92_0a, reset);
  tko0m3_1nm3b1 I41 (L94_0r, L94_0a, L100_0r0[2:0], L100_0r1[2:0], L100_0a, reset);
  tko0m3_1nm3b2 I42 (L96_0r, L96_0a, L101_0r0[2:0], L101_0r1[2:0], L101_0a, reset);
  tko0m3_1nm3b4 I43 (L98_0r, L98_0a, L102_0r0[2:0], L102_0r1[2:0], L102_0a, reset);
  tkm3x3b I44 (L100_0r0[2:0], L100_0r1[2:0], L100_0a, L101_0r0[2:0], L101_0r1[2:0], L101_0a, L102_0r0[2:0], L102_0r1[2:0], L102_0a, L103_0r0[2:0], L103_0r1[2:0], L103_0a, reset);
  tkj3m0_3 I45 (L93_0r, L93_0a, L103_0r0[2:0], L103_0r1[2:0], L103_0a, L104_0r0[2:0], L104_0r1[2:0], L104_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_4o0w0 I46 (L104_0r0[2:0], L104_0r1[2:0], L104_0a, L81_0r, L81_0a, L30_0r, L30_0a, L9_0r, L9_0a, reset);
  tkvnewStream1_wo0w1_ro0w1 I47 (L92_0r0, L92_0r1, L92_0a, L93_0r, L93_0a, L49_0r, L49_0a, L50_0r0, L50_0r1, L50_0a, reset);
  tkvpcTemp32_wo0w32_ro0w32 I48 (L70_0r0[31:0], L70_0r1[31:0], L70_0a, L71_0r, L71_0a, L74_0r, L74_0a, L76_0r0[31:0], L76_0r1[31:0], L76_0a, reset);
  tkf32mo0w0_o0w32 I49 (L76_0r0[31:0], L76_0r1[31:0], L76_0a, L107_0r, L107_0a, L108_0r0[31:0], L108_0r1[31:0], L108_0a, reset);
  tkf32mo0w0_o0w32 I50 (L19_0r0[31:0], L19_0r1[31:0], L19_0a, L109_0r, L109_0a, L110_0r0[31:0], L110_0r1[31:0], L110_0a, reset);
  tkf32mo0w0_o0w32 I51 (L4_0r0[31:0], L4_0r1[31:0], L4_0a, L111_0r, L111_0a, L112_0r0[31:0], L112_0r1[31:0], L112_0a, reset);
  tkm3x32b I52 (L108_0r0[31:0], L108_0r1[31:0], L108_0a, L110_0r0[31:0], L110_0r1[31:0], L110_0a, L112_0r0[31:0], L112_0r1[31:0], L112_0a, L105_0r0[31:0], L105_0r1[31:0], L105_0a, reset);
  tko0m3_1nm3b1 I53 (L107_0r, L107_0a, L113_0r0[2:0], L113_0r1[2:0], L113_0a, reset);
  tko0m3_1nm3b2 I54 (L109_0r, L109_0a, L114_0r0[2:0], L114_0r1[2:0], L114_0a, reset);
  tko0m3_1nm3b4 I55 (L111_0r, L111_0a, L115_0r0[2:0], L115_0r1[2:0], L115_0a, reset);
  tkm3x3b I56 (L113_0r0[2:0], L113_0r1[2:0], L113_0a, L114_0r0[2:0], L114_0r1[2:0], L114_0a, L115_0r0[2:0], L115_0r1[2:0], L115_0a, L116_0r0[2:0], L116_0r1[2:0], L116_0a, reset);
  tkj3m0_3 I57 (L106_0r, L106_0a, L116_0r0[2:0], L116_0r1[2:0], L116_0a, L117_0r0[2:0], L117_0r1[2:0], L117_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_4o0w0 I58 (L117_0r0[2:0], L117_0r1[2:0], L117_0a, L77_0r, L77_0a, L20_0r, L20_0a, L5_0r, L5_0a, reset);
  tkvpc32_wo0w32_ro0w32o0w32o0w32 I59 (L105_0r0[31:0], L105_0r1[31:0], L105_0a, L106_0r, L106_0a, L63_0r, L63_0a, L47_0r, L47_0a, L41_0r, L41_0a, L64_0r0[31:0], L64_0r1[31:0], L64_0a, L48_0r0[31:0], L48_0r1[31:0], L48_0a, L43_0r0[31:0], L43_0r1[31:0], L43_0a, reset);
  tkj1m1_0 I60 (doFetch_0r0, doFetch_0r1, doFetch_0a, L38_0r, L38_0a, L36_0r0, L36_0r1, L36_0a, reset);
  tkj32m32_0 I61 (newPc_0r0[31:0], newPc_0r1[31:0], newPc_0a, L26_0r, L26_0a, L24_0r0[31:0], L24_0r1[31:0], L24_0a, reset);
  tkf65mo0w0_o0w65 I62 (L54_0r0[64:0], L54_0r1[64:0], L54_0a, L55_0r, L55_0a, inst_0r0[64:0], inst_0r1[64:0], inst_0a, reset);
  tkf32mo0w0_o0w32 I63 (L43_0r0[31:0], L43_0r1[31:0], L43_0a, L44_0r, L44_0a, faddr_0r0[31:0], faddr_0r1[31:0], faddr_0a, reset);
  tkj32m32_0 I64 (finst_0r0[31:0], finst_0r1[31:0], finst_0a, L61_0r, L61_0a, L59_0r0[31:0], L59_0r1[31:0], L59_0a, reset);
  tkr I65 (L2_0r, L2_0a, reset);
  tkr I66 (L6_0r, L6_0a, reset);
endmodule

module teak_Decode (inst_0r0, inst_0r1, inst_0a, decoded_0r0, decoded_0r1, decoded_0a, pc_0r0, pc_0r1, pc_0a, reset);
  input [64:0] inst_0r0;
  input [64:0] inst_0r1;
  output inst_0a;
  output [73:0] decoded_0r0;
  output [73:0] decoded_0r1;
  input decoded_0a;
  output [32:0] pc_0r0;
  output [32:0] pc_0r1;
  input pc_0a;
  input reset;
  wire L3_0r;
  wire L3_0a;
  wire [64:0] L4_0r0;
  wire [64:0] L4_0r1;
  wire L4_0a;
  wire L6_0r;
  wire L6_0a;
  wire L7_0r;
  wire L7_0a;
  wire [32:0] L9_0r0;
  wire [32:0] L9_0r1;
  wire L9_0a;
  wire L10_0r;
  wire L10_0a;
  wire L11_0r;
  wire L11_0a;
  wire [1:0] L12_0r0;
  wire [1:0] L12_0r1;
  wire L12_0a;
  wire L14_0r;
  wire L14_0a;
  wire L15_0r;
  wire L15_0a;
  wire L16_0r;
  wire L16_0a;
  wire [5:0] L17_0r0;
  wire [5:0] L17_0r1;
  wire L17_0a;
  wire L18_0r;
  wire L18_0a;
  wire L19_0r;
  wire L19_0a;
  wire L20_0r;
  wire L20_0a;
  wire L21_0r;
  wire L21_0a;
  wire L22_0r;
  wire L22_0a;
  wire L23_0r;
  wire L23_0a;
  wire [2:0] L24_0r0;
  wire [2:0] L24_0r1;
  wire L24_0a;
  wire L25_0r;
  wire L25_0a;
  wire [3:0] L26_0r0;
  wire [3:0] L26_0r1;
  wire L26_0a;
  wire L27_0r;
  wire L27_0a;
  wire L28_0r0;
  wire L28_0r1;
  wire L28_0a;
  wire L29_0r0;
  wire L29_0r1;
  wire L29_0a;
  wire L30_0r;
  wire L30_0a;
  wire L31_0r0;
  wire L31_0r1;
  wire L31_0a;
  wire L32_0r;
  wire L32_0a;
  wire L33_0r0;
  wire L33_0r1;
  wire L33_0a;
  wire [2:0] L34_0r0;
  wire [2:0] L34_0r1;
  wire L34_0a;
  wire L35_0r;
  wire L35_0a;
  wire [4:0] L36_0r0;
  wire [4:0] L36_0r1;
  wire L36_0a;
  wire L37_0r;
  wire L37_0a;
  wire [4:0] L38_0r0;
  wire [4:0] L38_0r1;
  wire L38_0a;
  wire L39_0r;
  wire L39_0a;
  wire [4:0] L40_0r0;
  wire [4:0] L40_0r1;
  wire L40_0a;
  wire [14:0] L41_0r0;
  wire [14:0] L41_0r1;
  wire L41_0a;
  wire L42_0r;
  wire L42_0a;
  wire L43_0r0;
  wire L43_0r1;
  wire L43_0a;
  wire L44_0r;
  wire L44_0a;
  wire [4:0] L45_0r0;
  wire [4:0] L45_0r1;
  wire L45_0a;
  wire L46_0r;
  wire L46_0a;
  wire [5:0] L47_0r0;
  wire [5:0] L47_0r1;
  wire L47_0a;
  wire L48_0r;
  wire L48_0a;
  wire L49_0r0;
  wire L49_0r1;
  wire L49_0a;
  wire [31:0] L50_0r0;
  wire [31:0] L50_0r1;
  wire L50_0a;
  wire L51_0r;
  wire L51_0a;
  wire [12:0] L52_0r0;
  wire [12:0] L52_0r1;
  wire L52_0a;
  wire L53_0r;
  wire L53_0a;
  wire [3:0] L54_0r0;
  wire [3:0] L54_0r1;
  wire L54_0a;
  wire L56_0r;
  wire L56_0a;
  wire [73:0] L57_0r0;
  wire [73:0] L57_0r1;
  wire L57_0a;
  wire L58_0r;
  wire L58_0a;
  wire L59_0r0;
  wire L59_0r1;
  wire L59_0a;
  wire L61_0r;
  wire L61_0a;
  wire L62_0r;
  wire L62_0a;
  wire L63_0r0;
  wire L63_0r1;
  wire L63_0a;
  wire L64_0r;
  wire L64_0a;
  wire L66_0r0;
  wire L66_0r1;
  wire L66_0a;
  wire L67_0r;
  wire L67_0a;
  wire L68_0r;
  wire L68_0a;
  wire L70_0r0;
  wire L70_0r1;
  wire L70_0a;
  wire L71_0r;
  wire L71_0a;
  wire L72_0r;
  wire L72_0a;
  wire L73_0r;
  wire L73_0a;
  wire L74_0r;
  wire L74_0a;
  wire L75_0r;
  wire L75_0a;
  wire L76_0r;
  wire L76_0a;
  wire L77_0r0;
  wire L77_0r1;
  wire L77_0a;
  wire L78_0r;
  wire L78_0a;
  wire L79_0r0;
  wire L79_0r1;
  wire L79_0a;
  wire L80_0r0;
  wire L80_0r1;
  wire L80_0a;
  wire L81_0r;
  wire L81_0a;
  wire L82_0r0;
  wire L82_0r1;
  wire L82_0a;
  wire [1:0] L83_0r0;
  wire [1:0] L83_0r1;
  wire L83_0a;
  wire [1:0] L84_0r0;
  wire [1:0] L84_0r1;
  wire L84_0a;
  wire [1:0] L85_0r0;
  wire [1:0] L85_0r1;
  wire L85_0a;
  wire [1:0] L86_0r0;
  wire [1:0] L86_0r1;
  wire L86_0a;
  wire L87_0r;
  wire L87_0a;
  wire [2:0] L88_0r0;
  wire [2:0] L88_0r1;
  wire L88_0a;
  wire L90_0r;
  wire L90_0a;
  wire [2:0] L91_0r0;
  wire [2:0] L91_0r1;
  wire L91_0a;
  wire L92_0r;
  wire L92_0a;
  wire L94_0r0;
  wire L94_0r1;
  wire L94_0a;
  wire L95_0r;
  wire L95_0a;
  wire L96_0r;
  wire L96_0a;
  wire L98_0r0;
  wire L98_0r1;
  wire L98_0a;
  wire L99_0r;
  wire L99_0a;
  wire L101_0r;
  wire L101_0a;
  wire [2:0] L102_0r0;
  wire [2:0] L102_0r1;
  wire L102_0a;
  wire L103_0r;
  wire L103_0a;
  wire [3:0] L104_0r0;
  wire [3:0] L104_0r1;
  wire L104_0a;
  wire L105_0r;
  wire L105_0a;
  wire L106_0r0;
  wire L106_0r1;
  wire L106_0a;
  wire L107_0r0;
  wire L107_0r1;
  wire L107_0a;
  wire L108_0r;
  wire L108_0a;
  wire L109_0r0;
  wire L109_0r1;
  wire L109_0a;
  wire L110_0r;
  wire L110_0a;
  wire L111_0r0;
  wire L111_0r1;
  wire L111_0a;
  wire [2:0] L112_0r0;
  wire [2:0] L112_0r1;
  wire L112_0a;
  wire L113_0r;
  wire L113_0a;
  wire [4:0] L114_0r0;
  wire [4:0] L114_0r1;
  wire L114_0a;
  wire L115_0r;
  wire L115_0a;
  wire [4:0] L116_0r0;
  wire [4:0] L116_0r1;
  wire L116_0a;
  wire L117_0r;
  wire L117_0a;
  wire [4:0] L118_0r0;
  wire [4:0] L118_0r1;
  wire L118_0a;
  wire [14:0] L119_0r0;
  wire [14:0] L119_0r1;
  wire L119_0a;
  wire L120_0r0;
  wire L120_0r1;
  wire L120_0a;
  wire L121_0r;
  wire L121_0a;
  wire L122_0r0;
  wire L122_0r1;
  wire L122_0a;
  wire L123_0r;
  wire L123_0a;
  wire [4:0] L124_0r0;
  wire [4:0] L124_0r1;
  wire L124_0a;
  wire L125_0r;
  wire L125_0a;
  wire [5:0] L126_0r0;
  wire [5:0] L126_0r1;
  wire L126_0a;
  wire L127_0r;
  wire L127_0a;
  wire L128_0r0;
  wire L128_0r1;
  wire L128_0a;
  wire [31:0] L129_0r0;
  wire [31:0] L129_0r1;
  wire L129_0a;
  wire L130_0r;
  wire L130_0a;
  wire [12:0] L131_0r0;
  wire [12:0] L131_0r1;
  wire L131_0a;
  wire L132_0r;
  wire L132_0a;
  wire [3:0] L133_0r0;
  wire [3:0] L133_0r1;
  wire L133_0a;
  wire L135_0r;
  wire L135_0a;
  wire [73:0] L136_0r0;
  wire [73:0] L136_0r1;
  wire L136_0a;
  wire L137_0r;
  wire L137_0a;
  wire L138_0r;
  wire L138_0a;
  wire L139_0r;
  wire L139_0a;
  wire L140_0r;
  wire L140_0a;
  wire L141_0r0;
  wire L141_0r1;
  wire L141_0a;
  wire L142_0r;
  wire L142_0a;
  wire L143_0r;
  wire L143_0a;
  wire L144_0r0;
  wire L144_0r1;
  wire L144_0a;
  wire L145_0r;
  wire L145_0a;
  wire L146_0r0;
  wire L146_0r1;
  wire L146_0a;
  wire [1:0] L147_0r0;
  wire [1:0] L147_0r1;
  wire L147_0a;
  wire [1:0] L148_0r0;
  wire [1:0] L148_0r1;
  wire L148_0a;
  wire [1:0] L149_0r0;
  wire [1:0] L149_0r1;
  wire L149_0a;
  wire [1:0] L150_0r0;
  wire [1:0] L150_0r1;
  wire L150_0a;
  wire [3:0] L151_0r0;
  wire [3:0] L151_0r1;
  wire L151_0a;
  wire L152_0r;
  wire L152_0a;
  wire [2:0] L153_0r0;
  wire [2:0] L153_0r1;
  wire L153_0a;
  wire L154_0r;
  wire L154_0a;
  wire L155_0r0;
  wire L155_0r1;
  wire L155_0a;
  wire L156_0r;
  wire L156_0a;
  wire L158_0r;
  wire L158_0a;
  wire L159_0r;
  wire L159_0a;
  wire L160_0r;
  wire L160_0a;
  wire L161_0r;
  wire L161_0a;
  wire L162_0r;
  wire L162_0a;
  wire L163_0r0;
  wire L163_0r1;
  wire L163_0a;
  wire L164_0r;
  wire L164_0a;
  wire L166_0r0;
  wire L166_0r1;
  wire L166_0a;
  wire L167_0r;
  wire L167_0a;
  wire L168_0r;
  wire L168_0a;
  wire L170_0r0;
  wire L170_0r1;
  wire L170_0a;
  wire L171_0r;
  wire L171_0a;
  wire L172_0r;
  wire L172_0a;
  wire L173_0r;
  wire L173_0a;
  wire [5:0] L174_0r0;
  wire [5:0] L174_0r1;
  wire L174_0a;
  wire L176_0r;
  wire L176_0a;
  wire [3:0] L178_0r0;
  wire [3:0] L178_0r1;
  wire L178_0a;
  wire L179_0r;
  wire L179_0a;
  wire L180_0r;
  wire L180_0a;
  wire [2:0] L182_0r0;
  wire [2:0] L182_0r1;
  wire L182_0a;
  wire L183_0r;
  wire L183_0a;
  wire L184_0r;
  wire L184_0a;
  wire L185_0r;
  wire L185_0a;
  wire L186_0r;
  wire L186_0a;
  wire [3:0] L188_0r0;
  wire [3:0] L188_0r1;
  wire L188_0a;
  wire L189_0r;
  wire L189_0a;
  wire L190_0r;
  wire L190_0a;
  wire [2:0] L192_0r0;
  wire [2:0] L192_0r1;
  wire L192_0a;
  wire L193_0r;
  wire L193_0a;
  wire L194_0r;
  wire L194_0a;
  wire L195_0r;
  wire L195_0a;
  wire L196_0r;
  wire L196_0a;
  wire [3:0] L198_0r0;
  wire [3:0] L198_0r1;
  wire L198_0a;
  wire L199_0r;
  wire L199_0a;
  wire L200_0r;
  wire L200_0a;
  wire [2:0] L202_0r0;
  wire [2:0] L202_0r1;
  wire L202_0a;
  wire L203_0r;
  wire L203_0a;
  wire L204_0r;
  wire L204_0a;
  wire L205_0r;
  wire L205_0a;
  wire L206_0r;
  wire L206_0a;
  wire [3:0] L208_0r0;
  wire [3:0] L208_0r1;
  wire L208_0a;
  wire L209_0r;
  wire L209_0a;
  wire L210_0r;
  wire L210_0a;
  wire [2:0] L212_0r0;
  wire [2:0] L212_0r1;
  wire L212_0a;
  wire L213_0r;
  wire L213_0a;
  wire L214_0r;
  wire L214_0a;
  wire L215_0r;
  wire L215_0a;
  wire L216_0r;
  wire L216_0a;
  wire [3:0] L218_0r0;
  wire [3:0] L218_0r1;
  wire L218_0a;
  wire L219_0r;
  wire L219_0a;
  wire L220_0r;
  wire L220_0a;
  wire [2:0] L222_0r0;
  wire [2:0] L222_0r1;
  wire L222_0a;
  wire L223_0r;
  wire L223_0a;
  wire L224_0r;
  wire L224_0a;
  wire L225_0r;
  wire L225_0a;
  wire L226_0r;
  wire L226_0a;
  wire [3:0] L228_0r0;
  wire [3:0] L228_0r1;
  wire L228_0a;
  wire L229_0r;
  wire L229_0a;
  wire L230_0r;
  wire L230_0a;
  wire [2:0] L232_0r0;
  wire [2:0] L232_0r1;
  wire L232_0a;
  wire L233_0r;
  wire L233_0a;
  wire L234_0r;
  wire L234_0a;
  wire L235_0r;
  wire L235_0a;
  wire L236_0r;
  wire L236_0a;
  wire [3:0] L238_0r0;
  wire [3:0] L238_0r1;
  wire L238_0a;
  wire L239_0r;
  wire L239_0a;
  wire L240_0r;
  wire L240_0a;
  wire [2:0] L242_0r0;
  wire [2:0] L242_0r1;
  wire L242_0a;
  wire L243_0r;
  wire L243_0a;
  wire L244_0r;
  wire L244_0a;
  wire L245_0r;
  wire L245_0a;
  wire L246_0r;
  wire L246_0a;
  wire [3:0] L248_0r0;
  wire [3:0] L248_0r1;
  wire L248_0a;
  wire L249_0r;
  wire L249_0a;
  wire L250_0r;
  wire L250_0a;
  wire [2:0] L252_0r0;
  wire [2:0] L252_0r1;
  wire L252_0a;
  wire L253_0r;
  wire L253_0a;
  wire L254_0r;
  wire L254_0a;
  wire L255_0r;
  wire L255_0a;
  wire L256_0r;
  wire L256_0a;
  wire [3:0] L258_0r0;
  wire [3:0] L258_0r1;
  wire L258_0a;
  wire L259_0r;
  wire L259_0a;
  wire L260_0r;
  wire L260_0a;
  wire [2:0] L262_0r0;
  wire [2:0] L262_0r1;
  wire L262_0a;
  wire L263_0r;
  wire L263_0a;
  wire L264_0r;
  wire L264_0a;
  wire L265_0r;
  wire L265_0a;
  wire L266_0r;
  wire L266_0a;
  wire [3:0] L268_0r0;
  wire [3:0] L268_0r1;
  wire L268_0a;
  wire L269_0r;
  wire L269_0a;
  wire L270_0r;
  wire L270_0a;
  wire [2:0] L272_0r0;
  wire [2:0] L272_0r1;
  wire L272_0a;
  wire L273_0r;
  wire L273_0a;
  wire L274_0r;
  wire L274_0a;
  wire L275_0r;
  wire L275_0a;
  wire L276_0r;
  wire L276_0a;
  wire [3:0] L278_0r0;
  wire [3:0] L278_0r1;
  wire L278_0a;
  wire L279_0r;
  wire L279_0a;
  wire L280_0r;
  wire L280_0a;
  wire [2:0] L282_0r0;
  wire [2:0] L282_0r1;
  wire L282_0a;
  wire L283_0r;
  wire L283_0a;
  wire L284_0r;
  wire L284_0a;
  wire L285_0r;
  wire L285_0a;
  wire L286_0r;
  wire L286_0a;
  wire L287_0r;
  wire L287_0a;
  wire L288_0r;
  wire L288_0a;
  wire L289_0r;
  wire L289_0a;
  wire L290_0r0;
  wire L290_0r1;
  wire L290_0a;
  wire L291_0r;
  wire L291_0a;
  wire L292_0r0;
  wire L292_0r1;
  wire L292_0a;
  wire L293_0r0;
  wire L293_0r1;
  wire L293_0a;
  wire L294_0r;
  wire L294_0a;
  wire L295_0r0;
  wire L295_0r1;
  wire L295_0a;
  wire [1:0] L296_0r0;
  wire [1:0] L296_0r1;
  wire L296_0a;
  wire [1:0] L297_0r0;
  wire [1:0] L297_0r1;
  wire L297_0a;
  wire [1:0] L298_0r0;
  wire [1:0] L298_0r1;
  wire L298_0a;
  wire [1:0] L299_0r0;
  wire [1:0] L299_0r1;
  wire L299_0a;
  wire L300_0r;
  wire L300_0a;
  wire [2:0] L301_0r0;
  wire [2:0] L301_0r1;
  wire L301_0a;
  wire L302_0r;
  wire L302_0a;
  wire [2:0] L303_0r0;
  wire [2:0] L303_0r1;
  wire L303_0a;
  wire L304_0r;
  wire L304_0a;
  wire [2:0] L305_0r0;
  wire [2:0] L305_0r1;
  wire L305_0a;
  wire L306_0r;
  wire L306_0a;
  wire [2:0] L307_0r0;
  wire [2:0] L307_0r1;
  wire L307_0a;
  wire L308_0r;
  wire L308_0a;
  wire [2:0] L309_0r0;
  wire [2:0] L309_0r1;
  wire L309_0a;
  wire L310_0r;
  wire L310_0a;
  wire [2:0] L311_0r0;
  wire [2:0] L311_0r1;
  wire L311_0a;
  wire L312_0r;
  wire L312_0a;
  wire [2:0] L313_0r0;
  wire [2:0] L313_0r1;
  wire L313_0a;
  wire L314_0r;
  wire L314_0a;
  wire [2:0] L315_0r0;
  wire [2:0] L315_0r1;
  wire L315_0a;
  wire L316_0r;
  wire L316_0a;
  wire [2:0] L317_0r0;
  wire [2:0] L317_0r1;
  wire L317_0a;
  wire L318_0r;
  wire L318_0a;
  wire [2:0] L319_0r0;
  wire [2:0] L319_0r1;
  wire L319_0a;
  wire L320_0r;
  wire L320_0a;
  wire [2:0] L321_0r0;
  wire [2:0] L321_0r1;
  wire L321_0a;
  wire [2:0] L322_0r0;
  wire [2:0] L322_0r1;
  wire L322_0a;
  wire L323_0r;
  wire L323_0a;
  wire [2:0] L324_0r0;
  wire [2:0] L324_0r1;
  wire L324_0a;
  wire [10:0] L325_0r0;
  wire [10:0] L325_0r1;
  wire L325_0a;
  wire [10:0] L326_0r0;
  wire [10:0] L326_0r1;
  wire L326_0a;
  wire [10:0] L327_0r0;
  wire [10:0] L327_0r1;
  wire L327_0a;
  wire [10:0] L328_0r0;
  wire [10:0] L328_0r1;
  wire L328_0a;
  wire [10:0] L329_0r0;
  wire [10:0] L329_0r1;
  wire L329_0a;
  wire [10:0] L330_0r0;
  wire [10:0] L330_0r1;
  wire L330_0a;
  wire [10:0] L331_0r0;
  wire [10:0] L331_0r1;
  wire L331_0a;
  wire [10:0] L332_0r0;
  wire [10:0] L332_0r1;
  wire L332_0a;
  wire [10:0] L333_0r0;
  wire [10:0] L333_0r1;
  wire L333_0a;
  wire [10:0] L334_0r0;
  wire [10:0] L334_0r1;
  wire L334_0a;
  wire [10:0] L335_0r0;
  wire [10:0] L335_0r1;
  wire L335_0a;
  wire [10:0] L336_0r0;
  wire [10:0] L336_0r1;
  wire L336_0a;
  wire [10:0] L337_0r0;
  wire [10:0] L337_0r1;
  wire L337_0a;
  wire L338_0r;
  wire L338_0a;
  wire [3:0] L339_0r0;
  wire [3:0] L339_0r1;
  wire L339_0a;
  wire L340_0r;
  wire L340_0a;
  wire [3:0] L341_0r0;
  wire [3:0] L341_0r1;
  wire L341_0a;
  wire L342_0r;
  wire L342_0a;
  wire [3:0] L343_0r0;
  wire [3:0] L343_0r1;
  wire L343_0a;
  wire L344_0r;
  wire L344_0a;
  wire [3:0] L345_0r0;
  wire [3:0] L345_0r1;
  wire L345_0a;
  wire L346_0r;
  wire L346_0a;
  wire [3:0] L347_0r0;
  wire [3:0] L347_0r1;
  wire L347_0a;
  wire L348_0r;
  wire L348_0a;
  wire [3:0] L349_0r0;
  wire [3:0] L349_0r1;
  wire L349_0a;
  wire L350_0r;
  wire L350_0a;
  wire [3:0] L351_0r0;
  wire [3:0] L351_0r1;
  wire L351_0a;
  wire L352_0r;
  wire L352_0a;
  wire [3:0] L353_0r0;
  wire [3:0] L353_0r1;
  wire L353_0a;
  wire L354_0r;
  wire L354_0a;
  wire [3:0] L355_0r0;
  wire [3:0] L355_0r1;
  wire L355_0a;
  wire L356_0r;
  wire L356_0a;
  wire [3:0] L357_0r0;
  wire [3:0] L357_0r1;
  wire L357_0a;
  wire L358_0r;
  wire L358_0a;
  wire [3:0] L359_0r0;
  wire [3:0] L359_0r1;
  wire L359_0a;
  wire [3:0] L360_0r0;
  wire [3:0] L360_0r1;
  wire L360_0a;
  wire L361_0r;
  wire L361_0a;
  wire [3:0] L362_0r0;
  wire [3:0] L362_0r1;
  wire L362_0a;
  wire [10:0] L363_0r0;
  wire [10:0] L363_0r1;
  wire L363_0a;
  wire [10:0] L364_0r0;
  wire [10:0] L364_0r1;
  wire L364_0a;
  wire [10:0] L365_0r0;
  wire [10:0] L365_0r1;
  wire L365_0a;
  wire [10:0] L366_0r0;
  wire [10:0] L366_0r1;
  wire L366_0a;
  wire [10:0] L367_0r0;
  wire [10:0] L367_0r1;
  wire L367_0a;
  wire [10:0] L368_0r0;
  wire [10:0] L368_0r1;
  wire L368_0a;
  wire [10:0] L369_0r0;
  wire [10:0] L369_0r1;
  wire L369_0a;
  wire [10:0] L370_0r0;
  wire [10:0] L370_0r1;
  wire L370_0a;
  wire [10:0] L371_0r0;
  wire [10:0] L371_0r1;
  wire L371_0a;
  wire [10:0] L372_0r0;
  wire [10:0] L372_0r1;
  wire L372_0a;
  wire [10:0] L373_0r0;
  wire [10:0] L373_0r1;
  wire L373_0a;
  wire [10:0] L374_0r0;
  wire [10:0] L374_0r1;
  wire L374_0a;
  wire [10:0] L375_0r0;
  wire [10:0] L375_0r1;
  wire L375_0a;
  wire L376_0r;
  wire L376_0a;
  wire [2:0] L377_0r0;
  wire [2:0] L377_0r1;
  wire L377_0a;
  wire L379_0r;
  wire L379_0a;
  wire L380_0r;
  wire L380_0a;
  wire L381_0r;
  wire L381_0a;
  wire [2:0] L382_0r0;
  wire [2:0] L382_0r1;
  wire L382_0a;
  wire L383_0r;
  wire L383_0a;
  wire [3:0] L384_0r0;
  wire [3:0] L384_0r1;
  wire L384_0a;
  wire L385_0r;
  wire L385_0a;
  wire [2:0] L386_0r0;
  wire [2:0] L386_0r1;
  wire L386_0a;
  wire L387_0r;
  wire L387_0a;
  wire [14:0] L388_0r0;
  wire [14:0] L388_0r1;
  wire L388_0a;
  wire L389_0r;
  wire L389_0a;
  wire L390_0r0;
  wire L390_0r1;
  wire L390_0a;
  wire L391_0r;
  wire L391_0a;
  wire [4:0] L392_0r0;
  wire [4:0] L392_0r1;
  wire L392_0a;
  wire L393_0r;
  wire L393_0a;
  wire [5:0] L394_0r0;
  wire [5:0] L394_0r1;
  wire L394_0a;
  wire L395_0r;
  wire L395_0a;
  wire L396_0r0;
  wire L396_0r1;
  wire L396_0a;
  wire [31:0] L397_0r0;
  wire [31:0] L397_0r1;
  wire L397_0a;
  wire L398_0r;
  wire L398_0a;
  wire [1:0] L399_0r0;
  wire [1:0] L399_0r1;
  wire L399_0a;
  wire L400_0r;
  wire L400_0a;
  wire [21:0] L401_0r0;
  wire [21:0] L401_0r1;
  wire L401_0a;
  wire [23:0] L402_0r0;
  wire [23:0] L402_0r1;
  wire L402_0a;
  wire L403_0r;
  wire L403_0a;
  wire [3:0] L404_0r0;
  wire [3:0] L404_0r1;
  wire L404_0a;
  wire L406_0r;
  wire L406_0a;
  wire [73:0] L407_0r0;
  wire [73:0] L407_0r1;
  wire L407_0a;
  wire L408_0r;
  wire L408_0a;
  wire L409_0r;
  wire L409_0a;
  wire [2:0] L410_0r0;
  wire [2:0] L410_0r1;
  wire L410_0a;
  wire L411_0r;
  wire L411_0a;
  wire [3:0] L412_0r0;
  wire [3:0] L412_0r1;
  wire L412_0a;
  wire L413_0r;
  wire L413_0a;
  wire [2:0] L414_0r0;
  wire [2:0] L414_0r1;
  wire L414_0a;
  wire L415_0r;
  wire L415_0a;
  wire [14:0] L416_0r0;
  wire [14:0] L416_0r1;
  wire L416_0a;
  wire L417_0r;
  wire L417_0a;
  wire L418_0r0;
  wire L418_0r1;
  wire L418_0a;
  wire L419_0r;
  wire L419_0a;
  wire [4:0] L420_0r0;
  wire [4:0] L420_0r1;
  wire L420_0a;
  wire L421_0r;
  wire L421_0a;
  wire [5:0] L422_0r0;
  wire [5:0] L422_0r1;
  wire L422_0a;
  wire L423_0r;
  wire L423_0a;
  wire L424_0r0;
  wire L424_0r1;
  wire L424_0a;
  wire L425_0r;
  wire L425_0a;
  wire [9:0] L426_0r0;
  wire [9:0] L426_0r1;
  wire L426_0a;
  wire L427_0r;
  wire L427_0a;
  wire [21:0] L428_0r0;
  wire [21:0] L428_0r1;
  wire L428_0a;
  wire [31:0] L429_0r0;
  wire [31:0] L429_0r1;
  wire L429_0a;
  wire L430_0r;
  wire L430_0a;
  wire [3:0] L431_0r0;
  wire [3:0] L431_0r1;
  wire L431_0a;
  wire L433_0r;
  wire L433_0a;
  wire [73:0] L434_0r0;
  wire [73:0] L434_0r1;
  wire L434_0a;
  wire L435_0r;
  wire L435_0a;
  wire L436_0r;
  wire L436_0a;
  wire L437_0r;
  wire L437_0a;
  wire L438_0r;
  wire L438_0a;
  wire L439_0r;
  wire L439_0a;
  wire L441_0r;
  wire L441_0a;
  wire [73:0] L443_0r0;
  wire [73:0] L443_0r1;
  wire L443_0a;
  wire L444_0r;
  wire L444_0a;
  wire L445_0r;
  wire L445_0a;
  wire L446_0r;
  wire L446_0a;
  wire L447_0r;
  wire L447_0a;
  wire L448_0r;
  wire L448_0a;
  wire L449_0r;
  wire L449_0a;
  wire L450_0r;
  wire L450_0a;
  wire L451_0r;
  wire L451_0a;
  wire L452_0r;
  wire L452_0a;
  wire [3:0] L453_0r0;
  wire [3:0] L453_0r1;
  wire L453_0a;
  wire [3:0] L454_0r0;
  wire [3:0] L454_0r1;
  wire L454_0a;
  wire [3:0] L455_0r0;
  wire [3:0] L455_0r1;
  wire L455_0a;
  wire [3:0] L456_0r0;
  wire [3:0] L456_0r1;
  wire L456_0a;
  wire [3:0] L457_0r0;
  wire [3:0] L457_0r1;
  wire L457_0a;
  wire [3:0] L458_0r0;
  wire [3:0] L458_0r1;
  wire L458_0a;
  wire L460_0r;
  wire L460_0a;
  wire [73:0] L461_0r0;
  wire [73:0] L461_0r1;
  wire L461_0a;
  wire L462_0r;
  wire L462_0a;
  wire [73:0] L463_0r0;
  wire [73:0] L463_0r1;
  wire L463_0a;
  wire L464_0r;
  wire L464_0a;
  wire [73:0] L465_0r0;
  wire [73:0] L465_0r1;
  wire L465_0a;
  wire L466_0r;
  wire L466_0a;
  wire [73:0] L467_0r0;
  wire [73:0] L467_0r1;
  wire L467_0a;
  wire L468_0r;
  wire L468_0a;
  wire [73:0] L469_0r0;
  wire [73:0] L469_0r1;
  wire L469_0a;
  wire [73:0] L470_0r0;
  wire [73:0] L470_0r1;
  wire L470_0a;
  wire L471_0r;
  wire L471_0a;
  wire [4:0] L473_0r0;
  wire [4:0] L473_0r1;
  wire L473_0a;
  wire [4:0] L474_0r0;
  wire [4:0] L474_0r1;
  wire L474_0a;
  wire [4:0] L475_0r0;
  wire [4:0] L475_0r1;
  wire L475_0a;
  wire [4:0] L476_0r0;
  wire [4:0] L476_0r1;
  wire L476_0a;
  wire [4:0] L477_0r0;
  wire [4:0] L477_0r1;
  wire L477_0a;
  wire [4:0] L478_0r0;
  wire [4:0] L478_0r1;
  wire L478_0a;
  wire [4:0] L479_0r0;
  wire [4:0] L479_0r1;
  wire L479_0a;
  tkf0mo0w0_o0w0 I0 (L21_0r, L21_0a, L18_0r, L18_0a, L19_0r, L19_0a, reset);
  tkj0m0_0 I1 (L18_0r, L18_0a, L20_0r, L20_0a, L22_0r, L22_0a, reset);
  tko0m3_1nm3b2 I2 (L23_0r, L23_0a, L24_0r0[2:0], L24_0r1[2:0], L24_0a, reset);
  tko0m4_1nm4b8 I3 (L25_0r, L25_0a, L26_0r0[3:0], L26_0r1[3:0], L26_0a, reset);
  tko0m1_1nm1b1 I4 (L27_0r, L27_0a, L28_0r0, L28_0r1, L28_0a, reset);
  tko1m1_1noti0w1b I5 (L31_0r0, L31_0r1, L31_0a, L29_0r0, L29_0r1, L29_0a, reset);
  tko0m1_1nm1b0 I6 (L32_0r, L32_0a, L33_0r0, L33_0r1, L33_0a, reset);
  tkj3m1_1_1 I7 (L28_0r0, L28_0r1, L28_0a, L29_0r0, L29_0r1, L29_0a, L33_0r0, L33_0r1, L33_0a, L34_0r0[2:0], L34_0r1[2:0], L34_0a, reset);
  tko0m5_1nm5b0 I8 (L39_0r, L39_0a, L40_0r0[4:0], L40_0r1[4:0], L40_0a, reset);
  tkj15m5_5_5 I9 (L36_0r0[4:0], L36_0r1[4:0], L36_0a, L38_0r0[4:0], L38_0r1[4:0], L38_0a, L40_0r0[4:0], L40_0r1[4:0], L40_0a, L41_0r0[14:0], L41_0r1[14:0], L41_0a, reset);
  tko0m1_1nm1b1 I10 (L42_0r, L42_0a, L43_0r0, L43_0r1, L43_0a, reset);
  tko13m32_1ap19xi12w1b_2api0w13bt1o0w19b I11 (L52_0r0[12:0], L52_0r1[12:0], L52_0a, L50_0r0[31:0], L50_0r1[31:0], L50_0a, reset);
  tko0m4_1nm4b7 I12 (L53_0r, L53_0a, L54_0r0[3:0], L54_0r1[3:0], L54_0a, reset);
  tkj74m3_4_3_15_1_5_6_1_32_4 I13 (L24_0r0[2:0], L24_0r1[2:0], L24_0a, L26_0r0[3:0], L26_0r1[3:0], L26_0a, L34_0r0[2:0], L34_0r1[2:0], L34_0a, L41_0r0[14:0], L41_0r1[14:0], L41_0a, L43_0r0, L43_0r1, L43_0a, L45_0r0[4:0], L45_0r1[4:0], L45_0a, L47_0r0[5:0], L47_0r1[5:0], L47_0a, L49_0r0, L49_0r1, L49_0a, L50_0r0[31:0], L50_0r1[31:0], L50_0a, L54_0r0[3:0], L54_0r1[3:0], L54_0a, L57_0r0[73:0], L57_0r1[73:0], L57_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 I14 (L56_0r, L56_0a, L23_0r, L23_0a, L25_0r, L25_0a, L27_0r, L27_0a, L30_0r, L30_0a, L32_0r, L32_0a, L35_0r, L35_0a, L37_0r, L37_0a, L39_0r, L39_0a, L42_0r, L42_0a, L44_0r, L44_0a, L46_0r, L46_0a, L48_0r, L48_0a, L51_0r, L51_0a, L53_0r, L53_0a, reset);
  tkvimmOrReg1_wo0w1_ro0w1 I15 (L59_0r0, L59_0r1, L59_0a, L56_0r, L56_0a, L48_0r, L48_0a, L49_0r0, L49_0r1, L49_0a, reset);
  tko0m1_1nm1b0 I16 (L64_0r, L64_0a, L66_0r0, L66_0r1, L66_0a, reset);
  tko0m1_1nm1b1 I17 (L68_0r, L68_0a, L70_0r0, L70_0r1, L70_0a, reset);
  tks1_o0w1_1o0w0_0o0w0 I18 (L63_0r0, L63_0r1, L63_0a, L64_0r, L64_0a, L68_0r, L68_0a, reset);
  tkm2x0b I19 (L67_0r, L67_0a, L71_0r, L71_0a, L72_0r, L72_0a, reset);
  tkf0mo0w0_o0w0 I20 (L73_0r, L73_0a, L61_0r, L61_0a, L62_0r, L62_0a, reset);
  tkj0m0_0 I21 (L58_0r, L58_0a, L72_0r, L72_0a, L74_0r, L74_0a, reset);
  tks6_o0w6_9c30mac30mbc30mdc30mec30mfc30m20m21m22m23m24m28m2cm30m31m32m33m34m35m36m37m38m3co0w0_0m1m2m3m4m5m6m7m8mcm10m11m12m13m14m15m16m17m18m1cm25m26m27o0w0 I22 (L17_0r0[5:0], L17_0r1[5:0], L17_0a, L21_0r, L21_0a, L73_0r, L73_0a, reset);
  tkm2x0b I23 (L22_0r, L22_0a, L74_0r, L74_0a, L75_0r, L75_0a, reset);
  tkf1mo0w0_o0w1 I24 (L66_0r0, L66_0r1, L66_0a, L76_0r, L76_0a, L77_0r0, L77_0r1, L77_0a, reset);
  tkf1mo0w0_o0w1 I25 (L70_0r0, L70_0r1, L70_0a, L78_0r, L78_0a, L79_0r0, L79_0r1, L79_0a, reset);
  tkm2x1b I26 (L77_0r0, L77_0r1, L77_0a, L79_0r0, L79_0r1, L79_0a, L80_0r0, L80_0r1, L80_0a, reset);
  tkf1mo0w0_o0w1 I27 (L80_0r0, L80_0r1, L80_0a, L81_0r, L81_0a, L82_0r0, L82_0r1, L82_0a, reset);
  tko0m2_1nm2b1 I28 (L76_0r, L76_0a, L83_0r0[1:0], L83_0r1[1:0], L83_0a, reset);
  tko0m2_1nm2b2 I29 (L78_0r, L78_0a, L84_0r0[1:0], L84_0r1[1:0], L84_0a, reset);
  tkm2x2b I30 (L83_0r0[1:0], L83_0r1[1:0], L83_0a, L84_0r0[1:0], L84_0r1[1:0], L84_0a, L85_0r0[1:0], L85_0r1[1:0], L85_0a, reset);
  tkj2m0_2 I31 (L81_0r, L81_0a, L85_0r0[1:0], L85_0r1[1:0], L85_0a, L86_0r0[1:0], L86_0r1[1:0], L86_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I32 (L86_0r0[1:0], L86_0r1[1:0], L86_0a, L67_0r, L67_0a, L71_0r, L71_0a, reset);
  tkj1m1_0 I33 (L82_0r0, L82_0r1, L82_0a, L61_0r, L61_0a, L59_0r0, L59_0r1, L59_0a, reset);
  tko0m1_1nm1b0 I34 (L92_0r, L92_0a, L94_0r0, L94_0r1, L94_0a, reset);
  tko0m1_1nm1b1 I35 (L96_0r, L96_0a, L98_0r0, L98_0r1, L98_0a, reset);
  tks3_o0w3_0c4m1m2m3c4o0w0_5m6o0w0 I36 (L91_0r0[2:0], L91_0r1[2:0], L91_0a, L92_0r, L92_0a, L96_0r, L96_0a, reset);
  tkm2x0b I37 (L95_0r, L95_0a, L99_0r, L99_0a, L135_0r, L135_0a, reset);
  tko0m4_1nm4b8 I38 (L103_0r, L103_0a, L104_0r0[3:0], L104_0r1[3:0], L104_0a, reset);
  tko0m1_1nm1b1 I39 (L105_0r, L105_0a, L106_0r0, L106_0r1, L106_0a, reset);
  tko1m1_1noti0w1b I40 (L109_0r0, L109_0r1, L109_0a, L107_0r0, L107_0r1, L107_0a, reset);
  tkj3m1_1_1 I41 (L106_0r0, L106_0r1, L106_0a, L107_0r0, L107_0r1, L107_0a, L111_0r0, L111_0r1, L111_0a, L112_0r0[2:0], L112_0r1[2:0], L112_0a, reset);
  tkj15m5_5_5 I42 (L114_0r0[4:0], L114_0r1[4:0], L114_0a, L116_0r0[4:0], L116_0r1[4:0], L116_0a, L118_0r0[4:0], L118_0r1[4:0], L118_0a, L119_0r0[14:0], L119_0r1[14:0], L119_0a, reset);
  tko1m1_1noti0w1b I43 (L122_0r0, L122_0r1, L122_0a, L120_0r0, L120_0r1, L120_0a, reset);
  tko13m32_1ap19xi12w1b_2api0w13bt1o0w19b I44 (L131_0r0[12:0], L131_0r1[12:0], L131_0a, L129_0r0[31:0], L129_0r1[31:0], L129_0a, reset);
  tkj74m3_4_3_15_1_5_6_1_32_4 I45 (L102_0r0[2:0], L102_0r1[2:0], L102_0a, L104_0r0[3:0], L104_0r1[3:0], L104_0a, L112_0r0[2:0], L112_0r1[2:0], L112_0a, L119_0r0[14:0], L119_0r1[14:0], L119_0a, L120_0r0, L120_0r1, L120_0a, L124_0r0[4:0], L124_0r1[4:0], L124_0a, L126_0r0[5:0], L126_0r1[5:0], L126_0a, L128_0r0, L128_0r1, L128_0a, L129_0r0[31:0], L129_0r1[31:0], L129_0a, L133_0r0[3:0], L133_0r1[3:0], L133_0a, L136_0r0[73:0], L136_0r1[73:0], L136_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 I46 (L135_0r, L135_0a, L101_0r, L101_0a, L103_0r, L103_0a, L105_0r, L105_0a, L108_0r, L108_0a, L110_0r, L110_0a, L113_0r, L113_0a, L115_0r, L115_0a, L117_0r, L117_0a, L121_0r, L121_0a, L123_0r, L123_0a, L125_0r, L125_0a, L127_0r, L127_0a, L130_0r, L130_0a, L132_0r, L132_0a, reset);
  tks3_o0w3_1c6m2c4m4o0w0_0o0w0 I47 (L88_0r0[2:0], L88_0r1[2:0], L88_0a, L90_0r, L90_0a, L138_0r, L138_0a, reset);
  tkm2x0b I48 (L137_0r, L137_0a, L139_0r, L139_0a, L140_0r, L140_0a, reset);
  tkf1mo0w0_o0w1 I49 (L98_0r0, L98_0r1, L98_0a, L143_0r, L143_0a, L144_0r0, L144_0r1, L144_0a, reset);
  tkf1mo0w0_o0w1 I50 (L94_0r0, L94_0r1, L94_0a, L145_0r, L145_0a, L146_0r0, L146_0r1, L146_0a, reset);
  tkm2x1b I51 (L144_0r0, L144_0r1, L144_0a, L146_0r0, L146_0r1, L146_0a, L141_0r0, L141_0r1, L141_0a, reset);
  tko0m2_1nm2b1 I52 (L143_0r, L143_0a, L147_0r0[1:0], L147_0r1[1:0], L147_0a, reset);
  tko0m2_1nm2b2 I53 (L145_0r, L145_0a, L148_0r0[1:0], L148_0r1[1:0], L148_0a, reset);
  tkm2x2b I54 (L147_0r0[1:0], L147_0r1[1:0], L147_0a, L148_0r0[1:0], L148_0r1[1:0], L148_0a, L149_0r0[1:0], L149_0r1[1:0], L149_0a, reset);
  tkj2m0_2 I55 (L142_0r, L142_0a, L149_0r0[1:0], L149_0r1[1:0], L149_0a, L150_0r0[1:0], L150_0r1[1:0], L150_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I56 (L150_0r0[1:0], L150_0r1[1:0], L150_0a, L99_0r, L99_0a, L95_0r, L95_0a, reset);
  tkvstore1_wo0w1_ro0w1o0w1 I57 (L141_0r0, L141_0r1, L141_0a, L142_0r, L142_0a, L121_0r, L121_0a, L110_0r, L110_0a, L122_0r0, L122_0r1, L122_0a, L111_0r0, L111_0r1, L111_0a, reset);
  tkvmemAccess4_wo0w4_ro0w4 I58 (L151_0r0[3:0], L151_0r1[3:0], L151_0a, L152_0r, L152_0a, L132_0r, L132_0a, L133_0r0[3:0], L133_0r1[3:0], L133_0a, reset);
  tkvinstKind3_wo0w3_ro0w3o0w3o0w3 I59 (L153_0r0[2:0], L153_0r1[2:0], L153_0a, L154_0r, L154_0a, L87_0r, L87_0a, L90_0r, L90_0a, L101_0r, L101_0a, L88_0r0[2:0], L88_0r1[2:0], L88_0a, L91_0r0[2:0], L91_0r1[2:0], L91_0a, L102_0r0[2:0], L102_0r1[2:0], L102_0a, reset);
  tkvimmOrReg1_wo0w1_ro0w1 I60 (L155_0r0, L155_0r1, L155_0a, L156_0r, L156_0a, L127_0r, L127_0a, L128_0r0, L128_0r1, L128_0a, reset);
  tkj0m0_0_0 I61 (L152_0r, L152_0a, L154_0r, L154_0a, L156_0r, L156_0a, L87_0r, L87_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I62 (L161_0r, L161_0a, L158_0r, L158_0a, L159_0r, L159_0a, L160_0r, L160_0a, reset);
  tko0m1_1nm1b0 I63 (L164_0r, L164_0a, L166_0r0, L166_0r1, L166_0a, reset);
  tko0m1_1nm1b1 I64 (L168_0r, L168_0a, L170_0r0, L170_0r1, L170_0a, reset);
  tks1_o0w1_1o0w0_0o0w0 I65 (L163_0r0, L163_0r1, L163_0a, L164_0r, L164_0a, L168_0r, L168_0a, reset);
  tkm2x0b I66 (L167_0r, L167_0a, L171_0r, L171_0a, L172_0r, L172_0a, reset);
  tko0m4_1nm4b7 I67 (L176_0r, L176_0a, L178_0r0[3:0], L178_0r1[3:0], L178_0a, reset);
  tko0m3_1nm3b0 I68 (L180_0r, L180_0a, L182_0r0[2:0], L182_0r1[2:0], L182_0a, reset);
  tkf0mo0w0_o0w0 I69 (L184_0r, L184_0a, L176_0r, L176_0a, L180_0r, L180_0a, reset);
  tkj0m0_0 I70 (L179_0r, L179_0a, L183_0r, L183_0a, L185_0r, L185_0a, reset);
  tko0m4_1nm4b7 I71 (L186_0r, L186_0a, L188_0r0[3:0], L188_0r1[3:0], L188_0a, reset);
  tko0m3_1nm3b3 I72 (L190_0r, L190_0a, L192_0r0[2:0], L192_0r1[2:0], L192_0a, reset);
  tkf0mo0w0_o0w0 I73 (L194_0r, L194_0a, L186_0r, L186_0a, L190_0r, L190_0a, reset);
  tkj0m0_0 I74 (L189_0r, L189_0a, L193_0r, L193_0a, L195_0r, L195_0a, reset);
  tko0m4_1nm4b3 I75 (L196_0r, L196_0a, L198_0r0[3:0], L198_0r1[3:0], L198_0a, reset);
  tko0m3_1nm3b3 I76 (L200_0r, L200_0a, L202_0r0[2:0], L202_0r1[2:0], L202_0a, reset);
  tkf0mo0w0_o0w0 I77 (L204_0r, L204_0a, L196_0r, L196_0a, L200_0r, L200_0a, reset);
  tkj0m0_0 I78 (L199_0r, L199_0a, L203_0r, L203_0a, L205_0r, L205_0a, reset);
  tko0m4_1nm4b5 I79 (L206_0r, L206_0a, L208_0r0[3:0], L208_0r1[3:0], L208_0a, reset);
  tko0m3_1nm3b3 I80 (L210_0r, L210_0a, L212_0r0[2:0], L212_0r1[2:0], L212_0a, reset);
  tkf0mo0w0_o0w0 I81 (L214_0r, L214_0a, L206_0r, L206_0a, L210_0r, L210_0a, reset);
  tkj0m0_0 I82 (L209_0r, L209_0a, L213_0r, L213_0a, L215_0r, L215_0a, reset);
  tko0m4_1nm4b7 I83 (L216_0r, L216_0a, L218_0r0[3:0], L218_0r1[3:0], L218_0a, reset);
  tko0m3_1nm3b4 I84 (L220_0r, L220_0a, L222_0r0[2:0], L222_0r1[2:0], L222_0a, reset);
  tkf0mo0w0_o0w0 I85 (L224_0r, L224_0a, L216_0r, L216_0a, L220_0r, L220_0a, reset);
  tkj0m0_0 I86 (L219_0r, L219_0a, L223_0r, L223_0a, L225_0r, L225_0a, reset);
  tko0m4_1nm4b6 I87 (L226_0r, L226_0a, L228_0r0[3:0], L228_0r1[3:0], L228_0a, reset);
  tko0m3_1nm3b5 I88 (L230_0r, L230_0a, L232_0r0[2:0], L232_0r1[2:0], L232_0a, reset);
  tkf0mo0w0_o0w0 I89 (L234_0r, L234_0a, L226_0r, L226_0a, L230_0r, L230_0a, reset);
  tkj0m0_0 I90 (L229_0r, L229_0a, L233_0r, L233_0a, L235_0r, L235_0a, reset);
  tko0m4_1nm4b2 I91 (L236_0r, L236_0a, L238_0r0[3:0], L238_0r1[3:0], L238_0a, reset);
  tko0m3_1nm3b5 I92 (L240_0r, L240_0a, L242_0r0[2:0], L242_0r1[2:0], L242_0a, reset);
  tkf0mo0w0_o0w0 I93 (L244_0r, L244_0a, L236_0r, L236_0a, L240_0r, L240_0a, reset);
  tkj0m0_0 I94 (L239_0r, L239_0a, L243_0r, L243_0a, L245_0r, L245_0a, reset);
  tko0m4_1nm4b4 I95 (L246_0r, L246_0a, L248_0r0[3:0], L248_0r1[3:0], L248_0a, reset);
  tko0m3_1nm3b5 I96 (L250_0r, L250_0a, L252_0r0[2:0], L252_0r1[2:0], L252_0a, reset);
  tkf0mo0w0_o0w0 I97 (L254_0r, L254_0a, L246_0r, L246_0a, L250_0r, L250_0a, reset);
  tkj0m0_0 I98 (L249_0r, L249_0a, L253_0r, L253_0a, L255_0r, L255_0a, reset);
  tko0m4_1nm4b6 I99 (L256_0r, L256_0a, L258_0r0[3:0], L258_0r1[3:0], L258_0a, reset);
  tko0m3_1nm3b5 I100 (L260_0r, L260_0a, L262_0r0[2:0], L262_0r1[2:0], L262_0a, reset);
  tkf0mo0w0_o0w0 I101 (L264_0r, L264_0a, L256_0r, L256_0a, L260_0r, L260_0a, reset);
  tkj0m0_0 I102 (L259_0r, L259_0a, L263_0r, L263_0a, L265_0r, L265_0a, reset);
  tko0m4_1nm4bb I103 (L266_0r, L266_0a, L268_0r0[3:0], L268_0r1[3:0], L268_0a, reset);
  tko0m3_1nm3b3 I104 (L270_0r, L270_0a, L272_0r0[2:0], L272_0r1[2:0], L272_0a, reset);
  tkf0mo0w0_o0w0 I105 (L274_0r, L274_0a, L266_0r, L266_0a, L270_0r, L270_0a, reset);
  tkj0m0_0 I106 (L269_0r, L269_0a, L273_0r, L273_0a, L275_0r, L275_0a, reset);
  tko0m4_1nm4bd I107 (L276_0r, L276_0a, L278_0r0[3:0], L278_0r1[3:0], L278_0a, reset);
  tko0m3_1nm3b3 I108 (L280_0r, L280_0a, L282_0r0[2:0], L282_0r1[2:0], L282_0a, reset);
  tkf0mo0w0_o0w0 I109 (L284_0r, L284_0a, L276_0r, L276_0a, L280_0r, L280_0a, reset);
  tkj0m0_0 I110 (L279_0r, L279_0a, L283_0r, L283_0a, L285_0r, L285_0a, reset);
  tks6_o0w6_8c30mbc30mcc30mdc30mec30mfc30m10c20m11c20m12c20m13c20m14c20m15c20m16c20m17c20m19c20m1ac20m20m21m22m23m24m25m26m27m29m2ao0w0_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0_9o0w0_ao0w0 I111 (L174_0r0[5:0], L174_0r1[5:0], L174_0a, L184_0r, L184_0a, L194_0r, L194_0a, L204_0r, L204_0a, L214_0r, L214_0a, L224_0r, L224_0a, L234_0r, L234_0a, L244_0r, L244_0a, L254_0r, L254_0a, L264_0r, L264_0a, L274_0r, L274_0a, L284_0r, L284_0a, reset);
  tkm11x0b I112 (L185_0r, L185_0a, L195_0r, L195_0a, L205_0r, L205_0a, L215_0r, L215_0a, L225_0r, L225_0a, L235_0r, L235_0a, L245_0r, L245_0a, L255_0r, L255_0a, L265_0r, L265_0a, L275_0r, L275_0a, L285_0r, L285_0a, L286_0r, L286_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I113 (L287_0r, L287_0a, L161_0r, L161_0a, L162_0r, L162_0a, L173_0r, L173_0a, reset);
  tkj0m0_0_0 I114 (L140_0r, L140_0a, L172_0r, L172_0a, L286_0r, L286_0a, L288_0r, L288_0a, reset);
  tkf1mo0w0_o0w1 I115 (L166_0r0, L166_0r1, L166_0a, L289_0r, L289_0a, L290_0r0, L290_0r1, L290_0a, reset);
  tkf1mo0w0_o0w1 I116 (L170_0r0, L170_0r1, L170_0a, L291_0r, L291_0a, L292_0r0, L292_0r1, L292_0a, reset);
  tkm2x1b I117 (L290_0r0, L290_0r1, L290_0a, L292_0r0, L292_0r1, L292_0a, L293_0r0, L293_0r1, L293_0a, reset);
  tkf1mo0w0_o0w1 I118 (L293_0r0, L293_0r1, L293_0a, L294_0r, L294_0a, L295_0r0, L295_0r1, L295_0a, reset);
  tko0m2_1nm2b1 I119 (L289_0r, L289_0a, L296_0r0[1:0], L296_0r1[1:0], L296_0a, reset);
  tko0m2_1nm2b2 I120 (L291_0r, L291_0a, L297_0r0[1:0], L297_0r1[1:0], L297_0a, reset);
  tkm2x2b I121 (L296_0r0[1:0], L296_0r1[1:0], L296_0a, L297_0r0[1:0], L297_0r1[1:0], L297_0a, L298_0r0[1:0], L298_0r1[1:0], L298_0a, reset);
  tkj2m0_2 I122 (L294_0r, L294_0a, L298_0r0[1:0], L298_0r1[1:0], L298_0a, L299_0r0[1:0], L299_0r1[1:0], L299_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I123 (L299_0r0[1:0], L299_0r1[1:0], L299_0a, L167_0r, L167_0a, L171_0r, L171_0a, reset);
  tkj1m1_0 I124 (L295_0r0, L295_0r1, L295_0a, L160_0r, L160_0a, L155_0r0, L155_0r1, L155_0a, reset);
  tkf3mo0w0_o0w3 I125 (L182_0r0[2:0], L182_0r1[2:0], L182_0a, L300_0r, L300_0a, L301_0r0[2:0], L301_0r1[2:0], L301_0a, reset);
  tkf3mo0w0_o0w3 I126 (L192_0r0[2:0], L192_0r1[2:0], L192_0a, L302_0r, L302_0a, L303_0r0[2:0], L303_0r1[2:0], L303_0a, reset);
  tkf3mo0w0_o0w3 I127 (L202_0r0[2:0], L202_0r1[2:0], L202_0a, L304_0r, L304_0a, L305_0r0[2:0], L305_0r1[2:0], L305_0a, reset);
  tkf3mo0w0_o0w3 I128 (L212_0r0[2:0], L212_0r1[2:0], L212_0a, L306_0r, L306_0a, L307_0r0[2:0], L307_0r1[2:0], L307_0a, reset);
  tkf3mo0w0_o0w3 I129 (L222_0r0[2:0], L222_0r1[2:0], L222_0a, L308_0r, L308_0a, L309_0r0[2:0], L309_0r1[2:0], L309_0a, reset);
  tkf3mo0w0_o0w3 I130 (L232_0r0[2:0], L232_0r1[2:0], L232_0a, L310_0r, L310_0a, L311_0r0[2:0], L311_0r1[2:0], L311_0a, reset);
  tkf3mo0w0_o0w3 I131 (L242_0r0[2:0], L242_0r1[2:0], L242_0a, L312_0r, L312_0a, L313_0r0[2:0], L313_0r1[2:0], L313_0a, reset);
  tkf3mo0w0_o0w3 I132 (L252_0r0[2:0], L252_0r1[2:0], L252_0a, L314_0r, L314_0a, L315_0r0[2:0], L315_0r1[2:0], L315_0a, reset);
  tkf3mo0w0_o0w3 I133 (L262_0r0[2:0], L262_0r1[2:0], L262_0a, L316_0r, L316_0a, L317_0r0[2:0], L317_0r1[2:0], L317_0a, reset);
  tkf3mo0w0_o0w3 I134 (L272_0r0[2:0], L272_0r1[2:0], L272_0a, L318_0r, L318_0a, L319_0r0[2:0], L319_0r1[2:0], L319_0a, reset);
  tkf3mo0w0_o0w3 I135 (L282_0r0[2:0], L282_0r1[2:0], L282_0a, L320_0r, L320_0a, L321_0r0[2:0], L321_0r1[2:0], L321_0a, reset);
  tkm11x3b I136 (L301_0r0[2:0], L301_0r1[2:0], L301_0a, L303_0r0[2:0], L303_0r1[2:0], L303_0a, L305_0r0[2:0], L305_0r1[2:0], L305_0a, L307_0r0[2:0], L307_0r1[2:0], L307_0a, L309_0r0[2:0], L309_0r1[2:0], L309_0a, L311_0r0[2:0], L311_0r1[2:0], L311_0a, L313_0r0[2:0], L313_0r1[2:0], L313_0a, L315_0r0[2:0], L315_0r1[2:0], L315_0a, L317_0r0[2:0], L317_0r1[2:0], L317_0a, L319_0r0[2:0], L319_0r1[2:0], L319_0a, L321_0r0[2:0], L321_0r1[2:0], L321_0a, L322_0r0[2:0], L322_0r1[2:0], L322_0a, reset);
  tkf3mo0w0_o0w3 I137 (L322_0r0[2:0], L322_0r1[2:0], L322_0a, L323_0r, L323_0a, L324_0r0[2:0], L324_0r1[2:0], L324_0a, reset);
  tko0m11_1nm11b1 I138 (L300_0r, L300_0a, L325_0r0[10:0], L325_0r1[10:0], L325_0a, reset);
  tko0m11_1nm11b2 I139 (L302_0r, L302_0a, L326_0r0[10:0], L326_0r1[10:0], L326_0a, reset);
  tko0m11_1nm11b4 I140 (L304_0r, L304_0a, L327_0r0[10:0], L327_0r1[10:0], L327_0a, reset);
  tko0m11_1nm11b8 I141 (L306_0r, L306_0a, L328_0r0[10:0], L328_0r1[10:0], L328_0a, reset);
  tko0m11_1nm11b10 I142 (L308_0r, L308_0a, L329_0r0[10:0], L329_0r1[10:0], L329_0a, reset);
  tko0m11_1nm11b20 I143 (L310_0r, L310_0a, L330_0r0[10:0], L330_0r1[10:0], L330_0a, reset);
  tko0m11_1nm11b40 I144 (L312_0r, L312_0a, L331_0r0[10:0], L331_0r1[10:0], L331_0a, reset);
  tko0m11_1nm11b80 I145 (L314_0r, L314_0a, L332_0r0[10:0], L332_0r1[10:0], L332_0a, reset);
  tko0m11_1nm11b100 I146 (L316_0r, L316_0a, L333_0r0[10:0], L333_0r1[10:0], L333_0a, reset);
  tko0m11_1nm11b200 I147 (L318_0r, L318_0a, L334_0r0[10:0], L334_0r1[10:0], L334_0a, reset);
  tko0m11_1nm11b400 I148 (L320_0r, L320_0a, L335_0r0[10:0], L335_0r1[10:0], L335_0a, reset);
  tkm11x11b I149 (L325_0r0[10:0], L325_0r1[10:0], L325_0a, L326_0r0[10:0], L326_0r1[10:0], L326_0a, L327_0r0[10:0], L327_0r1[10:0], L327_0a, L328_0r0[10:0], L328_0r1[10:0], L328_0a, L329_0r0[10:0], L329_0r1[10:0], L329_0a, L330_0r0[10:0], L330_0r1[10:0], L330_0a, L331_0r0[10:0], L331_0r1[10:0], L331_0a, L332_0r0[10:0], L332_0r1[10:0], L332_0a, L333_0r0[10:0], L333_0r1[10:0], L333_0a, L334_0r0[10:0], L334_0r1[10:0], L334_0a, L335_0r0[10:0], L335_0r1[10:0], L335_0a, L336_0r0[10:0], L336_0r1[10:0], L336_0a, reset);
  tkj11m0_11 I150 (L323_0r, L323_0a, L336_0r0[10:0], L336_0r1[10:0], L336_0a, L337_0r0[10:0], L337_0r1[10:0], L337_0a, reset);
  tks11_o0w11_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0_20o0w0_40o0w0_80o0w0_100o0w0_200o0w0_400o0w0 I151 (L337_0r0[10:0], L337_0r1[10:0], L337_0a, L183_0r, L183_0a, L193_0r, L193_0a, L203_0r, L203_0a, L213_0r, L213_0a, L223_0r, L223_0a, L233_0r, L233_0a, L243_0r, L243_0a, L253_0r, L253_0a, L263_0r, L263_0a, L273_0r, L273_0a, L283_0r, L283_0a, reset);
  tkj3m3_0 I152 (L324_0r0[2:0], L324_0r1[2:0], L324_0a, L159_0r, L159_0a, L153_0r0[2:0], L153_0r1[2:0], L153_0a, reset);
  tkf4mo0w0_o0w4 I153 (L178_0r0[3:0], L178_0r1[3:0], L178_0a, L338_0r, L338_0a, L339_0r0[3:0], L339_0r1[3:0], L339_0a, reset);
  tkf4mo0w0_o0w4 I154 (L188_0r0[3:0], L188_0r1[3:0], L188_0a, L340_0r, L340_0a, L341_0r0[3:0], L341_0r1[3:0], L341_0a, reset);
  tkf4mo0w0_o0w4 I155 (L198_0r0[3:0], L198_0r1[3:0], L198_0a, L342_0r, L342_0a, L343_0r0[3:0], L343_0r1[3:0], L343_0a, reset);
  tkf4mo0w0_o0w4 I156 (L208_0r0[3:0], L208_0r1[3:0], L208_0a, L344_0r, L344_0a, L345_0r0[3:0], L345_0r1[3:0], L345_0a, reset);
  tkf4mo0w0_o0w4 I157 (L218_0r0[3:0], L218_0r1[3:0], L218_0a, L346_0r, L346_0a, L347_0r0[3:0], L347_0r1[3:0], L347_0a, reset);
  tkf4mo0w0_o0w4 I158 (L228_0r0[3:0], L228_0r1[3:0], L228_0a, L348_0r, L348_0a, L349_0r0[3:0], L349_0r1[3:0], L349_0a, reset);
  tkf4mo0w0_o0w4 I159 (L238_0r0[3:0], L238_0r1[3:0], L238_0a, L350_0r, L350_0a, L351_0r0[3:0], L351_0r1[3:0], L351_0a, reset);
  tkf4mo0w0_o0w4 I160 (L248_0r0[3:0], L248_0r1[3:0], L248_0a, L352_0r, L352_0a, L353_0r0[3:0], L353_0r1[3:0], L353_0a, reset);
  tkf4mo0w0_o0w4 I161 (L258_0r0[3:0], L258_0r1[3:0], L258_0a, L354_0r, L354_0a, L355_0r0[3:0], L355_0r1[3:0], L355_0a, reset);
  tkf4mo0w0_o0w4 I162 (L268_0r0[3:0], L268_0r1[3:0], L268_0a, L356_0r, L356_0a, L357_0r0[3:0], L357_0r1[3:0], L357_0a, reset);
  tkf4mo0w0_o0w4 I163 (L278_0r0[3:0], L278_0r1[3:0], L278_0a, L358_0r, L358_0a, L359_0r0[3:0], L359_0r1[3:0], L359_0a, reset);
  tkm11x4b I164 (L339_0r0[3:0], L339_0r1[3:0], L339_0a, L341_0r0[3:0], L341_0r1[3:0], L341_0a, L343_0r0[3:0], L343_0r1[3:0], L343_0a, L345_0r0[3:0], L345_0r1[3:0], L345_0a, L347_0r0[3:0], L347_0r1[3:0], L347_0a, L349_0r0[3:0], L349_0r1[3:0], L349_0a, L351_0r0[3:0], L351_0r1[3:0], L351_0a, L353_0r0[3:0], L353_0r1[3:0], L353_0a, L355_0r0[3:0], L355_0r1[3:0], L355_0a, L357_0r0[3:0], L357_0r1[3:0], L357_0a, L359_0r0[3:0], L359_0r1[3:0], L359_0a, L360_0r0[3:0], L360_0r1[3:0], L360_0a, reset);
  tkf4mo0w0_o0w4 I165 (L360_0r0[3:0], L360_0r1[3:0], L360_0a, L361_0r, L361_0a, L362_0r0[3:0], L362_0r1[3:0], L362_0a, reset);
  tko0m11_1nm11b1 I166 (L338_0r, L338_0a, L363_0r0[10:0], L363_0r1[10:0], L363_0a, reset);
  tko0m11_1nm11b2 I167 (L340_0r, L340_0a, L364_0r0[10:0], L364_0r1[10:0], L364_0a, reset);
  tko0m11_1nm11b4 I168 (L342_0r, L342_0a, L365_0r0[10:0], L365_0r1[10:0], L365_0a, reset);
  tko0m11_1nm11b8 I169 (L344_0r, L344_0a, L366_0r0[10:0], L366_0r1[10:0], L366_0a, reset);
  tko0m11_1nm11b10 I170 (L346_0r, L346_0a, L367_0r0[10:0], L367_0r1[10:0], L367_0a, reset);
  tko0m11_1nm11b20 I171 (L348_0r, L348_0a, L368_0r0[10:0], L368_0r1[10:0], L368_0a, reset);
  tko0m11_1nm11b40 I172 (L350_0r, L350_0a, L369_0r0[10:0], L369_0r1[10:0], L369_0a, reset);
  tko0m11_1nm11b80 I173 (L352_0r, L352_0a, L370_0r0[10:0], L370_0r1[10:0], L370_0a, reset);
  tko0m11_1nm11b100 I174 (L354_0r, L354_0a, L371_0r0[10:0], L371_0r1[10:0], L371_0a, reset);
  tko0m11_1nm11b200 I175 (L356_0r, L356_0a, L372_0r0[10:0], L372_0r1[10:0], L372_0a, reset);
  tko0m11_1nm11b400 I176 (L358_0r, L358_0a, L373_0r0[10:0], L373_0r1[10:0], L373_0a, reset);
  tkm11x11b I177 (L363_0r0[10:0], L363_0r1[10:0], L363_0a, L364_0r0[10:0], L364_0r1[10:0], L364_0a, L365_0r0[10:0], L365_0r1[10:0], L365_0a, L366_0r0[10:0], L366_0r1[10:0], L366_0a, L367_0r0[10:0], L367_0r1[10:0], L367_0a, L368_0r0[10:0], L368_0r1[10:0], L368_0a, L369_0r0[10:0], L369_0r1[10:0], L369_0a, L370_0r0[10:0], L370_0r1[10:0], L370_0a, L371_0r0[10:0], L371_0r1[10:0], L371_0a, L372_0r0[10:0], L372_0r1[10:0], L372_0a, L373_0r0[10:0], L373_0r1[10:0], L373_0a, L374_0r0[10:0], L374_0r1[10:0], L374_0a, reset);
  tkj11m0_11 I178 (L361_0r, L361_0a, L374_0r0[10:0], L374_0r1[10:0], L374_0a, L375_0r0[10:0], L375_0r1[10:0], L375_0a, reset);
  tks11_o0w11_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0_20o0w0_40o0w0_80o0w0_100o0w0_200o0w0_400o0w0 I179 (L375_0r0[10:0], L375_0r1[10:0], L375_0a, L179_0r, L179_0a, L189_0r, L189_0a, L199_0r, L199_0a, L209_0r, L209_0a, L219_0r, L219_0a, L229_0r, L229_0a, L239_0r, L239_0a, L249_0r, L249_0a, L259_0r, L259_0a, L269_0r, L269_0a, L279_0r, L279_0a, reset);
  tkj4m4_0 I180 (L362_0r0[3:0], L362_0r1[3:0], L362_0a, L158_0r, L158_0a, L151_0r0[3:0], L151_0r1[3:0], L151_0a, reset);
  tko0m3_1nm3b1 I181 (L381_0r, L381_0a, L382_0r0[2:0], L382_0r1[2:0], L382_0a, reset);
  tko0m3_1nm3b0 I182 (L385_0r, L385_0a, L386_0r0[2:0], L386_0r1[2:0], L386_0a, reset);
  tko0m15_1nm15b0 I183 (L387_0r, L387_0a, L388_0r0[14:0], L388_0r1[14:0], L388_0a, reset);
  tko0m1_1nm1b0 I184 (L389_0r, L389_0a, L390_0r0, L390_0r1, L390_0a, reset);
  tko0m5_1nm5b0 I185 (L391_0r, L391_0a, L392_0r0[4:0], L392_0r1[4:0], L392_0a, reset);
  tko0m6_1nm6b0 I186 (L393_0r, L393_0a, L394_0r0[5:0], L394_0r1[5:0], L394_0a, reset);
  tko0m1_1nm1b0 I187 (L395_0r, L395_0a, L396_0r0, L396_0r1, L396_0a, reset);
  tko0m2_1nm2b0 I188 (L398_0r, L398_0a, L399_0r0[1:0], L399_0r1[1:0], L399_0a, reset);
  tkj24m2_22 I189 (L399_0r0[1:0], L399_0r1[1:0], L399_0a, L401_0r0[21:0], L401_0r1[21:0], L401_0a, L402_0r0[23:0], L402_0r1[23:0], L402_0a, reset);
  tko24m32_1ap8xi23w1b_2api0w24bt1o0w8b I190 (L402_0r0[23:0], L402_0r1[23:0], L402_0a, L397_0r0[31:0], L397_0r1[31:0], L397_0a, reset);
  tko0m4_1nm4b7 I191 (L403_0r, L403_0a, L404_0r0[3:0], L404_0r1[3:0], L404_0a, reset);
  tkj74m3_4_3_15_1_5_6_1_32_4 I192 (L382_0r0[2:0], L382_0r1[2:0], L382_0a, L384_0r0[3:0], L384_0r1[3:0], L384_0a, L386_0r0[2:0], L386_0r1[2:0], L386_0a, L388_0r0[14:0], L388_0r1[14:0], L388_0a, L390_0r0, L390_0r1, L390_0a, L392_0r0[4:0], L392_0r1[4:0], L392_0a, L394_0r0[5:0], L394_0r1[5:0], L394_0a, L396_0r0, L396_0r1, L396_0a, L397_0r0[31:0], L397_0r1[31:0], L397_0a, L404_0r0[3:0], L404_0r1[3:0], L404_0a, L407_0r0[73:0], L407_0r1[73:0], L407_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 I193 (L406_0r, L406_0a, L381_0r, L381_0a, L383_0r, L383_0a, L385_0r, L385_0a, L387_0r, L387_0a, L389_0r, L389_0a, L391_0r, L391_0a, L393_0r, L393_0a, L395_0r, L395_0a, L398_0r, L398_0a, L400_0r, L400_0a, L403_0r, L403_0a, reset);
  tko0m3_1nm3b2 I194 (L409_0r, L409_0a, L410_0r0[2:0], L410_0r1[2:0], L410_0a, reset);
  tko0m4_1nm4b8 I195 (L411_0r, L411_0a, L412_0r0[3:0], L412_0r1[3:0], L412_0a, reset);
  tko0m3_1nm3b1 I196 (L413_0r, L413_0a, L414_0r0[2:0], L414_0r1[2:0], L414_0a, reset);
  tko0m15_1nm15b0 I197 (L415_0r, L415_0a, L416_0r0[14:0], L416_0r1[14:0], L416_0a, reset);
  tko0m1_1nm1b1 I198 (L417_0r, L417_0a, L418_0r0, L418_0r1, L418_0a, reset);
  tko0m6_1nm6b0 I199 (L421_0r, L421_0a, L422_0r0[5:0], L422_0r1[5:0], L422_0a, reset);
  tko0m1_1nm1b0 I200 (L423_0r, L423_0a, L424_0r0, L424_0r1, L424_0a, reset);
  tko0m10_1nm10b0 I201 (L425_0r, L425_0a, L426_0r0[9:0], L426_0r1[9:0], L426_0a, reset);
  tkj32m10_22 I202 (L426_0r0[9:0], L426_0r1[9:0], L426_0a, L428_0r0[21:0], L428_0r1[21:0], L428_0a, L429_0r0[31:0], L429_0r1[31:0], L429_0a, reset);
  tko0m4_1nm4b7 I203 (L430_0r, L430_0a, L431_0r0[3:0], L431_0r1[3:0], L431_0a, reset);
  tkj74m3_4_3_15_1_5_6_1_32_4 I204 (L410_0r0[2:0], L410_0r1[2:0], L410_0a, L412_0r0[3:0], L412_0r1[3:0], L412_0a, L414_0r0[2:0], L414_0r1[2:0], L414_0a, L416_0r0[14:0], L416_0r1[14:0], L416_0a, L418_0r0, L418_0r1, L418_0a, L420_0r0[4:0], L420_0r1[4:0], L420_0a, L422_0r0[5:0], L422_0r1[5:0], L422_0a, L424_0r0, L424_0r1, L424_0a, L429_0r0[31:0], L429_0r1[31:0], L429_0a, L431_0r0[3:0], L431_0r1[3:0], L431_0a, L434_0r0[73:0], L434_0r1[73:0], L434_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 I205 (L433_0r, L433_0a, L409_0r, L409_0a, L411_0r, L411_0a, L413_0r, L413_0a, L415_0r, L415_0a, L417_0r, L417_0a, L419_0r, L419_0a, L421_0r, L421_0a, L423_0r, L423_0a, L425_0r, L425_0a, L427_0r, L427_0a, L430_0r, L430_0a, reset);
  tks3_o0w3_0m1c6m6o0w0_2o0w0_4o0w0 I206 (L377_0r0[2:0], L377_0r1[2:0], L377_0a, L379_0r, L379_0a, L406_0r, L406_0a, L433_0r, L433_0a, reset);
  tkm3x0b I207 (L380_0r, L380_0a, L408_0r, L408_0a, L435_0r, L435_0a, L436_0r, L436_0a, reset);
  tks2_o0w2_1o0w0_2o0w0_3o0w0_0o0w0 I208 (L12_0r0[1:0], L12_0r1[1:0], L12_0a, L14_0r, L14_0a, L16_0r, L16_0a, L287_0r, L287_0a, L376_0r, L376_0a, reset);
  tkm4x0b I209 (L15_0r, L15_0a, L75_0r, L75_0a, L288_0r, L288_0a, L436_0r, L436_0a, L437_0r, L437_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I210 (L438_0r, L438_0a, L6_0r, L6_0a, L7_0r, L7_0a, L11_0r, L11_0a, reset);
  tkj0m0_0_0 I211 (L6_0r, L6_0a, L10_0r, L10_0a, L437_0r, L437_0a, L439_0r, L439_0a, reset);
  tko0m74_1nm74b1c00000000000000040 I212 (L441_0r, L441_0a, L443_0r0[73:0], L443_0r1[73:0], L443_0a, reset);
  tkf0mo0w0_o0w0 I213 (L14_0r, L14_0a, L445_0r, L445_0a, L446_0r, L446_0a, reset);
  tkf0mo0w0_o0w0 I214 (L19_0r, L19_0a, L447_0r, L447_0a, L448_0r, L448_0a, reset);
  tkf0mo0w0_o0w0 I215 (L138_0r, L138_0a, L449_0r, L449_0a, L450_0r, L450_0a, reset);
  tkf0mo0w0_o0w0 I216 (L379_0r, L379_0a, L451_0r, L451_0a, L452_0r, L452_0a, reset);
  tkm4x0b I217 (L445_0r, L445_0a, L447_0r, L447_0a, L449_0r, L449_0a, L451_0r, L451_0a, L441_0r, L441_0a, reset);
  tko0m4_1nm4b1 I218 (L446_0r, L446_0a, L453_0r0[3:0], L453_0r1[3:0], L453_0a, reset);
  tko0m4_1nm4b2 I219 (L448_0r, L448_0a, L454_0r0[3:0], L454_0r1[3:0], L454_0a, reset);
  tko0m4_1nm4b4 I220 (L450_0r, L450_0a, L455_0r0[3:0], L455_0r1[3:0], L455_0a, reset);
  tko0m4_1nm4b8 I221 (L452_0r, L452_0a, L456_0r0[3:0], L456_0r1[3:0], L456_0a, reset);
  tkm4x4b I222 (L453_0r0[3:0], L453_0r1[3:0], L453_0a, L454_0r0[3:0], L454_0r1[3:0], L454_0a, L455_0r0[3:0], L455_0r1[3:0], L455_0a, L456_0r0[3:0], L456_0r1[3:0], L456_0a, L457_0r0[3:0], L457_0r1[3:0], L457_0a, reset);
  tkj4m0_4 I223 (L444_0r, L444_0a, L457_0r0[3:0], L457_0r1[3:0], L457_0a, L458_0r0[3:0], L458_0r1[3:0], L458_0a, reset);
  tks4_o0w4_1o0w0_2o0w0_4o0w0_8o0w0 I224 (L458_0r0[3:0], L458_0r1[3:0], L458_0a, L15_0r, L15_0a, L20_0r, L20_0a, L139_0r, L139_0a, L380_0r, L380_0a, reset);
  tkvir65_wo0w65_ro0w22o25w5o0w22o25w4o22w3o19w6o13w1o0w13o19w6o25w5o25w5o0w5o14w5o13w1o13w1o0w13o19w6o25w5o0w5o14w5o13w1o19w6o30w2o32w33 I225 (L4_0r0[64:0], L4_0r1[64:0], L4_0a, L438_0r, L438_0a, L427_0r, L427_0a, L419_0r, L419_0a, L400_0r, L400_0a, L383_0r, L383_0a, L376_0r, L376_0a, L173_0r, L173_0a, L162_0r, L162_0a, L130_0r, L130_0a, L125_0r, L125_0a, L123_0r, L123_0a, L117_0r, L117_0a, L115_0r, L115_0a, L113_0r, L113_0a, L108_0r, L108_0a, L62_0r, L62_0a, L51_0r, L51_0a, L46_0r, L46_0a, L44_0r, L44_0a, L37_0r, L37_0a, L35_0r, L35_0a, L30_0r, L30_0a, L16_0r, L16_0a, L11_0r, L11_0a, L7_0r, L7_0a, L428_0r0[21:0], L428_0r1[21:0], L428_0a, L420_0r0[4:0], L420_0r1[4:0], L420_0a, L401_0r0[21:0], L401_0r1[21:0], L401_0a, L384_0r0[3:0], L384_0r1[3:0], L384_0a, L377_0r0[2:0], L377_0r1[2:0], L377_0a, L174_0r0[5:0], L174_0r1[5:0], L174_0a, L163_0r0, L163_0r1, L163_0a, L131_0r0[12:0], L131_0r1[12:0], L131_0a, L126_0r0[5:0], L126_0r1[5:0], L126_0a, L124_0r0[4:0], L124_0r1[4:0], L124_0a, L118_0r0[4:0], L118_0r1[4:0], L118_0a, L116_0r0[4:0], L116_0r1[4:0], L116_0a, L114_0r0[4:0], L114_0r1[4:0], L114_0a, L109_0r0, L109_0r1, L109_0a, L63_0r0, L63_0r1, L63_0a, L52_0r0[12:0], L52_0r1[12:0], L52_0a, L47_0r0[5:0], L47_0r1[5:0], L47_0a, L45_0r0[4:0], L45_0r1[4:0], L45_0a, L38_0r0[4:0], L38_0r1[4:0], L38_0a, L36_0r0[4:0], L36_0r1[4:0], L36_0a, L31_0r0, L31_0r1, L31_0a, L17_0r0[5:0], L17_0r1[5:0], L17_0a, L12_0r0[1:0], L12_0r1[1:0], L12_0a, L9_0r0[32:0], L9_0r1[32:0], L9_0a, reset);
  tkj65m65_0 I226 (inst_0r0[64:0], inst_0r1[64:0], inst_0a, L3_0r, L3_0a, L4_0r0[64:0], L4_0r1[64:0], L4_0a, reset);
  tkf74mo0w0_o0w74 I227 (L57_0r0[73:0], L57_0r1[73:0], L57_0a, L460_0r, L460_0a, L461_0r0[73:0], L461_0r1[73:0], L461_0a, reset);
  tkf74mo0w0_o0w74 I228 (L136_0r0[73:0], L136_0r1[73:0], L136_0a, L462_0r, L462_0a, L463_0r0[73:0], L463_0r1[73:0], L463_0a, reset);
  tkf74mo0w0_o0w74 I229 (L407_0r0[73:0], L407_0r1[73:0], L407_0a, L464_0r, L464_0a, L465_0r0[73:0], L465_0r1[73:0], L465_0a, reset);
  tkf74mo0w0_o0w74 I230 (L434_0r0[73:0], L434_0r1[73:0], L434_0a, L466_0r, L466_0a, L467_0r0[73:0], L467_0r1[73:0], L467_0a, reset);
  tkf74mo0w0_o0w74 I231 (L443_0r0[73:0], L443_0r1[73:0], L443_0a, L468_0r, L468_0a, L469_0r0[73:0], L469_0r1[73:0], L469_0a, reset);
  tkm5x74b I232 (L461_0r0[73:0], L461_0r1[73:0], L461_0a, L463_0r0[73:0], L463_0r1[73:0], L463_0a, L465_0r0[73:0], L465_0r1[73:0], L465_0a, L467_0r0[73:0], L467_0r1[73:0], L467_0a, L469_0r0[73:0], L469_0r1[73:0], L469_0a, L470_0r0[73:0], L470_0r1[73:0], L470_0a, reset);
  tkf74mo0w0_o0w74 I233 (L470_0r0[73:0], L470_0r1[73:0], L470_0a, L471_0r, L471_0a, decoded_0r0[73:0], decoded_0r1[73:0], decoded_0a, reset);
  tko0m5_1nm5b1 I234 (L460_0r, L460_0a, L473_0r0[4:0], L473_0r1[4:0], L473_0a, reset);
  tko0m5_1nm5b2 I235 (L462_0r, L462_0a, L474_0r0[4:0], L474_0r1[4:0], L474_0a, reset);
  tko0m5_1nm5b4 I236 (L464_0r, L464_0a, L475_0r0[4:0], L475_0r1[4:0], L475_0a, reset);
  tko0m5_1nm5b8 I237 (L466_0r, L466_0a, L476_0r0[4:0], L476_0r1[4:0], L476_0a, reset);
  tko0m5_1nm5b10 I238 (L468_0r, L468_0a, L477_0r0[4:0], L477_0r1[4:0], L477_0a, reset);
  tkm5x5b I239 (L473_0r0[4:0], L473_0r1[4:0], L473_0a, L474_0r0[4:0], L474_0r1[4:0], L474_0a, L475_0r0[4:0], L475_0r1[4:0], L475_0a, L476_0r0[4:0], L476_0r1[4:0], L476_0a, L477_0r0[4:0], L477_0r1[4:0], L477_0a, L478_0r0[4:0], L478_0r1[4:0], L478_0a, reset);
  tkj5m0_5 I240 (L471_0r, L471_0a, L478_0r0[4:0], L478_0r1[4:0], L478_0a, L479_0r0[4:0], L479_0r1[4:0], L479_0a, reset);
  tks5_o0w5_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0 I241 (L479_0r0[4:0], L479_0r1[4:0], L479_0a, L58_0r, L58_0a, L137_0r, L137_0a, L408_0r, L408_0a, L435_0r, L435_0a, L444_0r, L444_0a, reset);
  tkf33mo0w0_o0w33 I242 (L9_0r0[32:0], L9_0r1[32:0], L9_0a, L10_0r, L10_0a, pc_0r0[32:0], pc_0r1[32:0], pc_0a, reset);
  tki I243 (L439_0r, L439_0a, L3_0r, L3_0a, reset);
endmodule

module teak_Shifter (shift_0r0, shift_0r1, shift_0a, distanceI_0r0, distanceI_0r1, distanceI_0a, result_0r0, result_0r1, result_0a, arg_0r0, arg_0r1, arg_0a, reset);
  input [1:0] shift_0r0;
  input [1:0] shift_0r1;
  output shift_0a;
  input [4:0] distanceI_0r0;
  input [4:0] distanceI_0r1;
  output distanceI_0a;
  output [31:0] result_0r0;
  output [31:0] result_0r1;
  input result_0a;
  input [31:0] arg_0r0;
  input [31:0] arg_0r1;
  output arg_0a;
  input reset;
  wire L1_0r;
  wire L1_0a;
  wire L2_0r0;
  wire L2_0r1;
  wire L2_0a;
  wire L3_0r;
  wire L3_0a;
  wire [31:0] L5_0r0;
  wire [31:0] L5_0r1;
  wire L5_0a;
  wire L6_0r;
  wire L6_0a;
  wire L7_0r;
  wire L7_0a;
  wire [1:0] L8_0r0;
  wire [1:0] L8_0r1;
  wire L8_0a;
  wire L9_0r;
  wire L9_0a;
  wire L10_0r0;
  wire L10_0r1;
  wire L10_0a;
  wire L11_0r;
  wire L11_0a;
  wire [30:0] L12_0r0;
  wire [30:0] L12_0r1;
  wire L12_0a;
  wire L14_0r;
  wire L14_0a;
  wire [31:0] L15_0r0;
  wire [31:0] L15_0r1;
  wire L15_0a;
  wire L16_0r;
  wire L16_0a;
  wire L17_0r;
  wire L17_0a;
  wire [30:0] L18_0r0;
  wire [30:0] L18_0r1;
  wire L18_0a;
  wire L19_0r;
  wire L19_0a;
  wire L20_0r0;
  wire L20_0r1;
  wire L20_0a;
  wire L22_0r;
  wire L22_0a;
  wire [31:0] L23_0r0;
  wire [31:0] L23_0r1;
  wire L23_0a;
  wire L24_0r;
  wire L24_0a;
  wire L25_0r;
  wire L25_0a;
  wire [30:0] L26_0r0;
  wire [30:0] L26_0r1;
  wire L26_0a;
  wire L27_0r;
  wire L27_0a;
  wire L28_0r0;
  wire L28_0r1;
  wire L28_0a;
  wire L30_0r;
  wire L30_0a;
  wire [31:0] L31_0r0;
  wire [31:0] L31_0r1;
  wire L31_0a;
  wire L32_0r;
  wire L32_0a;
  wire L33_0r;
  wire L33_0a;
  wire L34_0r;
  wire L34_0a;
  wire [31:0] L35_0r0;
  wire [31:0] L35_0r1;
  wire L35_0a;
  wire L37_0r;
  wire L37_0a;
  wire L38_0r;
  wire L38_0a;
  wire L39_0r0;
  wire L39_0r1;
  wire L39_0a;
  wire L40_0r;
  wire L40_0a;
  wire [31:0] L42_0r0;
  wire [31:0] L42_0r1;
  wire L42_0a;
  wire L43_0r;
  wire L43_0a;
  wire L44_0r;
  wire L44_0a;
  wire [1:0] L45_0r0;
  wire [1:0] L45_0r1;
  wire L45_0a;
  wire L46_0r;
  wire L46_0a;
  wire [1:0] L47_0r0;
  wire [1:0] L47_0r1;
  wire L47_0a;
  wire L48_0r;
  wire L48_0a;
  wire [29:0] L49_0r0;
  wire [29:0] L49_0r1;
  wire L49_0a;
  wire L51_0r;
  wire L51_0a;
  wire [31:0] L52_0r0;
  wire [31:0] L52_0r1;
  wire L52_0a;
  wire L53_0r;
  wire L53_0a;
  wire L54_0r;
  wire L54_0a;
  wire [29:0] L55_0r0;
  wire [29:0] L55_0r1;
  wire L55_0a;
  wire L56_0r;
  wire L56_0a;
  wire [1:0] L57_0r0;
  wire [1:0] L57_0r1;
  wire L57_0a;
  wire L59_0r;
  wire L59_0a;
  wire [31:0] L60_0r0;
  wire [31:0] L60_0r1;
  wire L60_0a;
  wire L61_0r;
  wire L61_0a;
  wire L62_0r;
  wire L62_0a;
  wire [29:0] L63_0r0;
  wire [29:0] L63_0r1;
  wire L63_0a;
  wire L64_0r;
  wire L64_0a;
  wire [1:0] L65_0r0;
  wire [1:0] L65_0r1;
  wire L65_0a;
  wire L67_0r;
  wire L67_0a;
  wire [31:0] L68_0r0;
  wire [31:0] L68_0r1;
  wire L68_0a;
  wire L69_0r;
  wire L69_0a;
  wire L70_0r;
  wire L70_0a;
  wire L71_0r;
  wire L71_0a;
  wire [31:0] L72_0r0;
  wire [31:0] L72_0r1;
  wire L72_0a;
  wire L74_0r;
  wire L74_0a;
  wire L75_0r;
  wire L75_0a;
  wire L76_0r;
  wire L76_0a;
  wire L77_0r;
  wire L77_0a;
  wire [31:0] L78_0r0;
  wire [31:0] L78_0r1;
  wire L78_0a;
  wire L79_0r;
  wire L79_0a;
  wire [31:0] L80_0r0;
  wire [31:0] L80_0r1;
  wire L80_0a;
  wire L81_0r;
  wire L81_0a;
  wire [31:0] L82_0r0;
  wire [31:0] L82_0r1;
  wire L82_0a;
  wire L83_0r;
  wire L83_0a;
  wire [31:0] L84_0r0;
  wire [31:0] L84_0r1;
  wire L84_0a;
  wire [31:0] L85_0r0;
  wire [31:0] L85_0r1;
  wire L85_0a;
  wire L86_0r;
  wire L86_0a;
  wire [31:0] L87_0r0;
  wire [31:0] L87_0r1;
  wire L87_0a;
  wire [3:0] L88_0r0;
  wire [3:0] L88_0r1;
  wire L88_0a;
  wire [3:0] L89_0r0;
  wire [3:0] L89_0r1;
  wire L89_0a;
  wire [3:0] L90_0r0;
  wire [3:0] L90_0r1;
  wire L90_0a;
  wire [3:0] L91_0r0;
  wire [3:0] L91_0r1;
  wire L91_0a;
  wire [3:0] L92_0r0;
  wire [3:0] L92_0r1;
  wire L92_0a;
  wire [3:0] L93_0r0;
  wire [3:0] L93_0r1;
  wire L93_0a;
  wire L94_0r;
  wire L94_0a;
  wire L95_0r0;
  wire L95_0r1;
  wire L95_0a;
  wire L96_0r;
  wire L96_0a;
  wire [31:0] L98_0r0;
  wire [31:0] L98_0r1;
  wire L98_0a;
  wire L99_0r;
  wire L99_0a;
  wire L100_0r;
  wire L100_0a;
  wire [1:0] L101_0r0;
  wire [1:0] L101_0r1;
  wire L101_0a;
  wire L102_0r;
  wire L102_0a;
  wire [3:0] L103_0r0;
  wire [3:0] L103_0r1;
  wire L103_0a;
  wire L104_0r;
  wire L104_0a;
  wire [27:0] L105_0r0;
  wire [27:0] L105_0r1;
  wire L105_0a;
  wire L107_0r;
  wire L107_0a;
  wire [31:0] L108_0r0;
  wire [31:0] L108_0r1;
  wire L108_0a;
  wire L109_0r;
  wire L109_0a;
  wire L110_0r;
  wire L110_0a;
  wire [27:0] L111_0r0;
  wire [27:0] L111_0r1;
  wire L111_0a;
  wire L112_0r;
  wire L112_0a;
  wire [3:0] L113_0r0;
  wire [3:0] L113_0r1;
  wire L113_0a;
  wire L115_0r;
  wire L115_0a;
  wire [31:0] L116_0r0;
  wire [31:0] L116_0r1;
  wire L116_0a;
  wire L117_0r;
  wire L117_0a;
  wire L118_0r;
  wire L118_0a;
  wire [27:0] L119_0r0;
  wire [27:0] L119_0r1;
  wire L119_0a;
  wire L120_0r;
  wire L120_0a;
  wire [3:0] L121_0r0;
  wire [3:0] L121_0r1;
  wire L121_0a;
  wire L123_0r;
  wire L123_0a;
  wire [31:0] L124_0r0;
  wire [31:0] L124_0r1;
  wire L124_0a;
  wire L125_0r;
  wire L125_0a;
  wire L126_0r;
  wire L126_0a;
  wire L127_0r;
  wire L127_0a;
  wire [31:0] L128_0r0;
  wire [31:0] L128_0r1;
  wire L128_0a;
  wire L130_0r;
  wire L130_0a;
  wire L131_0r;
  wire L131_0a;
  wire L132_0r;
  wire L132_0a;
  wire L133_0r;
  wire L133_0a;
  wire [31:0] L134_0r0;
  wire [31:0] L134_0r1;
  wire L134_0a;
  wire L135_0r;
  wire L135_0a;
  wire [31:0] L136_0r0;
  wire [31:0] L136_0r1;
  wire L136_0a;
  wire L137_0r;
  wire L137_0a;
  wire [31:0] L138_0r0;
  wire [31:0] L138_0r1;
  wire L138_0a;
  wire L139_0r;
  wire L139_0a;
  wire [31:0] L140_0r0;
  wire [31:0] L140_0r1;
  wire L140_0a;
  wire [31:0] L141_0r0;
  wire [31:0] L141_0r1;
  wire L141_0a;
  wire L142_0r;
  wire L142_0a;
  wire [31:0] L143_0r0;
  wire [31:0] L143_0r1;
  wire L143_0a;
  wire [3:0] L144_0r0;
  wire [3:0] L144_0r1;
  wire L144_0a;
  wire [3:0] L145_0r0;
  wire [3:0] L145_0r1;
  wire L145_0a;
  wire [3:0] L146_0r0;
  wire [3:0] L146_0r1;
  wire L146_0a;
  wire [3:0] L147_0r0;
  wire [3:0] L147_0r1;
  wire L147_0a;
  wire [3:0] L148_0r0;
  wire [3:0] L148_0r1;
  wire L148_0a;
  wire [3:0] L149_0r0;
  wire [3:0] L149_0r1;
  wire L149_0a;
  wire L150_0r;
  wire L150_0a;
  wire L151_0r0;
  wire L151_0r1;
  wire L151_0a;
  wire L152_0r;
  wire L152_0a;
  wire [31:0] L154_0r0;
  wire [31:0] L154_0r1;
  wire L154_0a;
  wire L155_0r;
  wire L155_0a;
  wire L156_0r;
  wire L156_0a;
  wire [1:0] L157_0r0;
  wire [1:0] L157_0r1;
  wire L157_0a;
  wire L158_0r;
  wire L158_0a;
  wire [7:0] L159_0r0;
  wire [7:0] L159_0r1;
  wire L159_0a;
  wire L160_0r;
  wire L160_0a;
  wire [23:0] L161_0r0;
  wire [23:0] L161_0r1;
  wire L161_0a;
  wire L163_0r;
  wire L163_0a;
  wire [31:0] L164_0r0;
  wire [31:0] L164_0r1;
  wire L164_0a;
  wire L165_0r;
  wire L165_0a;
  wire L166_0r;
  wire L166_0a;
  wire [23:0] L167_0r0;
  wire [23:0] L167_0r1;
  wire L167_0a;
  wire L168_0r;
  wire L168_0a;
  wire [7:0] L169_0r0;
  wire [7:0] L169_0r1;
  wire L169_0a;
  wire L171_0r;
  wire L171_0a;
  wire [31:0] L172_0r0;
  wire [31:0] L172_0r1;
  wire L172_0a;
  wire L173_0r;
  wire L173_0a;
  wire L174_0r;
  wire L174_0a;
  wire [23:0] L175_0r0;
  wire [23:0] L175_0r1;
  wire L175_0a;
  wire L176_0r;
  wire L176_0a;
  wire [7:0] L177_0r0;
  wire [7:0] L177_0r1;
  wire L177_0a;
  wire L179_0r;
  wire L179_0a;
  wire [31:0] L180_0r0;
  wire [31:0] L180_0r1;
  wire L180_0a;
  wire L181_0r;
  wire L181_0a;
  wire L182_0r;
  wire L182_0a;
  wire L183_0r;
  wire L183_0a;
  wire [31:0] L184_0r0;
  wire [31:0] L184_0r1;
  wire L184_0a;
  wire L186_0r;
  wire L186_0a;
  wire L187_0r;
  wire L187_0a;
  wire L188_0r;
  wire L188_0a;
  wire L189_0r;
  wire L189_0a;
  wire [31:0] L190_0r0;
  wire [31:0] L190_0r1;
  wire L190_0a;
  wire L191_0r;
  wire L191_0a;
  wire [31:0] L192_0r0;
  wire [31:0] L192_0r1;
  wire L192_0a;
  wire L193_0r;
  wire L193_0a;
  wire [31:0] L194_0r0;
  wire [31:0] L194_0r1;
  wire L194_0a;
  wire L195_0r;
  wire L195_0a;
  wire [31:0] L196_0r0;
  wire [31:0] L196_0r1;
  wire L196_0a;
  wire [31:0] L197_0r0;
  wire [31:0] L197_0r1;
  wire L197_0a;
  wire L198_0r;
  wire L198_0a;
  wire [31:0] L199_0r0;
  wire [31:0] L199_0r1;
  wire L199_0a;
  wire [3:0] L200_0r0;
  wire [3:0] L200_0r1;
  wire L200_0a;
  wire [3:0] L201_0r0;
  wire [3:0] L201_0r1;
  wire L201_0a;
  wire [3:0] L202_0r0;
  wire [3:0] L202_0r1;
  wire L202_0a;
  wire [3:0] L203_0r0;
  wire [3:0] L203_0r1;
  wire L203_0a;
  wire [3:0] L204_0r0;
  wire [3:0] L204_0r1;
  wire L204_0a;
  wire [3:0] L205_0r0;
  wire [3:0] L205_0r1;
  wire L205_0a;
  wire L206_0r;
  wire L206_0a;
  wire L207_0r0;
  wire L207_0r1;
  wire L207_0a;
  wire L208_0r;
  wire L208_0a;
  wire [31:0] L210_0r0;
  wire [31:0] L210_0r1;
  wire L210_0a;
  wire L211_0r;
  wire L211_0a;
  wire L212_0r;
  wire L212_0a;
  wire [1:0] L213_0r0;
  wire [1:0] L213_0r1;
  wire L213_0a;
  wire L214_0r;
  wire L214_0a;
  wire [15:0] L215_0r0;
  wire [15:0] L215_0r1;
  wire L215_0a;
  wire L216_0r;
  wire L216_0a;
  wire [15:0] L217_0r0;
  wire [15:0] L217_0r1;
  wire L217_0a;
  wire L219_0r;
  wire L219_0a;
  wire [31:0] L220_0r0;
  wire [31:0] L220_0r1;
  wire L220_0a;
  wire L221_0r;
  wire L221_0a;
  wire L222_0r;
  wire L222_0a;
  wire [15:0] L223_0r0;
  wire [15:0] L223_0r1;
  wire L223_0a;
  wire L224_0r;
  wire L224_0a;
  wire [15:0] L225_0r0;
  wire [15:0] L225_0r1;
  wire L225_0a;
  wire L227_0r;
  wire L227_0a;
  wire [31:0] L228_0r0;
  wire [31:0] L228_0r1;
  wire L228_0a;
  wire L229_0r;
  wire L229_0a;
  wire L230_0r;
  wire L230_0a;
  wire [15:0] L231_0r0;
  wire [15:0] L231_0r1;
  wire L231_0a;
  wire L232_0r;
  wire L232_0a;
  wire [15:0] L233_0r0;
  wire [15:0] L233_0r1;
  wire L233_0a;
  wire L235_0r;
  wire L235_0a;
  wire [31:0] L236_0r0;
  wire [31:0] L236_0r1;
  wire L236_0a;
  wire L237_0r;
  wire L237_0a;
  wire L238_0r;
  wire L238_0a;
  wire L239_0r;
  wire L239_0a;
  wire [31:0] L240_0r0;
  wire [31:0] L240_0r1;
  wire L240_0a;
  wire L242_0r;
  wire L242_0a;
  wire L243_0r;
  wire L243_0a;
  wire L244_0r;
  wire L244_0a;
  wire L245_0r;
  wire L245_0a;
  wire [31:0] L246_0r0;
  wire [31:0] L246_0r1;
  wire L246_0a;
  wire L247_0r;
  wire L247_0a;
  wire [31:0] L248_0r0;
  wire [31:0] L248_0r1;
  wire L248_0a;
  wire L249_0r;
  wire L249_0a;
  wire [31:0] L250_0r0;
  wire [31:0] L250_0r1;
  wire L250_0a;
  wire L251_0r;
  wire L251_0a;
  wire [31:0] L252_0r0;
  wire [31:0] L252_0r1;
  wire L252_0a;
  wire [31:0] L253_0r0;
  wire [31:0] L253_0r1;
  wire L253_0a;
  wire L254_0r;
  wire L254_0a;
  wire [31:0] L255_0r0;
  wire [31:0] L255_0r1;
  wire L255_0a;
  wire [3:0] L256_0r0;
  wire [3:0] L256_0r1;
  wire L256_0a;
  wire [3:0] L257_0r0;
  wire [3:0] L257_0r1;
  wire L257_0a;
  wire [3:0] L258_0r0;
  wire [3:0] L258_0r1;
  wire L258_0a;
  wire [3:0] L259_0r0;
  wire [3:0] L259_0r1;
  wire L259_0a;
  wire [3:0] L260_0r0;
  wire [3:0] L260_0r1;
  wire L260_0a;
  wire [3:0] L261_0r0;
  wire [3:0] L261_0r1;
  wire L261_0a;
  wire [4:0] L262_0r0;
  wire [4:0] L262_0r1;
  wire L262_0a;
  wire L263_0r;
  wire L263_0a;
  wire [1:0] L264_0r0;
  wire [1:0] L264_0r1;
  wire L264_0a;
  wire L265_0r;
  wire L265_0a;
  wire L267_0r;
  wire L267_0a;
  wire L268_0r;
  wire L268_0a;
  wire L269_0r;
  wire L269_0a;
  wire L273_0r;
  wire L273_0a;
  wire [31:0] L274_0r0;
  wire [31:0] L274_0r1;
  wire L274_0a;
  wire L275_0r;
  wire L275_0a;
  wire [31:0] L276_0r0;
  wire [31:0] L276_0r1;
  wire L276_0a;
  wire L277_0r;
  wire L277_0a;
  wire [31:0] L278_0r0;
  wire [31:0] L278_0r1;
  wire L278_0a;
  wire L279_0r;
  wire L279_0a;
  wire [31:0] L280_0r0;
  wire [31:0] L280_0r1;
  wire L280_0a;
  wire [31:0] L281_0r0;
  wire [31:0] L281_0r1;
  wire L281_0a;
  wire L282_0r;
  wire L282_0a;
  wire [3:0] L284_0r0;
  wire [3:0] L284_0r1;
  wire L284_0a;
  wire [3:0] L285_0r0;
  wire [3:0] L285_0r1;
  wire L285_0a;
  wire [3:0] L286_0r0;
  wire [3:0] L286_0r1;
  wire L286_0a;
  wire [3:0] L287_0r0;
  wire [3:0] L287_0r1;
  wire L287_0a;
  wire [3:0] L288_0r0;
  wire [3:0] L288_0r1;
  wire L288_0a;
  wire [3:0] L289_0r0;
  wire [3:0] L289_0r1;
  wire L289_0a;
  tko0m1_1nm1b0 I0 (L9_0r, L9_0a, L10_0r0, L10_0r1, L10_0a, reset);
  tkj32m1_31 I1 (L10_0r0, L10_0r1, L10_0a, L12_0r0[30:0], L12_0r1[30:0], L12_0a, L15_0r0[31:0], L15_0r1[31:0], L15_0a, reset);
  tkf0mo0w0_o0w0 I2 (L14_0r, L14_0a, L9_0r, L9_0a, L11_0r, L11_0a, reset);
  tko0m1_1nm1b0 I3 (L19_0r, L19_0a, L20_0r0, L20_0r1, L20_0a, reset);
  tkj32m31_1 I4 (L18_0r0[30:0], L18_0r1[30:0], L18_0a, L20_0r0, L20_0r1, L20_0a, L23_0r0[31:0], L23_0r1[31:0], L23_0a, reset);
  tkf0mo0w0_o0w0 I5 (L22_0r, L22_0a, L17_0r, L17_0a, L19_0r, L19_0a, reset);
  tko0m1_1nm1b1 I6 (L27_0r, L27_0a, L28_0r0, L28_0r1, L28_0a, reset);
  tkj32m31_1 I7 (L26_0r0[30:0], L26_0r1[30:0], L26_0a, L28_0r0, L28_0r1, L28_0a, L31_0r0[31:0], L31_0r1[31:0], L31_0a, reset);
  tkf0mo0w0_o0w0 I8 (L30_0r, L30_0a, L25_0r, L25_0a, L27_0r, L27_0a, reset);
  tks2_o0w2_0c2o0w0_1o0w0_3o0w0 I9 (L8_0r0[1:0], L8_0r1[1:0], L8_0a, L14_0r, L14_0a, L22_0r, L22_0a, L30_0r, L30_0a, reset);
  tkm3x0b I10 (L16_0r, L16_0a, L24_0r, L24_0a, L32_0r, L32_0a, L33_0r, L33_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I11 (L2_0r0, L2_0r1, L2_0a, L3_0r, L3_0a, L7_0r, L7_0a, reset);
  tkm2x0b I12 (L6_0r, L6_0a, L33_0r, L33_0a, L34_0r, L34_0a, reset);
  tkvi32_wo0w32_ro0w32o0w31o1w31o1w31 I13 (L35_0r0[31:0], L35_0r1[31:0], L35_0a, L1_0r, L1_0a, L3_0r, L3_0a, L11_0r, L11_0a, L17_0r, L17_0a, L25_0r, L25_0a, L5_0r0[31:0], L5_0r1[31:0], L5_0a, L12_0r0[30:0], L12_0r1[30:0], L12_0a, L18_0r0[30:0], L18_0r1[30:0], L18_0a, L26_0r0[30:0], L26_0r1[30:0], L26_0a, reset);
  tko0m2_1nm2b0 I14 (L46_0r, L46_0a, L47_0r0[1:0], L47_0r1[1:0], L47_0a, reset);
  tkj32m2_30 I15 (L47_0r0[1:0], L47_0r1[1:0], L47_0a, L49_0r0[29:0], L49_0r1[29:0], L49_0a, L52_0r0[31:0], L52_0r1[31:0], L52_0a, reset);
  tkf0mo0w0_o0w0 I16 (L51_0r, L51_0a, L46_0r, L46_0a, L48_0r, L48_0a, reset);
  tko0m2_1nm2b0 I17 (L56_0r, L56_0a, L57_0r0[1:0], L57_0r1[1:0], L57_0a, reset);
  tkj32m30_2 I18 (L55_0r0[29:0], L55_0r1[29:0], L55_0a, L57_0r0[1:0], L57_0r1[1:0], L57_0a, L60_0r0[31:0], L60_0r1[31:0], L60_0a, reset);
  tkf0mo0w0_o0w0 I19 (L59_0r, L59_0a, L54_0r, L54_0a, L56_0r, L56_0a, reset);
  tko0m2_1nm2b3 I20 (L64_0r, L64_0a, L65_0r0[1:0], L65_0r1[1:0], L65_0a, reset);
  tkj32m30_2 I21 (L63_0r0[29:0], L63_0r1[29:0], L63_0a, L65_0r0[1:0], L65_0r1[1:0], L65_0a, L68_0r0[31:0], L68_0r1[31:0], L68_0a, reset);
  tkf0mo0w0_o0w0 I22 (L67_0r, L67_0a, L62_0r, L62_0a, L64_0r, L64_0a, reset);
  tks2_o0w2_0c2o0w0_1o0w0_3o0w0 I23 (L45_0r0[1:0], L45_0r1[1:0], L45_0a, L51_0r, L51_0a, L59_0r, L59_0a, L67_0r, L67_0a, reset);
  tkm3x0b I24 (L53_0r, L53_0a, L61_0r, L61_0a, L69_0r, L69_0a, L70_0r, L70_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I25 (L39_0r0, L39_0r1, L39_0a, L40_0r, L40_0a, L44_0r, L44_0a, reset);
  tkm2x0b I26 (L43_0r, L43_0a, L70_0r, L70_0a, L71_0r, L71_0a, reset);
  tkvi32_wo0w32_ro0w32o0w30o2w30o2w30 I27 (L72_0r0[31:0], L72_0r1[31:0], L72_0a, L38_0r, L38_0a, L40_0r, L40_0a, L48_0r, L48_0a, L54_0r, L54_0a, L62_0r, L62_0a, L42_0r0[31:0], L42_0r1[31:0], L42_0a, L49_0r0[29:0], L49_0r1[29:0], L49_0a, L55_0r0[29:0], L55_0r1[29:0], L55_0a, L63_0r0[29:0], L63_0r1[29:0], L63_0a, reset);
  tkf0mo0w0_o0w0 I28 (L75_0r, L75_0a, L37_0r, L37_0a, L74_0r, L74_0a, reset);
  tkj0m0_0 I29 (L34_0r, L34_0a, L71_0r, L71_0a, L76_0r, L76_0a, reset);
  tkf32mo0w0_o0w32 I30 (L42_0r0[31:0], L42_0r1[31:0], L42_0a, L77_0r, L77_0a, L78_0r0[31:0], L78_0r1[31:0], L78_0a, reset);
  tkf32mo0w0_o0w32 I31 (L52_0r0[31:0], L52_0r1[31:0], L52_0a, L79_0r, L79_0a, L80_0r0[31:0], L80_0r1[31:0], L80_0a, reset);
  tkf32mo0w0_o0w32 I32 (L60_0r0[31:0], L60_0r1[31:0], L60_0a, L81_0r, L81_0a, L82_0r0[31:0], L82_0r1[31:0], L82_0a, reset);
  tkf32mo0w0_o0w32 I33 (L68_0r0[31:0], L68_0r1[31:0], L68_0a, L83_0r, L83_0a, L84_0r0[31:0], L84_0r1[31:0], L84_0a, reset);
  tkm4x32b I34 (L78_0r0[31:0], L78_0r1[31:0], L78_0a, L80_0r0[31:0], L80_0r1[31:0], L80_0a, L82_0r0[31:0], L82_0r1[31:0], L82_0a, L84_0r0[31:0], L84_0r1[31:0], L84_0a, L85_0r0[31:0], L85_0r1[31:0], L85_0a, reset);
  tkf32mo0w0_o0w32 I35 (L85_0r0[31:0], L85_0r1[31:0], L85_0a, L86_0r, L86_0a, L87_0r0[31:0], L87_0r1[31:0], L87_0a, reset);
  tko0m4_1nm4b1 I36 (L77_0r, L77_0a, L88_0r0[3:0], L88_0r1[3:0], L88_0a, reset);
  tko0m4_1nm4b2 I37 (L79_0r, L79_0a, L89_0r0[3:0], L89_0r1[3:0], L89_0a, reset);
  tko0m4_1nm4b4 I38 (L81_0r, L81_0a, L90_0r0[3:0], L90_0r1[3:0], L90_0a, reset);
  tko0m4_1nm4b8 I39 (L83_0r, L83_0a, L91_0r0[3:0], L91_0r1[3:0], L91_0a, reset);
  tkm4x4b I40 (L88_0r0[3:0], L88_0r1[3:0], L88_0a, L89_0r0[3:0], L89_0r1[3:0], L89_0a, L90_0r0[3:0], L90_0r1[3:0], L90_0a, L91_0r0[3:0], L91_0r1[3:0], L91_0a, L92_0r0[3:0], L92_0r1[3:0], L92_0a, reset);
  tkj4m0_4 I41 (L86_0r, L86_0a, L92_0r0[3:0], L92_0r1[3:0], L92_0a, L93_0r0[3:0], L93_0r1[3:0], L93_0a, reset);
  tks4_o0w4_1o0w0_2o0w0_4o0w0_8o0w0 I42 (L93_0r0[3:0], L93_0r1[3:0], L93_0a, L43_0r, L43_0a, L53_0r, L53_0a, L61_0r, L61_0a, L69_0r, L69_0a, reset);
  tkj32m32_0 I43 (L87_0r0[31:0], L87_0r1[31:0], L87_0a, L37_0r, L37_0a, L35_0r0[31:0], L35_0r1[31:0], L35_0a, reset);
  tko0m4_1nm4b0 I44 (L102_0r, L102_0a, L103_0r0[3:0], L103_0r1[3:0], L103_0a, reset);
  tkj32m4_28 I45 (L103_0r0[3:0], L103_0r1[3:0], L103_0a, L105_0r0[27:0], L105_0r1[27:0], L105_0a, L108_0r0[31:0], L108_0r1[31:0], L108_0a, reset);
  tkf0mo0w0_o0w0 I46 (L107_0r, L107_0a, L102_0r, L102_0a, L104_0r, L104_0a, reset);
  tko0m4_1nm4b0 I47 (L112_0r, L112_0a, L113_0r0[3:0], L113_0r1[3:0], L113_0a, reset);
  tkj32m28_4 I48 (L111_0r0[27:0], L111_0r1[27:0], L111_0a, L113_0r0[3:0], L113_0r1[3:0], L113_0a, L116_0r0[31:0], L116_0r1[31:0], L116_0a, reset);
  tkf0mo0w0_o0w0 I49 (L115_0r, L115_0a, L110_0r, L110_0a, L112_0r, L112_0a, reset);
  tko0m4_1nm4bf I50 (L120_0r, L120_0a, L121_0r0[3:0], L121_0r1[3:0], L121_0a, reset);
  tkj32m28_4 I51 (L119_0r0[27:0], L119_0r1[27:0], L119_0a, L121_0r0[3:0], L121_0r1[3:0], L121_0a, L124_0r0[31:0], L124_0r1[31:0], L124_0a, reset);
  tkf0mo0w0_o0w0 I52 (L123_0r, L123_0a, L118_0r, L118_0a, L120_0r, L120_0a, reset);
  tks2_o0w2_0c2o0w0_1o0w0_3o0w0 I53 (L101_0r0[1:0], L101_0r1[1:0], L101_0a, L107_0r, L107_0a, L115_0r, L115_0a, L123_0r, L123_0a, reset);
  tkm3x0b I54 (L109_0r, L109_0a, L117_0r, L117_0a, L125_0r, L125_0a, L126_0r, L126_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I55 (L95_0r0, L95_0r1, L95_0a, L96_0r, L96_0a, L100_0r, L100_0a, reset);
  tkm2x0b I56 (L99_0r, L99_0a, L126_0r, L126_0a, L127_0r, L127_0a, reset);
  tkvi32_wo0w32_ro0w32o0w28o4w28o4w28 I57 (L128_0r0[31:0], L128_0r1[31:0], L128_0a, L94_0r, L94_0a, L96_0r, L96_0a, L104_0r, L104_0a, L110_0r, L110_0a, L118_0r, L118_0a, L98_0r0[31:0], L98_0r1[31:0], L98_0a, L105_0r0[27:0], L105_0r1[27:0], L105_0a, L111_0r0[27:0], L111_0r1[27:0], L111_0a, L119_0r0[27:0], L119_0r1[27:0], L119_0a, reset);
  tkf0mo0w0_o0w0 I58 (L131_0r, L131_0a, L75_0r, L75_0a, L130_0r, L130_0a, reset);
  tkj0m0_0 I59 (L76_0r, L76_0a, L127_0r, L127_0a, L132_0r, L132_0a, reset);
  tkf32mo0w0_o0w32 I60 (L98_0r0[31:0], L98_0r1[31:0], L98_0a, L133_0r, L133_0a, L134_0r0[31:0], L134_0r1[31:0], L134_0a, reset);
  tkf32mo0w0_o0w32 I61 (L108_0r0[31:0], L108_0r1[31:0], L108_0a, L135_0r, L135_0a, L136_0r0[31:0], L136_0r1[31:0], L136_0a, reset);
  tkf32mo0w0_o0w32 I62 (L116_0r0[31:0], L116_0r1[31:0], L116_0a, L137_0r, L137_0a, L138_0r0[31:0], L138_0r1[31:0], L138_0a, reset);
  tkf32mo0w0_o0w32 I63 (L124_0r0[31:0], L124_0r1[31:0], L124_0a, L139_0r, L139_0a, L140_0r0[31:0], L140_0r1[31:0], L140_0a, reset);
  tkm4x32b I64 (L134_0r0[31:0], L134_0r1[31:0], L134_0a, L136_0r0[31:0], L136_0r1[31:0], L136_0a, L138_0r0[31:0], L138_0r1[31:0], L138_0a, L140_0r0[31:0], L140_0r1[31:0], L140_0a, L141_0r0[31:0], L141_0r1[31:0], L141_0a, reset);
  tkf32mo0w0_o0w32 I65 (L141_0r0[31:0], L141_0r1[31:0], L141_0a, L142_0r, L142_0a, L143_0r0[31:0], L143_0r1[31:0], L143_0a, reset);
  tko0m4_1nm4b1 I66 (L133_0r, L133_0a, L144_0r0[3:0], L144_0r1[3:0], L144_0a, reset);
  tko0m4_1nm4b2 I67 (L135_0r, L135_0a, L145_0r0[3:0], L145_0r1[3:0], L145_0a, reset);
  tko0m4_1nm4b4 I68 (L137_0r, L137_0a, L146_0r0[3:0], L146_0r1[3:0], L146_0a, reset);
  tko0m4_1nm4b8 I69 (L139_0r, L139_0a, L147_0r0[3:0], L147_0r1[3:0], L147_0a, reset);
  tkm4x4b I70 (L144_0r0[3:0], L144_0r1[3:0], L144_0a, L145_0r0[3:0], L145_0r1[3:0], L145_0a, L146_0r0[3:0], L146_0r1[3:0], L146_0a, L147_0r0[3:0], L147_0r1[3:0], L147_0a, L148_0r0[3:0], L148_0r1[3:0], L148_0a, reset);
  tkj4m0_4 I71 (L142_0r, L142_0a, L148_0r0[3:0], L148_0r1[3:0], L148_0a, L149_0r0[3:0], L149_0r1[3:0], L149_0a, reset);
  tks4_o0w4_1o0w0_2o0w0_4o0w0_8o0w0 I72 (L149_0r0[3:0], L149_0r1[3:0], L149_0a, L99_0r, L99_0a, L109_0r, L109_0a, L117_0r, L117_0a, L125_0r, L125_0a, reset);
  tkj32m32_0 I73 (L143_0r0[31:0], L143_0r1[31:0], L143_0a, L74_0r, L74_0a, L72_0r0[31:0], L72_0r1[31:0], L72_0a, reset);
  tko0m8_1nm8b0 I74 (L158_0r, L158_0a, L159_0r0[7:0], L159_0r1[7:0], L159_0a, reset);
  tkj32m8_24 I75 (L159_0r0[7:0], L159_0r1[7:0], L159_0a, L161_0r0[23:0], L161_0r1[23:0], L161_0a, L164_0r0[31:0], L164_0r1[31:0], L164_0a, reset);
  tkf0mo0w0_o0w0 I76 (L163_0r, L163_0a, L158_0r, L158_0a, L160_0r, L160_0a, reset);
  tko0m8_1nm8b0 I77 (L168_0r, L168_0a, L169_0r0[7:0], L169_0r1[7:0], L169_0a, reset);
  tkj32m24_8 I78 (L167_0r0[23:0], L167_0r1[23:0], L167_0a, L169_0r0[7:0], L169_0r1[7:0], L169_0a, L172_0r0[31:0], L172_0r1[31:0], L172_0a, reset);
  tkf0mo0w0_o0w0 I79 (L171_0r, L171_0a, L166_0r, L166_0a, L168_0r, L168_0a, reset);
  tko0m8_1nm8bff I80 (L176_0r, L176_0a, L177_0r0[7:0], L177_0r1[7:0], L177_0a, reset);
  tkj32m24_8 I81 (L175_0r0[23:0], L175_0r1[23:0], L175_0a, L177_0r0[7:0], L177_0r1[7:0], L177_0a, L180_0r0[31:0], L180_0r1[31:0], L180_0a, reset);
  tkf0mo0w0_o0w0 I82 (L179_0r, L179_0a, L174_0r, L174_0a, L176_0r, L176_0a, reset);
  tks2_o0w2_0c2o0w0_1o0w0_3o0w0 I83 (L157_0r0[1:0], L157_0r1[1:0], L157_0a, L163_0r, L163_0a, L171_0r, L171_0a, L179_0r, L179_0a, reset);
  tkm3x0b I84 (L165_0r, L165_0a, L173_0r, L173_0a, L181_0r, L181_0a, L182_0r, L182_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I85 (L151_0r0, L151_0r1, L151_0a, L152_0r, L152_0a, L156_0r, L156_0a, reset);
  tkm2x0b I86 (L155_0r, L155_0a, L182_0r, L182_0a, L183_0r, L183_0a, reset);
  tkvi32_wo0w32_ro0w32o0w24o8w24o8w24 I87 (L184_0r0[31:0], L184_0r1[31:0], L184_0a, L150_0r, L150_0a, L152_0r, L152_0a, L160_0r, L160_0a, L166_0r, L166_0a, L174_0r, L174_0a, L154_0r0[31:0], L154_0r1[31:0], L154_0a, L161_0r0[23:0], L161_0r1[23:0], L161_0a, L167_0r0[23:0], L167_0r1[23:0], L167_0a, L175_0r0[23:0], L175_0r1[23:0], L175_0a, reset);
  tkf0mo0w0_o0w0 I88 (L187_0r, L187_0a, L131_0r, L131_0a, L186_0r, L186_0a, reset);
  tkj0m0_0 I89 (L132_0r, L132_0a, L183_0r, L183_0a, L188_0r, L188_0a, reset);
  tkf32mo0w0_o0w32 I90 (L154_0r0[31:0], L154_0r1[31:0], L154_0a, L189_0r, L189_0a, L190_0r0[31:0], L190_0r1[31:0], L190_0a, reset);
  tkf32mo0w0_o0w32 I91 (L164_0r0[31:0], L164_0r1[31:0], L164_0a, L191_0r, L191_0a, L192_0r0[31:0], L192_0r1[31:0], L192_0a, reset);
  tkf32mo0w0_o0w32 I92 (L172_0r0[31:0], L172_0r1[31:0], L172_0a, L193_0r, L193_0a, L194_0r0[31:0], L194_0r1[31:0], L194_0a, reset);
  tkf32mo0w0_o0w32 I93 (L180_0r0[31:0], L180_0r1[31:0], L180_0a, L195_0r, L195_0a, L196_0r0[31:0], L196_0r1[31:0], L196_0a, reset);
  tkm4x32b I94 (L190_0r0[31:0], L190_0r1[31:0], L190_0a, L192_0r0[31:0], L192_0r1[31:0], L192_0a, L194_0r0[31:0], L194_0r1[31:0], L194_0a, L196_0r0[31:0], L196_0r1[31:0], L196_0a, L197_0r0[31:0], L197_0r1[31:0], L197_0a, reset);
  tkf32mo0w0_o0w32 I95 (L197_0r0[31:0], L197_0r1[31:0], L197_0a, L198_0r, L198_0a, L199_0r0[31:0], L199_0r1[31:0], L199_0a, reset);
  tko0m4_1nm4b1 I96 (L189_0r, L189_0a, L200_0r0[3:0], L200_0r1[3:0], L200_0a, reset);
  tko0m4_1nm4b2 I97 (L191_0r, L191_0a, L201_0r0[3:0], L201_0r1[3:0], L201_0a, reset);
  tko0m4_1nm4b4 I98 (L193_0r, L193_0a, L202_0r0[3:0], L202_0r1[3:0], L202_0a, reset);
  tko0m4_1nm4b8 I99 (L195_0r, L195_0a, L203_0r0[3:0], L203_0r1[3:0], L203_0a, reset);
  tkm4x4b I100 (L200_0r0[3:0], L200_0r1[3:0], L200_0a, L201_0r0[3:0], L201_0r1[3:0], L201_0a, L202_0r0[3:0], L202_0r1[3:0], L202_0a, L203_0r0[3:0], L203_0r1[3:0], L203_0a, L204_0r0[3:0], L204_0r1[3:0], L204_0a, reset);
  tkj4m0_4 I101 (L198_0r, L198_0a, L204_0r0[3:0], L204_0r1[3:0], L204_0a, L205_0r0[3:0], L205_0r1[3:0], L205_0a, reset);
  tks4_o0w4_1o0w0_2o0w0_4o0w0_8o0w0 I102 (L205_0r0[3:0], L205_0r1[3:0], L205_0a, L155_0r, L155_0a, L165_0r, L165_0a, L173_0r, L173_0a, L181_0r, L181_0a, reset);
  tkj32m32_0 I103 (L199_0r0[31:0], L199_0r1[31:0], L199_0a, L130_0r, L130_0a, L128_0r0[31:0], L128_0r1[31:0], L128_0a, reset);
  tko0m16_1nm16b0 I104 (L214_0r, L214_0a, L215_0r0[15:0], L215_0r1[15:0], L215_0a, reset);
  tkj32m16_16 I105 (L215_0r0[15:0], L215_0r1[15:0], L215_0a, L217_0r0[15:0], L217_0r1[15:0], L217_0a, L220_0r0[31:0], L220_0r1[31:0], L220_0a, reset);
  tkf0mo0w0_o0w0 I106 (L219_0r, L219_0a, L214_0r, L214_0a, L216_0r, L216_0a, reset);
  tko0m16_1nm16b0 I107 (L224_0r, L224_0a, L225_0r0[15:0], L225_0r1[15:0], L225_0a, reset);
  tkj32m16_16 I108 (L223_0r0[15:0], L223_0r1[15:0], L223_0a, L225_0r0[15:0], L225_0r1[15:0], L225_0a, L228_0r0[31:0], L228_0r1[31:0], L228_0a, reset);
  tkf0mo0w0_o0w0 I109 (L227_0r, L227_0a, L222_0r, L222_0a, L224_0r, L224_0a, reset);
  tko0m16_1nm16bffff I110 (L232_0r, L232_0a, L233_0r0[15:0], L233_0r1[15:0], L233_0a, reset);
  tkj32m16_16 I111 (L231_0r0[15:0], L231_0r1[15:0], L231_0a, L233_0r0[15:0], L233_0r1[15:0], L233_0a, L236_0r0[31:0], L236_0r1[31:0], L236_0a, reset);
  tkf0mo0w0_o0w0 I112 (L235_0r, L235_0a, L230_0r, L230_0a, L232_0r, L232_0a, reset);
  tks2_o0w2_0c2o0w0_1o0w0_3o0w0 I113 (L213_0r0[1:0], L213_0r1[1:0], L213_0a, L219_0r, L219_0a, L227_0r, L227_0a, L235_0r, L235_0a, reset);
  tkm3x0b I114 (L221_0r, L221_0a, L229_0r, L229_0a, L237_0r, L237_0a, L238_0r, L238_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I115 (L207_0r0, L207_0r1, L207_0a, L208_0r, L208_0a, L212_0r, L212_0a, reset);
  tkm2x0b I116 (L211_0r, L211_0a, L238_0r, L238_0a, L239_0r, L239_0a, reset);
  tkvi32_wo0w32_ro0w32o0w16o16w16o16w16 I117 (L240_0r0[31:0], L240_0r1[31:0], L240_0a, L206_0r, L206_0a, L208_0r, L208_0a, L216_0r, L216_0a, L222_0r, L222_0a, L230_0r, L230_0a, L210_0r0[31:0], L210_0r1[31:0], L210_0a, L217_0r0[15:0], L217_0r1[15:0], L217_0a, L223_0r0[15:0], L223_0r1[15:0], L223_0a, L231_0r0[15:0], L231_0r1[15:0], L231_0a, reset);
  tkf0mo0w0_o0w0 I118 (L243_0r, L243_0a, L187_0r, L187_0a, L242_0r, L242_0a, reset);
  tkj0m0_0 I119 (L188_0r, L188_0a, L239_0r, L239_0a, L244_0r, L244_0a, reset);
  tkf32mo0w0_o0w32 I120 (L210_0r0[31:0], L210_0r1[31:0], L210_0a, L245_0r, L245_0a, L246_0r0[31:0], L246_0r1[31:0], L246_0a, reset);
  tkf32mo0w0_o0w32 I121 (L220_0r0[31:0], L220_0r1[31:0], L220_0a, L247_0r, L247_0a, L248_0r0[31:0], L248_0r1[31:0], L248_0a, reset);
  tkf32mo0w0_o0w32 I122 (L228_0r0[31:0], L228_0r1[31:0], L228_0a, L249_0r, L249_0a, L250_0r0[31:0], L250_0r1[31:0], L250_0a, reset);
  tkf32mo0w0_o0w32 I123 (L236_0r0[31:0], L236_0r1[31:0], L236_0a, L251_0r, L251_0a, L252_0r0[31:0], L252_0r1[31:0], L252_0a, reset);
  tkm4x32b I124 (L246_0r0[31:0], L246_0r1[31:0], L246_0a, L248_0r0[31:0], L248_0r1[31:0], L248_0a, L250_0r0[31:0], L250_0r1[31:0], L250_0a, L252_0r0[31:0], L252_0r1[31:0], L252_0a, L253_0r0[31:0], L253_0r1[31:0], L253_0a, reset);
  tkf32mo0w0_o0w32 I125 (L253_0r0[31:0], L253_0r1[31:0], L253_0a, L254_0r, L254_0a, L255_0r0[31:0], L255_0r1[31:0], L255_0a, reset);
  tko0m4_1nm4b1 I126 (L245_0r, L245_0a, L256_0r0[3:0], L256_0r1[3:0], L256_0a, reset);
  tko0m4_1nm4b2 I127 (L247_0r, L247_0a, L257_0r0[3:0], L257_0r1[3:0], L257_0a, reset);
  tko0m4_1nm4b4 I128 (L249_0r, L249_0a, L258_0r0[3:0], L258_0r1[3:0], L258_0a, reset);
  tko0m4_1nm4b8 I129 (L251_0r, L251_0a, L259_0r0[3:0], L259_0r1[3:0], L259_0a, reset);
  tkm4x4b I130 (L256_0r0[3:0], L256_0r1[3:0], L256_0a, L257_0r0[3:0], L257_0r1[3:0], L257_0a, L258_0r0[3:0], L258_0r1[3:0], L258_0a, L259_0r0[3:0], L259_0r1[3:0], L259_0a, L260_0r0[3:0], L260_0r1[3:0], L260_0a, reset);
  tkj4m0_4 I131 (L254_0r, L254_0a, L260_0r0[3:0], L260_0r1[3:0], L260_0a, L261_0r0[3:0], L261_0r1[3:0], L261_0a, reset);
  tks4_o0w4_1o0w0_2o0w0_4o0w0_8o0w0 I132 (L261_0r0[3:0], L261_0r1[3:0], L261_0a, L211_0r, L211_0a, L221_0r, L221_0a, L229_0r, L229_0a, L237_0r, L237_0a, reset);
  tkj32m32_0 I133 (L255_0r0[31:0], L255_0r1[31:0], L255_0a, L186_0r, L186_0a, L184_0r0[31:0], L184_0r1[31:0], L184_0a, reset);
  tkvdistanceI5_wo0w5_ro0w1o1w1o2w1o3w1o4w1 I134 (L262_0r0[4:0], L262_0r1[4:0], L262_0a, L263_0r, L263_0a, L1_0r, L1_0a, L38_0r, L38_0a, L94_0r, L94_0a, L150_0r, L150_0a, L206_0r, L206_0a, L2_0r0, L2_0r1, L2_0a, L39_0r0, L39_0r1, L39_0a, L95_0r0, L95_0r1, L95_0a, L151_0r0, L151_0r1, L151_0a, L207_0r0, L207_0r1, L207_0a, reset);
  tkvshift2_wo0w2_ro0w2o0w2o0w2o0w2o0w2 I135 (L264_0r0[1:0], L264_0r1[1:0], L264_0a, L265_0r, L265_0a, L7_0r, L7_0a, L44_0r, L44_0a, L100_0r, L100_0a, L156_0r, L156_0a, L212_0r, L212_0a, L8_0r0[1:0], L8_0r1[1:0], L8_0a, L45_0r0[1:0], L45_0r1[1:0], L45_0a, L101_0r0[1:0], L101_0r1[1:0], L101_0a, L157_0r0[1:0], L157_0r1[1:0], L157_0a, L213_0r0[1:0], L213_0r1[1:0], L213_0a, reset);
  tkj0m0_0 I136 (L263_0r, L263_0a, L265_0r, L265_0a, L243_0r, L243_0a, reset);
  tkf0mo0w0_o0w0 I137 (L269_0r, L269_0a, L267_0r, L267_0a, L268_0r, L268_0a, reset);
  tkj2m2_0 I138 (shift_0r0[1:0], shift_0r1[1:0], shift_0a, L268_0r, L268_0a, L264_0r0[1:0], L264_0r1[1:0], L264_0a, reset);
  tkj5m5_0 I139 (distanceI_0r0[4:0], distanceI_0r1[4:0], distanceI_0a, L267_0r, L267_0a, L262_0r0[4:0], L262_0r1[4:0], L262_0a, reset);
  tkf32mo0w0_o0w32 I140 (L5_0r0[31:0], L5_0r1[31:0], L5_0a, L273_0r, L273_0a, L274_0r0[31:0], L274_0r1[31:0], L274_0a, reset);
  tkf32mo0w0_o0w32 I141 (L15_0r0[31:0], L15_0r1[31:0], L15_0a, L275_0r, L275_0a, L276_0r0[31:0], L276_0r1[31:0], L276_0a, reset);
  tkf32mo0w0_o0w32 I142 (L23_0r0[31:0], L23_0r1[31:0], L23_0a, L277_0r, L277_0a, L278_0r0[31:0], L278_0r1[31:0], L278_0a, reset);
  tkf32mo0w0_o0w32 I143 (L31_0r0[31:0], L31_0r1[31:0], L31_0a, L279_0r, L279_0a, L280_0r0[31:0], L280_0r1[31:0], L280_0a, reset);
  tkm4x32b I144 (L274_0r0[31:0], L274_0r1[31:0], L274_0a, L276_0r0[31:0], L276_0r1[31:0], L276_0a, L278_0r0[31:0], L278_0r1[31:0], L278_0a, L280_0r0[31:0], L280_0r1[31:0], L280_0a, L281_0r0[31:0], L281_0r1[31:0], L281_0a, reset);
  tkf32mo0w0_o0w32 I145 (L281_0r0[31:0], L281_0r1[31:0], L281_0a, L282_0r, L282_0a, result_0r0[31:0], result_0r1[31:0], result_0a, reset);
  tko0m4_1nm4b1 I146 (L273_0r, L273_0a, L284_0r0[3:0], L284_0r1[3:0], L284_0a, reset);
  tko0m4_1nm4b2 I147 (L275_0r, L275_0a, L285_0r0[3:0], L285_0r1[3:0], L285_0a, reset);
  tko0m4_1nm4b4 I148 (L277_0r, L277_0a, L286_0r0[3:0], L286_0r1[3:0], L286_0a, reset);
  tko0m4_1nm4b8 I149 (L279_0r, L279_0a, L287_0r0[3:0], L287_0r1[3:0], L287_0a, reset);
  tkm4x4b I150 (L284_0r0[3:0], L284_0r1[3:0], L284_0a, L285_0r0[3:0], L285_0r1[3:0], L285_0a, L286_0r0[3:0], L286_0r1[3:0], L286_0a, L287_0r0[3:0], L287_0r1[3:0], L287_0a, L288_0r0[3:0], L288_0r1[3:0], L288_0a, reset);
  tkj4m0_4 I151 (L282_0r, L282_0a, L288_0r0[3:0], L288_0r1[3:0], L288_0a, L289_0r0[3:0], L289_0r1[3:0], L289_0a, reset);
  tks4_o0w4_1o0w0_2o0w0_4o0w0_8o0w0 I152 (L289_0r0[3:0], L289_0r1[3:0], L289_0a, L6_0r, L6_0a, L16_0r, L16_0a, L24_0r, L24_0a, L32_0r, L32_0a, reset);
  tkj32m32_0 I153 (arg_0r0[31:0], arg_0r1[31:0], arg_0a, L242_0r, L242_0a, L240_0r0[31:0], L240_0r1[31:0], L240_0a, reset);
  tki I154 (L244_0r, L244_0a, L269_0r, L269_0a, reset);
endmodule

module teak_Alu (op_0r0, op_0r1, op_0a, result_0r0, result_0r1, result_0a, flags_0r0, flags_0r1, flags_0a, lhs_0r0, lhs_0r1, lhs_0a, rhs_0r0, rhs_0r1, rhs_0a, reset);
  input [6:0] op_0r0;
  input [6:0] op_0r1;
  output op_0a;
  output [31:0] result_0r0;
  output [31:0] result_0r1;
  input result_0a;
  output [3:0] flags_0r0;
  output [3:0] flags_0r1;
  input flags_0a;
  input [31:0] lhs_0r0;
  input [31:0] lhs_0r1;
  output lhs_0a;
  input [31:0] rhs_0r0;
  input [31:0] rhs_0r1;
  output rhs_0a;
  input reset;
  wire [1:0] L1_0r0;
  wire [1:0] L1_0r1;
  wire L1_0a;
  wire [4:0] L2_0r0;
  wire [4:0] L2_0r1;
  wire L2_0a;
  wire [31:0] L4_0r0;
  wire [31:0] L4_0r1;
  wire L4_0a;
  wire L6_0r;
  wire L6_0a;
  wire [5:0] L7_0r0;
  wire [5:0] L7_0r1;
  wire L7_0a;
  wire L8_0r;
  wire L8_0a;
  wire [31:0] L10_0r0;
  wire [31:0] L10_0r1;
  wire L10_0a;
  wire L11_0r;
  wire L11_0a;
  wire L13_0r;
  wire L13_0a;
  wire [31:0] L14_0r0;
  wire [31:0] L14_0r1;
  wire L14_0a;
  wire [31:0] L15_0r0;
  wire [31:0] L15_0r1;
  wire L15_0a;
  wire L16_0r;
  wire L16_0a;
  wire L17_0r;
  wire L17_0a;
  wire L18_0r;
  wire L18_0a;
  wire [5:0] L19_0r0;
  wire [5:0] L19_0r1;
  wire L19_0a;
  wire L20_0r;
  wire L20_0a;
  wire L22_0r0;
  wire L22_0r1;
  wire L22_0a;
  wire L23_0r;
  wire L23_0a;
  wire L24_0r;
  wire L24_0a;
  wire L26_0r0;
  wire L26_0r1;
  wire L26_0a;
  wire L27_0r;
  wire L27_0a;
  wire L28_0r;
  wire L28_0a;
  wire L30_0r0;
  wire L30_0r1;
  wire L30_0a;
  wire L31_0r;
  wire L31_0a;
  wire L33_0r;
  wire L33_0a;
  wire L34_0r0;
  wire L34_0r1;
  wire L34_0a;
  wire L35_0r0;
  wire L35_0r1;
  wire L35_0a;
  wire L36_0r;
  wire L36_0a;
  wire L37_0r;
  wire L37_0a;
  wire L39_0r;
  wire L39_0a;
  wire [5:0] L40_0r0;
  wire [5:0] L40_0r1;
  wire L40_0a;
  wire L41_0r;
  wire L41_0a;
  wire L43_0r;
  wire L43_0a;
  wire L44_0r0;
  wire L44_0r1;
  wire L44_0a;
  wire L45_0r;
  wire L45_0a;
  wire [31:0] L46_0r0;
  wire [31:0] L46_0r1;
  wire L46_0a;
  wire [32:0] L47_0r0;
  wire [32:0] L47_0r1;
  wire L47_0a;
  wire L48_0r;
  wire L48_0a;
  wire L49_0r0;
  wire L49_0r1;
  wire L49_0a;
  wire L50_0r;
  wire L50_0a;
  wire [31:0] L51_0r0;
  wire [31:0] L51_0r1;
  wire L51_0a;
  wire [32:0] L52_0r0;
  wire [32:0] L52_0r1;
  wire L52_0a;
  wire [65:0] L53_0r0;
  wire [65:0] L53_0r1;
  wire L53_0a;
  wire [33:0] L54_0r0;
  wire [33:0] L54_0r1;
  wire L54_0a;
  wire L55_0r;
  wire L55_0a;
  wire [32:0] L56_0r0;
  wire [32:0] L56_0r1;
  wire L56_0a;
  wire L57_0r;
  wire L57_0a;
  wire L58_0r;
  wire L58_0a;
  wire [31:0] L59_0r0;
  wire [31:0] L59_0r1;
  wire L59_0a;
  wire L60_0r;
  wire L60_0a;
  wire [31:0] L61_0r0;
  wire [31:0] L61_0r1;
  wire L61_0a;
  wire [63:0] L62_0r0;
  wire [63:0] L62_0r1;
  wire L62_0a;
  wire L64_0r;
  wire L64_0a;
  wire [31:0] L65_0r0;
  wire [31:0] L65_0r1;
  wire L65_0a;
  wire L66_0r;
  wire L66_0a;
  wire L67_0r;
  wire L67_0a;
  wire [31:0] L68_0r0;
  wire [31:0] L68_0r1;
  wire L68_0a;
  wire L69_0r;
  wire L69_0a;
  wire [31:0] L70_0r0;
  wire [31:0] L70_0r1;
  wire L70_0a;
  wire [63:0] L71_0r0;
  wire [63:0] L71_0r1;
  wire L71_0a;
  wire L73_0r;
  wire L73_0a;
  wire [31:0] L74_0r0;
  wire [31:0] L74_0r1;
  wire L74_0a;
  wire L75_0r;
  wire L75_0a;
  wire L76_0r;
  wire L76_0a;
  wire [31:0] L77_0r0;
  wire [31:0] L77_0r1;
  wire L77_0a;
  wire L78_0r;
  wire L78_0a;
  wire [31:0] L79_0r0;
  wire [31:0] L79_0r1;
  wire L79_0a;
  wire [63:0] L80_0r0;
  wire [63:0] L80_0r1;
  wire L80_0a;
  wire L82_0r;
  wire L82_0a;
  wire [31:0] L83_0r0;
  wire [31:0] L83_0r1;
  wire L83_0a;
  wire L84_0r;
  wire L84_0a;
  wire L85_0r;
  wire L85_0a;
  wire [1:0] L87_0r0;
  wire [1:0] L87_0r1;
  wire L87_0a;
  wire L88_0r;
  wire L88_0a;
  wire L89_0r;
  wire L89_0a;
  wire [1:0] L91_0r0;
  wire [1:0] L91_0r1;
  wire L91_0a;
  wire L92_0r;
  wire L92_0a;
  wire L93_0r;
  wire L93_0a;
  wire L94_0r0;
  wire L94_0r1;
  wire L94_0a;
  wire L95_0r;
  wire L95_0a;
  wire L96_0r0;
  wire L96_0r1;
  wire L96_0a;
  wire L98_0r;
  wire L98_0a;
  wire [1:0] L99_0r0;
  wire [1:0] L99_0r1;
  wire L99_0a;
  wire L100_0r;
  wire L100_0a;
  wire L101_0r;
  wire L101_0a;
  wire L102_0r;
  wire L102_0a;
  wire [5:0] L103_0r0;
  wire [5:0] L103_0r1;
  wire L103_0a;
  wire L104_0r;
  wire L104_0a;
  wire L105_0r;
  wire L105_0a;
  wire [4:0] L107_0r0;
  wire [4:0] L107_0r1;
  wire L107_0a;
  wire L108_0r;
  wire L108_0a;
  wire L109_0r;
  wire L109_0a;
  wire [31:0] L111_0r0;
  wire [31:0] L111_0r1;
  wire L111_0a;
  wire L112_0r;
  wire L112_0a;
  wire L113_0r;
  wire L113_0a;
  wire L114_0r;
  wire L114_0a;
  wire L115_0r;
  wire L115_0a;
  wire L116_0r;
  wire L116_0a;
  wire L117_0r;
  wire L117_0a;
  wire L118_0r;
  wire L118_0a;
  wire [32:0] L120_0r0;
  wire [32:0] L120_0r1;
  wire L120_0a;
  wire L121_0r;
  wire L121_0a;
  wire [32:0] L122_0r0;
  wire [32:0] L122_0r1;
  wire L122_0a;
  wire L124_0r;
  wire L124_0a;
  wire [32:0] L125_0r0;
  wire [32:0] L125_0r1;
  wire L125_0a;
  wire [32:0] L126_0r0;
  wire [32:0] L126_0r1;
  wire L126_0a;
  wire L127_0r;
  wire L127_0a;
  wire L128_0r;
  wire L128_0a;
  wire [31:0] L129_0r0;
  wire [31:0] L129_0r1;
  wire L129_0a;
  wire L130_0r;
  wire L130_0a;
  wire L131_0r0;
  wire L131_0r1;
  wire L131_0a;
  wire L133_0r;
  wire L133_0a;
  wire [32:0] L134_0r0;
  wire [32:0] L134_0r1;
  wire L134_0a;
  wire L135_0r;
  wire L135_0a;
  wire [31:0] L136_0r0;
  wire [31:0] L136_0r1;
  wire L136_0a;
  wire L138_0r;
  wire L138_0a;
  wire [31:0] L139_0r0;
  wire [31:0] L139_0r1;
  wire L139_0a;
  wire [31:0] L140_0r0;
  wire [31:0] L140_0r1;
  wire L140_0a;
  wire L141_0r;
  wire L141_0a;
  wire L142_0r;
  wire L142_0a;
  wire [31:0] L143_0r0;
  wire [31:0] L143_0r1;
  wire L143_0a;
  wire L144_0r;
  wire L144_0a;
  wire L145_0r0;
  wire L145_0r1;
  wire L145_0a;
  wire L147_0r;
  wire L147_0a;
  wire [32:0] L148_0r0;
  wire [32:0] L148_0r1;
  wire L148_0a;
  wire L149_0r;
  wire L149_0a;
  wire [31:0] L150_0r0;
  wire [31:0] L150_0r1;
  wire L150_0a;
  wire L152_0r;
  wire L152_0a;
  wire [31:0] L153_0r0;
  wire [31:0] L153_0r1;
  wire L153_0a;
  wire [31:0] L154_0r0;
  wire [31:0] L154_0r1;
  wire L154_0a;
  wire L155_0r;
  wire L155_0a;
  wire L156_0r;
  wire L156_0a;
  wire [2:0] L157_0r0;
  wire [2:0] L157_0r1;
  wire L157_0a;
  wire [2:0] L158_0r0;
  wire [2:0] L158_0r1;
  wire L158_0a;
  wire [2:0] L159_0r0;
  wire [2:0] L159_0r1;
  wire L159_0a;
  wire [2:0] L160_0r0;
  wire [2:0] L160_0r1;
  wire L160_0a;
  wire [2:0] L161_0r0;
  wire [2:0] L161_0r1;
  wire L161_0a;
  wire L162_0r;
  wire L162_0a;
  wire L163_0r;
  wire L163_0a;
  wire [31:0] L165_0r0;
  wire [31:0] L165_0r1;
  wire L165_0a;
  wire L166_0r;
  wire L166_0a;
  wire L167_0r;
  wire L167_0a;
  wire L168_0r;
  wire L168_0a;
  wire [31:0] L169_0r0;
  wire [31:0] L169_0r1;
  wire L169_0a;
  wire L170_0r;
  wire L170_0a;
  wire L171_0r0;
  wire L171_0r1;
  wire L171_0a;
  wire [32:0] L172_0r0;
  wire [32:0] L172_0r1;
  wire L172_0a;
  wire L173_0r0;
  wire L173_0r1;
  wire L173_0a;
  wire L174_0r;
  wire L174_0a;
  wire L175_0r0;
  wire L175_0r1;
  wire L175_0a;
  wire L176_0r;
  wire L176_0a;
  wire L177_0r0;
  wire L177_0r1;
  wire L177_0a;
  wire L178_0r;
  wire L178_0a;
  wire L179_0r0;
  wire L179_0r1;
  wire L179_0a;
  wire L180_0r;
  wire L180_0a;
  wire L181_0r0;
  wire L181_0r1;
  wire L181_0a;
  wire L182_0r;
  wire L182_0a;
  wire L183_0r0;
  wire L183_0r1;
  wire L183_0a;
  wire [1:0] L184_0r0;
  wire [1:0] L184_0r1;
  wire L184_0a;
  wire L185_0r0;
  wire L185_0r1;
  wire L185_0a;
  wire [1:0] L186_0r0;
  wire [1:0] L186_0r1;
  wire L186_0a;
  wire L187_0r0;
  wire L187_0r1;
  wire L187_0a;
  wire [1:0] L188_0r0;
  wire [1:0] L188_0r1;
  wire L188_0a;
  wire L189_0r0;
  wire L189_0r1;
  wire L189_0a;
  wire L190_0r;
  wire L190_0a;
  wire L191_0r0;
  wire L191_0r1;
  wire L191_0a;
  wire L192_0r;
  wire L192_0a;
  wire [5:0] L193_0r0;
  wire [5:0] L193_0r1;
  wire L193_0a;
  wire L194_0r;
  wire L194_0a;
  wire [5:0] L195_0r0;
  wire [5:0] L195_0r1;
  wire L195_0a;
  wire [11:0] L196_0r0;
  wire [11:0] L196_0r1;
  wire L196_0a;
  wire L197_0r0;
  wire L197_0r1;
  wire L197_0a;
  wire [1:0] L198_0r0;
  wire [1:0] L198_0r1;
  wire L198_0a;
  wire L199_0r0;
  wire L199_0r1;
  wire L199_0a;
  wire L201_0r;
  wire L201_0a;
  wire [3:0] L202_0r0;
  wire [3:0] L202_0r1;
  wire L202_0a;
  wire L203_0r;
  wire L203_0a;
  wire L204_0r;
  wire L204_0a;
  wire L205_0r;
  wire L205_0a;
  wire [32:0] L206_0r0;
  wire [32:0] L206_0r1;
  wire L206_0a;
  wire L208_0r;
  wire L208_0a;
  wire L209_0r;
  wire L209_0a;
  wire L210_0r;
  wire L210_0a;
  wire L211_0r;
  wire L211_0a;
  wire [32:0] L212_0r0;
  wire [32:0] L212_0r1;
  wire L212_0a;
  wire L213_0r;
  wire L213_0a;
  wire [32:0] L214_0r0;
  wire [32:0] L214_0r1;
  wire L214_0a;
  wire L215_0r;
  wire L215_0a;
  wire [32:0] L216_0r0;
  wire [32:0] L216_0r1;
  wire L216_0a;
  wire [32:0] L217_0r0;
  wire [32:0] L217_0r1;
  wire L217_0a;
  wire L218_0r;
  wire L218_0a;
  wire [32:0] L219_0r0;
  wire [32:0] L219_0r1;
  wire L219_0a;
  wire [2:0] L220_0r0;
  wire [2:0] L220_0r1;
  wire L220_0a;
  wire [2:0] L221_0r0;
  wire [2:0] L221_0r1;
  wire L221_0a;
  wire [2:0] L222_0r0;
  wire [2:0] L222_0r1;
  wire L222_0a;
  wire [2:0] L223_0r0;
  wire [2:0] L223_0r1;
  wire L223_0a;
  wire [2:0] L224_0r0;
  wire [2:0] L224_0r1;
  wire L224_0a;
  wire L226_0r;
  wire L226_0a;
  wire [31:0] L227_0r0;
  wire [31:0] L227_0r1;
  wire L227_0a;
  wire L228_0r;
  wire L228_0a;
  wire [31:0] L229_0r0;
  wire [31:0] L229_0r1;
  wire L229_0a;
  wire L230_0r;
  wire L230_0a;
  wire [31:0] L231_0r0;
  wire [31:0] L231_0r1;
  wire L231_0a;
  wire [31:0] L232_0r0;
  wire [31:0] L232_0r1;
  wire L232_0a;
  wire L233_0r;
  wire L233_0a;
  wire [2:0] L235_0r0;
  wire [2:0] L235_0r1;
  wire L235_0a;
  wire [2:0] L236_0r0;
  wire [2:0] L236_0r1;
  wire L236_0a;
  wire [2:0] L237_0r0;
  wire [2:0] L237_0r1;
  wire L237_0a;
  wire [2:0] L238_0r0;
  wire [2:0] L238_0r1;
  wire L238_0a;
  wire [2:0] L239_0r0;
  wire [2:0] L239_0r1;
  wire L239_0a;
  wire [31:0] L240_0r0;
  wire [31:0] L240_0r1;
  wire L240_0a;
  wire L241_0r;
  wire L241_0a;
  wire L242_0r0;
  wire L242_0r1;
  wire L242_0a;
  wire L243_0r;
  wire L243_0a;
  wire L245_0r;
  wire L245_0a;
  wire L246_0r;
  wire L246_0a;
  wire L247_0r;
  wire L247_0a;
  wire L248_0r;
  wire L248_0a;
  wire L249_0r;
  wire L249_0a;
  wire [6:0] L250_0r0;
  wire [6:0] L250_0r1;
  wire L250_0a;
  wire L251_0r;
  wire L251_0a;
  wire [31:0] L252_0r0;
  wire [31:0] L252_0r1;
  wire L252_0a;
  wire L253_0r;
  wire L253_0a;
  wire [31:0] L254_0r0;
  wire [31:0] L254_0r1;
  wire L254_0a;
  wire L255_0r;
  wire L255_0a;
  wire L257_0r;
  wire L257_0a;
  wire L258_0r;
  wire L258_0a;
  wire L259_0r;
  wire L259_0a;
  wire L260_0r;
  wire L260_0a;
  wire L265_0r;
  wire L265_0a;
  wire [1:0] L266_0r0;
  wire [1:0] L266_0r1;
  wire L266_0a;
  wire L267_0r;
  wire L267_0a;
  wire [1:0] L268_0r0;
  wire [1:0] L268_0r1;
  wire L268_0a;
  wire L269_0r;
  wire L269_0a;
  wire [1:0] L270_0r0;
  wire [1:0] L270_0r1;
  wire L270_0a;
  wire [1:0] L271_0r0;
  wire [1:0] L271_0r1;
  wire L271_0a;
  wire L272_0r;
  wire L272_0a;
  wire [2:0] L274_0r0;
  wire [2:0] L274_0r1;
  wire L274_0a;
  wire [2:0] L275_0r0;
  wire [2:0] L275_0r1;
  wire L275_0a;
  wire [2:0] L276_0r0;
  wire [2:0] L276_0r1;
  wire L276_0a;
  wire [2:0] L277_0r0;
  wire [2:0] L277_0r1;
  wire L277_0a;
  wire [2:0] L278_0r0;
  wire [2:0] L278_0r1;
  wire L278_0a;
  wire L279_0r;
  wire L279_0a;
  wire L280_0r0;
  wire L280_0r1;
  wire L280_0a;
  wire L281_0r;
  wire L281_0a;
  wire L282_0r0;
  wire L282_0r1;
  wire L282_0a;
  wire L283_0r;
  wire L283_0a;
  wire L284_0r0;
  wire L284_0r1;
  wire L284_0a;
  wire L285_0r;
  wire L285_0a;
  wire L286_0r0;
  wire L286_0r1;
  wire L286_0a;
  wire L287_0r0;
  wire L287_0r1;
  wire L287_0a;
  wire L288_0r;
  wire L288_0a;
  wire L289_0r0;
  wire L289_0r1;
  wire L289_0a;
  wire [3:0] L290_0r0;
  wire [3:0] L290_0r1;
  wire L290_0a;
  wire [3:0] L291_0r0;
  wire [3:0] L291_0r1;
  wire L291_0a;
  wire [3:0] L292_0r0;
  wire [3:0] L292_0r1;
  wire L292_0a;
  wire [3:0] L293_0r0;
  wire [3:0] L293_0r1;
  wire L293_0a;
  wire [3:0] L294_0r0;
  wire [3:0] L294_0r1;
  wire L294_0a;
  wire [3:0] L295_0r0;
  wire [3:0] L295_0r1;
  wire L295_0a;
  wire L296_0r;
  wire L296_0a;
  wire [31:0] L297_0r0;
  wire [31:0] L297_0r1;
  wire L297_0a;
  wire L298_0r;
  wire L298_0a;
  wire [31:0] L299_0r0;
  wire [31:0] L299_0r1;
  wire L299_0a;
  wire [31:0] L300_0r0;
  wire [31:0] L300_0r1;
  wire L300_0a;
  wire L301_0r;
  wire L301_0a;
  wire [31:0] L302_0r0;
  wire [31:0] L302_0r1;
  wire L302_0a;
  wire [1:0] L303_0r0;
  wire [1:0] L303_0r1;
  wire L303_0a;
  wire [1:0] L304_0r0;
  wire [1:0] L304_0r1;
  wire L304_0a;
  wire [1:0] L305_0r0;
  wire [1:0] L305_0r1;
  wire L305_0a;
  wire [1:0] L306_0r0;
  wire [1:0] L306_0r1;
  wire L306_0a;
  teak_Shifter I0 (L1_0r0[1:0], L1_0r1[1:0], L1_0a, L2_0r0[4:0], L2_0r1[4:0], L2_0a, L153_0r0[31:0], L153_0r1[31:0], L153_0a, L4_0r0[31:0], L4_0r1[31:0], L4_0a, reset);
  tko32m32_1noti0w32b I1 (L14_0r0[31:0], L14_0r1[31:0], L14_0a, L15_0r0[31:0], L15_0r1[31:0], L15_0a, reset);
  tks6_o0w6_0c38m1c3em2c3cm24m2cm34m3co0w0_4mcm14m1co0w0 I2 (L7_0r0[5:0], L7_0r1[5:0], L7_0a, L8_0r, L8_0a, L13_0r, L13_0a, reset);
  tkm2x0b I3 (L11_0r, L11_0a, L16_0r, L16_0a, L17_0r, L17_0a, reset);
  tko0m1_1nm1b0 I4 (L20_0r, L20_0a, L22_0r0, L22_0r1, L22_0a, reset);
  tko0m1_1nm1b1 I5 (L24_0r, L24_0a, L26_0r0, L26_0r1, L26_0a, reset);
  tko1m1_1noti0w1b I6 (L34_0r0, L34_0r1, L34_0a, L35_0r0, L35_0r1, L35_0a, reset);
  tks6_o0w6_0c30m1c3em2c3cm24m28m2cm34m38m3co0w0_4m14o0w0_8m18o0w0_cm1co0w0 I7 (L19_0r0[5:0], L19_0r1[5:0], L19_0a, L20_0r, L20_0a, L24_0r, L24_0a, L28_0r, L28_0a, L33_0r, L33_0a, reset);
  tkm4x0b I8 (L23_0r, L23_0a, L27_0r, L27_0a, L31_0r, L31_0a, L36_0r, L36_0a, L37_0r, L37_0a, reset);
  tkj33m1_32 I9 (L44_0r0, L44_0r1, L44_0a, L46_0r0[31:0], L46_0r1[31:0], L46_0a, L47_0r0[32:0], L47_0r1[32:0], L47_0a, reset);
  tkj33m1_32 I10 (L49_0r0, L49_0r1, L49_0a, L51_0r0[31:0], L51_0r1[31:0], L51_0a, L52_0r0[32:0], L52_0r1[32:0], L52_0a, reset);
  tkj66m33_33 I11 (L47_0r0[32:0], L47_0r1[32:0], L47_0a, L52_0r0[32:0], L52_0r1[32:0], L52_0a, L53_0r0[65:0], L53_0r1[65:0], L53_0a, reset);
  tko66m34_1api0w33b_2api33w33b_3nm1b0_4apt1o0w33bt3o0w1b_5nm1b0_6apt2o0w33bt5o0w1b_7addt4o0w34bt6o0w34b I12 (L53_0r0[65:0], L53_0r1[65:0], L53_0a, L54_0r0[33:0], L54_0r1[33:0], L54_0a, reset);
  tkf34mo1w33 I13 (L54_0r0[33:0], L54_0r1[33:0], L54_0a, L56_0r0[32:0], L56_0r1[32:0], L56_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0 I14 (L55_0r, L55_0a, L43_0r, L43_0a, L45_0r, L45_0a, L48_0r, L48_0a, L50_0r, L50_0a, reset);
  tkj64m32_32 I15 (L59_0r0[31:0], L59_0r1[31:0], L59_0a, L61_0r0[31:0], L61_0r1[31:0], L61_0a, L62_0r0[63:0], L62_0r1[63:0], L62_0a, reset);
  tko64m32_1api0w32b_2api32w32b_3andt1o0w32bt2o0w32b I16 (L62_0r0[63:0], L62_0r1[63:0], L62_0a, L65_0r0[31:0], L65_0r1[31:0], L65_0a, reset);
  tkf0mo0w0_o0w0 I17 (L64_0r, L64_0a, L58_0r, L58_0a, L60_0r, L60_0a, reset);
  tkj64m32_32 I18 (L68_0r0[31:0], L68_0r1[31:0], L68_0a, L70_0r0[31:0], L70_0r1[31:0], L70_0a, L71_0r0[63:0], L71_0r1[63:0], L71_0a, reset);
  tko64m32_1api0w32b_2api32w32b_3ort1o0w32bt2o0w32b I19 (L71_0r0[63:0], L71_0r1[63:0], L71_0a, L74_0r0[31:0], L74_0r1[31:0], L74_0a, reset);
  tkf0mo0w0_o0w0 I20 (L73_0r, L73_0a, L67_0r, L67_0a, L69_0r, L69_0a, reset);
  tkj64m32_32 I21 (L77_0r0[31:0], L77_0r1[31:0], L77_0a, L79_0r0[31:0], L79_0r1[31:0], L79_0a, L80_0r0[63:0], L80_0r1[63:0], L80_0a, reset);
  tko64m32_1api0w32b_2api32w32b_3xort1o0w32bt2o0w32b I22 (L80_0r0[63:0], L80_0r1[63:0], L80_0a, L83_0r0[31:0], L83_0r1[31:0], L83_0a, reset);
  tkf0mo0w0_o0w0 I23 (L82_0r, L82_0a, L76_0r, L76_0a, L78_0r, L78_0a, reset);
  tko0m2_1nm2b0 I24 (L85_0r, L85_0a, L87_0r0[1:0], L87_0r1[1:0], L87_0a, reset);
  tko0m2_1nm2b1 I25 (L89_0r, L89_0a, L91_0r0[1:0], L91_0r1[1:0], L91_0a, reset);
  tko0m1_1nm1b1 I26 (L93_0r, L93_0a, L94_0r0, L94_0r1, L94_0a, reset);
  tkj2m1_1 I27 (L94_0r0, L94_0r1, L94_0a, L96_0r0, L96_0r1, L96_0a, L99_0r0[1:0], L99_0r1[1:0], L99_0a, reset);
  tkf0mo0w0_o0w0 I28 (L98_0r, L98_0a, L93_0r, L93_0a, L95_0r, L95_0a, reset);
  tks6_o0w6_4c20m9c30mac30mbc30mdc30mec30mfc30m20m21m22m23m28m2cm30m31m32m33m34m35m36m37m38m3co0w0_0m8mcm10m14m18m1co0w0_1m5m11m15o0w0_2m6m12m16o0w0_3m7m13m17o0w0_25o0w0_26o0w0_27o0w0 I29 (L40_0r0[5:0], L40_0r1[5:0], L40_0a, L41_0r, L41_0a, L55_0r, L55_0a, L64_0r, L64_0a, L73_0r, L73_0a, L82_0r, L82_0a, L85_0r, L85_0a, L89_0r, L89_0a, L98_0r, L98_0a, reset);
  tkm8x0b I30 (L41_0r, L41_0a, L57_0r, L57_0a, L66_0r, L66_0a, L75_0r, L75_0a, L84_0r, L84_0a, L88_0r, L88_0a, L92_0r, L92_0a, L100_0r, L100_0a, L101_0r, L101_0a, reset);
  tkf0mo0w0_o0w0 I31 (L113_0r, L113_0a, L105_0r, L105_0a, L109_0r, L109_0a, reset);
  tkj0m0_0 I32 (L108_0r, L108_0a, L112_0r, L112_0a, L114_0r, L114_0a, reset);
  tks6_o0w6_0c3cm1c38m2c38m3c38m5m6m7mdc30mec30mfc30m15c20m16c20m17c20o0w0_25m26m27o0w0 I33 (L103_0r0[5:0], L103_0r1[5:0], L103_0a, L104_0r, L104_0a, L113_0r, L113_0a, reset);
  tkm2x0b I34 (L104_0r, L104_0a, L114_0r, L114_0a, L115_0r, L115_0a, reset);
  tkf0mo0w0_o0w0 I35 (L116_0r, L116_0a, L39_0r, L39_0a, L102_0r, L102_0a, reset);
  tkj0m0_0 I36 (L101_0r, L101_0a, L115_0r, L115_0a, L117_0r, L117_0a, reset);
  tkvaddResult33_wo0w33_ro0w33 I37 (L122_0r0[32:0], L122_0r1[32:0], L122_0a, L118_0r, L118_0a, L118_0r, L118_0a, L120_0r0[32:0], L120_0r1[32:0], L120_0a, reset);
  tkf33mo0w0_o0w33 I38 (L125_0r0[32:0], L125_0r1[32:0], L125_0a, L124_0r, L124_0a, L126_0r0[32:0], L126_0r1[32:0], L126_0a, reset);
  tkj33m0_33 I39 (L127_0r, L127_0a, L126_0r0[32:0], L126_0r1[32:0], L126_0a, L122_0r0[32:0], L122_0r1[32:0], L122_0a, reset);
  tko0m1_1nm1b0 I40 (L130_0r, L130_0a, L131_0r0, L131_0r1, L131_0a, reset);
  tkj33m32_1 I41 (L129_0r0[31:0], L129_0r1[31:0], L129_0a, L131_0r0, L131_0r1, L131_0a, L134_0r0[32:0], L134_0r1[32:0], L134_0a, reset);
  tkf0mo0w0_o0w0 I42 (L133_0r, L133_0a, L128_0r, L128_0a, L130_0r, L130_0a, reset);
  tkvlogicResult32_wo0w32_ro0w32 I43 (L136_0r0[31:0], L136_0r1[31:0], L136_0a, L133_0r, L133_0a, L128_0r, L128_0a, L129_0r0[31:0], L129_0r1[31:0], L129_0a, reset);
  tkf32mo0w0_o0w32 I44 (L139_0r0[31:0], L139_0r1[31:0], L139_0a, L138_0r, L138_0a, L140_0r0[31:0], L140_0r1[31:0], L140_0a, reset);
  tkj32m0_32 I45 (L141_0r, L141_0a, L140_0r0[31:0], L140_0r1[31:0], L140_0a, L136_0r0[31:0], L136_0r1[31:0], L136_0a, reset);
  tko0m1_1nm1b0 I46 (L144_0r, L144_0a, L145_0r0, L145_0r1, L145_0a, reset);
  tkj33m32_1 I47 (L143_0r0[31:0], L143_0r1[31:0], L143_0a, L145_0r0, L145_0r1, L145_0a, L148_0r0[32:0], L148_0r1[32:0], L148_0a, reset);
  tkf0mo0w0_o0w0 I48 (L147_0r, L147_0a, L142_0r, L142_0a, L144_0r, L144_0a, reset);
  tkvshiftResult32_wo0w32_ro0w32 I49 (L150_0r0[31:0], L150_0r1[31:0], L150_0a, L147_0r, L147_0a, L142_0r, L142_0a, L143_0r0[31:0], L143_0r1[31:0], L143_0a, reset);
  tkf32mo0w0_o0w32 I50 (L153_0r0[31:0], L153_0r1[31:0], L153_0a, L152_0r, L152_0a, L154_0r0[31:0], L154_0r1[31:0], L154_0a, reset);
  tkj32m0_32 I51 (L155_0r, L155_0a, L154_0r0[31:0], L154_0r1[31:0], L154_0a, L150_0r0[31:0], L150_0r1[31:0], L150_0a, reset);
  tko0m3_1nm3b1 I52 (L124_0r, L124_0a, L157_0r0[2:0], L157_0r1[2:0], L157_0a, reset);
  tko0m3_1nm3b2 I53 (L138_0r, L138_0a, L158_0r0[2:0], L158_0r1[2:0], L158_0a, reset);
  tko0m3_1nm3b4 I54 (L152_0r, L152_0a, L159_0r0[2:0], L159_0r1[2:0], L159_0a, reset);
  tkm3x3b I55 (L157_0r0[2:0], L157_0r1[2:0], L157_0a, L158_0r0[2:0], L158_0r1[2:0], L158_0a, L159_0r0[2:0], L159_0r1[2:0], L159_0a, L160_0r0[2:0], L160_0r1[2:0], L160_0a, reset);
  tkj3m0_3 I56 (L156_0r, L156_0a, L160_0r0[2:0], L160_0r1[2:0], L160_0a, L161_0r0[2:0], L161_0r1[2:0], L161_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_4o0w0 I57 (L161_0r0[2:0], L161_0r1[2:0], L161_0a, L127_0r, L127_0a, L141_0r, L141_0a, L155_0r, L155_0a, reset);
  tkm3x0b I58 (L121_0r, L121_0a, L135_0r, L135_0a, L149_0r, L149_0a, L162_0r, L162_0a, reset);
  tko0m1_1nm1b0 I59 (L170_0r, L170_0a, L171_0r0, L171_0r1, L171_0a, reset);
  tkj33m32_1 I60 (L169_0r0[31:0], L169_0r1[31:0], L169_0a, L171_0r0, L171_0r1, L171_0a, L172_0r0[32:0], L172_0r1[32:0], L172_0a, reset);
  tko33m1_1api0w32b_2api32w1b_3nm31b0_4apt2o0w1bt3o0w31b_5eqt1o0w32bt4o0w32b I61 (L172_0r0[32:0], L172_0r1[32:0], L172_0a, L173_0r0, L173_0r1, L173_0a, reset);
  tkj2m1_1 I62 (L181_0r0, L181_0r1, L181_0a, L183_0r0, L183_0r1, L183_0a, L184_0r0[1:0], L184_0r1[1:0], L184_0a, reset);
  tko2m1_1api0w1b_2api1w1b_3xort1o0w1bt2o0w1b I63 (L184_0r0[1:0], L184_0r1[1:0], L184_0a, L185_0r0, L185_0r1, L185_0a, reset);
  tkj2m1_1 I64 (L179_0r0, L179_0r1, L179_0a, L185_0r0, L185_0r1, L185_0a, L186_0r0[1:0], L186_0r1[1:0], L186_0a, reset);
  tko2m1_1api0w1b_2api1w1b_3xort1o0w1bt2o0w1b I65 (L186_0r0[1:0], L186_0r1[1:0], L186_0a, L187_0r0, L187_0r1, L187_0a, reset);
  tkj2m1_1 I66 (L177_0r0, L177_0r1, L177_0a, L187_0r0, L187_0r1, L187_0a, L188_0r0[1:0], L188_0r1[1:0], L188_0a, reset);
  tko2m1_1api0w1b_2api1w1b_3xort1o0w1bt2o0w1b I67 (L188_0r0[1:0], L188_0r1[1:0], L188_0a, L189_0r0, L189_0r1, L189_0a, reset);
  tko0m6_1nm6b4 I68 (L194_0r, L194_0a, L195_0r0[5:0], L195_0r1[5:0], L195_0a, reset);
  tkj12m6_6 I69 (L193_0r0[5:0], L193_0r1[5:0], L193_0a, L195_0r0[5:0], L195_0r1[5:0], L195_0a, L196_0r0[11:0], L196_0r1[11:0], L196_0a, reset);
  tko12m1_1api0w6b_2api6w6b_3eqt1o0w6bt2o0w6b I70 (L196_0r0[11:0], L196_0r1[11:0], L196_0a, L197_0r0, L197_0r1, L197_0a, reset);
  tkj2m1_1 I71 (L191_0r0, L191_0r1, L191_0a, L197_0r0, L197_0r1, L197_0a, L198_0r0[1:0], L198_0r1[1:0], L198_0a, reset);
  tko2m1_1api0w1b_2api1w1b_3net1o0w1bt2o0w1b I72 (L198_0r0[1:0], L198_0r1[1:0], L198_0a, L199_0r0, L199_0r1, L199_0a, reset);
  tkj4m1_1_1_1 I73 (L173_0r0, L173_0r1, L173_0a, L175_0r0, L175_0r1, L175_0a, L189_0r0, L189_0r1, L189_0a, L199_0r0, L199_0r1, L199_0a, L202_0r0[3:0], L202_0r1[3:0], L202_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 I74 (L201_0r, L201_0a, L168_0r, L168_0a, L170_0r, L170_0a, L174_0r, L174_0a, L176_0r, L176_0a, L178_0r, L178_0a, L180_0r, L180_0a, L182_0r, L182_0a, L190_0r, L190_0a, L192_0r, L192_0a, L194_0r, L194_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I75 (L204_0r, L204_0a, L163_0r, L163_0a, L167_0r, L167_0a, L201_0r, L201_0a, reset);
  tkj0m0_0_0 I76 (L166_0r, L166_0a, L167_0r, L167_0a, L203_0r, L203_0a, L205_0r, L205_0a, reset);
  tkvmergedResult33_wo0w33_ro0w32o0w32o31w1o32w1o31w1o32w1 I77 (L206_0r0[32:0], L206_0r1[32:0], L206_0a, L204_0r, L204_0a, L163_0r, L163_0a, L168_0r, L168_0a, L174_0r, L174_0a, L176_0r, L176_0a, L178_0r, L178_0a, L190_0r, L190_0a, L165_0r0[31:0], L165_0r1[31:0], L165_0a, L169_0r0[31:0], L169_0r1[31:0], L169_0a, L175_0r0, L175_0r1, L175_0a, L177_0r0, L177_0r1, L177_0a, L179_0r0, L179_0r1, L179_0a, L191_0r0, L191_0r1, L191_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I78 (L209_0r, L209_0a, L116_0r, L116_0a, L156_0r, L156_0a, L208_0r, L208_0a, reset);
  tkj0m0_0_0 I79 (L117_0r, L117_0a, L162_0r, L162_0a, L205_0r, L205_0a, L210_0r, L210_0a, reset);
  tkf33mo0w0_o0w33 I80 (L120_0r0[32:0], L120_0r1[32:0], L120_0a, L211_0r, L211_0a, L212_0r0[32:0], L212_0r1[32:0], L212_0a, reset);
  tkf33mo0w0_o0w33 I81 (L134_0r0[32:0], L134_0r1[32:0], L134_0a, L213_0r, L213_0a, L214_0r0[32:0], L214_0r1[32:0], L214_0a, reset);
  tkf33mo0w0_o0w33 I82 (L148_0r0[32:0], L148_0r1[32:0], L148_0a, L215_0r, L215_0a, L216_0r0[32:0], L216_0r1[32:0], L216_0a, reset);
  tkm3x33b I83 (L212_0r0[32:0], L212_0r1[32:0], L212_0a, L214_0r0[32:0], L214_0r1[32:0], L214_0a, L216_0r0[32:0], L216_0r1[32:0], L216_0a, L217_0r0[32:0], L217_0r1[32:0], L217_0a, reset);
  tkf33mo0w0_o0w33 I84 (L217_0r0[32:0], L217_0r1[32:0], L217_0a, L218_0r, L218_0a, L219_0r0[32:0], L219_0r1[32:0], L219_0a, reset);
  tko0m3_1nm3b1 I85 (L211_0r, L211_0a, L220_0r0[2:0], L220_0r1[2:0], L220_0a, reset);
  tko0m3_1nm3b2 I86 (L213_0r, L213_0a, L221_0r0[2:0], L221_0r1[2:0], L221_0a, reset);
  tko0m3_1nm3b4 I87 (L215_0r, L215_0a, L222_0r0[2:0], L222_0r1[2:0], L222_0a, reset);
  tkm3x3b I88 (L220_0r0[2:0], L220_0r1[2:0], L220_0a, L221_0r0[2:0], L221_0r1[2:0], L221_0a, L222_0r0[2:0], L222_0r1[2:0], L222_0a, L223_0r0[2:0], L223_0r1[2:0], L223_0a, reset);
  tkj3m0_3 I89 (L218_0r, L218_0a, L223_0r0[2:0], L223_0r1[2:0], L223_0a, L224_0r0[2:0], L224_0r1[2:0], L224_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_4o0w0 I90 (L224_0r0[2:0], L224_0r1[2:0], L224_0a, L121_0r, L121_0a, L135_0r, L135_0a, L149_0r, L149_0a, reset);
  tkj33m33_0 I91 (L219_0r0[32:0], L219_0r1[32:0], L219_0a, L208_0r, L208_0a, L206_0r0[32:0], L206_0r1[32:0], L206_0a, reset);
  tkf33mo0w0_o0w33 I92 (L56_0r0[32:0], L56_0r1[32:0], L56_0a, L57_0r, L57_0a, L125_0r0[32:0], L125_0r1[32:0], L125_0a, reset);
  tkf32mo0w0_o0w32 I93 (L65_0r0[31:0], L65_0r1[31:0], L65_0a, L226_0r, L226_0a, L227_0r0[31:0], L227_0r1[31:0], L227_0a, reset);
  tkf32mo0w0_o0w32 I94 (L74_0r0[31:0], L74_0r1[31:0], L74_0a, L228_0r, L228_0a, L229_0r0[31:0], L229_0r1[31:0], L229_0a, reset);
  tkf32mo0w0_o0w32 I95 (L83_0r0[31:0], L83_0r1[31:0], L83_0a, L230_0r, L230_0a, L231_0r0[31:0], L231_0r1[31:0], L231_0a, reset);
  tkm3x32b I96 (L227_0r0[31:0], L227_0r1[31:0], L227_0a, L229_0r0[31:0], L229_0r1[31:0], L229_0a, L231_0r0[31:0], L231_0r1[31:0], L231_0a, L232_0r0[31:0], L232_0r1[31:0], L232_0a, reset);
  tkf32mo0w0_o0w32 I97 (L232_0r0[31:0], L232_0r1[31:0], L232_0a, L233_0r, L233_0a, L139_0r0[31:0], L139_0r1[31:0], L139_0a, reset);
  tko0m3_1nm3b1 I98 (L226_0r, L226_0a, L235_0r0[2:0], L235_0r1[2:0], L235_0a, reset);
  tko0m3_1nm3b2 I99 (L228_0r, L228_0a, L236_0r0[2:0], L236_0r1[2:0], L236_0a, reset);
  tko0m3_1nm3b4 I100 (L230_0r, L230_0a, L237_0r0[2:0], L237_0r1[2:0], L237_0a, reset);
  tkm3x3b I101 (L235_0r0[2:0], L235_0r1[2:0], L235_0a, L236_0r0[2:0], L236_0r1[2:0], L236_0a, L237_0r0[2:0], L237_0r1[2:0], L237_0a, L238_0r0[2:0], L238_0r1[2:0], L238_0a, reset);
  tkj3m0_3 I102 (L233_0r, L233_0a, L238_0r0[2:0], L238_0r1[2:0], L238_0a, L239_0r0[2:0], L239_0r1[2:0], L239_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_4o0w0 I103 (L239_0r0[2:0], L239_0r1[2:0], L239_0a, L66_0r, L66_0a, L75_0r, L75_0a, L84_0r, L84_0a, reset);
  tkvpostRhs32_wo0w32_ro0w32o31w1o0w5o31w1 I104 (L240_0r0[31:0], L240_0r1[31:0], L240_0a, L241_0r, L241_0a, L50_0r, L50_0a, L95_0r, L95_0a, L105_0r, L105_0a, L182_0r, L182_0a, L51_0r0[31:0], L51_0r1[31:0], L51_0a, L96_0r0, L96_0r1, L96_0a, L107_0r0[4:0], L107_0r1[4:0], L107_0a, L183_0r0, L183_0r1, L183_0a, reset);
  tkvaddCarryIn1_wo0w1_ro0w1o0w1 I105 (L242_0r0, L242_0r1, L242_0a, L243_0r, L243_0a, L43_0r, L43_0a, L48_0r, L48_0a, L44_0r0, L44_0r1, L44_0a, L49_0r0, L49_0r1, L49_0a, reset);
  tkj0m0_0 I106 (L241_0r, L241_0a, L243_0r, L243_0a, L209_0r, L209_0a, reset);
  tkf0mo0w0_o0w0 I107 (L247_0r, L247_0a, L245_0r, L245_0a, L246_0r, L246_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I108 (L248_0r, L248_0a, L6_0r, L6_0a, L18_0r, L18_0a, L247_0r, L247_0a, reset);
  tkj0m0_0_0 I109 (L17_0r, L17_0a, L37_0r, L37_0a, L210_0r, L210_0a, L249_0r, L249_0a, reset);
  tkvop7_wo0w7_ro0w6o0w6o6w1o6w1o0w6o0w6o0w6 I110 (L250_0r0[6:0], L250_0r1[6:0], L250_0a, L251_0r, L251_0a, L6_0r, L6_0a, L18_0r, L18_0a, L28_0r, L28_0a, L33_0r, L33_0a, L39_0r, L39_0a, L102_0r, L102_0a, L192_0r, L192_0a, L7_0r0[5:0], L7_0r1[5:0], L7_0a, L19_0r0[5:0], L19_0r1[5:0], L19_0a, L30_0r0, L30_0r1, L30_0a, L34_0r0, L34_0r1, L34_0a, L40_0r0[5:0], L40_0r1[5:0], L40_0a, L103_0r0[5:0], L103_0r1[5:0], L103_0a, L193_0r0[5:0], L193_0r1[5:0], L193_0a, reset);
  tkvlhs32_wo0w32_ro0w32o0w32o0w32o0w32o0w32o31w1 I111 (L252_0r0[31:0], L252_0r1[31:0], L252_0a, L253_0r, L253_0a, L45_0r, L45_0a, L58_0r, L58_0a, L67_0r, L67_0a, L76_0r, L76_0a, L109_0r, L109_0a, L180_0r, L180_0a, L46_0r0[31:0], L46_0r1[31:0], L46_0a, L59_0r0[31:0], L59_0r1[31:0], L59_0a, L68_0r0[31:0], L68_0r1[31:0], L68_0a, L77_0r0[31:0], L77_0r1[31:0], L77_0a, L111_0r0[31:0], L111_0r1[31:0], L111_0a, L181_0r0, L181_0r1, L181_0a, reset);
  tkvrhs32_wo0w32_ro0w32o0w32o0w32o0w32o0w32 I112 (L254_0r0[31:0], L254_0r1[31:0], L254_0a, L255_0r, L255_0a, L8_0r, L8_0a, L13_0r, L13_0a, L60_0r, L60_0a, L69_0r, L69_0a, L78_0r, L78_0a, L10_0r0[31:0], L10_0r1[31:0], L10_0a, L14_0r0[31:0], L14_0r1[31:0], L14_0a, L61_0r0[31:0], L61_0r1[31:0], L61_0a, L70_0r0[31:0], L70_0r1[31:0], L70_0a, L79_0r0[31:0], L79_0r1[31:0], L79_0a, reset);
  tkj0m0_0_0 I113 (L251_0r, L251_0a, L253_0r, L253_0a, L255_0r, L255_0a, L248_0r, L248_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I114 (L260_0r, L260_0a, L257_0r, L257_0a, L258_0r, L258_0a, L259_0r, L259_0a, reset);
  tkf32mo0w0_o0w32 I115 (L111_0r0[31:0], L111_0r1[31:0], L111_0a, L112_0r, L112_0a, L4_0r0[31:0], L4_0r1[31:0], L4_0a, reset);
  tkf5mo0w0_o0w5 I116 (L107_0r0[4:0], L107_0r1[4:0], L107_0a, L108_0r, L108_0a, L2_0r0[4:0], L2_0r1[4:0], L2_0a, reset);
  tkf2mo0w0_o0w2 I117 (L87_0r0[1:0], L87_0r1[1:0], L87_0a, L265_0r, L265_0a, L266_0r0[1:0], L266_0r1[1:0], L266_0a, reset);
  tkf2mo0w0_o0w2 I118 (L91_0r0[1:0], L91_0r1[1:0], L91_0a, L267_0r, L267_0a, L268_0r0[1:0], L268_0r1[1:0], L268_0a, reset);
  tkf2mo0w0_o0w2 I119 (L99_0r0[1:0], L99_0r1[1:0], L99_0a, L269_0r, L269_0a, L270_0r0[1:0], L270_0r1[1:0], L270_0a, reset);
  tkm3x2b I120 (L266_0r0[1:0], L266_0r1[1:0], L266_0a, L268_0r0[1:0], L268_0r1[1:0], L268_0a, L270_0r0[1:0], L270_0r1[1:0], L270_0a, L271_0r0[1:0], L271_0r1[1:0], L271_0a, reset);
  tkf2mo0w0_o0w2 I121 (L271_0r0[1:0], L271_0r1[1:0], L271_0a, L272_0r, L272_0a, L1_0r0[1:0], L1_0r1[1:0], L1_0a, reset);
  tko0m3_1nm3b1 I122 (L265_0r, L265_0a, L274_0r0[2:0], L274_0r1[2:0], L274_0a, reset);
  tko0m3_1nm3b2 I123 (L267_0r, L267_0a, L275_0r0[2:0], L275_0r1[2:0], L275_0a, reset);
  tko0m3_1nm3b4 I124 (L269_0r, L269_0a, L276_0r0[2:0], L276_0r1[2:0], L276_0a, reset);
  tkm3x3b I125 (L274_0r0[2:0], L274_0r1[2:0], L274_0a, L275_0r0[2:0], L275_0r1[2:0], L275_0a, L276_0r0[2:0], L276_0r1[2:0], L276_0a, L277_0r0[2:0], L277_0r1[2:0], L277_0a, reset);
  tkj3m0_3 I126 (L272_0r, L272_0a, L277_0r0[2:0], L277_0r1[2:0], L277_0a, L278_0r0[2:0], L278_0r1[2:0], L278_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_4o0w0 I127 (L278_0r0[2:0], L278_0r1[2:0], L278_0a, L88_0r, L88_0a, L92_0r, L92_0a, L100_0r, L100_0a, reset);
  tkf1mo0w0_o0w1 I128 (L22_0r0, L22_0r1, L22_0a, L279_0r, L279_0a, L280_0r0, L280_0r1, L280_0a, reset);
  tkf1mo0w0_o0w1 I129 (L26_0r0, L26_0r1, L26_0a, L281_0r, L281_0a, L282_0r0, L282_0r1, L282_0a, reset);
  tkf1mo0w0_o0w1 I130 (L30_0r0, L30_0r1, L30_0a, L283_0r, L283_0a, L284_0r0, L284_0r1, L284_0a, reset);
  tkf1mo0w0_o0w1 I131 (L35_0r0, L35_0r1, L35_0a, L285_0r, L285_0a, L286_0r0, L286_0r1, L286_0a, reset);
  tkm4x1b I132 (L280_0r0, L280_0r1, L280_0a, L282_0r0, L282_0r1, L282_0a, L284_0r0, L284_0r1, L284_0a, L286_0r0, L286_0r1, L286_0a, L287_0r0, L287_0r1, L287_0a, reset);
  tkf1mo0w0_o0w1 I133 (L287_0r0, L287_0r1, L287_0a, L288_0r, L288_0a, L289_0r0, L289_0r1, L289_0a, reset);
  tko0m4_1nm4b1 I134 (L279_0r, L279_0a, L290_0r0[3:0], L290_0r1[3:0], L290_0a, reset);
  tko0m4_1nm4b2 I135 (L281_0r, L281_0a, L291_0r0[3:0], L291_0r1[3:0], L291_0a, reset);
  tko0m4_1nm4b4 I136 (L283_0r, L283_0a, L292_0r0[3:0], L292_0r1[3:0], L292_0a, reset);
  tko0m4_1nm4b8 I137 (L285_0r, L285_0a, L293_0r0[3:0], L293_0r1[3:0], L293_0a, reset);
  tkm4x4b I138 (L290_0r0[3:0], L290_0r1[3:0], L290_0a, L291_0r0[3:0], L291_0r1[3:0], L291_0a, L292_0r0[3:0], L292_0r1[3:0], L292_0a, L293_0r0[3:0], L293_0r1[3:0], L293_0a, L294_0r0[3:0], L294_0r1[3:0], L294_0a, reset);
  tkj4m0_4 I139 (L288_0r, L288_0a, L294_0r0[3:0], L294_0r1[3:0], L294_0a, L295_0r0[3:0], L295_0r1[3:0], L295_0a, reset);
  tks4_o0w4_1o0w0_2o0w0_4o0w0_8o0w0 I140 (L295_0r0[3:0], L295_0r1[3:0], L295_0a, L23_0r, L23_0a, L27_0r, L27_0a, L31_0r, L31_0a, L36_0r, L36_0a, reset);
  tkj1m1_0 I141 (L289_0r0, L289_0r1, L289_0a, L246_0r, L246_0a, L242_0r0, L242_0r1, L242_0a, reset);
  tkf32mo0w0_o0w32 I142 (L10_0r0[31:0], L10_0r1[31:0], L10_0a, L296_0r, L296_0a, L297_0r0[31:0], L297_0r1[31:0], L297_0a, reset);
  tkf32mo0w0_o0w32 I143 (L15_0r0[31:0], L15_0r1[31:0], L15_0a, L298_0r, L298_0a, L299_0r0[31:0], L299_0r1[31:0], L299_0a, reset);
  tkm2x32b I144 (L297_0r0[31:0], L297_0r1[31:0], L297_0a, L299_0r0[31:0], L299_0r1[31:0], L299_0a, L300_0r0[31:0], L300_0r1[31:0], L300_0a, reset);
  tkf32mo0w0_o0w32 I145 (L300_0r0[31:0], L300_0r1[31:0], L300_0a, L301_0r, L301_0a, L302_0r0[31:0], L302_0r1[31:0], L302_0a, reset);
  tko0m2_1nm2b1 I146 (L296_0r, L296_0a, L303_0r0[1:0], L303_0r1[1:0], L303_0a, reset);
  tko0m2_1nm2b2 I147 (L298_0r, L298_0a, L304_0r0[1:0], L304_0r1[1:0], L304_0a, reset);
  tkm2x2b I148 (L303_0r0[1:0], L303_0r1[1:0], L303_0a, L304_0r0[1:0], L304_0r1[1:0], L304_0a, L305_0r0[1:0], L305_0r1[1:0], L305_0a, reset);
  tkj2m0_2 I149 (L301_0r, L301_0a, L305_0r0[1:0], L305_0r1[1:0], L305_0a, L306_0r0[1:0], L306_0r1[1:0], L306_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I150 (L306_0r0[1:0], L306_0r1[1:0], L306_0a, L11_0r, L11_0a, L16_0r, L16_0a, reset);
  tkj32m32_0 I151 (L302_0r0[31:0], L302_0r1[31:0], L302_0a, L245_0r, L245_0a, L240_0r0[31:0], L240_0r1[31:0], L240_0a, reset);
  tkj7m7_0 I152 (op_0r0[6:0], op_0r1[6:0], op_0a, L257_0r, L257_0a, L250_0r0[6:0], L250_0r1[6:0], L250_0a, reset);
  tkf32mo0w0_o0w32 I153 (L165_0r0[31:0], L165_0r1[31:0], L165_0a, L166_0r, L166_0a, result_0r0[31:0], result_0r1[31:0], result_0a, reset);
  tkf4mo0w0_o0w4 I154 (L202_0r0[3:0], L202_0r1[3:0], L202_0a, L203_0r, L203_0a, flags_0r0[3:0], flags_0r1[3:0], flags_0a, reset);
  tkj32m32_0 I155 (lhs_0r0[31:0], lhs_0r1[31:0], lhs_0a, L258_0r, L258_0a, L252_0r0[31:0], L252_0r1[31:0], L252_0a, reset);
  tkj32m32_0 I156 (rhs_0r0[31:0], rhs_0r1[31:0], rhs_0a, L259_0r, L259_0a, L254_0r0[31:0], L254_0r1[31:0], L254_0a, reset);
  tki I157 (L249_0r, L249_0a, L260_0r, L260_0a, reset);
endmodule

module teak_RegBank (wEn_0r0, wEn_0r1, wEn_0a, rEn_0r0, rEn_0r1, rEn_0a, wSel_0r0, wSel_0r1, wSel_0a, r0Sel_0r0, r0Sel_0r1, r0Sel_0a, r1Sel_0r0, r1Sel_0r1, r1Sel_0a, r2Sel_0r0, r2Sel_0r1, r2Sel_0a, window_0r0, window_0r1, window_0a, w_0r0, w_0r1, w_0a, r0_0r0, r0_0r1, r0_0a, r1_0r0, r1_0r1, r1_0a, r2_0r0, r2_0r1, r2_0a, reset);
  input wEn_0r0;
  input wEn_0r1;
  output wEn_0a;
  input [2:0] rEn_0r0;
  input [2:0] rEn_0r1;
  output rEn_0a;
  input [4:0] wSel_0r0;
  input [4:0] wSel_0r1;
  output wSel_0a;
  input [4:0] r0Sel_0r0;
  input [4:0] r0Sel_0r1;
  output r0Sel_0a;
  input [4:0] r1Sel_0r0;
  input [4:0] r1Sel_0r1;
  output r1Sel_0a;
  input [4:0] r2Sel_0r0;
  input [4:0] r2Sel_0r1;
  output r2Sel_0a;
  input window_0r0;
  input window_0r1;
  output window_0a;
  input [31:0] w_0r0;
  input [31:0] w_0r1;
  output w_0a;
  output [31:0] r0_0r0;
  output [31:0] r0_0r1;
  input r0_0a;
  output [31:0] r1_0r0;
  output [31:0] r1_0r1;
  input r1_0a;
  output [31:0] r2_0r0;
  output [31:0] r2_0r1;
  input r2_0a;
  input reset;
  wire L2_0r;
  wire L2_0a;
  wire L3_0r0;
  wire L3_0r1;
  wire L3_0a;
  wire L4_0r;
  wire L4_0a;
  wire L5_0r;
  wire L5_0a;
  wire [4:0] L6_0r0;
  wire [4:0] L6_0r1;
  wire L6_0a;
  wire L7_0r;
  wire L7_0a;
  wire [31:0] L9_0r0;
  wire [31:0] L9_0r1;
  wire L9_0a;
  wire L10_0r;
  wire L10_0a;
  wire L11_0r;
  wire L11_0a;
  wire [31:0] L12_0r0;
  wire [31:0] L12_0r1;
  wire L12_0a;
  wire L13_0r;
  wire L13_0a;
  wire [31:0] L14_0r0;
  wire [31:0] L14_0r1;
  wire L14_0a;
  wire L15_0r;
  wire L15_0a;
  wire [31:0] L16_0r0;
  wire [31:0] L16_0r1;
  wire L16_0a;
  wire L17_0r;
  wire L17_0a;
  wire [31:0] L18_0r0;
  wire [31:0] L18_0r1;
  wire L18_0a;
  wire L19_0r;
  wire L19_0a;
  wire [31:0] L20_0r0;
  wire [31:0] L20_0r1;
  wire L20_0a;
  wire L21_0r;
  wire L21_0a;
  wire [31:0] L22_0r0;
  wire [31:0] L22_0r1;
  wire L22_0a;
  wire L23_0r;
  wire L23_0a;
  wire [31:0] L24_0r0;
  wire [31:0] L24_0r1;
  wire L24_0a;
  wire L25_0r;
  wire L25_0a;
  wire [2:0] L26_0r0;
  wire [2:0] L26_0r1;
  wire L26_0a;
  wire [31:0] L28_0r0;
  wire [31:0] L28_0r1;
  wire L28_0a;
  wire L29_0r;
  wire L29_0a;
  wire L30_0r;
  wire L30_0a;
  wire [31:0] L31_0r0;
  wire [31:0] L31_0r1;
  wire L31_0a;
  wire L32_0r;
  wire L32_0a;
  wire [31:0] L33_0r0;
  wire [31:0] L33_0r1;
  wire L33_0a;
  wire L34_0r;
  wire L34_0a;
  wire [31:0] L35_0r0;
  wire [31:0] L35_0r1;
  wire L35_0a;
  wire L36_0r;
  wire L36_0a;
  wire [31:0] L37_0r0;
  wire [31:0] L37_0r1;
  wire L37_0a;
  wire L38_0r;
  wire L38_0a;
  wire [31:0] L39_0r0;
  wire [31:0] L39_0r1;
  wire L39_0a;
  wire L40_0r;
  wire L40_0a;
  wire [31:0] L41_0r0;
  wire [31:0] L41_0r1;
  wire L41_0a;
  wire L42_0r;
  wire L42_0a;
  wire [31:0] L43_0r0;
  wire [31:0] L43_0r1;
  wire L43_0a;
  wire L44_0r;
  wire L44_0a;
  wire [31:0] L45_0r0;
  wire [31:0] L45_0r1;
  wire L45_0a;
  wire [2:0] L46_0r0;
  wire [2:0] L46_0r1;
  wire L46_0a;
  wire L47_0r;
  wire L47_0a;
  wire [2:0] L48_0r0;
  wire [2:0] L48_0r1;
  wire L48_0a;
  wire L49_0r;
  wire L49_0a;
  wire L50_0r0;
  wire L50_0r1;
  wire L50_0a;
  wire [3:0] L51_0r0;
  wire [3:0] L51_0r1;
  wire L51_0a;
  wire L53_0r;
  wire L53_0a;
  wire [31:0] L54_0r0;
  wire [31:0] L54_0r1;
  wire L54_0a;
  wire L55_0r;
  wire L55_0a;
  wire L56_0r;
  wire L56_0a;
  wire [31:0] L57_0r0;
  wire [31:0] L57_0r1;
  wire L57_0a;
  wire L58_0r;
  wire L58_0a;
  wire [31:0] L59_0r0;
  wire [31:0] L59_0r1;
  wire L59_0a;
  wire L60_0r;
  wire L60_0a;
  wire [31:0] L61_0r0;
  wire [31:0] L61_0r1;
  wire L61_0a;
  wire L62_0r;
  wire L62_0a;
  wire [31:0] L63_0r0;
  wire [31:0] L63_0r1;
  wire L63_0a;
  wire L64_0r;
  wire L64_0a;
  wire [31:0] L65_0r0;
  wire [31:0] L65_0r1;
  wire L65_0a;
  wire L66_0r;
  wire L66_0a;
  wire [31:0] L67_0r0;
  wire [31:0] L67_0r1;
  wire L67_0a;
  wire L68_0r;
  wire L68_0a;
  wire [31:0] L69_0r0;
  wire [31:0] L69_0r1;
  wire L69_0a;
  wire L70_0r;
  wire L70_0a;
  wire [31:0] L71_0r0;
  wire [31:0] L71_0r1;
  wire L71_0a;
  wire [2:0] L72_0r0;
  wire [2:0] L72_0r1;
  wire L72_0a;
  wire L73_0r;
  wire L73_0a;
  wire [2:0] L74_0r0;
  wire [2:0] L74_0r1;
  wire L74_0a;
  wire L75_0r;
  wire L75_0a;
  wire L76_0r0;
  wire L76_0r1;
  wire L76_0a;
  wire [3:0] L77_0r0;
  wire [3:0] L77_0r1;
  wire L77_0a;
  wire L79_0r;
  wire L79_0a;
  wire [31:0] L80_0r0;
  wire [31:0] L80_0r1;
  wire L80_0a;
  wire L81_0r;
  wire L81_0a;
  wire L82_0r;
  wire L82_0a;
  wire [31:0] L83_0r0;
  wire [31:0] L83_0r1;
  wire L83_0a;
  wire L84_0r;
  wire L84_0a;
  wire [31:0] L85_0r0;
  wire [31:0] L85_0r1;
  wire L85_0a;
  wire L86_0r;
  wire L86_0a;
  wire [31:0] L87_0r0;
  wire [31:0] L87_0r1;
  wire L87_0a;
  wire L88_0r;
  wire L88_0a;
  wire [31:0] L89_0r0;
  wire [31:0] L89_0r1;
  wire L89_0a;
  wire L90_0r;
  wire L90_0a;
  wire [31:0] L91_0r0;
  wire [31:0] L91_0r1;
  wire L91_0a;
  wire L92_0r;
  wire L92_0a;
  wire [31:0] L93_0r0;
  wire [31:0] L93_0r1;
  wire L93_0a;
  wire L94_0r;
  wire L94_0a;
  wire [31:0] L95_0r0;
  wire [31:0] L95_0r1;
  wire L95_0a;
  wire L96_0r;
  wire L96_0a;
  wire [31:0] L97_0r0;
  wire [31:0] L97_0r1;
  wire L97_0a;
  wire [2:0] L98_0r0;
  wire [2:0] L98_0r1;
  wire L98_0a;
  wire L99_0r;
  wire L99_0a;
  wire [2:0] L100_0r0;
  wire [2:0] L100_0r1;
  wire L100_0a;
  wire L101_0r0;
  wire L101_0r1;
  wire L101_0a;
  wire L102_0r;
  wire L102_0a;
  wire L103_0r0;
  wire L103_0r1;
  wire L103_0a;
  wire L104_0r;
  wire L104_0a;
  wire L105_0r0;
  wire L105_0r1;
  wire L105_0a;
  wire [1:0] L106_0r0;
  wire [1:0] L106_0r1;
  wire L106_0a;
  wire [1:0] L107_0r0;
  wire [1:0] L107_0r1;
  wire L107_0a;
  wire [3:0] L108_0r0;
  wire [3:0] L108_0r1;
  wire L108_0a;
  wire L110_0r;
  wire L110_0a;
  wire [31:0] L111_0r0;
  wire [31:0] L111_0r1;
  wire L111_0a;
  wire L112_0r;
  wire L112_0a;
  wire L113_0r;
  wire L113_0a;
  wire [4:0] L114_0r0;
  wire [4:0] L114_0r1;
  wire L114_0a;
  wire L116_0r;
  wire L116_0a;
  wire L117_0r;
  wire L117_0a;
  wire L118_0r;
  wire L118_0a;
  wire L119_0r0;
  wire L119_0r1;
  wire L119_0a;
  wire L120_0r;
  wire L120_0a;
  wire L121_0r;
  wire L121_0a;
  wire [4:0] L122_0r0;
  wire [4:0] L122_0r1;
  wire L122_0a;
  wire L123_0r;
  wire L123_0a;
  wire [31:0] L125_0r0;
  wire [31:0] L125_0r1;
  wire L125_0a;
  wire L126_0r;
  wire L126_0a;
  wire L127_0r;
  wire L127_0a;
  wire [31:0] L128_0r0;
  wire [31:0] L128_0r1;
  wire L128_0a;
  wire L129_0r;
  wire L129_0a;
  wire [31:0] L130_0r0;
  wire [31:0] L130_0r1;
  wire L130_0a;
  wire L131_0r;
  wire L131_0a;
  wire [31:0] L132_0r0;
  wire [31:0] L132_0r1;
  wire L132_0a;
  wire L133_0r;
  wire L133_0a;
  wire [31:0] L134_0r0;
  wire [31:0] L134_0r1;
  wire L134_0a;
  wire L135_0r;
  wire L135_0a;
  wire [31:0] L136_0r0;
  wire [31:0] L136_0r1;
  wire L136_0a;
  wire L137_0r;
  wire L137_0a;
  wire [31:0] L138_0r0;
  wire [31:0] L138_0r1;
  wire L138_0a;
  wire L139_0r;
  wire L139_0a;
  wire [31:0] L140_0r0;
  wire [31:0] L140_0r1;
  wire L140_0a;
  wire L141_0r;
  wire L141_0a;
  wire [2:0] L142_0r0;
  wire [2:0] L142_0r1;
  wire L142_0a;
  wire [31:0] L144_0r0;
  wire [31:0] L144_0r1;
  wire L144_0a;
  wire L145_0r;
  wire L145_0a;
  wire L146_0r;
  wire L146_0a;
  wire [31:0] L147_0r0;
  wire [31:0] L147_0r1;
  wire L147_0a;
  wire L148_0r;
  wire L148_0a;
  wire [31:0] L149_0r0;
  wire [31:0] L149_0r1;
  wire L149_0a;
  wire L150_0r;
  wire L150_0a;
  wire [31:0] L151_0r0;
  wire [31:0] L151_0r1;
  wire L151_0a;
  wire L152_0r;
  wire L152_0a;
  wire [31:0] L153_0r0;
  wire [31:0] L153_0r1;
  wire L153_0a;
  wire L154_0r;
  wire L154_0a;
  wire [31:0] L155_0r0;
  wire [31:0] L155_0r1;
  wire L155_0a;
  wire L156_0r;
  wire L156_0a;
  wire [31:0] L157_0r0;
  wire [31:0] L157_0r1;
  wire L157_0a;
  wire L158_0r;
  wire L158_0a;
  wire [31:0] L159_0r0;
  wire [31:0] L159_0r1;
  wire L159_0a;
  wire L160_0r;
  wire L160_0a;
  wire [31:0] L161_0r0;
  wire [31:0] L161_0r1;
  wire L161_0a;
  wire [2:0] L162_0r0;
  wire [2:0] L162_0r1;
  wire L162_0a;
  wire L163_0r;
  wire L163_0a;
  wire [2:0] L164_0r0;
  wire [2:0] L164_0r1;
  wire L164_0a;
  wire L165_0r;
  wire L165_0a;
  wire L166_0r0;
  wire L166_0r1;
  wire L166_0a;
  wire [3:0] L167_0r0;
  wire [3:0] L167_0r1;
  wire L167_0a;
  wire L169_0r;
  wire L169_0a;
  wire [31:0] L170_0r0;
  wire [31:0] L170_0r1;
  wire L170_0a;
  wire L171_0r;
  wire L171_0a;
  wire L172_0r;
  wire L172_0a;
  wire [31:0] L173_0r0;
  wire [31:0] L173_0r1;
  wire L173_0a;
  wire L174_0r;
  wire L174_0a;
  wire [31:0] L175_0r0;
  wire [31:0] L175_0r1;
  wire L175_0a;
  wire L176_0r;
  wire L176_0a;
  wire [31:0] L177_0r0;
  wire [31:0] L177_0r1;
  wire L177_0a;
  wire L178_0r;
  wire L178_0a;
  wire [31:0] L179_0r0;
  wire [31:0] L179_0r1;
  wire L179_0a;
  wire L180_0r;
  wire L180_0a;
  wire [31:0] L181_0r0;
  wire [31:0] L181_0r1;
  wire L181_0a;
  wire L182_0r;
  wire L182_0a;
  wire [31:0] L183_0r0;
  wire [31:0] L183_0r1;
  wire L183_0a;
  wire L184_0r;
  wire L184_0a;
  wire [31:0] L185_0r0;
  wire [31:0] L185_0r1;
  wire L185_0a;
  wire L186_0r;
  wire L186_0a;
  wire [31:0] L187_0r0;
  wire [31:0] L187_0r1;
  wire L187_0a;
  wire [2:0] L188_0r0;
  wire [2:0] L188_0r1;
  wire L188_0a;
  wire L189_0r;
  wire L189_0a;
  wire [2:0] L190_0r0;
  wire [2:0] L190_0r1;
  wire L190_0a;
  wire L191_0r;
  wire L191_0a;
  wire L192_0r0;
  wire L192_0r1;
  wire L192_0a;
  wire [3:0] L193_0r0;
  wire [3:0] L193_0r1;
  wire L193_0a;
  wire L195_0r;
  wire L195_0a;
  wire [31:0] L196_0r0;
  wire [31:0] L196_0r1;
  wire L196_0a;
  wire L197_0r;
  wire L197_0a;
  wire L198_0r;
  wire L198_0a;
  wire [31:0] L199_0r0;
  wire [31:0] L199_0r1;
  wire L199_0a;
  wire L200_0r;
  wire L200_0a;
  wire [31:0] L201_0r0;
  wire [31:0] L201_0r1;
  wire L201_0a;
  wire L202_0r;
  wire L202_0a;
  wire [31:0] L203_0r0;
  wire [31:0] L203_0r1;
  wire L203_0a;
  wire L204_0r;
  wire L204_0a;
  wire [31:0] L205_0r0;
  wire [31:0] L205_0r1;
  wire L205_0a;
  wire L206_0r;
  wire L206_0a;
  wire [31:0] L207_0r0;
  wire [31:0] L207_0r1;
  wire L207_0a;
  wire L208_0r;
  wire L208_0a;
  wire [31:0] L209_0r0;
  wire [31:0] L209_0r1;
  wire L209_0a;
  wire L210_0r;
  wire L210_0a;
  wire [31:0] L211_0r0;
  wire [31:0] L211_0r1;
  wire L211_0a;
  wire L212_0r;
  wire L212_0a;
  wire [31:0] L213_0r0;
  wire [31:0] L213_0r1;
  wire L213_0a;
  wire [2:0] L214_0r0;
  wire [2:0] L214_0r1;
  wire L214_0a;
  wire L215_0r;
  wire L215_0a;
  wire [2:0] L216_0r0;
  wire [2:0] L216_0r1;
  wire L216_0a;
  wire L217_0r0;
  wire L217_0r1;
  wire L217_0a;
  wire L218_0r;
  wire L218_0a;
  wire L219_0r0;
  wire L219_0r1;
  wire L219_0a;
  wire L220_0r;
  wire L220_0a;
  wire L221_0r0;
  wire L221_0r1;
  wire L221_0a;
  wire [1:0] L222_0r0;
  wire [1:0] L222_0r1;
  wire L222_0a;
  wire [1:0] L223_0r0;
  wire [1:0] L223_0r1;
  wire L223_0a;
  wire [3:0] L224_0r0;
  wire [3:0] L224_0r1;
  wire L224_0a;
  wire L226_0r;
  wire L226_0a;
  wire [31:0] L227_0r0;
  wire [31:0] L227_0r1;
  wire L227_0a;
  wire L228_0r;
  wire L228_0a;
  wire L229_0r;
  wire L229_0a;
  wire [4:0] L230_0r0;
  wire [4:0] L230_0r1;
  wire L230_0a;
  wire L232_0r;
  wire L232_0a;
  wire L233_0r;
  wire L233_0a;
  wire L234_0r;
  wire L234_0a;
  wire L235_0r0;
  wire L235_0r1;
  wire L235_0a;
  wire L236_0r;
  wire L236_0a;
  wire L237_0r;
  wire L237_0a;
  wire [4:0] L238_0r0;
  wire [4:0] L238_0r1;
  wire L238_0a;
  wire L239_0r;
  wire L239_0a;
  wire [31:0] L241_0r0;
  wire [31:0] L241_0r1;
  wire L241_0a;
  wire L242_0r;
  wire L242_0a;
  wire L243_0r;
  wire L243_0a;
  wire [31:0] L244_0r0;
  wire [31:0] L244_0r1;
  wire L244_0a;
  wire L245_0r;
  wire L245_0a;
  wire [31:0] L246_0r0;
  wire [31:0] L246_0r1;
  wire L246_0a;
  wire L247_0r;
  wire L247_0a;
  wire [31:0] L248_0r0;
  wire [31:0] L248_0r1;
  wire L248_0a;
  wire L249_0r;
  wire L249_0a;
  wire [31:0] L250_0r0;
  wire [31:0] L250_0r1;
  wire L250_0a;
  wire L251_0r;
  wire L251_0a;
  wire [31:0] L252_0r0;
  wire [31:0] L252_0r1;
  wire L252_0a;
  wire L253_0r;
  wire L253_0a;
  wire [31:0] L254_0r0;
  wire [31:0] L254_0r1;
  wire L254_0a;
  wire L255_0r;
  wire L255_0a;
  wire [31:0] L256_0r0;
  wire [31:0] L256_0r1;
  wire L256_0a;
  wire L257_0r;
  wire L257_0a;
  wire [2:0] L258_0r0;
  wire [2:0] L258_0r1;
  wire L258_0a;
  wire [31:0] L260_0r0;
  wire [31:0] L260_0r1;
  wire L260_0a;
  wire L261_0r;
  wire L261_0a;
  wire L262_0r;
  wire L262_0a;
  wire [31:0] L263_0r0;
  wire [31:0] L263_0r1;
  wire L263_0a;
  wire L264_0r;
  wire L264_0a;
  wire [31:0] L265_0r0;
  wire [31:0] L265_0r1;
  wire L265_0a;
  wire L266_0r;
  wire L266_0a;
  wire [31:0] L267_0r0;
  wire [31:0] L267_0r1;
  wire L267_0a;
  wire L268_0r;
  wire L268_0a;
  wire [31:0] L269_0r0;
  wire [31:0] L269_0r1;
  wire L269_0a;
  wire L270_0r;
  wire L270_0a;
  wire [31:0] L271_0r0;
  wire [31:0] L271_0r1;
  wire L271_0a;
  wire L272_0r;
  wire L272_0a;
  wire [31:0] L273_0r0;
  wire [31:0] L273_0r1;
  wire L273_0a;
  wire L274_0r;
  wire L274_0a;
  wire [31:0] L275_0r0;
  wire [31:0] L275_0r1;
  wire L275_0a;
  wire L276_0r;
  wire L276_0a;
  wire [31:0] L277_0r0;
  wire [31:0] L277_0r1;
  wire L277_0a;
  wire [2:0] L278_0r0;
  wire [2:0] L278_0r1;
  wire L278_0a;
  wire L279_0r;
  wire L279_0a;
  wire [2:0] L280_0r0;
  wire [2:0] L280_0r1;
  wire L280_0a;
  wire L281_0r;
  wire L281_0a;
  wire L282_0r0;
  wire L282_0r1;
  wire L282_0a;
  wire [3:0] L283_0r0;
  wire [3:0] L283_0r1;
  wire L283_0a;
  wire L285_0r;
  wire L285_0a;
  wire [31:0] L286_0r0;
  wire [31:0] L286_0r1;
  wire L286_0a;
  wire L287_0r;
  wire L287_0a;
  wire L288_0r;
  wire L288_0a;
  wire [31:0] L289_0r0;
  wire [31:0] L289_0r1;
  wire L289_0a;
  wire L290_0r;
  wire L290_0a;
  wire [31:0] L291_0r0;
  wire [31:0] L291_0r1;
  wire L291_0a;
  wire L292_0r;
  wire L292_0a;
  wire [31:0] L293_0r0;
  wire [31:0] L293_0r1;
  wire L293_0a;
  wire L294_0r;
  wire L294_0a;
  wire [31:0] L295_0r0;
  wire [31:0] L295_0r1;
  wire L295_0a;
  wire L296_0r;
  wire L296_0a;
  wire [31:0] L297_0r0;
  wire [31:0] L297_0r1;
  wire L297_0a;
  wire L298_0r;
  wire L298_0a;
  wire [31:0] L299_0r0;
  wire [31:0] L299_0r1;
  wire L299_0a;
  wire L300_0r;
  wire L300_0a;
  wire [31:0] L301_0r0;
  wire [31:0] L301_0r1;
  wire L301_0a;
  wire L302_0r;
  wire L302_0a;
  wire [31:0] L303_0r0;
  wire [31:0] L303_0r1;
  wire L303_0a;
  wire [2:0] L304_0r0;
  wire [2:0] L304_0r1;
  wire L304_0a;
  wire L305_0r;
  wire L305_0a;
  wire [2:0] L306_0r0;
  wire [2:0] L306_0r1;
  wire L306_0a;
  wire L307_0r;
  wire L307_0a;
  wire L308_0r0;
  wire L308_0r1;
  wire L308_0a;
  wire [3:0] L309_0r0;
  wire [3:0] L309_0r1;
  wire L309_0a;
  wire L311_0r;
  wire L311_0a;
  wire [31:0] L312_0r0;
  wire [31:0] L312_0r1;
  wire L312_0a;
  wire L313_0r;
  wire L313_0a;
  wire L314_0r;
  wire L314_0a;
  wire [31:0] L315_0r0;
  wire [31:0] L315_0r1;
  wire L315_0a;
  wire L316_0r;
  wire L316_0a;
  wire [31:0] L317_0r0;
  wire [31:0] L317_0r1;
  wire L317_0a;
  wire L318_0r;
  wire L318_0a;
  wire [31:0] L319_0r0;
  wire [31:0] L319_0r1;
  wire L319_0a;
  wire L320_0r;
  wire L320_0a;
  wire [31:0] L321_0r0;
  wire [31:0] L321_0r1;
  wire L321_0a;
  wire L322_0r;
  wire L322_0a;
  wire [31:0] L323_0r0;
  wire [31:0] L323_0r1;
  wire L323_0a;
  wire L324_0r;
  wire L324_0a;
  wire [31:0] L325_0r0;
  wire [31:0] L325_0r1;
  wire L325_0a;
  wire L326_0r;
  wire L326_0a;
  wire [31:0] L327_0r0;
  wire [31:0] L327_0r1;
  wire L327_0a;
  wire L328_0r;
  wire L328_0a;
  wire [31:0] L329_0r0;
  wire [31:0] L329_0r1;
  wire L329_0a;
  wire [2:0] L330_0r0;
  wire [2:0] L330_0r1;
  wire L330_0a;
  wire L331_0r;
  wire L331_0a;
  wire [2:0] L332_0r0;
  wire [2:0] L332_0r1;
  wire L332_0a;
  wire L333_0r0;
  wire L333_0r1;
  wire L333_0a;
  wire L334_0r;
  wire L334_0a;
  wire L335_0r0;
  wire L335_0r1;
  wire L335_0a;
  wire L336_0r;
  wire L336_0a;
  wire L337_0r0;
  wire L337_0r1;
  wire L337_0a;
  wire [1:0] L338_0r0;
  wire [1:0] L338_0r1;
  wire L338_0a;
  wire [1:0] L339_0r0;
  wire [1:0] L339_0r1;
  wire L339_0a;
  wire [3:0] L340_0r0;
  wire [3:0] L340_0r1;
  wire L340_0a;
  wire L342_0r;
  wire L342_0a;
  wire [31:0] L343_0r0;
  wire [31:0] L343_0r1;
  wire L343_0a;
  wire L344_0r;
  wire L344_0a;
  wire L345_0r;
  wire L345_0a;
  wire [4:0] L346_0r0;
  wire [4:0] L346_0r1;
  wire L346_0a;
  wire L348_0r;
  wire L348_0a;
  wire L349_0r;
  wire L349_0a;
  wire L350_0r;
  wire L350_0a;
  wire L352_0r;
  wire L352_0a;
  wire L353_0r0;
  wire L353_0r1;
  wire L353_0a;
  wire L354_0r;
  wire L354_0a;
  wire L355_0r;
  wire L355_0a;
  wire [4:0] L356_0r0;
  wire [4:0] L356_0r1;
  wire L356_0a;
  wire L357_0r;
  wire L357_0a;
  wire L358_0r;
  wire L358_0a;
  wire [31:0] L360_0r0;
  wire [31:0] L360_0r1;
  wire L360_0a;
  wire L361_0r;
  wire L361_0a;
  wire [2:0] L362_0r0;
  wire [2:0] L362_0r1;
  wire L362_0a;
  wire [31:0] L363_0r0;
  wire [31:0] L363_0r1;
  wire L363_0a;
  wire L364_0r;
  wire L364_0a;
  wire [31:0] L365_0r0;
  wire [31:0] L365_0r1;
  wire L365_0a;
  wire L366_0r;
  wire L366_0a;
  wire [31:0] L367_0r0;
  wire [31:0] L367_0r1;
  wire L367_0a;
  wire L368_0r;
  wire L368_0a;
  wire [31:0] L369_0r0;
  wire [31:0] L369_0r1;
  wire L369_0a;
  wire L370_0r;
  wire L370_0a;
  wire [31:0] L371_0r0;
  wire [31:0] L371_0r1;
  wire L371_0a;
  wire L372_0r;
  wire L372_0a;
  wire [31:0] L373_0r0;
  wire [31:0] L373_0r1;
  wire L373_0a;
  wire L374_0r;
  wire L374_0a;
  wire [31:0] L375_0r0;
  wire [31:0] L375_0r1;
  wire L375_0a;
  wire L376_0r;
  wire L376_0a;
  wire [31:0] L377_0r0;
  wire [31:0] L377_0r1;
  wire L377_0a;
  wire [34:0] L378_0r0;
  wire [34:0] L378_0r1;
  wire L378_0a;
  wire L379_0r;
  wire L379_0a;
  wire L380_0r;
  wire L380_0a;
  wire [31:0] L382_0r0;
  wire [31:0] L382_0r1;
  wire L382_0a;
  wire [2:0] L383_0r0;
  wire [2:0] L383_0r1;
  wire L383_0a;
  wire L384_0r;
  wire L384_0a;
  wire [2:0] L385_0r0;
  wire [2:0] L385_0r1;
  wire L385_0a;
  wire L386_0r;
  wire L386_0a;
  wire L387_0r0;
  wire L387_0r1;
  wire L387_0a;
  wire [3:0] L388_0r0;
  wire [3:0] L388_0r1;
  wire L388_0a;
  wire L389_0r;
  wire L389_0a;
  wire [31:0] L390_0r0;
  wire [31:0] L390_0r1;
  wire L390_0a;
  wire L391_0r;
  wire L391_0a;
  wire [31:0] L392_0r0;
  wire [31:0] L392_0r1;
  wire L392_0a;
  wire L393_0r;
  wire L393_0a;
  wire [31:0] L394_0r0;
  wire [31:0] L394_0r1;
  wire L394_0a;
  wire L395_0r;
  wire L395_0a;
  wire [31:0] L396_0r0;
  wire [31:0] L396_0r1;
  wire L396_0a;
  wire L397_0r;
  wire L397_0a;
  wire [31:0] L398_0r0;
  wire [31:0] L398_0r1;
  wire L398_0a;
  wire L399_0r;
  wire L399_0a;
  wire [31:0] L400_0r0;
  wire [31:0] L400_0r1;
  wire L400_0a;
  wire L401_0r;
  wire L401_0a;
  wire [31:0] L402_0r0;
  wire [31:0] L402_0r1;
  wire L402_0a;
  wire L403_0r;
  wire L403_0a;
  wire [31:0] L404_0r0;
  wire [31:0] L404_0r1;
  wire L404_0a;
  wire L405_0r;
  wire L405_0a;
  wire [31:0] L406_0r0;
  wire [31:0] L406_0r1;
  wire L406_0a;
  wire [34:0] L407_0r0;
  wire [34:0] L407_0r1;
  wire L407_0a;
  wire L408_0r;
  wire L408_0a;
  wire L409_0r;
  wire L409_0a;
  wire [31:0] L411_0r0;
  wire [31:0] L411_0r1;
  wire L411_0a;
  wire [2:0] L412_0r0;
  wire [2:0] L412_0r1;
  wire L412_0a;
  wire L413_0r;
  wire L413_0a;
  wire [2:0] L414_0r0;
  wire [2:0] L414_0r1;
  wire L414_0a;
  wire L415_0r;
  wire L415_0a;
  wire L416_0r0;
  wire L416_0r1;
  wire L416_0a;
  wire [3:0] L417_0r0;
  wire [3:0] L417_0r1;
  wire L417_0a;
  wire L418_0r;
  wire L418_0a;
  wire [31:0] L419_0r0;
  wire [31:0] L419_0r1;
  wire L419_0a;
  wire L420_0r;
  wire L420_0a;
  wire [31:0] L421_0r0;
  wire [31:0] L421_0r1;
  wire L421_0a;
  wire L422_0r;
  wire L422_0a;
  wire [31:0] L423_0r0;
  wire [31:0] L423_0r1;
  wire L423_0a;
  wire L424_0r;
  wire L424_0a;
  wire [31:0] L425_0r0;
  wire [31:0] L425_0r1;
  wire L425_0a;
  wire L426_0r;
  wire L426_0a;
  wire [31:0] L427_0r0;
  wire [31:0] L427_0r1;
  wire L427_0a;
  wire L428_0r;
  wire L428_0a;
  wire [31:0] L429_0r0;
  wire [31:0] L429_0r1;
  wire L429_0a;
  wire L430_0r;
  wire L430_0a;
  wire [31:0] L431_0r0;
  wire [31:0] L431_0r1;
  wire L431_0a;
  wire L432_0r;
  wire L432_0a;
  wire [31:0] L433_0r0;
  wire [31:0] L433_0r1;
  wire L433_0a;
  wire L434_0r;
  wire L434_0a;
  wire [31:0] L435_0r0;
  wire [31:0] L435_0r1;
  wire L435_0a;
  wire [34:0] L436_0r0;
  wire [34:0] L436_0r1;
  wire L436_0a;
  wire L437_0r;
  wire L437_0a;
  wire L438_0r;
  wire L438_0a;
  wire [31:0] L440_0r0;
  wire [31:0] L440_0r1;
  wire L440_0a;
  wire [2:0] L441_0r0;
  wire [2:0] L441_0r1;
  wire L441_0a;
  wire L442_0r;
  wire L442_0a;
  wire [2:0] L443_0r0;
  wire [2:0] L443_0r1;
  wire L443_0a;
  wire L444_0r0;
  wire L444_0r1;
  wire L444_0a;
  wire L445_0r;
  wire L445_0a;
  wire L446_0r0;
  wire L446_0r1;
  wire L446_0a;
  wire L447_0r;
  wire L447_0a;
  wire L448_0r0;
  wire L448_0r1;
  wire L448_0a;
  wire [1:0] L449_0r0;
  wire [1:0] L449_0r1;
  wire L449_0a;
  wire [1:0] L450_0r0;
  wire [1:0] L450_0r1;
  wire L450_0a;
  wire [3:0] L451_0r0;
  wire [3:0] L451_0r1;
  wire L451_0a;
  wire L452_0r;
  wire L452_0a;
  wire [31:0] L453_0r0;
  wire [31:0] L453_0r1;
  wire L453_0a;
  wire L454_0r;
  wire L454_0a;
  wire [31:0] L455_0r0;
  wire [31:0] L455_0r1;
  wire L455_0a;
  wire L456_0r;
  wire L456_0a;
  wire [31:0] L457_0r0;
  wire [31:0] L457_0r1;
  wire L457_0a;
  wire L458_0r;
  wire L458_0a;
  wire [31:0] L459_0r0;
  wire [31:0] L459_0r1;
  wire L459_0a;
  wire L460_0r;
  wire L460_0a;
  wire [31:0] L461_0r0;
  wire [31:0] L461_0r1;
  wire L461_0a;
  wire L462_0r;
  wire L462_0a;
  wire [31:0] L463_0r0;
  wire [31:0] L463_0r1;
  wire L463_0a;
  wire L464_0r;
  wire L464_0a;
  wire [31:0] L465_0r0;
  wire [31:0] L465_0r1;
  wire L465_0a;
  wire L466_0r;
  wire L466_0a;
  wire [31:0] L467_0r0;
  wire [31:0] L467_0r1;
  wire L467_0a;
  wire L468_0r;
  wire L468_0a;
  wire [31:0] L469_0r0;
  wire [31:0] L469_0r1;
  wire L469_0a;
  wire [34:0] L470_0r0;
  wire [34:0] L470_0r1;
  wire L470_0a;
  wire L471_0r;
  wire L471_0a;
  wire L472_0r;
  wire L472_0a;
  wire [4:0] L473_0r0;
  wire [4:0] L473_0r1;
  wire L473_0a;
  wire L474_0r;
  wire L474_0a;
  wire [31:0] L475_0r0;
  wire [31:0] L475_0r1;
  wire L475_0a;
  wire L476_0r;
  wire L476_0a;
  wire L478_0r;
  wire L478_0a;
  wire L479_0r;
  wire L479_0a;
  wire L480_0r;
  wire L480_0a;
  wire L481_0r;
  wire L481_0a;
  wire L482_0r0;
  wire L482_0r1;
  wire L482_0a;
  wire L483_0r;
  wire L483_0a;
  wire [2:0] L484_0r0;
  wire [2:0] L484_0r1;
  wire L484_0a;
  wire L485_0r;
  wire L485_0a;
  wire L486_0r0;
  wire L486_0r1;
  wire L486_0a;
  wire L487_0r;
  wire L487_0a;
  wire L489_0r;
  wire L489_0a;
  wire L490_0r;
  wire L490_0a;
  wire L491_0r;
  wire L491_0a;
  wire L492_0r;
  wire L492_0a;
  wire [31:0] L494_0r0;
  wire [31:0] L494_0r1;
  wire L494_0a;
  wire L495_0r;
  wire L495_0a;
  wire L496_0r;
  wire L496_0a;
  wire [31:0] L497_0r0;
  wire [31:0] L497_0r1;
  wire L497_0a;
  wire L498_0r;
  wire L498_0a;
  wire [31:0] L499_0r0;
  wire [31:0] L499_0r1;
  wire L499_0a;
  wire [1:0] L500_0r0;
  wire [1:0] L500_0r1;
  wire L500_0a;
  wire [1:0] L501_0r0;
  wire [1:0] L501_0r1;
  wire L501_0a;
  wire [1:0] L502_0r0;
  wire [1:0] L502_0r1;
  wire L502_0a;
  wire [1:0] L503_0r0;
  wire [1:0] L503_0r1;
  wire L503_0a;
  wire [31:0] L504_0r0;
  wire [31:0] L504_0r1;
  wire L504_0a;
  wire L505_0r;
  wire L505_0a;
  wire L506_0r;
  wire L506_0a;
  wire [31:0] L507_0r0;
  wire [31:0] L507_0r1;
  wire L507_0a;
  wire L508_0r;
  wire L508_0a;
  wire [31:0] L509_0r0;
  wire [31:0] L509_0r1;
  wire L509_0a;
  wire [1:0] L510_0r0;
  wire [1:0] L510_0r1;
  wire L510_0a;
  wire [1:0] L511_0r0;
  wire [1:0] L511_0r1;
  wire L511_0a;
  wire [1:0] L512_0r0;
  wire [1:0] L512_0r1;
  wire L512_0a;
  wire [1:0] L513_0r0;
  wire [1:0] L513_0r1;
  wire L513_0a;
  wire [31:0] L514_0r0;
  wire [31:0] L514_0r1;
  wire L514_0a;
  wire L515_0r;
  wire L515_0a;
  wire L516_0r;
  wire L516_0a;
  wire [31:0] L517_0r0;
  wire [31:0] L517_0r1;
  wire L517_0a;
  wire L518_0r;
  wire L518_0a;
  wire [31:0] L519_0r0;
  wire [31:0] L519_0r1;
  wire L519_0a;
  wire [1:0] L520_0r0;
  wire [1:0] L520_0r1;
  wire L520_0a;
  wire [1:0] L521_0r0;
  wire [1:0] L521_0r1;
  wire L521_0a;
  wire [1:0] L522_0r0;
  wire [1:0] L522_0r1;
  wire L522_0a;
  wire [1:0] L523_0r0;
  wire [1:0] L523_0r1;
  wire L523_0a;
  wire [31:0] L524_0r0;
  wire [31:0] L524_0r1;
  wire L524_0a;
  wire L525_0r;
  wire L525_0a;
  wire L526_0r;
  wire L526_0a;
  wire [31:0] L527_0r0;
  wire [31:0] L527_0r1;
  wire L527_0a;
  wire L528_0r;
  wire L528_0a;
  wire [31:0] L529_0r0;
  wire [31:0] L529_0r1;
  wire L529_0a;
  wire [1:0] L530_0r0;
  wire [1:0] L530_0r1;
  wire L530_0a;
  wire [1:0] L531_0r0;
  wire [1:0] L531_0r1;
  wire L531_0a;
  wire [1:0] L532_0r0;
  wire [1:0] L532_0r1;
  wire L532_0a;
  wire [1:0] L533_0r0;
  wire [1:0] L533_0r1;
  wire L533_0a;
  wire [31:0] L534_0r0;
  wire [31:0] L534_0r1;
  wire L534_0a;
  wire L535_0r;
  wire L535_0a;
  wire L536_0r;
  wire L536_0a;
  wire [31:0] L537_0r0;
  wire [31:0] L537_0r1;
  wire L537_0a;
  wire L538_0r;
  wire L538_0a;
  wire [31:0] L539_0r0;
  wire [31:0] L539_0r1;
  wire L539_0a;
  wire [1:0] L540_0r0;
  wire [1:0] L540_0r1;
  wire L540_0a;
  wire [1:0] L541_0r0;
  wire [1:0] L541_0r1;
  wire L541_0a;
  wire [1:0] L542_0r0;
  wire [1:0] L542_0r1;
  wire L542_0a;
  wire [1:0] L543_0r0;
  wire [1:0] L543_0r1;
  wire L543_0a;
  wire [31:0] L544_0r0;
  wire [31:0] L544_0r1;
  wire L544_0a;
  wire L545_0r;
  wire L545_0a;
  wire L546_0r;
  wire L546_0a;
  wire [31:0] L547_0r0;
  wire [31:0] L547_0r1;
  wire L547_0a;
  wire L548_0r;
  wire L548_0a;
  wire [31:0] L549_0r0;
  wire [31:0] L549_0r1;
  wire L549_0a;
  wire [1:0] L550_0r0;
  wire [1:0] L550_0r1;
  wire L550_0a;
  wire [1:0] L551_0r0;
  wire [1:0] L551_0r1;
  wire L551_0a;
  wire [1:0] L552_0r0;
  wire [1:0] L552_0r1;
  wire L552_0a;
  wire [1:0] L553_0r0;
  wire [1:0] L553_0r1;
  wire L553_0a;
  wire [31:0] L554_0r0;
  wire [31:0] L554_0r1;
  wire L554_0a;
  wire L555_0r;
  wire L555_0a;
  wire L556_0r;
  wire L556_0a;
  wire [31:0] L557_0r0;
  wire [31:0] L557_0r1;
  wire L557_0a;
  wire L558_0r;
  wire L558_0a;
  wire [31:0] L559_0r0;
  wire [31:0] L559_0r1;
  wire L559_0a;
  wire [1:0] L560_0r0;
  wire [1:0] L560_0r1;
  wire L560_0a;
  wire [1:0] L561_0r0;
  wire [1:0] L561_0r1;
  wire L561_0a;
  wire [1:0] L562_0r0;
  wire [1:0] L562_0r1;
  wire L562_0a;
  wire [1:0] L563_0r0;
  wire [1:0] L563_0r1;
  wire L563_0a;
  wire [31:0] L564_0r0;
  wire [31:0] L564_0r1;
  wire L564_0a;
  wire L565_0r;
  wire L565_0a;
  wire L566_0r;
  wire L566_0a;
  wire [31:0] L567_0r0;
  wire [31:0] L567_0r1;
  wire L567_0a;
  wire L568_0r;
  wire L568_0a;
  wire [31:0] L569_0r0;
  wire [31:0] L569_0r1;
  wire L569_0a;
  wire [1:0] L570_0r0;
  wire [1:0] L570_0r1;
  wire L570_0a;
  wire [1:0] L571_0r0;
  wire [1:0] L571_0r1;
  wire L571_0a;
  wire [1:0] L572_0r0;
  wire [1:0] L572_0r1;
  wire L572_0a;
  wire [1:0] L573_0r0;
  wire [1:0] L573_0r1;
  wire L573_0a;
  wire L582_0r;
  wire L582_0a;
  wire [31:0] L583_0r0;
  wire [31:0] L583_0r1;
  wire L583_0a;
  wire L584_0r;
  wire L584_0a;
  wire [31:0] L585_0r0;
  wire [31:0] L585_0r1;
  wire L585_0a;
  wire L586_0r;
  wire L586_0a;
  wire [31:0] L587_0r0;
  wire [31:0] L587_0r1;
  wire L587_0a;
  wire L588_0r;
  wire L588_0a;
  wire [31:0] L589_0r0;
  wire [31:0] L589_0r1;
  wire L589_0a;
  wire L590_0r;
  wire L590_0a;
  wire [31:0] L591_0r0;
  wire [31:0] L591_0r1;
  wire L591_0a;
  wire [31:0] L592_0r0;
  wire [31:0] L592_0r1;
  wire L592_0a;
  wire L593_0r;
  wire L593_0a;
  wire [4:0] L595_0r0;
  wire [4:0] L595_0r1;
  wire L595_0a;
  wire [4:0] L596_0r0;
  wire [4:0] L596_0r1;
  wire L596_0a;
  wire [4:0] L597_0r0;
  wire [4:0] L597_0r1;
  wire L597_0a;
  wire [4:0] L598_0r0;
  wire [4:0] L598_0r1;
  wire L598_0a;
  wire [4:0] L599_0r0;
  wire [4:0] L599_0r1;
  wire L599_0a;
  wire [4:0] L600_0r0;
  wire [4:0] L600_0r1;
  wire L600_0a;
  wire [4:0] L601_0r0;
  wire [4:0] L601_0r1;
  wire L601_0a;
  wire L602_0r;
  wire L602_0a;
  wire [31:0] L603_0r0;
  wire [31:0] L603_0r1;
  wire L603_0a;
  wire L604_0r;
  wire L604_0a;
  wire [31:0] L605_0r0;
  wire [31:0] L605_0r1;
  wire L605_0a;
  wire L606_0r;
  wire L606_0a;
  wire [31:0] L607_0r0;
  wire [31:0] L607_0r1;
  wire L607_0a;
  wire L608_0r;
  wire L608_0a;
  wire [31:0] L609_0r0;
  wire [31:0] L609_0r1;
  wire L609_0a;
  wire L610_0r;
  wire L610_0a;
  wire [31:0] L611_0r0;
  wire [31:0] L611_0r1;
  wire L611_0a;
  wire [31:0] L612_0r0;
  wire [31:0] L612_0r1;
  wire L612_0a;
  wire L613_0r;
  wire L613_0a;
  wire [4:0] L615_0r0;
  wire [4:0] L615_0r1;
  wire L615_0a;
  wire [4:0] L616_0r0;
  wire [4:0] L616_0r1;
  wire L616_0a;
  wire [4:0] L617_0r0;
  wire [4:0] L617_0r1;
  wire L617_0a;
  wire [4:0] L618_0r0;
  wire [4:0] L618_0r1;
  wire L618_0a;
  wire [4:0] L619_0r0;
  wire [4:0] L619_0r1;
  wire L619_0a;
  wire [4:0] L620_0r0;
  wire [4:0] L620_0r1;
  wire L620_0a;
  wire [4:0] L621_0r0;
  wire [4:0] L621_0r1;
  wire L621_0a;
  wire L622_0r;
  wire L622_0a;
  wire [31:0] L623_0r0;
  wire [31:0] L623_0r1;
  wire L623_0a;
  wire L624_0r;
  wire L624_0a;
  wire [31:0] L625_0r0;
  wire [31:0] L625_0r1;
  wire L625_0a;
  wire L626_0r;
  wire L626_0a;
  wire [31:0] L627_0r0;
  wire [31:0] L627_0r1;
  wire L627_0a;
  wire L628_0r;
  wire L628_0a;
  wire [31:0] L629_0r0;
  wire [31:0] L629_0r1;
  wire L629_0a;
  wire L630_0r;
  wire L630_0a;
  wire [31:0] L631_0r0;
  wire [31:0] L631_0r1;
  wire L631_0a;
  wire [31:0] L632_0r0;
  wire [31:0] L632_0r1;
  wire L632_0a;
  wire L633_0r;
  wire L633_0a;
  wire [4:0] L635_0r0;
  wire [4:0] L635_0r1;
  wire L635_0a;
  wire [4:0] L636_0r0;
  wire [4:0] L636_0r1;
  wire L636_0a;
  wire [4:0] L637_0r0;
  wire [4:0] L637_0r1;
  wire L637_0a;
  wire [4:0] L638_0r0;
  wire [4:0] L638_0r1;
  wire L638_0a;
  wire [4:0] L639_0r0;
  wire [4:0] L639_0r1;
  wire L639_0a;
  wire [4:0] L640_0r0;
  wire [4:0] L640_0r1;
  wire L640_0a;
  wire [4:0] L641_0r0;
  wire [4:0] L641_0r1;
  wire L641_0a;
  tko0m32_1nm32b0 I0 (L7_0r, L7_0a, L9_0r0[31:0], L9_0r1[31:0], L9_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0 I1 (L26_0r0[2:0], L26_0r1[2:0], L26_0a, L11_0r, L11_0a, L13_0r, L13_0a, L15_0r, L15_0a, L17_0r, L17_0a, L19_0r, L19_0a, L21_0r, L21_0a, L23_0r, L23_0a, reset);
  tkm7x32b I2 (L12_0r0[31:0], L12_0r1[31:0], L12_0a, L14_0r0[31:0], L14_0r1[31:0], L14_0a, L16_0r0[31:0], L16_0r1[31:0], L16_0a, L18_0r0[31:0], L18_0r1[31:0], L18_0a, L20_0r0[31:0], L20_0r1[31:0], L20_0a, L22_0r0[31:0], L22_0r1[31:0], L22_0a, L24_0r0[31:0], L24_0r1[31:0], L24_0a, L28_0r0[31:0], L28_0r1[31:0], L28_0a, reset);
  tkj4m3_1 I3 (L48_0r0[2:0], L48_0r1[2:0], L48_0a, L50_0r0, L50_0r1, L50_0a, L51_0r0[3:0], L51_0r1[3:0], L51_0a, reset);
  tkf4mo0w3 I4 (L51_0r0[3:0], L51_0r1[3:0], L51_0a, L46_0r0[2:0], L46_0r1[2:0], L46_0a, reset);
  tks3_o0w3_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0 I5 (L46_0r0[2:0], L46_0r1[2:0], L46_0a, L30_0r, L30_0a, L32_0r, L32_0a, L34_0r, L34_0a, L36_0r, L36_0a, L38_0r, L38_0a, L40_0r, L40_0a, L42_0r, L42_0a, L44_0r, L44_0a, reset);
  tkm8x32b I6 (L31_0r0[31:0], L31_0r1[31:0], L31_0a, L33_0r0[31:0], L33_0r1[31:0], L33_0a, L35_0r0[31:0], L35_0r1[31:0], L35_0a, L37_0r0[31:0], L37_0r1[31:0], L37_0a, L39_0r0[31:0], L39_0r1[31:0], L39_0a, L41_0r0[31:0], L41_0r1[31:0], L41_0a, L43_0r0[31:0], L43_0r1[31:0], L43_0a, L45_0r0[31:0], L45_0r1[31:0], L45_0a, L54_0r0[31:0], L54_0r1[31:0], L54_0a, reset);
  tkf0mo0w0_o0w0 I7 (L53_0r, L53_0a, L47_0r, L47_0a, L49_0r, L49_0a, reset);
  tkj4m3_1 I8 (L74_0r0[2:0], L74_0r1[2:0], L74_0a, L76_0r0, L76_0r1, L76_0a, L77_0r0[3:0], L77_0r1[3:0], L77_0a, reset);
  tkf4mo0w3 I9 (L77_0r0[3:0], L77_0r1[3:0], L77_0a, L72_0r0[2:0], L72_0r1[2:0], L72_0a, reset);
  tks3_o0w3_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0 I10 (L72_0r0[2:0], L72_0r1[2:0], L72_0a, L56_0r, L56_0a, L58_0r, L58_0a, L60_0r, L60_0a, L62_0r, L62_0a, L64_0r, L64_0a, L66_0r, L66_0a, L68_0r, L68_0a, L70_0r, L70_0a, reset);
  tkm8x32b I11 (L57_0r0[31:0], L57_0r1[31:0], L57_0a, L59_0r0[31:0], L59_0r1[31:0], L59_0a, L61_0r0[31:0], L61_0r1[31:0], L61_0a, L63_0r0[31:0], L63_0r1[31:0], L63_0a, L65_0r0[31:0], L65_0r1[31:0], L65_0a, L67_0r0[31:0], L67_0r1[31:0], L67_0a, L69_0r0[31:0], L69_0r1[31:0], L69_0a, L71_0r0[31:0], L71_0r1[31:0], L71_0a, L80_0r0[31:0], L80_0r1[31:0], L80_0a, reset);
  tkf0mo0w0_o0w0 I12 (L79_0r, L79_0a, L73_0r, L73_0a, L75_0r, L75_0a, reset);
  tko0m1_1nm1b1 I13 (L104_0r, L104_0a, L105_0r0, L105_0r1, L105_0a, reset);
  tkj2m1_1 I14 (L103_0r0, L103_0r1, L103_0a, L105_0r0, L105_0r1, L105_0a, L106_0r0[1:0], L106_0r1[1:0], L106_0a, reset);
  tko2m2_1api0w1b_2api1w1b_3nm1b0_4apt1o0w1bt3o0w1b_5nm1b0_6apt2o0w1bt5o0w1b_7addt4o0w2bt6o0w2b I15 (L106_0r0[1:0], L106_0r1[1:0], L106_0a, L107_0r0[1:0], L107_0r1[1:0], L107_0a, reset);
  tkf2mo0w1 I16 (L107_0r0[1:0], L107_0r1[1:0], L107_0a, L101_0r0, L101_0r1, L101_0a, reset);
  tkj4m3_1 I17 (L100_0r0[2:0], L100_0r1[2:0], L100_0a, L101_0r0, L101_0r1, L101_0a, L108_0r0[3:0], L108_0r1[3:0], L108_0a, reset);
  tkf4mo0w3 I18 (L108_0r0[3:0], L108_0r1[3:0], L108_0a, L98_0r0[2:0], L98_0r1[2:0], L98_0a, reset);
  tks3_o0w3_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0 I19 (L98_0r0[2:0], L98_0r1[2:0], L98_0a, L82_0r, L82_0a, L84_0r, L84_0a, L86_0r, L86_0a, L88_0r, L88_0a, L90_0r, L90_0a, L92_0r, L92_0a, L94_0r, L94_0a, L96_0r, L96_0a, reset);
  tkm8x32b I20 (L83_0r0[31:0], L83_0r1[31:0], L83_0a, L85_0r0[31:0], L85_0r1[31:0], L85_0a, L87_0r0[31:0], L87_0r1[31:0], L87_0a, L89_0r0[31:0], L89_0r1[31:0], L89_0a, L91_0r0[31:0], L91_0r1[31:0], L91_0a, L93_0r0[31:0], L93_0r1[31:0], L93_0a, L95_0r0[31:0], L95_0r1[31:0], L95_0a, L97_0r0[31:0], L97_0r1[31:0], L97_0a, L111_0r0[31:0], L111_0r1[31:0], L111_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I21 (L110_0r, L110_0a, L99_0r, L99_0a, L102_0r, L102_0a, L104_0r, L104_0a, reset);
  tks5_o0w5_0o0w0_1m2c1m4c3o0w0_8c7o0w0_10c7o0w0_18c7o0w0 I22 (L6_0r0[4:0], L6_0r1[4:0], L6_0a, L7_0r, L7_0a, L25_0r, L25_0a, L53_0r, L53_0a, L79_0r, L79_0a, L110_0r, L110_0a, reset);
  tkm5x0b I23 (L10_0r, L10_0a, L29_0r, L29_0a, L55_0r, L55_0a, L81_0r, L81_0a, L112_0r, L112_0a, L113_0r, L113_0a, reset);
  tkvsel5_wo0w5_ro0w5o0w3o0w3o0w3o0w3 I24 (L114_0r0[4:0], L114_0r1[4:0], L114_0a, L5_0r, L5_0a, L5_0r, L5_0a, L25_0r, L25_0a, L47_0r, L47_0a, L73_0r, L73_0a, L99_0r, L99_0a, L6_0r0[4:0], L6_0r1[4:0], L6_0a, L26_0r0[2:0], L26_0r1[2:0], L26_0a, L48_0r0[2:0], L48_0r1[2:0], L48_0a, L74_0r0[2:0], L74_0r1[2:0], L74_0a, L100_0r0[2:0], L100_0r1[2:0], L100_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I25 (L3_0r0, L3_0r1, L3_0a, L4_0r, L4_0a, L116_0r, L116_0a, reset);
  tkm2x0b I26 (L4_0r, L4_0a, L113_0r, L113_0a, L117_0r, L117_0a, reset);
  tko0m32_1nm32b0 I27 (L123_0r, L123_0a, L125_0r0[31:0], L125_0r1[31:0], L125_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0 I28 (L142_0r0[2:0], L142_0r1[2:0], L142_0a, L127_0r, L127_0a, L129_0r, L129_0a, L131_0r, L131_0a, L133_0r, L133_0a, L135_0r, L135_0a, L137_0r, L137_0a, L139_0r, L139_0a, reset);
  tkm7x32b I29 (L128_0r0[31:0], L128_0r1[31:0], L128_0a, L130_0r0[31:0], L130_0r1[31:0], L130_0a, L132_0r0[31:0], L132_0r1[31:0], L132_0a, L134_0r0[31:0], L134_0r1[31:0], L134_0a, L136_0r0[31:0], L136_0r1[31:0], L136_0a, L138_0r0[31:0], L138_0r1[31:0], L138_0a, L140_0r0[31:0], L140_0r1[31:0], L140_0a, L144_0r0[31:0], L144_0r1[31:0], L144_0a, reset);
  tkj4m3_1 I30 (L164_0r0[2:0], L164_0r1[2:0], L164_0a, L166_0r0, L166_0r1, L166_0a, L167_0r0[3:0], L167_0r1[3:0], L167_0a, reset);
  tkf4mo0w3 I31 (L167_0r0[3:0], L167_0r1[3:0], L167_0a, L162_0r0[2:0], L162_0r1[2:0], L162_0a, reset);
  tks3_o0w3_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0 I32 (L162_0r0[2:0], L162_0r1[2:0], L162_0a, L146_0r, L146_0a, L148_0r, L148_0a, L150_0r, L150_0a, L152_0r, L152_0a, L154_0r, L154_0a, L156_0r, L156_0a, L158_0r, L158_0a, L160_0r, L160_0a, reset);
  tkm8x32b I33 (L147_0r0[31:0], L147_0r1[31:0], L147_0a, L149_0r0[31:0], L149_0r1[31:0], L149_0a, L151_0r0[31:0], L151_0r1[31:0], L151_0a, L153_0r0[31:0], L153_0r1[31:0], L153_0a, L155_0r0[31:0], L155_0r1[31:0], L155_0a, L157_0r0[31:0], L157_0r1[31:0], L157_0a, L159_0r0[31:0], L159_0r1[31:0], L159_0a, L161_0r0[31:0], L161_0r1[31:0], L161_0a, L170_0r0[31:0], L170_0r1[31:0], L170_0a, reset);
  tkf0mo0w0_o0w0 I34 (L169_0r, L169_0a, L163_0r, L163_0a, L165_0r, L165_0a, reset);
  tkj4m3_1 I35 (L190_0r0[2:0], L190_0r1[2:0], L190_0a, L192_0r0, L192_0r1, L192_0a, L193_0r0[3:0], L193_0r1[3:0], L193_0a, reset);
  tkf4mo0w3 I36 (L193_0r0[3:0], L193_0r1[3:0], L193_0a, L188_0r0[2:0], L188_0r1[2:0], L188_0a, reset);
  tks3_o0w3_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0 I37 (L188_0r0[2:0], L188_0r1[2:0], L188_0a, L172_0r, L172_0a, L174_0r, L174_0a, L176_0r, L176_0a, L178_0r, L178_0a, L180_0r, L180_0a, L182_0r, L182_0a, L184_0r, L184_0a, L186_0r, L186_0a, reset);
  tkm8x32b I38 (L173_0r0[31:0], L173_0r1[31:0], L173_0a, L175_0r0[31:0], L175_0r1[31:0], L175_0a, L177_0r0[31:0], L177_0r1[31:0], L177_0a, L179_0r0[31:0], L179_0r1[31:0], L179_0a, L181_0r0[31:0], L181_0r1[31:0], L181_0a, L183_0r0[31:0], L183_0r1[31:0], L183_0a, L185_0r0[31:0], L185_0r1[31:0], L185_0a, L187_0r0[31:0], L187_0r1[31:0], L187_0a, L196_0r0[31:0], L196_0r1[31:0], L196_0a, reset);
  tkf0mo0w0_o0w0 I39 (L195_0r, L195_0a, L189_0r, L189_0a, L191_0r, L191_0a, reset);
  tko0m1_1nm1b1 I40 (L220_0r, L220_0a, L221_0r0, L221_0r1, L221_0a, reset);
  tkj2m1_1 I41 (L219_0r0, L219_0r1, L219_0a, L221_0r0, L221_0r1, L221_0a, L222_0r0[1:0], L222_0r1[1:0], L222_0a, reset);
  tko2m2_1api0w1b_2api1w1b_3nm1b0_4apt1o0w1bt3o0w1b_5nm1b0_6apt2o0w1bt5o0w1b_7addt4o0w2bt6o0w2b I42 (L222_0r0[1:0], L222_0r1[1:0], L222_0a, L223_0r0[1:0], L223_0r1[1:0], L223_0a, reset);
  tkf2mo0w1 I43 (L223_0r0[1:0], L223_0r1[1:0], L223_0a, L217_0r0, L217_0r1, L217_0a, reset);
  tkj4m3_1 I44 (L216_0r0[2:0], L216_0r1[2:0], L216_0a, L217_0r0, L217_0r1, L217_0a, L224_0r0[3:0], L224_0r1[3:0], L224_0a, reset);
  tkf4mo0w3 I45 (L224_0r0[3:0], L224_0r1[3:0], L224_0a, L214_0r0[2:0], L214_0r1[2:0], L214_0a, reset);
  tks3_o0w3_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0 I46 (L214_0r0[2:0], L214_0r1[2:0], L214_0a, L198_0r, L198_0a, L200_0r, L200_0a, L202_0r, L202_0a, L204_0r, L204_0a, L206_0r, L206_0a, L208_0r, L208_0a, L210_0r, L210_0a, L212_0r, L212_0a, reset);
  tkm8x32b I47 (L199_0r0[31:0], L199_0r1[31:0], L199_0a, L201_0r0[31:0], L201_0r1[31:0], L201_0a, L203_0r0[31:0], L203_0r1[31:0], L203_0a, L205_0r0[31:0], L205_0r1[31:0], L205_0a, L207_0r0[31:0], L207_0r1[31:0], L207_0a, L209_0r0[31:0], L209_0r1[31:0], L209_0a, L211_0r0[31:0], L211_0r1[31:0], L211_0a, L213_0r0[31:0], L213_0r1[31:0], L213_0a, L227_0r0[31:0], L227_0r1[31:0], L227_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I48 (L226_0r, L226_0a, L215_0r, L215_0a, L218_0r, L218_0a, L220_0r, L220_0a, reset);
  tks5_o0w5_0o0w0_1m2c1m4c3o0w0_8c7o0w0_10c7o0w0_18c7o0w0 I49 (L122_0r0[4:0], L122_0r1[4:0], L122_0a, L123_0r, L123_0a, L141_0r, L141_0a, L169_0r, L169_0a, L195_0r, L195_0a, L226_0r, L226_0a, reset);
  tkm5x0b I50 (L126_0r, L126_0a, L145_0r, L145_0a, L171_0r, L171_0a, L197_0r, L197_0a, L228_0r, L228_0a, L229_0r, L229_0a, reset);
  tkvsel5_wo0w5_ro0w5o0w3o0w3o0w3o0w3 I51 (L230_0r0[4:0], L230_0r1[4:0], L230_0a, L121_0r, L121_0a, L121_0r, L121_0a, L141_0r, L141_0a, L163_0r, L163_0a, L189_0r, L189_0a, L215_0r, L215_0a, L122_0r0[4:0], L122_0r1[4:0], L122_0a, L142_0r0[2:0], L142_0r1[2:0], L142_0a, L164_0r0[2:0], L164_0r1[2:0], L164_0a, L190_0r0[2:0], L190_0r1[2:0], L190_0a, L216_0r0[2:0], L216_0r1[2:0], L216_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I52 (L119_0r0, L119_0r1, L119_0a, L120_0r, L120_0a, L232_0r, L232_0a, reset);
  tkm2x0b I53 (L120_0r, L120_0a, L229_0r, L229_0a, L233_0r, L233_0a, reset);
  tko0m32_1nm32b0 I54 (L239_0r, L239_0a, L241_0r0[31:0], L241_0r1[31:0], L241_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0 I55 (L258_0r0[2:0], L258_0r1[2:0], L258_0a, L243_0r, L243_0a, L245_0r, L245_0a, L247_0r, L247_0a, L249_0r, L249_0a, L251_0r, L251_0a, L253_0r, L253_0a, L255_0r, L255_0a, reset);
  tkm7x32b I56 (L244_0r0[31:0], L244_0r1[31:0], L244_0a, L246_0r0[31:0], L246_0r1[31:0], L246_0a, L248_0r0[31:0], L248_0r1[31:0], L248_0a, L250_0r0[31:0], L250_0r1[31:0], L250_0a, L252_0r0[31:0], L252_0r1[31:0], L252_0a, L254_0r0[31:0], L254_0r1[31:0], L254_0a, L256_0r0[31:0], L256_0r1[31:0], L256_0a, L260_0r0[31:0], L260_0r1[31:0], L260_0a, reset);
  tkj4m3_1 I57 (L280_0r0[2:0], L280_0r1[2:0], L280_0a, L282_0r0, L282_0r1, L282_0a, L283_0r0[3:0], L283_0r1[3:0], L283_0a, reset);
  tkf4mo0w3 I58 (L283_0r0[3:0], L283_0r1[3:0], L283_0a, L278_0r0[2:0], L278_0r1[2:0], L278_0a, reset);
  tks3_o0w3_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0 I59 (L278_0r0[2:0], L278_0r1[2:0], L278_0a, L262_0r, L262_0a, L264_0r, L264_0a, L266_0r, L266_0a, L268_0r, L268_0a, L270_0r, L270_0a, L272_0r, L272_0a, L274_0r, L274_0a, L276_0r, L276_0a, reset);
  tkm8x32b I60 (L263_0r0[31:0], L263_0r1[31:0], L263_0a, L265_0r0[31:0], L265_0r1[31:0], L265_0a, L267_0r0[31:0], L267_0r1[31:0], L267_0a, L269_0r0[31:0], L269_0r1[31:0], L269_0a, L271_0r0[31:0], L271_0r1[31:0], L271_0a, L273_0r0[31:0], L273_0r1[31:0], L273_0a, L275_0r0[31:0], L275_0r1[31:0], L275_0a, L277_0r0[31:0], L277_0r1[31:0], L277_0a, L286_0r0[31:0], L286_0r1[31:0], L286_0a, reset);
  tkf0mo0w0_o0w0 I61 (L285_0r, L285_0a, L279_0r, L279_0a, L281_0r, L281_0a, reset);
  tkj4m3_1 I62 (L306_0r0[2:0], L306_0r1[2:0], L306_0a, L308_0r0, L308_0r1, L308_0a, L309_0r0[3:0], L309_0r1[3:0], L309_0a, reset);
  tkf4mo0w3 I63 (L309_0r0[3:0], L309_0r1[3:0], L309_0a, L304_0r0[2:0], L304_0r1[2:0], L304_0a, reset);
  tks3_o0w3_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0 I64 (L304_0r0[2:0], L304_0r1[2:0], L304_0a, L288_0r, L288_0a, L290_0r, L290_0a, L292_0r, L292_0a, L294_0r, L294_0a, L296_0r, L296_0a, L298_0r, L298_0a, L300_0r, L300_0a, L302_0r, L302_0a, reset);
  tkm8x32b I65 (L289_0r0[31:0], L289_0r1[31:0], L289_0a, L291_0r0[31:0], L291_0r1[31:0], L291_0a, L293_0r0[31:0], L293_0r1[31:0], L293_0a, L295_0r0[31:0], L295_0r1[31:0], L295_0a, L297_0r0[31:0], L297_0r1[31:0], L297_0a, L299_0r0[31:0], L299_0r1[31:0], L299_0a, L301_0r0[31:0], L301_0r1[31:0], L301_0a, L303_0r0[31:0], L303_0r1[31:0], L303_0a, L312_0r0[31:0], L312_0r1[31:0], L312_0a, reset);
  tkf0mo0w0_o0w0 I66 (L311_0r, L311_0a, L305_0r, L305_0a, L307_0r, L307_0a, reset);
  tko0m1_1nm1b1 I67 (L336_0r, L336_0a, L337_0r0, L337_0r1, L337_0a, reset);
  tkj2m1_1 I68 (L335_0r0, L335_0r1, L335_0a, L337_0r0, L337_0r1, L337_0a, L338_0r0[1:0], L338_0r1[1:0], L338_0a, reset);
  tko2m2_1api0w1b_2api1w1b_3nm1b0_4apt1o0w1bt3o0w1b_5nm1b0_6apt2o0w1bt5o0w1b_7addt4o0w2bt6o0w2b I69 (L338_0r0[1:0], L338_0r1[1:0], L338_0a, L339_0r0[1:0], L339_0r1[1:0], L339_0a, reset);
  tkf2mo0w1 I70 (L339_0r0[1:0], L339_0r1[1:0], L339_0a, L333_0r0, L333_0r1, L333_0a, reset);
  tkj4m3_1 I71 (L332_0r0[2:0], L332_0r1[2:0], L332_0a, L333_0r0, L333_0r1, L333_0a, L340_0r0[3:0], L340_0r1[3:0], L340_0a, reset);
  tkf4mo0w3 I72 (L340_0r0[3:0], L340_0r1[3:0], L340_0a, L330_0r0[2:0], L330_0r1[2:0], L330_0a, reset);
  tks3_o0w3_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0 I73 (L330_0r0[2:0], L330_0r1[2:0], L330_0a, L314_0r, L314_0a, L316_0r, L316_0a, L318_0r, L318_0a, L320_0r, L320_0a, L322_0r, L322_0a, L324_0r, L324_0a, L326_0r, L326_0a, L328_0r, L328_0a, reset);
  tkm8x32b I74 (L315_0r0[31:0], L315_0r1[31:0], L315_0a, L317_0r0[31:0], L317_0r1[31:0], L317_0a, L319_0r0[31:0], L319_0r1[31:0], L319_0a, L321_0r0[31:0], L321_0r1[31:0], L321_0a, L323_0r0[31:0], L323_0r1[31:0], L323_0a, L325_0r0[31:0], L325_0r1[31:0], L325_0a, L327_0r0[31:0], L327_0r1[31:0], L327_0a, L329_0r0[31:0], L329_0r1[31:0], L329_0a, L343_0r0[31:0], L343_0r1[31:0], L343_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I75 (L342_0r, L342_0a, L331_0r, L331_0a, L334_0r, L334_0a, L336_0r, L336_0a, reset);
  tks5_o0w5_0o0w0_1m2c1m4c3o0w0_8c7o0w0_10c7o0w0_18c7o0w0 I76 (L238_0r0[4:0], L238_0r1[4:0], L238_0a, L239_0r, L239_0a, L257_0r, L257_0a, L285_0r, L285_0a, L311_0r, L311_0a, L342_0r, L342_0a, reset);
  tkm5x0b I77 (L242_0r, L242_0a, L261_0r, L261_0a, L287_0r, L287_0a, L313_0r, L313_0a, L344_0r, L344_0a, L345_0r, L345_0a, reset);
  tkvsel5_wo0w5_ro0w5o0w3o0w3o0w3o0w3 I78 (L346_0r0[4:0], L346_0r1[4:0], L346_0a, L237_0r, L237_0a, L237_0r, L237_0a, L257_0r, L257_0a, L279_0r, L279_0a, L305_0r, L305_0a, L331_0r, L331_0a, L238_0r0[4:0], L238_0r1[4:0], L238_0a, L258_0r0[2:0], L258_0r1[2:0], L258_0a, L280_0r0[2:0], L280_0r1[2:0], L280_0a, L306_0r0[2:0], L306_0r1[2:0], L306_0a, L332_0r0[2:0], L332_0r1[2:0], L332_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I79 (L235_0r0, L235_0r1, L235_0a, L236_0r, L236_0a, L348_0r, L348_0a, reset);
  tkm2x0b I80 (L236_0r, L236_0a, L345_0r, L345_0a, L349_0r, L349_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I81 (L350_0r, L350_0a, L2_0r, L2_0a, L118_0r, L118_0a, L234_0r, L234_0a, reset);
  tkj0m0_0_0 I82 (L117_0r, L117_0a, L233_0r, L233_0a, L349_0r, L349_0a, L352_0r, L352_0a, reset);
  tkf32mo0w0_o0w32 I83 (L360_0r0[31:0], L360_0r1[31:0], L360_0a, L361_0r, L361_0a, L377_0r0[31:0], L377_0r1[31:0], L377_0a, reset);
  tkj35m32_3 I84 (L377_0r0[31:0], L377_0r1[31:0], L377_0a, L362_0r0[2:0], L362_0r1[2:0], L362_0a, L378_0r0[34:0], L378_0r1[34:0], L378_0a, reset);
  tks35_o32w3_1o0w32_2o0w32_3o0w32_4o0w32_5o0w32_6o0w32_7o0w32 I85 (L378_0r0[34:0], L378_0r1[34:0], L378_0a, L363_0r0[31:0], L363_0r1[31:0], L363_0a, L365_0r0[31:0], L365_0r1[31:0], L365_0a, L367_0r0[31:0], L367_0r1[31:0], L367_0a, L369_0r0[31:0], L369_0r1[31:0], L369_0a, L371_0r0[31:0], L371_0r1[31:0], L371_0a, L373_0r0[31:0], L373_0r1[31:0], L373_0a, L375_0r0[31:0], L375_0r1[31:0], L375_0a, reset);
  tkm7x0b I86 (L364_0r, L364_0a, L366_0r, L366_0a, L368_0r, L368_0a, L370_0r, L370_0a, L372_0r, L372_0a, L374_0r, L374_0a, L376_0r, L376_0a, L379_0r, L379_0a, reset);
  tkj4m3_1 I87 (L385_0r0[2:0], L385_0r1[2:0], L385_0a, L387_0r0, L387_0r1, L387_0a, L388_0r0[3:0], L388_0r1[3:0], L388_0a, reset);
  tkf4mo0w3 I88 (L388_0r0[3:0], L388_0r1[3:0], L388_0a, L383_0r0[2:0], L383_0r1[2:0], L383_0a, reset);
  tkf0mo0w0_o0w0 I89 (L389_0r, L389_0a, L384_0r, L384_0a, L386_0r, L386_0a, reset);
  tkf32mo0w0_o0w32 I90 (L382_0r0[31:0], L382_0r1[31:0], L382_0a, L389_0r, L389_0a, L406_0r0[31:0], L406_0r1[31:0], L406_0a, reset);
  tkj35m32_3 I91 (L406_0r0[31:0], L406_0r1[31:0], L406_0a, L383_0r0[2:0], L383_0r1[2:0], L383_0a, L407_0r0[34:0], L407_0r1[34:0], L407_0a, reset);
  tks35_o32w3_0o0w32_1o0w32_2o0w32_3o0w32_4o0w32_5o0w32_6o0w32_7o0w32 I92 (L407_0r0[34:0], L407_0r1[34:0], L407_0a, L390_0r0[31:0], L390_0r1[31:0], L390_0a, L392_0r0[31:0], L392_0r1[31:0], L392_0a, L394_0r0[31:0], L394_0r1[31:0], L394_0a, L396_0r0[31:0], L396_0r1[31:0], L396_0a, L398_0r0[31:0], L398_0r1[31:0], L398_0a, L400_0r0[31:0], L400_0r1[31:0], L400_0a, L402_0r0[31:0], L402_0r1[31:0], L402_0a, L404_0r0[31:0], L404_0r1[31:0], L404_0a, reset);
  tkm8x0b I93 (L391_0r, L391_0a, L393_0r, L393_0a, L395_0r, L395_0a, L397_0r, L397_0a, L399_0r, L399_0a, L401_0r, L401_0a, L403_0r, L403_0a, L405_0r, L405_0a, L408_0r, L408_0a, reset);
  tkj4m3_1 I94 (L414_0r0[2:0], L414_0r1[2:0], L414_0a, L416_0r0, L416_0r1, L416_0a, L417_0r0[3:0], L417_0r1[3:0], L417_0a, reset);
  tkf4mo0w3 I95 (L417_0r0[3:0], L417_0r1[3:0], L417_0a, L412_0r0[2:0], L412_0r1[2:0], L412_0a, reset);
  tkf0mo0w0_o0w0 I96 (L418_0r, L418_0a, L413_0r, L413_0a, L415_0r, L415_0a, reset);
  tkf32mo0w0_o0w32 I97 (L411_0r0[31:0], L411_0r1[31:0], L411_0a, L418_0r, L418_0a, L435_0r0[31:0], L435_0r1[31:0], L435_0a, reset);
  tkj35m32_3 I98 (L435_0r0[31:0], L435_0r1[31:0], L435_0a, L412_0r0[2:0], L412_0r1[2:0], L412_0a, L436_0r0[34:0], L436_0r1[34:0], L436_0a, reset);
  tks35_o32w3_0o0w32_1o0w32_2o0w32_3o0w32_4o0w32_5o0w32_6o0w32_7o0w32 I99 (L436_0r0[34:0], L436_0r1[34:0], L436_0a, L419_0r0[31:0], L419_0r1[31:0], L419_0a, L421_0r0[31:0], L421_0r1[31:0], L421_0a, L423_0r0[31:0], L423_0r1[31:0], L423_0a, L425_0r0[31:0], L425_0r1[31:0], L425_0a, L427_0r0[31:0], L427_0r1[31:0], L427_0a, L429_0r0[31:0], L429_0r1[31:0], L429_0a, L431_0r0[31:0], L431_0r1[31:0], L431_0a, L433_0r0[31:0], L433_0r1[31:0], L433_0a, reset);
  tkm8x0b I100 (L420_0r, L420_0a, L422_0r, L422_0a, L424_0r, L424_0a, L426_0r, L426_0a, L428_0r, L428_0a, L430_0r, L430_0a, L432_0r, L432_0a, L434_0r, L434_0a, L437_0r, L437_0a, reset);
  tko0m1_1nm1b1 I101 (L447_0r, L447_0a, L448_0r0, L448_0r1, L448_0a, reset);
  tkj2m1_1 I102 (L446_0r0, L446_0r1, L446_0a, L448_0r0, L448_0r1, L448_0a, L449_0r0[1:0], L449_0r1[1:0], L449_0a, reset);
  tko2m2_1api0w1b_2api1w1b_3nm1b0_4apt1o0w1bt3o0w1b_5nm1b0_6apt2o0w1bt5o0w1b_7addt4o0w2bt6o0w2b I103 (L449_0r0[1:0], L449_0r1[1:0], L449_0a, L450_0r0[1:0], L450_0r1[1:0], L450_0a, reset);
  tkf2mo0w1 I104 (L450_0r0[1:0], L450_0r1[1:0], L450_0a, L444_0r0, L444_0r1, L444_0a, reset);
  tkj4m3_1 I105 (L443_0r0[2:0], L443_0r1[2:0], L443_0a, L444_0r0, L444_0r1, L444_0a, L451_0r0[3:0], L451_0r1[3:0], L451_0a, reset);
  tkf4mo0w3 I106 (L451_0r0[3:0], L451_0r1[3:0], L451_0a, L441_0r0[2:0], L441_0r1[2:0], L441_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I107 (L452_0r, L452_0a, L442_0r, L442_0a, L445_0r, L445_0a, L447_0r, L447_0a, reset);
  tkf32mo0w0_o0w32 I108 (L440_0r0[31:0], L440_0r1[31:0], L440_0a, L452_0r, L452_0a, L469_0r0[31:0], L469_0r1[31:0], L469_0a, reset);
  tkj35m32_3 I109 (L469_0r0[31:0], L469_0r1[31:0], L469_0a, L441_0r0[2:0], L441_0r1[2:0], L441_0a, L470_0r0[34:0], L470_0r1[34:0], L470_0a, reset);
  tks35_o32w3_0o0w32_1o0w32_2o0w32_3o0w32_4o0w32_5o0w32_6o0w32_7o0w32 I110 (L470_0r0[34:0], L470_0r1[34:0], L470_0a, L453_0r0[31:0], L453_0r1[31:0], L453_0a, L455_0r0[31:0], L455_0r1[31:0], L455_0a, L457_0r0[31:0], L457_0r1[31:0], L457_0a, L459_0r0[31:0], L459_0r1[31:0], L459_0a, L461_0r0[31:0], L461_0r1[31:0], L461_0a, L463_0r0[31:0], L463_0r1[31:0], L463_0a, L465_0r0[31:0], L465_0r1[31:0], L465_0a, L467_0r0[31:0], L467_0r1[31:0], L467_0a, reset);
  tkm8x0b I111 (L454_0r, L454_0a, L456_0r, L456_0a, L458_0r, L458_0a, L460_0r, L460_0a, L462_0r, L462_0a, L464_0r, L464_0a, L466_0r, L466_0a, L468_0r, L468_0a, L471_0r, L471_0a, reset);
  tks5_o0w5_0o0w0_1m2c1m4c3o0w0_8c7o0w0_10c7o0w0_18c7o0w0 I112 (L356_0r0[4:0], L356_0r1[4:0], L356_0a, L357_0r, L357_0a, L358_0r, L358_0a, L380_0r, L380_0a, L409_0r, L409_0a, L438_0r, L438_0a, reset);
  tkm5x0b I113 (L357_0r, L357_0a, L379_0r, L379_0a, L408_0r, L408_0a, L437_0r, L437_0a, L471_0r, L471_0a, L472_0r, L472_0a, reset);
  tkvsel5_wo0w5_ro0w5o0w3o0w3o0w3o0w3 I114 (L473_0r0[4:0], L473_0r1[4:0], L473_0a, L474_0r, L474_0a, L355_0r, L355_0a, L361_0r, L361_0a, L384_0r, L384_0a, L413_0r, L413_0a, L442_0r, L442_0a, L356_0r0[4:0], L356_0r1[4:0], L356_0a, L362_0r0[2:0], L362_0r1[2:0], L362_0a, L385_0r0[2:0], L385_0r1[2:0], L385_0a, L414_0r0[2:0], L414_0r1[2:0], L414_0a, L443_0r0[2:0], L443_0r1[2:0], L443_0a, reset);
  tkvw32_wo0w32_ro0w32o0w32o0w32o0w32 I115 (L475_0r0[31:0], L475_0r1[31:0], L475_0a, L476_0r, L476_0a, L358_0r, L358_0a, L380_0r, L380_0a, L409_0r, L409_0a, L438_0r, L438_0a, L360_0r0[31:0], L360_0r1[31:0], L360_0a, L382_0r0[31:0], L382_0r1[31:0], L382_0a, L411_0r0[31:0], L411_0r1[31:0], L411_0a, L440_0r0[31:0], L440_0r1[31:0], L440_0a, reset);
  tkj0m0_0 I116 (L474_0r, L474_0a, L476_0r, L476_0a, L355_0r, L355_0a, reset);
  tkf0mo0w0_o0w0 I117 (L480_0r, L480_0a, L478_0r, L478_0a, L479_0r, L479_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I118 (L353_0r0, L353_0r1, L353_0a, L354_0r, L354_0a, L480_0r, L480_0a, reset);
  tkm2x0b I119 (L354_0r, L354_0a, L472_0r, L472_0a, L481_0r, L481_0a, reset);
  tkvwindow1_wo0w1_ro0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1 I120 (L482_0r0, L482_0r1, L482_0a, L483_0r, L483_0a, L49_0r, L49_0a, L75_0r, L75_0a, L102_0r, L102_0a, L165_0r, L165_0a, L191_0r, L191_0a, L218_0r, L218_0a, L281_0r, L281_0a, L307_0r, L307_0a, L334_0r, L334_0a, L386_0r, L386_0a, L415_0r, L415_0a, L445_0r, L445_0a, L50_0r0, L50_0r1, L50_0a, L76_0r0, L76_0r1, L76_0a, L103_0r0, L103_0r1, L103_0a, L166_0r0, L166_0r1, L166_0a, L192_0r0, L192_0r1, L192_0a, L219_0r0, L219_0r1, L219_0a, L282_0r0, L282_0r1, L282_0a, L308_0r0, L308_0r1, L308_0a, L335_0r0, L335_0r1, L335_0a, L387_0r0, L387_0r1, L387_0a, L416_0r0, L416_0r1, L416_0a, L446_0r0, L446_0r1, L446_0a, reset);
  tkvrEn3_wo0w3_ro0w1o1w1o2w1 I121 (L484_0r0[2:0], L484_0r1[2:0], L484_0a, L485_0r, L485_0a, L2_0r, L2_0a, L118_0r, L118_0a, L234_0r, L234_0a, L3_0r0, L3_0r1, L3_0a, L119_0r0, L119_0r1, L119_0a, L235_0r0, L235_0r1, L235_0a, reset);
  tkvwEn1_wo0w1_ro0w1 I122 (L486_0r0, L486_0r1, L486_0a, L487_0r, L487_0a, L352_0r, L352_0a, L353_0r0, L353_0r1, L353_0a, reset);
  tkj0m0_0_0 I123 (L483_0r, L483_0a, L485_0r, L485_0a, L487_0r, L487_0a, L350_0r, L350_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I124 (L492_0r, L492_0a, L489_0r, L489_0a, L490_0r, L490_0a, L491_0r, L491_0a, reset);
  tkf32mo0w0_o0w32 I125 (L453_0r0[31:0], L453_0r1[31:0], L453_0a, L496_0r, L496_0a, L497_0r0[31:0], L497_0r1[31:0], L497_0a, reset);
  tkf32mo0w0_o0w32 I126 (L390_0r0[31:0], L390_0r1[31:0], L390_0a, L498_0r, L498_0a, L499_0r0[31:0], L499_0r1[31:0], L499_0a, reset);
  tkm2x32b I127 (L497_0r0[31:0], L497_0r1[31:0], L497_0a, L499_0r0[31:0], L499_0r1[31:0], L499_0a, L494_0r0[31:0], L494_0r1[31:0], L494_0a, reset);
  tko0m2_1nm2b1 I128 (L496_0r, L496_0a, L500_0r0[1:0], L500_0r1[1:0], L500_0a, reset);
  tko0m2_1nm2b2 I129 (L498_0r, L498_0a, L501_0r0[1:0], L501_0r1[1:0], L501_0a, reset);
  tkm2x2b I130 (L500_0r0[1:0], L500_0r1[1:0], L500_0a, L501_0r0[1:0], L501_0r1[1:0], L501_0a, L502_0r0[1:0], L502_0r1[1:0], L502_0a, reset);
  tkj2m0_2 I131 (L495_0r, L495_0a, L502_0r0[1:0], L502_0r1[1:0], L502_0a, L503_0r0[1:0], L503_0r1[1:0], L503_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I132 (L503_0r0[1:0], L503_0r1[1:0], L503_0a, L454_0r, L454_0a, L391_0r, L391_0a, reset);
  tkvinouts_31032_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 I133 (L494_0r0[31:0], L494_0r1[31:0], L494_0a, L495_0r, L495_0a, L314_0r, L314_0a, L262_0r, L262_0a, L198_0r, L198_0a, L146_0r, L146_0a, L82_0r, L82_0a, L30_0r, L30_0a, L315_0r0[31:0], L315_0r1[31:0], L315_0a, L263_0r0[31:0], L263_0r1[31:0], L263_0a, L199_0r0[31:0], L199_0r1[31:0], L199_0a, L147_0r0[31:0], L147_0r1[31:0], L147_0a, L83_0r0[31:0], L83_0r1[31:0], L83_0a, L31_0r0[31:0], L31_0r1[31:0], L31_0a, reset);
  tkf32mo0w0_o0w32 I134 (L455_0r0[31:0], L455_0r1[31:0], L455_0a, L506_0r, L506_0a, L507_0r0[31:0], L507_0r1[31:0], L507_0a, reset);
  tkf32mo0w0_o0w32 I135 (L392_0r0[31:0], L392_0r1[31:0], L392_0a, L508_0r, L508_0a, L509_0r0[31:0], L509_0r1[31:0], L509_0a, reset);
  tkm2x32b I136 (L507_0r0[31:0], L507_0r1[31:0], L507_0a, L509_0r0[31:0], L509_0r1[31:0], L509_0a, L504_0r0[31:0], L504_0r1[31:0], L504_0a, reset);
  tko0m2_1nm2b1 I137 (L506_0r, L506_0a, L510_0r0[1:0], L510_0r1[1:0], L510_0a, reset);
  tko0m2_1nm2b2 I138 (L508_0r, L508_0a, L511_0r0[1:0], L511_0r1[1:0], L511_0a, reset);
  tkm2x2b I139 (L510_0r0[1:0], L510_0r1[1:0], L510_0a, L511_0r0[1:0], L511_0r1[1:0], L511_0a, L512_0r0[1:0], L512_0r1[1:0], L512_0a, reset);
  tkj2m0_2 I140 (L505_0r, L505_0a, L512_0r0[1:0], L512_0r1[1:0], L512_0a, L513_0r0[1:0], L513_0r1[1:0], L513_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I141 (L513_0r0[1:0], L513_0r1[1:0], L513_0a, L456_0r, L456_0a, L393_0r, L393_0a, reset);
  tkvinouts_633232_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 I142 (L504_0r0[31:0], L504_0r1[31:0], L504_0a, L505_0r, L505_0a, L316_0r, L316_0a, L264_0r, L264_0a, L200_0r, L200_0a, L148_0r, L148_0a, L84_0r, L84_0a, L32_0r, L32_0a, L317_0r0[31:0], L317_0r1[31:0], L317_0a, L265_0r0[31:0], L265_0r1[31:0], L265_0a, L201_0r0[31:0], L201_0r1[31:0], L201_0a, L149_0r0[31:0], L149_0r1[31:0], L149_0a, L85_0r0[31:0], L85_0r1[31:0], L85_0a, L33_0r0[31:0], L33_0r1[31:0], L33_0a, reset);
  tkf32mo0w0_o0w32 I143 (L457_0r0[31:0], L457_0r1[31:0], L457_0a, L516_0r, L516_0a, L517_0r0[31:0], L517_0r1[31:0], L517_0a, reset);
  tkf32mo0w0_o0w32 I144 (L394_0r0[31:0], L394_0r1[31:0], L394_0a, L518_0r, L518_0a, L519_0r0[31:0], L519_0r1[31:0], L519_0a, reset);
  tkm2x32b I145 (L517_0r0[31:0], L517_0r1[31:0], L517_0a, L519_0r0[31:0], L519_0r1[31:0], L519_0a, L514_0r0[31:0], L514_0r1[31:0], L514_0a, reset);
  tko0m2_1nm2b1 I146 (L516_0r, L516_0a, L520_0r0[1:0], L520_0r1[1:0], L520_0a, reset);
  tko0m2_1nm2b2 I147 (L518_0r, L518_0a, L521_0r0[1:0], L521_0r1[1:0], L521_0a, reset);
  tkm2x2b I148 (L520_0r0[1:0], L520_0r1[1:0], L520_0a, L521_0r0[1:0], L521_0r1[1:0], L521_0a, L522_0r0[1:0], L522_0r1[1:0], L522_0a, reset);
  tkj2m0_2 I149 (L515_0r, L515_0a, L522_0r0[1:0], L522_0r1[1:0], L522_0a, L523_0r0[1:0], L523_0r1[1:0], L523_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I150 (L523_0r0[1:0], L523_0r1[1:0], L523_0a, L458_0r, L458_0a, L395_0r, L395_0a, reset);
  tkvinouts_956432_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 I151 (L514_0r0[31:0], L514_0r1[31:0], L514_0a, L515_0r, L515_0a, L318_0r, L318_0a, L266_0r, L266_0a, L202_0r, L202_0a, L150_0r, L150_0a, L86_0r, L86_0a, L34_0r, L34_0a, L319_0r0[31:0], L319_0r1[31:0], L319_0a, L267_0r0[31:0], L267_0r1[31:0], L267_0a, L203_0r0[31:0], L203_0r1[31:0], L203_0a, L151_0r0[31:0], L151_0r1[31:0], L151_0a, L87_0r0[31:0], L87_0r1[31:0], L87_0a, L35_0r0[31:0], L35_0r1[31:0], L35_0a, reset);
  tkf32mo0w0_o0w32 I152 (L459_0r0[31:0], L459_0r1[31:0], L459_0a, L526_0r, L526_0a, L527_0r0[31:0], L527_0r1[31:0], L527_0a, reset);
  tkf32mo0w0_o0w32 I153 (L396_0r0[31:0], L396_0r1[31:0], L396_0a, L528_0r, L528_0a, L529_0r0[31:0], L529_0r1[31:0], L529_0a, reset);
  tkm2x32b I154 (L527_0r0[31:0], L527_0r1[31:0], L527_0a, L529_0r0[31:0], L529_0r1[31:0], L529_0a, L524_0r0[31:0], L524_0r1[31:0], L524_0a, reset);
  tko0m2_1nm2b1 I155 (L526_0r, L526_0a, L530_0r0[1:0], L530_0r1[1:0], L530_0a, reset);
  tko0m2_1nm2b2 I156 (L528_0r, L528_0a, L531_0r0[1:0], L531_0r1[1:0], L531_0a, reset);
  tkm2x2b I157 (L530_0r0[1:0], L530_0r1[1:0], L530_0a, L531_0r0[1:0], L531_0r1[1:0], L531_0a, L532_0r0[1:0], L532_0r1[1:0], L532_0a, reset);
  tkj2m0_2 I158 (L525_0r, L525_0a, L532_0r0[1:0], L532_0r1[1:0], L532_0a, L533_0r0[1:0], L533_0r1[1:0], L533_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I159 (L533_0r0[1:0], L533_0r1[1:0], L533_0a, L460_0r, L460_0a, L397_0r, L397_0a, reset);
  tkvinouts_1279632_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 I160 (L524_0r0[31:0], L524_0r1[31:0], L524_0a, L525_0r, L525_0a, L320_0r, L320_0a, L268_0r, L268_0a, L204_0r, L204_0a, L152_0r, L152_0a, L88_0r, L88_0a, L36_0r, L36_0a, L321_0r0[31:0], L321_0r1[31:0], L321_0a, L269_0r0[31:0], L269_0r1[31:0], L269_0a, L205_0r0[31:0], L205_0r1[31:0], L205_0a, L153_0r0[31:0], L153_0r1[31:0], L153_0a, L89_0r0[31:0], L89_0r1[31:0], L89_0a, L37_0r0[31:0], L37_0r1[31:0], L37_0a, reset);
  tkf32mo0w0_o0w32 I161 (L461_0r0[31:0], L461_0r1[31:0], L461_0a, L536_0r, L536_0a, L537_0r0[31:0], L537_0r1[31:0], L537_0a, reset);
  tkf32mo0w0_o0w32 I162 (L398_0r0[31:0], L398_0r1[31:0], L398_0a, L538_0r, L538_0a, L539_0r0[31:0], L539_0r1[31:0], L539_0a, reset);
  tkm2x32b I163 (L537_0r0[31:0], L537_0r1[31:0], L537_0a, L539_0r0[31:0], L539_0r1[31:0], L539_0a, L534_0r0[31:0], L534_0r1[31:0], L534_0a, reset);
  tko0m2_1nm2b1 I164 (L536_0r, L536_0a, L540_0r0[1:0], L540_0r1[1:0], L540_0a, reset);
  tko0m2_1nm2b2 I165 (L538_0r, L538_0a, L541_0r0[1:0], L541_0r1[1:0], L541_0a, reset);
  tkm2x2b I166 (L540_0r0[1:0], L540_0r1[1:0], L540_0a, L541_0r0[1:0], L541_0r1[1:0], L541_0a, L542_0r0[1:0], L542_0r1[1:0], L542_0a, reset);
  tkj2m0_2 I167 (L535_0r, L535_0a, L542_0r0[1:0], L542_0r1[1:0], L542_0a, L543_0r0[1:0], L543_0r1[1:0], L543_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I168 (L543_0r0[1:0], L543_0r1[1:0], L543_0a, L462_0r, L462_0a, L399_0r, L399_0a, reset);
  tkvinouts_15912832_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 I169 (L534_0r0[31:0], L534_0r1[31:0], L534_0a, L535_0r, L535_0a, L322_0r, L322_0a, L270_0r, L270_0a, L206_0r, L206_0a, L154_0r, L154_0a, L90_0r, L90_0a, L38_0r, L38_0a, L323_0r0[31:0], L323_0r1[31:0], L323_0a, L271_0r0[31:0], L271_0r1[31:0], L271_0a, L207_0r0[31:0], L207_0r1[31:0], L207_0a, L155_0r0[31:0], L155_0r1[31:0], L155_0a, L91_0r0[31:0], L91_0r1[31:0], L91_0a, L39_0r0[31:0], L39_0r1[31:0], L39_0a, reset);
  tkf32mo0w0_o0w32 I170 (L463_0r0[31:0], L463_0r1[31:0], L463_0a, L546_0r, L546_0a, L547_0r0[31:0], L547_0r1[31:0], L547_0a, reset);
  tkf32mo0w0_o0w32 I171 (L400_0r0[31:0], L400_0r1[31:0], L400_0a, L548_0r, L548_0a, L549_0r0[31:0], L549_0r1[31:0], L549_0a, reset);
  tkm2x32b I172 (L547_0r0[31:0], L547_0r1[31:0], L547_0a, L549_0r0[31:0], L549_0r1[31:0], L549_0a, L544_0r0[31:0], L544_0r1[31:0], L544_0a, reset);
  tko0m2_1nm2b1 I173 (L546_0r, L546_0a, L550_0r0[1:0], L550_0r1[1:0], L550_0a, reset);
  tko0m2_1nm2b2 I174 (L548_0r, L548_0a, L551_0r0[1:0], L551_0r1[1:0], L551_0a, reset);
  tkm2x2b I175 (L550_0r0[1:0], L550_0r1[1:0], L550_0a, L551_0r0[1:0], L551_0r1[1:0], L551_0a, L552_0r0[1:0], L552_0r1[1:0], L552_0a, reset);
  tkj2m0_2 I176 (L545_0r, L545_0a, L552_0r0[1:0], L552_0r1[1:0], L552_0a, L553_0r0[1:0], L553_0r1[1:0], L553_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I177 (L553_0r0[1:0], L553_0r1[1:0], L553_0a, L464_0r, L464_0a, L401_0r, L401_0a, reset);
  tkvinouts_19116032_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 I178 (L544_0r0[31:0], L544_0r1[31:0], L544_0a, L545_0r, L545_0a, L324_0r, L324_0a, L272_0r, L272_0a, L208_0r, L208_0a, L156_0r, L156_0a, L92_0r, L92_0a, L40_0r, L40_0a, L325_0r0[31:0], L325_0r1[31:0], L325_0a, L273_0r0[31:0], L273_0r1[31:0], L273_0a, L209_0r0[31:0], L209_0r1[31:0], L209_0a, L157_0r0[31:0], L157_0r1[31:0], L157_0a, L93_0r0[31:0], L93_0r1[31:0], L93_0a, L41_0r0[31:0], L41_0r1[31:0], L41_0a, reset);
  tkf32mo0w0_o0w32 I179 (L465_0r0[31:0], L465_0r1[31:0], L465_0a, L556_0r, L556_0a, L557_0r0[31:0], L557_0r1[31:0], L557_0a, reset);
  tkf32mo0w0_o0w32 I180 (L402_0r0[31:0], L402_0r1[31:0], L402_0a, L558_0r, L558_0a, L559_0r0[31:0], L559_0r1[31:0], L559_0a, reset);
  tkm2x32b I181 (L557_0r0[31:0], L557_0r1[31:0], L557_0a, L559_0r0[31:0], L559_0r1[31:0], L559_0a, L554_0r0[31:0], L554_0r1[31:0], L554_0a, reset);
  tko0m2_1nm2b1 I182 (L556_0r, L556_0a, L560_0r0[1:0], L560_0r1[1:0], L560_0a, reset);
  tko0m2_1nm2b2 I183 (L558_0r, L558_0a, L561_0r0[1:0], L561_0r1[1:0], L561_0a, reset);
  tkm2x2b I184 (L560_0r0[1:0], L560_0r1[1:0], L560_0a, L561_0r0[1:0], L561_0r1[1:0], L561_0a, L562_0r0[1:0], L562_0r1[1:0], L562_0a, reset);
  tkj2m0_2 I185 (L555_0r, L555_0a, L562_0r0[1:0], L562_0r1[1:0], L562_0a, L563_0r0[1:0], L563_0r1[1:0], L563_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I186 (L563_0r0[1:0], L563_0r1[1:0], L563_0a, L466_0r, L466_0a, L403_0r, L403_0a, reset);
  tkvinouts_22319232_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 I187 (L554_0r0[31:0], L554_0r1[31:0], L554_0a, L555_0r, L555_0a, L326_0r, L326_0a, L274_0r, L274_0a, L210_0r, L210_0a, L158_0r, L158_0a, L94_0r, L94_0a, L42_0r, L42_0a, L327_0r0[31:0], L327_0r1[31:0], L327_0a, L275_0r0[31:0], L275_0r1[31:0], L275_0a, L211_0r0[31:0], L211_0r1[31:0], L211_0a, L159_0r0[31:0], L159_0r1[31:0], L159_0a, L95_0r0[31:0], L95_0r1[31:0], L95_0a, L43_0r0[31:0], L43_0r1[31:0], L43_0a, reset);
  tkf32mo0w0_o0w32 I188 (L467_0r0[31:0], L467_0r1[31:0], L467_0a, L566_0r, L566_0a, L567_0r0[31:0], L567_0r1[31:0], L567_0a, reset);
  tkf32mo0w0_o0w32 I189 (L404_0r0[31:0], L404_0r1[31:0], L404_0a, L568_0r, L568_0a, L569_0r0[31:0], L569_0r1[31:0], L569_0a, reset);
  tkm2x32b I190 (L567_0r0[31:0], L567_0r1[31:0], L567_0a, L569_0r0[31:0], L569_0r1[31:0], L569_0a, L564_0r0[31:0], L564_0r1[31:0], L564_0a, reset);
  tko0m2_1nm2b1 I191 (L566_0r, L566_0a, L570_0r0[1:0], L570_0r1[1:0], L570_0a, reset);
  tko0m2_1nm2b2 I192 (L568_0r, L568_0a, L571_0r0[1:0], L571_0r1[1:0], L571_0a, reset);
  tkm2x2b I193 (L570_0r0[1:0], L570_0r1[1:0], L570_0a, L571_0r0[1:0], L571_0r1[1:0], L571_0a, L572_0r0[1:0], L572_0r1[1:0], L572_0a, reset);
  tkj2m0_2 I194 (L565_0r, L565_0a, L572_0r0[1:0], L572_0r1[1:0], L572_0a, L573_0r0[1:0], L573_0r1[1:0], L573_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I195 (L573_0r0[1:0], L573_0r1[1:0], L573_0a, L468_0r, L468_0a, L405_0r, L405_0a, reset);
  tkvinouts_25522432_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32 I196 (L564_0r0[31:0], L564_0r1[31:0], L564_0a, L565_0r, L565_0a, L328_0r, L328_0a, L276_0r, L276_0a, L212_0r, L212_0a, L160_0r, L160_0a, L96_0r, L96_0a, L44_0r, L44_0a, L329_0r0[31:0], L329_0r1[31:0], L329_0a, L277_0r0[31:0], L277_0r1[31:0], L277_0a, L213_0r0[31:0], L213_0r1[31:0], L213_0a, L161_0r0[31:0], L161_0r1[31:0], L161_0a, L97_0r0[31:0], L97_0r1[31:0], L97_0a, L45_0r0[31:0], L45_0r1[31:0], L45_0a, reset);
  tkvlocals_31032_wo0w32_ro0w32o0w32o0w32 I197 (L419_0r0[31:0], L419_0r1[31:0], L419_0a, L420_0r, L420_0a, L288_0r, L288_0a, L172_0r, L172_0a, L56_0r, L56_0a, L289_0r0[31:0], L289_0r1[31:0], L289_0a, L173_0r0[31:0], L173_0r1[31:0], L173_0a, L57_0r0[31:0], L57_0r1[31:0], L57_0a, reset);
  tkvlocals_633232_wo0w32_ro0w32o0w32o0w32 I198 (L421_0r0[31:0], L421_0r1[31:0], L421_0a, L422_0r, L422_0a, L290_0r, L290_0a, L174_0r, L174_0a, L58_0r, L58_0a, L291_0r0[31:0], L291_0r1[31:0], L291_0a, L175_0r0[31:0], L175_0r1[31:0], L175_0a, L59_0r0[31:0], L59_0r1[31:0], L59_0a, reset);
  tkvlocals_956432_wo0w32_ro0w32o0w32o0w32 I199 (L423_0r0[31:0], L423_0r1[31:0], L423_0a, L424_0r, L424_0a, L292_0r, L292_0a, L176_0r, L176_0a, L60_0r, L60_0a, L293_0r0[31:0], L293_0r1[31:0], L293_0a, L177_0r0[31:0], L177_0r1[31:0], L177_0a, L61_0r0[31:0], L61_0r1[31:0], L61_0a, reset);
  tkvlocals_1279632_wo0w32_ro0w32o0w32o0w32 I200 (L425_0r0[31:0], L425_0r1[31:0], L425_0a, L426_0r, L426_0a, L294_0r, L294_0a, L178_0r, L178_0a, L62_0r, L62_0a, L295_0r0[31:0], L295_0r1[31:0], L295_0a, L179_0r0[31:0], L179_0r1[31:0], L179_0a, L63_0r0[31:0], L63_0r1[31:0], L63_0a, reset);
  tkvlocals_15912832_wo0w32_ro0w32o0w32o0w32 I201 (L427_0r0[31:0], L427_0r1[31:0], L427_0a, L428_0r, L428_0a, L296_0r, L296_0a, L180_0r, L180_0a, L64_0r, L64_0a, L297_0r0[31:0], L297_0r1[31:0], L297_0a, L181_0r0[31:0], L181_0r1[31:0], L181_0a, L65_0r0[31:0], L65_0r1[31:0], L65_0a, reset);
  tkvlocals_19116032_wo0w32_ro0w32o0w32o0w32 I202 (L429_0r0[31:0], L429_0r1[31:0], L429_0a, L430_0r, L430_0a, L298_0r, L298_0a, L182_0r, L182_0a, L66_0r, L66_0a, L299_0r0[31:0], L299_0r1[31:0], L299_0a, L183_0r0[31:0], L183_0r1[31:0], L183_0a, L67_0r0[31:0], L67_0r1[31:0], L67_0a, reset);
  tkvlocals_22319232_wo0w32_ro0w32o0w32o0w32 I203 (L431_0r0[31:0], L431_0r1[31:0], L431_0a, L432_0r, L432_0a, L300_0r, L300_0a, L184_0r, L184_0a, L68_0r, L68_0a, L301_0r0[31:0], L301_0r1[31:0], L301_0a, L185_0r0[31:0], L185_0r1[31:0], L185_0a, L69_0r0[31:0], L69_0r1[31:0], L69_0a, reset);
  tkvlocals_25522432_wo0w32_ro0w32o0w32o0w32 I204 (L433_0r0[31:0], L433_0r1[31:0], L433_0a, L434_0r, L434_0a, L302_0r, L302_0a, L186_0r, L186_0a, L70_0r, L70_0a, L303_0r0[31:0], L303_0r1[31:0], L303_0a, L187_0r0[31:0], L187_0r1[31:0], L187_0a, L71_0r0[31:0], L71_0r1[31:0], L71_0a, reset);
  tkvglobals_31032_wo0w32_ro0w32o0w32o0w32 I205 (L363_0r0[31:0], L363_0r1[31:0], L363_0a, L364_0r, L364_0a, L243_0r, L243_0a, L127_0r, L127_0a, L11_0r, L11_0a, L244_0r0[31:0], L244_0r1[31:0], L244_0a, L128_0r0[31:0], L128_0r1[31:0], L128_0a, L12_0r0[31:0], L12_0r1[31:0], L12_0a, reset);
  tkvglobals_633232_wo0w32_ro0w32o0w32o0w32 I206 (L365_0r0[31:0], L365_0r1[31:0], L365_0a, L366_0r, L366_0a, L245_0r, L245_0a, L129_0r, L129_0a, L13_0r, L13_0a, L246_0r0[31:0], L246_0r1[31:0], L246_0a, L130_0r0[31:0], L130_0r1[31:0], L130_0a, L14_0r0[31:0], L14_0r1[31:0], L14_0a, reset);
  tkvglobals_956432_wo0w32_ro0w32o0w32o0w32 I207 (L367_0r0[31:0], L367_0r1[31:0], L367_0a, L368_0r, L368_0a, L247_0r, L247_0a, L131_0r, L131_0a, L15_0r, L15_0a, L248_0r0[31:0], L248_0r1[31:0], L248_0a, L132_0r0[31:0], L132_0r1[31:0], L132_0a, L16_0r0[31:0], L16_0r1[31:0], L16_0a, reset);
  tkvglobals_1279632_wo0w32_ro0w32o0w32o0w32 I208 (L369_0r0[31:0], L369_0r1[31:0], L369_0a, L370_0r, L370_0a, L249_0r, L249_0a, L133_0r, L133_0a, L17_0r, L17_0a, L250_0r0[31:0], L250_0r1[31:0], L250_0a, L134_0r0[31:0], L134_0r1[31:0], L134_0a, L18_0r0[31:0], L18_0r1[31:0], L18_0a, reset);
  tkvglobals_15912832_wo0w32_ro0w32o0w32o0w32 I209 (L371_0r0[31:0], L371_0r1[31:0], L371_0a, L372_0r, L372_0a, L251_0r, L251_0a, L135_0r, L135_0a, L19_0r, L19_0a, L252_0r0[31:0], L252_0r1[31:0], L252_0a, L136_0r0[31:0], L136_0r1[31:0], L136_0a, L20_0r0[31:0], L20_0r1[31:0], L20_0a, reset);
  tkvglobals_19116032_wo0w32_ro0w32o0w32o0w32 I210 (L373_0r0[31:0], L373_0r1[31:0], L373_0a, L374_0r, L374_0a, L253_0r, L253_0a, L137_0r, L137_0a, L21_0r, L21_0a, L254_0r0[31:0], L254_0r1[31:0], L254_0a, L138_0r0[31:0], L138_0r1[31:0], L138_0a, L22_0r0[31:0], L22_0r1[31:0], L22_0a, reset);
  tkvglobals_22319232_wo0w32_ro0w32o0w32o0w32 I211 (L375_0r0[31:0], L375_0r1[31:0], L375_0a, L376_0r, L376_0a, L255_0r, L255_0a, L139_0r, L139_0a, L23_0r, L23_0a, L256_0r0[31:0], L256_0r1[31:0], L256_0a, L140_0r0[31:0], L140_0r1[31:0], L140_0a, L24_0r0[31:0], L24_0r1[31:0], L24_0a, reset);
  tkj1m1_0 I212 (wEn_0r0, wEn_0r1, wEn_0a, L491_0r, L491_0a, L486_0r0, L486_0r1, L486_0a, reset);
  tkj3m3_0 I213 (rEn_0r0[2:0], rEn_0r1[2:0], rEn_0a, L490_0r, L490_0a, L484_0r0[2:0], L484_0r1[2:0], L484_0a, reset);
  tkj5m5_0 I214 (wSel_0r0[4:0], wSel_0r1[4:0], wSel_0a, L478_0r, L478_0a, L473_0r0[4:0], L473_0r1[4:0], L473_0a, reset);
  tkj5m5_0 I215 (r0Sel_0r0[4:0], r0Sel_0r1[4:0], r0Sel_0a, L116_0r, L116_0a, L114_0r0[4:0], L114_0r1[4:0], L114_0a, reset);
  tkj5m5_0 I216 (r1Sel_0r0[4:0], r1Sel_0r1[4:0], r1Sel_0a, L232_0r, L232_0a, L230_0r0[4:0], L230_0r1[4:0], L230_0a, reset);
  tkj5m5_0 I217 (r2Sel_0r0[4:0], r2Sel_0r1[4:0], r2Sel_0a, L348_0r, L348_0a, L346_0r0[4:0], L346_0r1[4:0], L346_0a, reset);
  tkj1m1_0 I218 (window_0r0, window_0r1, window_0a, L489_0r, L489_0a, L482_0r0, L482_0r1, L482_0a, reset);
  tkj32m32_0 I219 (w_0r0[31:0], w_0r1[31:0], w_0a, L479_0r, L479_0a, L475_0r0[31:0], L475_0r1[31:0], L475_0a, reset);
  tkf32mo0w0_o0w32 I220 (L9_0r0[31:0], L9_0r1[31:0], L9_0a, L582_0r, L582_0a, L583_0r0[31:0], L583_0r1[31:0], L583_0a, reset);
  tkf32mo0w0_o0w32 I221 (L28_0r0[31:0], L28_0r1[31:0], L28_0a, L584_0r, L584_0a, L585_0r0[31:0], L585_0r1[31:0], L585_0a, reset);
  tkf32mo0w0_o0w32 I222 (L54_0r0[31:0], L54_0r1[31:0], L54_0a, L586_0r, L586_0a, L587_0r0[31:0], L587_0r1[31:0], L587_0a, reset);
  tkf32mo0w0_o0w32 I223 (L80_0r0[31:0], L80_0r1[31:0], L80_0a, L588_0r, L588_0a, L589_0r0[31:0], L589_0r1[31:0], L589_0a, reset);
  tkf32mo0w0_o0w32 I224 (L111_0r0[31:0], L111_0r1[31:0], L111_0a, L590_0r, L590_0a, L591_0r0[31:0], L591_0r1[31:0], L591_0a, reset);
  tkm5x32b I225 (L583_0r0[31:0], L583_0r1[31:0], L583_0a, L585_0r0[31:0], L585_0r1[31:0], L585_0a, L587_0r0[31:0], L587_0r1[31:0], L587_0a, L589_0r0[31:0], L589_0r1[31:0], L589_0a, L591_0r0[31:0], L591_0r1[31:0], L591_0a, L592_0r0[31:0], L592_0r1[31:0], L592_0a, reset);
  tkf32mo0w0_o0w32 I226 (L592_0r0[31:0], L592_0r1[31:0], L592_0a, L593_0r, L593_0a, r0_0r0[31:0], r0_0r1[31:0], r0_0a, reset);
  tko0m5_1nm5b1 I227 (L582_0r, L582_0a, L595_0r0[4:0], L595_0r1[4:0], L595_0a, reset);
  tko0m5_1nm5b2 I228 (L584_0r, L584_0a, L596_0r0[4:0], L596_0r1[4:0], L596_0a, reset);
  tko0m5_1nm5b4 I229 (L586_0r, L586_0a, L597_0r0[4:0], L597_0r1[4:0], L597_0a, reset);
  tko0m5_1nm5b8 I230 (L588_0r, L588_0a, L598_0r0[4:0], L598_0r1[4:0], L598_0a, reset);
  tko0m5_1nm5b10 I231 (L590_0r, L590_0a, L599_0r0[4:0], L599_0r1[4:0], L599_0a, reset);
  tkm5x5b I232 (L595_0r0[4:0], L595_0r1[4:0], L595_0a, L596_0r0[4:0], L596_0r1[4:0], L596_0a, L597_0r0[4:0], L597_0r1[4:0], L597_0a, L598_0r0[4:0], L598_0r1[4:0], L598_0a, L599_0r0[4:0], L599_0r1[4:0], L599_0a, L600_0r0[4:0], L600_0r1[4:0], L600_0a, reset);
  tkj5m0_5 I233 (L593_0r, L593_0a, L600_0r0[4:0], L600_0r1[4:0], L600_0a, L601_0r0[4:0], L601_0r1[4:0], L601_0a, reset);
  tks5_o0w5_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0 I234 (L601_0r0[4:0], L601_0r1[4:0], L601_0a, L10_0r, L10_0a, L29_0r, L29_0a, L55_0r, L55_0a, L81_0r, L81_0a, L112_0r, L112_0a, reset);
  tkf32mo0w0_o0w32 I235 (L125_0r0[31:0], L125_0r1[31:0], L125_0a, L602_0r, L602_0a, L603_0r0[31:0], L603_0r1[31:0], L603_0a, reset);
  tkf32mo0w0_o0w32 I236 (L144_0r0[31:0], L144_0r1[31:0], L144_0a, L604_0r, L604_0a, L605_0r0[31:0], L605_0r1[31:0], L605_0a, reset);
  tkf32mo0w0_o0w32 I237 (L170_0r0[31:0], L170_0r1[31:0], L170_0a, L606_0r, L606_0a, L607_0r0[31:0], L607_0r1[31:0], L607_0a, reset);
  tkf32mo0w0_o0w32 I238 (L196_0r0[31:0], L196_0r1[31:0], L196_0a, L608_0r, L608_0a, L609_0r0[31:0], L609_0r1[31:0], L609_0a, reset);
  tkf32mo0w0_o0w32 I239 (L227_0r0[31:0], L227_0r1[31:0], L227_0a, L610_0r, L610_0a, L611_0r0[31:0], L611_0r1[31:0], L611_0a, reset);
  tkm5x32b I240 (L603_0r0[31:0], L603_0r1[31:0], L603_0a, L605_0r0[31:0], L605_0r1[31:0], L605_0a, L607_0r0[31:0], L607_0r1[31:0], L607_0a, L609_0r0[31:0], L609_0r1[31:0], L609_0a, L611_0r0[31:0], L611_0r1[31:0], L611_0a, L612_0r0[31:0], L612_0r1[31:0], L612_0a, reset);
  tkf32mo0w0_o0w32 I241 (L612_0r0[31:0], L612_0r1[31:0], L612_0a, L613_0r, L613_0a, r1_0r0[31:0], r1_0r1[31:0], r1_0a, reset);
  tko0m5_1nm5b1 I242 (L602_0r, L602_0a, L615_0r0[4:0], L615_0r1[4:0], L615_0a, reset);
  tko0m5_1nm5b2 I243 (L604_0r, L604_0a, L616_0r0[4:0], L616_0r1[4:0], L616_0a, reset);
  tko0m5_1nm5b4 I244 (L606_0r, L606_0a, L617_0r0[4:0], L617_0r1[4:0], L617_0a, reset);
  tko0m5_1nm5b8 I245 (L608_0r, L608_0a, L618_0r0[4:0], L618_0r1[4:0], L618_0a, reset);
  tko0m5_1nm5b10 I246 (L610_0r, L610_0a, L619_0r0[4:0], L619_0r1[4:0], L619_0a, reset);
  tkm5x5b I247 (L615_0r0[4:0], L615_0r1[4:0], L615_0a, L616_0r0[4:0], L616_0r1[4:0], L616_0a, L617_0r0[4:0], L617_0r1[4:0], L617_0a, L618_0r0[4:0], L618_0r1[4:0], L618_0a, L619_0r0[4:0], L619_0r1[4:0], L619_0a, L620_0r0[4:0], L620_0r1[4:0], L620_0a, reset);
  tkj5m0_5 I248 (L613_0r, L613_0a, L620_0r0[4:0], L620_0r1[4:0], L620_0a, L621_0r0[4:0], L621_0r1[4:0], L621_0a, reset);
  tks5_o0w5_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0 I249 (L621_0r0[4:0], L621_0r1[4:0], L621_0a, L126_0r, L126_0a, L145_0r, L145_0a, L171_0r, L171_0a, L197_0r, L197_0a, L228_0r, L228_0a, reset);
  tkf32mo0w0_o0w32 I250 (L241_0r0[31:0], L241_0r1[31:0], L241_0a, L622_0r, L622_0a, L623_0r0[31:0], L623_0r1[31:0], L623_0a, reset);
  tkf32mo0w0_o0w32 I251 (L260_0r0[31:0], L260_0r1[31:0], L260_0a, L624_0r, L624_0a, L625_0r0[31:0], L625_0r1[31:0], L625_0a, reset);
  tkf32mo0w0_o0w32 I252 (L286_0r0[31:0], L286_0r1[31:0], L286_0a, L626_0r, L626_0a, L627_0r0[31:0], L627_0r1[31:0], L627_0a, reset);
  tkf32mo0w0_o0w32 I253 (L312_0r0[31:0], L312_0r1[31:0], L312_0a, L628_0r, L628_0a, L629_0r0[31:0], L629_0r1[31:0], L629_0a, reset);
  tkf32mo0w0_o0w32 I254 (L343_0r0[31:0], L343_0r1[31:0], L343_0a, L630_0r, L630_0a, L631_0r0[31:0], L631_0r1[31:0], L631_0a, reset);
  tkm5x32b I255 (L623_0r0[31:0], L623_0r1[31:0], L623_0a, L625_0r0[31:0], L625_0r1[31:0], L625_0a, L627_0r0[31:0], L627_0r1[31:0], L627_0a, L629_0r0[31:0], L629_0r1[31:0], L629_0a, L631_0r0[31:0], L631_0r1[31:0], L631_0a, L632_0r0[31:0], L632_0r1[31:0], L632_0a, reset);
  tkf32mo0w0_o0w32 I256 (L632_0r0[31:0], L632_0r1[31:0], L632_0a, L633_0r, L633_0a, r2_0r0[31:0], r2_0r1[31:0], r2_0a, reset);
  tko0m5_1nm5b1 I257 (L622_0r, L622_0a, L635_0r0[4:0], L635_0r1[4:0], L635_0a, reset);
  tko0m5_1nm5b2 I258 (L624_0r, L624_0a, L636_0r0[4:0], L636_0r1[4:0], L636_0a, reset);
  tko0m5_1nm5b4 I259 (L626_0r, L626_0a, L637_0r0[4:0], L637_0r1[4:0], L637_0a, reset);
  tko0m5_1nm5b8 I260 (L628_0r, L628_0a, L638_0r0[4:0], L638_0r1[4:0], L638_0a, reset);
  tko0m5_1nm5b10 I261 (L630_0r, L630_0a, L639_0r0[4:0], L639_0r1[4:0], L639_0a, reset);
  tkm5x5b I262 (L635_0r0[4:0], L635_0r1[4:0], L635_0a, L636_0r0[4:0], L636_0r1[4:0], L636_0a, L637_0r0[4:0], L637_0r1[4:0], L637_0a, L638_0r0[4:0], L638_0r1[4:0], L638_0a, L639_0r0[4:0], L639_0r1[4:0], L639_0a, L640_0r0[4:0], L640_0r1[4:0], L640_0a, reset);
  tkj5m0_5 I263 (L633_0r, L633_0a, L640_0r0[4:0], L640_0r1[4:0], L640_0a, L641_0r0[4:0], L641_0r1[4:0], L641_0a, reset);
  tks5_o0w5_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0 I264 (L641_0r0[4:0], L641_0r1[4:0], L641_0a, L242_0r, L242_0a, L261_0r, L261_0a, L287_0r, L287_0a, L313_0r, L313_0a, L344_0r, L344_0a, reset);
  tki I265 (L481_0r, L481_0a, L492_0r, L492_0a, reset);
endmodule

module teak_ExecuteCtrl (op_0r0, op_0r1, op_0a, pc_0r0, pc_0r1, pc_0a, doFetch_0r0, doFetch_0r1, doFetch_0a, newPc_0r0, newPc_0r1, newPc_0a, wEn_0r0, wEn_0r1, wEn_0a, rEn_0r0, rEn_0r1, rEn_0a, wSel_0r0, wSel_0r1, wSel_0a, r0Sel_0r0, r0Sel_0r1, r0Sel_0a, r1Sel_0r0, r1Sel_0r1, r1Sel_0a, r2Sel_0r0, r2Sel_0r1, r2Sel_0a, window_0r0, window_0r1, window_0a, w_0r0, w_0r1, w_0a, r0_0r0, r0_0r1, r0_0a, r1_0r0, r1_0r1, r1_0a, r2_0r0, r2_0r1, r2_0a, aluOp_0r0, aluOp_0r1, aluOp_0a, aluResult_0r0, aluResult_0r1, aluResult_0a, aluFlags_0r0, aluFlags_0r1, aluFlags_0a, aluLhs_0r0, aluLhs_0r1, aluLhs_0a, aluRhs_0r0, aluRhs_0r1, aluRhs_0a, daddr_0r0, daddr_0r1, daddr_0a, daccess_0r0, daccess_0r1, daccess_0a, dread_0r0, dread_0r1, dread_0a, dwrite_0r0, dwrite_0r1, dwrite_0a, reset);
  input [73:0] op_0r0;
  input [73:0] op_0r1;
  output op_0a;
  input [32:0] pc_0r0;
  input [32:0] pc_0r1;
  output pc_0a;
  output doFetch_0r0;
  output doFetch_0r1;
  input doFetch_0a;
  output [31:0] newPc_0r0;
  output [31:0] newPc_0r1;
  input newPc_0a;
  output wEn_0r0;
  output wEn_0r1;
  input wEn_0a;
  output [2:0] rEn_0r0;
  output [2:0] rEn_0r1;
  input rEn_0a;
  output [4:0] wSel_0r0;
  output [4:0] wSel_0r1;
  input wSel_0a;
  output [4:0] r0Sel_0r0;
  output [4:0] r0Sel_0r1;
  input r0Sel_0a;
  output [4:0] r1Sel_0r0;
  output [4:0] r1Sel_0r1;
  input r1Sel_0a;
  output [4:0] r2Sel_0r0;
  output [4:0] r2Sel_0r1;
  input r2Sel_0a;
  output window_0r0;
  output window_0r1;
  input window_0a;
  output [31:0] w_0r0;
  output [31:0] w_0r1;
  input w_0a;
  input [31:0] r0_0r0;
  input [31:0] r0_0r1;
  output r0_0a;
  input [31:0] r1_0r0;
  input [31:0] r1_0r1;
  output r1_0a;
  input [31:0] r2_0r0;
  input [31:0] r2_0r1;
  output r2_0a;
  output [6:0] aluOp_0r0;
  output [6:0] aluOp_0r1;
  input aluOp_0a;
  input [31:0] aluResult_0r0;
  input [31:0] aluResult_0r1;
  output aluResult_0a;
  input [3:0] aluFlags_0r0;
  input [3:0] aluFlags_0r1;
  output aluFlags_0a;
  output [31:0] aluLhs_0r0;
  output [31:0] aluLhs_0r1;
  input aluLhs_0a;
  output [31:0] aluRhs_0r0;
  output [31:0] aluRhs_0r1;
  input aluRhs_0a;
  output [31:0] daddr_0r0;
  output [31:0] daddr_0r1;
  input daddr_0a;
  output [2:0] daccess_0r0;
  output [2:0] daccess_0r1;
  input daccess_0a;
  input [31:0] dread_0r0;
  input [31:0] dread_0r1;
  output dread_0a;
  output [31:0] dwrite_0r0;
  output [31:0] dwrite_0r1;
  input dwrite_0a;
  input reset;
  wire L2_0r;
  wire L2_0a;
  wire L4_0r0;
  wire L4_0r1;
  wire L4_0a;
  wire L5_0r;
  wire L5_0a;
  wire L6_0r;
  wire L6_0a;
  wire [3:0] L8_0r0;
  wire [3:0] L8_0r1;
  wire L8_0a;
  wire L9_0r;
  wire L9_0a;
  wire L10_0r;
  wire L10_0a;
  wire L12_0r0;
  wire L12_0r1;
  wire L12_0a;
  wire L13_0r;
  wire L13_0a;
  wire L14_0r;
  wire L14_0a;
  wire L16_0r0;
  wire L16_0r1;
  wire L16_0a;
  wire L17_0r;
  wire L17_0a;
  wire L23_0r;
  wire L23_0a;
  wire L25_0r;
  wire L25_0a;
  wire L26_0r;
  wire L26_0a;
  wire L27_0r0;
  wire L27_0r1;
  wire L27_0a;
  wire L28_0r0;
  wire L28_0r1;
  wire L28_0a;
  wire L29_0r;
  wire L29_0a;
  wire L30_0r0;
  wire L30_0r1;
  wire L30_0a;
  wire [1:0] L31_0r0;
  wire [1:0] L31_0r1;
  wire L31_0a;
  wire L32_0r0;
  wire L32_0r1;
  wire L32_0a;
  wire L33_0r;
  wire L33_0a;
  wire L34_0r;
  wire L34_0a;
  wire L36_0r0;
  wire L36_0r1;
  wire L36_0a;
  wire L37_0r;
  wire L37_0a;
  wire L38_0r;
  wire L38_0a;
  wire L40_0r0;
  wire L40_0r1;
  wire L40_0a;
  wire L41_0r;
  wire L41_0a;
  wire L42_0r;
  wire L42_0a;
  wire L44_0r;
  wire L44_0a;
  wire L46_0r0;
  wire L46_0r1;
  wire L46_0a;
  wire L48_0r;
  wire L48_0a;
  wire [2:0] L49_0r0;
  wire [2:0] L49_0r1;
  wire L49_0a;
  wire L50_0r;
  wire L50_0a;
  wire L51_0r;
  wire L51_0a;
  wire L52_0r;
  wire L52_0a;
  wire L53_0r;
  wire L53_0a;
  wire L54_0r;
  wire L54_0a;
  wire L55_0r;
  wire L55_0a;
  wire L57_0r;
  wire L57_0a;
  wire [3:0] L58_0r0;
  wire [3:0] L58_0r1;
  wire L58_0a;
  wire L59_0r;
  wire L59_0a;
  wire L61_0r0;
  wire L61_0r1;
  wire L61_0a;
  wire L62_0r;
  wire L62_0a;
  wire L63_0r;
  wire L63_0a;
  wire L65_0r0;
  wire L65_0r1;
  wire L65_0a;
  wire L66_0r;
  wire L66_0a;
  wire L67_0r;
  wire L67_0a;
  wire L68_0r0;
  wire L68_0r1;
  wire L68_0a;
  wire L69_0r;
  wire L69_0a;
  wire L70_0r0;
  wire L70_0r1;
  wire L70_0a;
  wire L71_0r;
  wire L71_0a;
  wire L72_0r0;
  wire L72_0r1;
  wire L72_0a;
  wire [1:0] L73_0r0;
  wire [1:0] L73_0r1;
  wire L73_0a;
  wire L74_0r0;
  wire L74_0r1;
  wire L74_0a;
  wire [1:0] L75_0r0;
  wire [1:0] L75_0r1;
  wire L75_0a;
  wire L77_0r;
  wire L77_0a;
  wire L78_0r0;
  wire L78_0r1;
  wire L78_0a;
  wire L79_0r;
  wire L79_0a;
  wire L80_0r;
  wire L80_0a;
  wire L81_0r0;
  wire L81_0r1;
  wire L81_0a;
  wire L82_0r;
  wire L82_0a;
  wire L83_0r0;
  wire L83_0r1;
  wire L83_0a;
  wire [1:0] L84_0r0;
  wire [1:0] L84_0r1;
  wire L84_0a;
  wire L86_0r;
  wire L86_0a;
  wire L87_0r0;
  wire L87_0r1;
  wire L87_0a;
  wire L88_0r;
  wire L88_0a;
  wire L89_0r;
  wire L89_0a;
  wire L90_0r0;
  wire L90_0r1;
  wire L90_0a;
  wire L91_0r;
  wire L91_0a;
  wire L92_0r0;
  wire L92_0r1;
  wire L92_0a;
  wire [1:0] L93_0r0;
  wire [1:0] L93_0r1;
  wire L93_0a;
  wire L95_0r;
  wire L95_0a;
  wire L96_0r0;
  wire L96_0r1;
  wire L96_0a;
  wire L97_0r;
  wire L97_0a;
  wire L98_0r;
  wire L98_0a;
  wire L100_0r0;
  wire L100_0r1;
  wire L100_0a;
  wire L101_0r;
  wire L101_0a;
  wire L102_0r;
  wire L102_0a;
  wire L104_0r0;
  wire L104_0r1;
  wire L104_0a;
  wire L105_0r;
  wire L105_0a;
  wire L106_0r;
  wire L106_0a;
  wire L108_0r0;
  wire L108_0r1;
  wire L108_0a;
  wire L109_0r;
  wire L109_0a;
  wire L110_0r;
  wire L110_0a;
  wire L112_0r;
  wire L112_0a;
  wire L113_0r0;
  wire L113_0r1;
  wire L113_0a;
  wire L114_0r;
  wire L114_0a;
  wire L115_0r0;
  wire L115_0r1;
  wire L115_0a;
  wire [1:0] L116_0r0;
  wire [1:0] L116_0r1;
  wire L116_0a;
  wire L118_0r;
  wire L118_0a;
  wire L119_0r0;
  wire L119_0r1;
  wire L119_0a;
  wire L121_0r;
  wire L121_0a;
  wire L122_0r0;
  wire L122_0r1;
  wire L122_0a;
  wire L123_0r;
  wire L123_0a;
  wire L124_0r;
  wire L124_0a;
  wire L127_0r;
  wire L127_0a;
  wire [31:0] L128_0r0;
  wire [31:0] L128_0r1;
  wire L128_0a;
  wire L129_0r;
  wire L129_0a;
  wire [31:0] L130_0r0;
  wire [31:0] L130_0r1;
  wire L130_0a;
  wire [63:0] L131_0r0;
  wire [63:0] L131_0r1;
  wire L131_0a;
  wire [32:0] L132_0r0;
  wire [32:0] L132_0r1;
  wire L132_0a;
  wire L133_0r;
  wire L133_0a;
  wire [31:0] L134_0r0;
  wire [31:0] L134_0r1;
  wire L134_0a;
  wire L135_0r;
  wire L135_0a;
  wire L136_0r;
  wire L136_0a;
  wire L138_0r0;
  wire L138_0r1;
  wire L138_0a;
  wire L139_0r;
  wire L139_0a;
  wire L140_0r;
  wire L140_0a;
  wire L141_0r;
  wire L141_0a;
  wire L142_0r;
  wire L142_0a;
  wire L143_0r0;
  wire L143_0r1;
  wire L143_0a;
  wire L145_0r;
  wire L145_0a;
  wire L146_0r;
  wire L146_0a;
  wire L147_0r;
  wire L147_0a;
  wire L148_0r;
  wire L148_0a;
  wire L149_0r0;
  wire L149_0r1;
  wire L149_0a;
  wire L150_0r;
  wire L150_0a;
  wire L151_0r0;
  wire L151_0r1;
  wire L151_0a;
  wire L152_0r;
  wire L152_0a;
  wire L153_0r0;
  wire L153_0r1;
  wire L153_0a;
  wire L154_0r;
  wire L154_0a;
  wire L155_0r0;
  wire L155_0r1;
  wire L155_0a;
  wire L156_0r;
  wire L156_0a;
  wire L157_0r0;
  wire L157_0r1;
  wire L157_0a;
  wire L158_0r;
  wire L158_0a;
  wire L159_0r0;
  wire L159_0r1;
  wire L159_0a;
  wire L160_0r;
  wire L160_0a;
  wire L161_0r0;
  wire L161_0r1;
  wire L161_0a;
  wire L162_0r;
  wire L162_0a;
  wire L163_0r0;
  wire L163_0r1;
  wire L163_0a;
  wire L164_0r0;
  wire L164_0r1;
  wire L164_0a;
  wire L165_0r;
  wire L165_0a;
  wire L166_0r0;
  wire L166_0r1;
  wire L166_0a;
  wire [7:0] L167_0r0;
  wire [7:0] L167_0r1;
  wire L167_0a;
  wire [7:0] L168_0r0;
  wire [7:0] L168_0r1;
  wire L168_0a;
  wire [7:0] L169_0r0;
  wire [7:0] L169_0r1;
  wire L169_0a;
  wire [7:0] L170_0r0;
  wire [7:0] L170_0r1;
  wire L170_0a;
  wire [7:0] L171_0r0;
  wire [7:0] L171_0r1;
  wire L171_0a;
  wire [7:0] L172_0r0;
  wire [7:0] L172_0r1;
  wire L172_0a;
  wire [7:0] L173_0r0;
  wire [7:0] L173_0r1;
  wire L173_0a;
  wire [7:0] L174_0r0;
  wire [7:0] L174_0r1;
  wire L174_0a;
  wire [7:0] L175_0r0;
  wire [7:0] L175_0r1;
  wire L175_0a;
  wire [7:0] L176_0r0;
  wire [7:0] L176_0r1;
  wire L176_0a;
  wire L178_0r;
  wire L178_0a;
  wire L179_0r;
  wire L179_0a;
  wire L180_0r;
  wire L180_0a;
  wire L181_0r;
  wire L181_0a;
  wire L182_0r;
  wire L182_0a;
  wire [5:0] L183_0r0;
  wire [5:0] L183_0r1;
  wire L183_0a;
  wire L184_0r;
  wire L184_0a;
  wire L185_0r0;
  wire L185_0r1;
  wire L185_0a;
  wire L187_0r;
  wire L187_0a;
  wire [6:0] L188_0r0;
  wire [6:0] L188_0r1;
  wire L188_0a;
  wire L189_0r;
  wire L189_0a;
  wire L191_0r;
  wire L191_0a;
  wire [3:0] L192_0r0;
  wire [3:0] L192_0r1;
  wire L192_0a;
  wire L193_0r;
  wire L193_0a;
  wire L194_0r;
  wire L194_0a;
  wire L195_0r;
  wire L195_0a;
  wire L196_0r0;
  wire L196_0r1;
  wire L196_0a;
  wire L197_0r;
  wire L197_0a;
  wire L198_0r;
  wire L198_0a;
  wire [31:0] L200_0r0;
  wire [31:0] L200_0r1;
  wire L200_0a;
  wire L201_0r;
  wire L201_0a;
  wire L202_0r;
  wire L202_0a;
  wire L203_0r;
  wire L203_0a;
  wire L204_0r;
  wire L204_0a;
  wire [31:0] L205_0r0;
  wire [31:0] L205_0r1;
  wire L205_0a;
  wire L207_0r;
  wire L207_0a;
  wire L208_0r;
  wire L208_0a;
  wire L209_0r;
  wire L209_0a;
  wire L210_0r;
  wire L210_0a;
  wire L211_0r;
  wire L211_0a;
  wire L213_0r;
  wire L213_0a;
  wire L214_0r;
  wire L214_0a;
  wire L215_0r;
  wire L215_0a;
  wire L216_0r;
  wire L216_0a;
  wire L217_0r;
  wire L217_0a;
  wire [5:0] L218_0r0;
  wire [5:0] L218_0r1;
  wire L218_0a;
  wire L219_0r;
  wire L219_0a;
  wire L220_0r0;
  wire L220_0r1;
  wire L220_0a;
  wire L222_0r;
  wire L222_0a;
  wire [6:0] L223_0r0;
  wire [6:0] L223_0r1;
  wire L223_0a;
  wire L224_0r;
  wire L224_0a;
  wire L226_0r;
  wire L226_0a;
  wire [31:0] L228_0r0;
  wire [31:0] L228_0r1;
  wire L228_0a;
  wire L229_0r;
  wire L229_0a;
  wire [31:0] L230_0r0;
  wire [31:0] L230_0r1;
  wire L230_0a;
  wire L232_0r;
  wire L232_0a;
  wire L233_0r;
  wire L233_0a;
  wire L234_0r0;
  wire L234_0r1;
  wire L234_0a;
  wire L235_0r;
  wire L235_0a;
  wire [1:0] L236_0r0;
  wire [1:0] L236_0r1;
  wire L236_0a;
  wire L238_0r;
  wire L238_0a;
  wire [2:0] L239_0r0;
  wire [2:0] L239_0r1;
  wire L239_0a;
  wire L240_0r;
  wire L240_0a;
  wire L241_0r;
  wire L241_0a;
  wire [3:0] L242_0r0;
  wire [3:0] L242_0r1;
  wire L242_0a;
  wire L244_0r;
  wire L244_0a;
  wire L245_0r;
  wire L245_0a;
  wire [31:0] L247_0r0;
  wire [31:0] L247_0r1;
  wire L247_0a;
  wire L248_0r;
  wire L248_0a;
  wire [31:0] L249_0r0;
  wire [31:0] L249_0r1;
  wire L249_0a;
  wire L251_0r;
  wire L251_0a;
  wire L252_0r;
  wire L252_0a;
  wire L253_0r;
  wire L253_0a;
  wire L254_0r;
  wire L254_0a;
  wire L255_0r;
  wire L255_0a;
  wire L257_0r;
  wire L257_0a;
  wire L258_0r;
  wire L258_0a;
  wire L260_0r;
  wire L260_0a;
  wire L261_0r;
  wire L261_0a;
  wire L262_0r;
  wire L262_0a;
  wire L263_0r;
  wire L263_0a;
  wire L264_0r;
  wire L264_0a;
  wire [5:0] L265_0r0;
  wire [5:0] L265_0r1;
  wire L265_0a;
  wire L266_0r;
  wire L266_0a;
  wire L267_0r0;
  wire L267_0r1;
  wire L267_0a;
  wire L269_0r;
  wire L269_0a;
  wire [6:0] L270_0r0;
  wire [6:0] L270_0r1;
  wire L270_0a;
  wire L271_0r;
  wire L271_0a;
  wire L273_0r;
  wire L273_0a;
  wire [31:0] L275_0r0;
  wire [31:0] L275_0r1;
  wire L275_0a;
  wire L276_0r;
  wire L276_0a;
  wire [31:0] L277_0r0;
  wire [31:0] L277_0r1;
  wire L277_0a;
  wire L279_0r;
  wire L279_0a;
  wire L280_0r;
  wire L280_0a;
  wire L281_0r0;
  wire L281_0r1;
  wire L281_0a;
  wire L282_0r;
  wire L282_0a;
  wire [1:0] L283_0r0;
  wire [1:0] L283_0r1;
  wire L283_0a;
  wire L285_0r;
  wire L285_0a;
  wire [2:0] L286_0r0;
  wire [2:0] L286_0r1;
  wire L286_0a;
  wire L287_0r;
  wire L287_0a;
  wire L288_0r;
  wire L288_0a;
  wire [3:0] L289_0r0;
  wire [3:0] L289_0r1;
  wire L289_0a;
  wire L291_0r;
  wire L291_0a;
  wire L293_0r;
  wire L293_0a;
  wire [31:0] L295_0r0;
  wire [31:0] L295_0r1;
  wire L295_0a;
  wire L296_0r;
  wire L296_0a;
  wire [31:0] L297_0r0;
  wire [31:0] L297_0r1;
  wire L297_0a;
  wire L299_0r;
  wire L299_0a;
  wire L300_0r;
  wire L300_0a;
  wire L301_0r;
  wire L301_0a;
  wire L302_0r;
  wire L302_0a;
  wire L303_0r;
  wire L303_0a;
  wire L305_0r;
  wire L305_0a;
  wire L306_0r;
  wire L306_0a;
  wire L307_0r;
  wire L307_0a;
  wire L308_0r;
  wire L308_0a;
  wire L310_0r;
  wire L310_0a;
  wire [73:0] L311_0r0;
  wire [73:0] L311_0r1;
  wire L311_0a;
  wire L312_0r;
  wire L312_0a;
  wire L314_0r;
  wire L314_0a;
  wire [32:0] L315_0r0;
  wire [32:0] L315_0r1;
  wire L315_0a;
  wire L316_0r;
  wire L316_0a;
  wire L317_0r;
  wire L317_0a;
  wire L319_0r;
  wire L319_0a;
  wire L321_0r0;
  wire L321_0r1;
  wire L321_0a;
  wire L322_0r;
  wire L322_0a;
  wire L323_0r;
  wire L323_0a;
  wire L324_0r;
  wire L324_0a;
  wire L325_0r;
  wire L325_0a;
  wire L326_0r;
  wire L326_0a;
  wire L327_0r;
  wire L327_0a;
  wire L328_0r;
  wire L328_0a;
  wire L329_0r;
  wire L329_0a;
  wire L330_0r;
  wire L330_0a;
  wire L331_0r;
  wire L331_0a;
  wire L332_0r;
  wire L332_0a;
  wire L333_0r;
  wire L333_0a;
  wire L334_0r;
  wire L334_0a;
  wire L335_0r;
  wire L335_0a;
  wire L336_0r;
  wire L336_0a;
  wire [6:0] L337_0r0;
  wire [6:0] L337_0r1;
  wire L337_0a;
  wire [6:0] L338_0r0;
  wire [6:0] L338_0r1;
  wire L338_0a;
  wire [6:0] L339_0r0;
  wire [6:0] L339_0r1;
  wire L339_0a;
  wire [6:0] L340_0r0;
  wire [6:0] L340_0r1;
  wire L340_0a;
  wire [6:0] L341_0r0;
  wire [6:0] L341_0r1;
  wire L341_0a;
  wire [6:0] L342_0r0;
  wire [6:0] L342_0r1;
  wire L342_0a;
  wire [6:0] L343_0r0;
  wire [6:0] L343_0r1;
  wire L343_0a;
  wire [6:0] L344_0r0;
  wire [6:0] L344_0r1;
  wire L344_0a;
  wire [6:0] L345_0r0;
  wire [6:0] L345_0r1;
  wire L345_0a;
  wire L347_0r;
  wire L347_0a;
  wire L348_0r0;
  wire L348_0r1;
  wire L348_0a;
  wire L349_0r;
  wire L349_0a;
  wire [31:0] L351_0r0;
  wire [31:0] L351_0r1;
  wire L351_0a;
  wire L352_0r;
  wire L352_0a;
  wire L353_0r;
  wire L353_0a;
  wire [31:0] L355_0r0;
  wire [31:0] L355_0r1;
  wire L355_0a;
  wire L356_0r;
  wire L356_0a;
  wire [31:0] L357_0r0;
  wire [31:0] L357_0r1;
  wire L357_0a;
  wire L359_0r;
  wire L359_0a;
  wire L360_0r;
  wire L360_0a;
  wire L361_0r;
  wire L361_0a;
  wire [31:0] L363_0r0;
  wire [31:0] L363_0r1;
  wire L363_0a;
  wire L364_0r;
  wire L364_0a;
  wire [31:0] L365_0r0;
  wire [31:0] L365_0r1;
  wire L365_0a;
  wire L367_0r;
  wire L367_0a;
  wire L368_0r;
  wire L368_0a;
  wire L369_0r;
  wire L369_0a;
  wire L370_0r;
  wire L370_0a;
  wire L371_0r;
  wire L371_0a;
  wire L372_0r;
  wire L372_0a;
  wire L373_0r;
  wire L373_0a;
  wire L374_0r;
  wire L374_0a;
  wire L375_0r;
  wire L375_0a;
  wire [2:0] L376_0r0;
  wire [2:0] L376_0r1;
  wire L376_0a;
  wire [2:0] L377_0r0;
  wire [2:0] L377_0r1;
  wire L377_0a;
  wire [2:0] L378_0r0;
  wire [2:0] L378_0r1;
  wire L378_0a;
  wire [2:0] L379_0r0;
  wire [2:0] L379_0r1;
  wire L379_0a;
  wire [2:0] L380_0r0;
  wire [2:0] L380_0r1;
  wire L380_0a;
  wire L382_0r;
  wire L382_0a;
  wire [2:0] L384_0r0;
  wire [2:0] L384_0r1;
  wire L384_0a;
  wire L385_0r;
  wire L385_0a;
  wire L386_0r;
  wire L386_0a;
  wire L387_0r0;
  wire L387_0r1;
  wire L387_0a;
  wire L388_0r;
  wire L388_0a;
  wire L389_0r;
  wire L389_0a;
  wire [4:0] L391_0r0;
  wire [4:0] L391_0r1;
  wire L391_0a;
  wire L392_0r;
  wire L392_0a;
  wire L393_0r;
  wire L393_0a;
  wire L394_0r;
  wire L394_0a;
  wire L395_0r0;
  wire L395_0r1;
  wire L395_0a;
  wire L396_0r;
  wire L396_0a;
  wire L397_0r;
  wire L397_0a;
  wire [4:0] L399_0r0;
  wire [4:0] L399_0r1;
  wire L399_0a;
  wire L400_0r;
  wire L400_0a;
  wire L401_0r;
  wire L401_0a;
  wire L402_0r;
  wire L402_0a;
  wire L403_0r0;
  wire L403_0r1;
  wire L403_0a;
  wire L404_0r;
  wire L404_0a;
  wire L405_0r;
  wire L405_0a;
  wire [4:0] L407_0r0;
  wire [4:0] L407_0r1;
  wire L407_0a;
  wire L408_0r;
  wire L408_0a;
  wire L409_0r;
  wire L409_0a;
  wire L410_0r;
  wire L410_0a;
  wire L412_0r0;
  wire L412_0r1;
  wire L412_0a;
  wire L413_0r;
  wire L413_0a;
  wire L414_0r;
  wire L414_0a;
  wire L415_0r0;
  wire L415_0r1;
  wire L415_0a;
  wire L416_0r;
  wire L416_0a;
  wire L417_0r;
  wire L417_0a;
  wire [4:0] L419_0r0;
  wire [4:0] L419_0r1;
  wire L419_0a;
  wire L420_0r;
  wire L420_0a;
  wire L421_0r;
  wire L421_0a;
  wire L422_0r;
  wire L422_0a;
  wire L424_0r0;
  wire L424_0r1;
  wire L424_0a;
  wire L425_0r;
  wire L425_0a;
  wire L426_0r;
  wire L426_0a;
  wire L427_0r;
  wire L427_0a;
  wire L428_0r;
  wire L428_0a;
  wire L429_0r;
  wire L429_0a;
  wire L430_0r;
  wire L430_0a;
  wire L431_0r;
  wire L431_0a;
  wire L432_0r;
  wire L432_0a;
  wire L433_0r;
  wire L433_0a;
  wire [2:0] L434_0r0;
  wire [2:0] L434_0r1;
  wire L434_0a;
  wire [2:0] L435_0r0;
  wire [2:0] L435_0r1;
  wire L435_0a;
  wire [2:0] L436_0r0;
  wire [2:0] L436_0r1;
  wire L436_0a;
  wire [2:0] L437_0r0;
  wire [2:0] L437_0r1;
  wire L437_0a;
  wire [2:0] L438_0r0;
  wire [2:0] L438_0r1;
  wire L438_0a;
  wire L439_0r0;
  wire L439_0r1;
  wire L439_0a;
  wire L440_0r;
  wire L440_0a;
  wire L441_0r;
  wire L441_0a;
  wire L442_0r0;
  wire L442_0r1;
  wire L442_0a;
  wire L443_0r;
  wire L443_0a;
  wire L444_0r0;
  wire L444_0r1;
  wire L444_0a;
  wire [1:0] L445_0r0;
  wire [1:0] L445_0r1;
  wire L445_0a;
  wire [1:0] L446_0r0;
  wire [1:0] L446_0r1;
  wire L446_0a;
  wire [1:0] L447_0r0;
  wire [1:0] L447_0r1;
  wire L447_0a;
  wire [1:0] L448_0r0;
  wire [1:0] L448_0r1;
  wire L448_0a;
  wire L449_0r0;
  wire L449_0r1;
  wire L449_0a;
  wire L450_0r;
  wire L450_0a;
  wire L451_0r;
  wire L451_0a;
  wire L452_0r0;
  wire L452_0r1;
  wire L452_0a;
  wire L453_0r;
  wire L453_0a;
  wire L454_0r0;
  wire L454_0r1;
  wire L454_0a;
  wire L455_0r;
  wire L455_0a;
  wire L456_0r0;
  wire L456_0r1;
  wire L456_0a;
  wire [2:0] L457_0r0;
  wire [2:0] L457_0r1;
  wire L457_0a;
  wire [2:0] L458_0r0;
  wire [2:0] L458_0r1;
  wire L458_0a;
  wire [2:0] L459_0r0;
  wire [2:0] L459_0r1;
  wire L459_0a;
  wire [2:0] L460_0r0;
  wire [2:0] L460_0r1;
  wire L460_0a;
  wire [2:0] L461_0r0;
  wire [2:0] L461_0r1;
  wire L461_0a;
  wire [3:0] L462_0r0;
  wire [3:0] L462_0r1;
  wire L462_0a;
  wire L463_0r;
  wire L463_0a;
  wire L464_0r;
  wire L464_0a;
  wire [3:0] L465_0r0;
  wire [3:0] L465_0r1;
  wire L465_0a;
  wire L466_0r;
  wire L466_0a;
  wire [3:0] L467_0r0;
  wire [3:0] L467_0r1;
  wire L467_0a;
  wire [1:0] L468_0r0;
  wire [1:0] L468_0r1;
  wire L468_0a;
  wire [1:0] L469_0r0;
  wire [1:0] L469_0r1;
  wire L469_0a;
  wire [1:0] L470_0r0;
  wire [1:0] L470_0r1;
  wire L470_0a;
  wire [1:0] L471_0r0;
  wire [1:0] L471_0r1;
  wire L471_0a;
  wire L474_0r;
  wire L474_0a;
  wire L475_0r0;
  wire L475_0r1;
  wire L475_0a;
  wire L476_0r;
  wire L476_0a;
  wire L477_0r0;
  wire L477_0r1;
  wire L477_0a;
  wire L478_0r0;
  wire L478_0r1;
  wire L478_0a;
  wire L479_0r;
  wire L479_0a;
  wire [1:0] L481_0r0;
  wire [1:0] L481_0r1;
  wire L481_0a;
  wire [1:0] L482_0r0;
  wire [1:0] L482_0r1;
  wire L482_0a;
  wire [1:0] L483_0r0;
  wire [1:0] L483_0r1;
  wire L483_0a;
  wire [1:0] L484_0r0;
  wire [1:0] L484_0r1;
  wire L484_0a;
  wire L493_0r;
  wire L493_0a;
  wire [31:0] L494_0r0;
  wire [31:0] L494_0r1;
  wire L494_0a;
  wire L495_0r;
  wire L495_0a;
  wire [31:0] L496_0r0;
  wire [31:0] L496_0r1;
  wire L496_0a;
  wire [31:0] L497_0r0;
  wire [31:0] L497_0r1;
  wire L497_0a;
  wire L498_0r;
  wire L498_0a;
  wire [1:0] L500_0r0;
  wire [1:0] L500_0r1;
  wire L500_0a;
  wire [1:0] L501_0r0;
  wire [1:0] L501_0r1;
  wire L501_0a;
  wire [1:0] L502_0r0;
  wire [1:0] L502_0r1;
  wire L502_0a;
  wire [1:0] L503_0r0;
  wire [1:0] L503_0r1;
  wire L503_0a;
  wire L507_0r;
  wire L507_0a;
  wire [6:0] L508_0r0;
  wire [6:0] L508_0r1;
  wire L508_0a;
  wire L509_0r;
  wire L509_0a;
  wire [6:0] L510_0r0;
  wire [6:0] L510_0r1;
  wire L510_0a;
  wire L511_0r;
  wire L511_0a;
  wire [6:0] L512_0r0;
  wire [6:0] L512_0r1;
  wire L512_0a;
  wire [6:0] L513_0r0;
  wire [6:0] L513_0r1;
  wire L513_0a;
  wire L514_0r;
  wire L514_0a;
  wire [2:0] L516_0r0;
  wire [2:0] L516_0r1;
  wire L516_0a;
  wire [2:0] L517_0r0;
  wire [2:0] L517_0r1;
  wire L517_0a;
  wire [2:0] L518_0r0;
  wire [2:0] L518_0r1;
  wire L518_0a;
  wire [2:0] L519_0r0;
  wire [2:0] L519_0r1;
  wire L519_0a;
  wire [2:0] L520_0r0;
  wire [2:0] L520_0r1;
  wire L520_0a;
  wire [2:0] L522_0r0;
  wire [2:0] L522_0r1;
  wire L522_0a;
  wire [2:0] L523_0r0;
  wire [2:0] L523_0r1;
  wire L523_0a;
  wire [2:0] L524_0r0;
  wire [2:0] L524_0r1;
  wire L524_0a;
  wire [2:0] L525_0r0;
  wire [2:0] L525_0r1;
  wire L525_0a;
  wire [34:0] L526_0r0;
  wire [34:0] L526_0r1;
  wire L526_0a;
  wire [2:0] L528_0r0;
  wire [2:0] L528_0r1;
  wire L528_0a;
  wire [2:0] L529_0r0;
  wire [2:0] L529_0r1;
  wire L529_0a;
  wire [2:0] L530_0r0;
  wire [2:0] L530_0r1;
  wire L530_0a;
  wire [2:0] L531_0r0;
  wire [2:0] L531_0r1;
  wire L531_0a;
  wire [6:0] L532_0r0;
  wire [6:0] L532_0r1;
  wire L532_0a;
  wire L534_0r;
  wire L534_0a;
  wire [31:0] L535_0r0;
  wire [31:0] L535_0r1;
  wire L535_0a;
  wire L536_0r;
  wire L536_0a;
  wire [31:0] L537_0r0;
  wire [31:0] L537_0r1;
  wire L537_0a;
  wire [31:0] L538_0r0;
  wire [31:0] L538_0r1;
  wire L538_0a;
  wire L539_0r;
  wire L539_0a;
  wire [1:0] L541_0r0;
  wire [1:0] L541_0r1;
  wire L541_0a;
  wire [1:0] L542_0r0;
  wire [1:0] L542_0r1;
  wire L542_0a;
  wire [1:0] L543_0r0;
  wire [1:0] L543_0r1;
  wire L543_0a;
  wire [1:0] L544_0r0;
  wire [1:0] L544_0r1;
  wire L544_0a;
  wire L545_0r;
  wire L545_0a;
  wire [31:0] L546_0r0;
  wire [31:0] L546_0r1;
  wire L546_0a;
  wire L547_0r;
  wire L547_0a;
  wire [31:0] L548_0r0;
  wire [31:0] L548_0r1;
  wire L548_0a;
  wire [31:0] L549_0r0;
  wire [31:0] L549_0r1;
  wire L549_0a;
  wire L550_0r;
  wire L550_0a;
  wire [1:0] L552_0r0;
  wire [1:0] L552_0r1;
  wire L552_0a;
  wire [1:0] L553_0r0;
  wire [1:0] L553_0r1;
  wire L553_0a;
  wire [1:0] L554_0r0;
  wire [1:0] L554_0r1;
  wire L554_0a;
  wire [1:0] L555_0r0;
  wire [1:0] L555_0r1;
  wire L555_0a;
  wire L556_0r;
  wire L556_0a;
  wire [2:0] L557_0r0;
  wire [2:0] L557_0r1;
  wire L557_0a;
  wire L558_0r;
  wire L558_0a;
  wire [2:0] L559_0r0;
  wire [2:0] L559_0r1;
  wire L559_0a;
  wire [2:0] L560_0r0;
  wire [2:0] L560_0r1;
  wire L560_0a;
  wire L561_0r;
  wire L561_0a;
  wire [1:0] L563_0r0;
  wire [1:0] L563_0r1;
  wire L563_0a;
  wire [1:0] L564_0r0;
  wire [1:0] L564_0r1;
  wire L564_0a;
  wire [1:0] L565_0r0;
  wire [1:0] L565_0r1;
  wire L565_0a;
  wire [1:0] L566_0r0;
  wire [1:0] L566_0r1;
  wire L566_0a;
  tko0m1_1nm1b0 I0 (L2_0r, L2_0a, L4_0r0, L4_0r1, L4_0a, reset);
  tko0m4_1nm4b0 I1 (L6_0r, L6_0a, L8_0r0[3:0], L8_0r1[3:0], L8_0a, reset);
  tko0m1_1nm1b0 I2 (L10_0r, L10_0a, L12_0r0, L12_0r1, L12_0a, reset);
  tko0m1_1nm1b0 I3 (L14_0r, L14_0a, L16_0r0, L16_0r1, L16_0a, reset);
  tkj0m0_0_0_0 I4 (L5_0r, L5_0a, L9_0r, L9_0a, L13_0r, L13_0a, L17_0r, L17_0a, L308_0r, L308_0a, reset);
  tko1m1_1noti0w1b I5 (L30_0r0, L30_0r1, L30_0a, L28_0r0, L28_0r1, L28_0a, reset);
  tkj2m1_1 I6 (L27_0r0, L27_0r1, L27_0a, L28_0r0, L28_0r1, L28_0a, L31_0r0[1:0], L31_0r1[1:0], L31_0a, reset);
  tko2m1_1api0w1b_2api1w1b_3andt1o0w1bt2o0w1b I7 (L31_0r0[1:0], L31_0r1[1:0], L31_0a, L32_0r0, L32_0r1, L32_0a, reset);
  tkf0mo0w0_o0w0 I8 (L33_0r, L33_0a, L26_0r, L26_0a, L29_0r, L29_0a, reset);
  tkm2x0b I9 (L23_0r, L23_0a, L25_0r, L25_0a, L317_0r, L317_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I10 (L32_0r0, L32_0r1, L32_0a, L42_0r, L42_0a, L25_0r, L25_0a, reset);
  tkf0mo0w0_o0w0 I11 (L42_0r, L42_0a, L34_0r, L34_0a, L38_0r, L38_0a, reset);
  tkj0m0_0 I12 (L37_0r, L37_0a, L41_0r, L41_0a, L44_0r, L44_0a, reset);
  tko0m1_1nm1b0 I13 (L44_0r, L44_0a, L46_0r0, L46_0r1, L46_0a, reset);
  tkf0mo0w0_o0w0 I14 (L54_0r, L54_0a, L51_0r, L51_0a, L52_0r, L52_0a, reset);
  tkj0m0_0 I15 (L51_0r, L51_0a, L53_0r, L53_0a, L55_0r, L55_0a, reset);
  tko0m1_1nm1b0 I16 (L59_0r, L59_0a, L61_0r0, L61_0r1, L61_0a, reset);
  tkj2m1_1 I17 (L70_0r0, L70_0r1, L70_0a, L72_0r0, L72_0r1, L72_0a, L73_0r0[1:0], L73_0r1[1:0], L73_0a, reset);
  tko2m1_1api0w1b_2api1w1b_3net1o0w1bt2o0w1b I18 (L73_0r0[1:0], L73_0r1[1:0], L73_0a, L74_0r0, L74_0r1, L74_0a, reset);
  tkj2m1_1 I19 (L68_0r0, L68_0r1, L68_0a, L74_0r0, L74_0r1, L74_0a, L75_0r0[1:0], L75_0r1[1:0], L75_0a, reset);
  tko2m1_1api0w1b_2api1w1b_3ort1o0w1bt2o0w1b I20 (L75_0r0[1:0], L75_0r1[1:0], L75_0a, L78_0r0, L78_0r1, L78_0a, reset);
  tkf0mo0w0_o0w0_o0w0 I21 (L77_0r, L77_0a, L67_0r, L67_0a, L69_0r, L69_0a, L71_0r, L71_0a, reset);
  tkj2m1_1 I22 (L81_0r0, L81_0r1, L81_0a, L83_0r0, L83_0r1, L83_0a, L84_0r0[1:0], L84_0r1[1:0], L84_0a, reset);
  tko2m1_1api0w1b_2api1w1b_3net1o0w1bt2o0w1b I23 (L84_0r0[1:0], L84_0r1[1:0], L84_0a, L87_0r0, L87_0r1, L87_0a, reset);
  tkf0mo0w0_o0w0 I24 (L86_0r, L86_0a, L80_0r, L80_0a, L82_0r, L82_0a, reset);
  tkj2m1_1 I25 (L90_0r0, L90_0r1, L90_0a, L92_0r0, L92_0r1, L92_0a, L93_0r0[1:0], L93_0r1[1:0], L93_0a, reset);
  tko2m1_1api0w1b_2api1w1b_3ort1o0w1bt2o0w1b I26 (L93_0r0[1:0], L93_0r1[1:0], L93_0a, L96_0r0, L96_0r1, L96_0a, reset);
  tkf0mo0w0_o0w0 I27 (L95_0r, L95_0a, L89_0r, L89_0a, L91_0r, L91_0a, reset);
  tks4_o0w4_0m8o0w0_1m9o0w0_2mao0w0_3mbo0w0_4mco0w0_5mdo0w0_6meo0w0_7mfo0w0 I28 (L58_0r0[3:0], L58_0r1[3:0], L58_0a, L59_0r, L59_0a, L63_0r, L63_0a, L77_0r, L77_0a, L86_0r, L86_0a, L95_0r, L95_0a, L98_0r, L98_0a, L102_0r, L102_0a, L106_0r, L106_0a, reset);
  tkm8x0b I29 (L62_0r, L62_0a, L66_0r, L66_0a, L79_0r, L79_0a, L88_0r, L88_0a, L97_0r, L97_0a, L101_0r, L101_0a, L105_0r, L105_0a, L109_0r, L109_0a, L110_0r, L110_0a, reset);
  tkj2m1_1 I30 (L113_0r0, L113_0r1, L113_0a, L115_0r0, L115_0r1, L115_0a, L116_0r0[1:0], L116_0r1[1:0], L116_0a, reset);
  tko2m1_1api0w1b_2api1w1b_3net1o0w1bt2o0w1b I31 (L116_0r0[1:0], L116_0r1[1:0], L116_0a, L119_0r0, L119_0r1, L119_0a, reset);
  tkf0mo0w0_o0w0 I32 (L118_0r, L118_0a, L112_0r, L112_0a, L114_0r, L114_0a, reset);
  tkj64m32_32 I33 (L128_0r0[31:0], L128_0r1[31:0], L128_0a, L130_0r0[31:0], L130_0r1[31:0], L130_0a, L131_0r0[63:0], L131_0r1[63:0], L131_0a, reset);
  tko64m33_1api0w32b_2api32w32b_3nm1b0_4apt1o0w32bt3o0w1b_5nm1b0_6apt2o0w32bt5o0w1b_7addt4o0w33bt6o0w33b I34 (L131_0r0[63:0], L131_0r1[63:0], L131_0a, L132_0r0[32:0], L132_0r1[32:0], L132_0a, reset);
  tkf33mo0w32 I35 (L132_0r0[32:0], L132_0r1[32:0], L132_0a, L134_0r0[31:0], L134_0r1[31:0], L134_0a, reset);
  tkf0mo0w0_o0w0 I36 (L133_0r, L133_0a, L127_0r, L127_0a, L129_0r, L129_0a, reset);
  tko0m1_1nm1b1 I37 (L136_0r, L136_0a, L138_0r0, L138_0r1, L138_0a, reset);
  tkf0mo0w0_o0w0 I38 (L140_0r, L140_0a, L133_0r, L133_0a, L136_0r, L136_0a, reset);
  tkj0m0_0 I39 (L135_0r, L135_0a, L139_0r, L139_0a, L141_0r, L141_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I40 (L122_0r0, L122_0r1, L122_0a, L123_0r, L123_0a, L140_0r, L140_0a, reset);
  tkm2x0b I41 (L124_0r, L124_0a, L141_0r, L141_0a, L142_0r, L142_0a, reset);
  tkvtake1_wo0w1_ro0w1 I42 (L143_0r0, L143_0r1, L143_0a, L118_0r, L118_0a, L112_0r, L112_0a, L113_0r0, L113_0r1, L113_0a, reset);
  tkf0mo0w0_o0w0 I43 (L146_0r, L146_0a, L57_0r, L57_0a, L145_0r, L145_0a, reset);
  tkj0m0_0 I44 (L110_0r, L110_0a, L142_0r, L142_0a, L147_0r, L147_0a, reset);
  tkf1mo0w0_o0w1 I45 (L61_0r0, L61_0r1, L61_0a, L148_0r, L148_0a, L149_0r0, L149_0r1, L149_0a, reset);
  tkf1mo0w0_o0w1 I46 (L65_0r0, L65_0r1, L65_0a, L150_0r, L150_0a, L151_0r0, L151_0r1, L151_0a, reset);
  tkf1mo0w0_o0w1 I47 (L78_0r0, L78_0r1, L78_0a, L152_0r, L152_0a, L153_0r0, L153_0r1, L153_0a, reset);
  tkf1mo0w0_o0w1 I48 (L87_0r0, L87_0r1, L87_0a, L154_0r, L154_0a, L155_0r0, L155_0r1, L155_0a, reset);
  tkf1mo0w0_o0w1 I49 (L96_0r0, L96_0r1, L96_0a, L156_0r, L156_0a, L157_0r0, L157_0r1, L157_0a, reset);
  tkf1mo0w0_o0w1 I50 (L100_0r0, L100_0r1, L100_0a, L158_0r, L158_0a, L159_0r0, L159_0r1, L159_0a, reset);
  tkf1mo0w0_o0w1 I51 (L104_0r0, L104_0r1, L104_0a, L160_0r, L160_0a, L161_0r0, L161_0r1, L161_0a, reset);
  tkf1mo0w0_o0w1 I52 (L108_0r0, L108_0r1, L108_0a, L162_0r, L162_0a, L163_0r0, L163_0r1, L163_0a, reset);
  tkm8x1b I53 (L149_0r0, L149_0r1, L149_0a, L151_0r0, L151_0r1, L151_0a, L153_0r0, L153_0r1, L153_0a, L155_0r0, L155_0r1, L155_0a, L157_0r0, L157_0r1, L157_0a, L159_0r0, L159_0r1, L159_0a, L161_0r0, L161_0r1, L161_0a, L163_0r0, L163_0r1, L163_0a, L164_0r0, L164_0r1, L164_0a, reset);
  tkf1mo0w0_o0w1 I54 (L164_0r0, L164_0r1, L164_0a, L165_0r, L165_0a, L166_0r0, L166_0r1, L166_0a, reset);
  tko0m8_1nm8b1 I55 (L148_0r, L148_0a, L167_0r0[7:0], L167_0r1[7:0], L167_0a, reset);
  tko0m8_1nm8b2 I56 (L150_0r, L150_0a, L168_0r0[7:0], L168_0r1[7:0], L168_0a, reset);
  tko0m8_1nm8b4 I57 (L152_0r, L152_0a, L169_0r0[7:0], L169_0r1[7:0], L169_0a, reset);
  tko0m8_1nm8b8 I58 (L154_0r, L154_0a, L170_0r0[7:0], L170_0r1[7:0], L170_0a, reset);
  tko0m8_1nm8b10 I59 (L156_0r, L156_0a, L171_0r0[7:0], L171_0r1[7:0], L171_0a, reset);
  tko0m8_1nm8b20 I60 (L158_0r, L158_0a, L172_0r0[7:0], L172_0r1[7:0], L172_0a, reset);
  tko0m8_1nm8b40 I61 (L160_0r, L160_0a, L173_0r0[7:0], L173_0r1[7:0], L173_0a, reset);
  tko0m8_1nm8b80 I62 (L162_0r, L162_0a, L174_0r0[7:0], L174_0r1[7:0], L174_0a, reset);
  tkm8x8b I63 (L167_0r0[7:0], L167_0r1[7:0], L167_0a, L168_0r0[7:0], L168_0r1[7:0], L168_0a, L169_0r0[7:0], L169_0r1[7:0], L169_0a, L170_0r0[7:0], L170_0r1[7:0], L170_0a, L171_0r0[7:0], L171_0r1[7:0], L171_0a, L172_0r0[7:0], L172_0r1[7:0], L172_0a, L173_0r0[7:0], L173_0r1[7:0], L173_0a, L174_0r0[7:0], L174_0r1[7:0], L174_0a, L175_0r0[7:0], L175_0r1[7:0], L175_0a, reset);
  tkj8m0_8 I64 (L165_0r, L165_0a, L175_0r0[7:0], L175_0r1[7:0], L175_0a, L176_0r0[7:0], L176_0r1[7:0], L176_0a, reset);
  tks8_o0w8_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0_20o0w0_40o0w0_80o0w0 I65 (L176_0r0[7:0], L176_0r1[7:0], L176_0a, L62_0r, L62_0a, L66_0r, L66_0a, L79_0r, L79_0a, L88_0r, L88_0a, L97_0r, L97_0a, L101_0r, L101_0a, L105_0r, L105_0a, L109_0r, L109_0a, reset);
  tkj1m1_0 I66 (L166_0r0, L166_0r1, L166_0a, L145_0r, L145_0a, L143_0r0, L143_0r1, L143_0a, reset);
  tkj7m6_1 I67 (L183_0r0[5:0], L183_0r1[5:0], L183_0a, L185_0r0, L185_0r1, L185_0a, L188_0r0[6:0], L188_0r1[6:0], L188_0a, reset);
  tkf0mo0w0_o0w0 I68 (L187_0r, L187_0a, L182_0r, L182_0a, L184_0r, L184_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I69 (L196_0r0, L196_0r1, L196_0a, L197_0r, L197_0a, L198_0r, L198_0a, reset);
  tkm2x0b I70 (L197_0r, L197_0a, L201_0r, L201_0a, L202_0r, L202_0a, reset);
  tkf0mo0w0_o0w0 I71 (L203_0r, L203_0a, L194_0r, L194_0a, L195_0r, L195_0a, reset);
  tkj0m0_0 I72 (L194_0r, L194_0a, L202_0r, L202_0a, L204_0r, L204_0a, reset);
  tkvaluResult32_wo0w32_ro0w32 I73 (L205_0r0[31:0], L205_0r1[31:0], L205_0a, L203_0r, L203_0a, L198_0r, L198_0a, L200_0r0[31:0], L200_0r1[31:0], L200_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0 I74 (L210_0r, L210_0a, L178_0r, L178_0a, L180_0r, L180_0a, L187_0r, L187_0a, L191_0r, L191_0a, L207_0r, L207_0a, L208_0r, L208_0a, reset);
  tkj0m0_0_0_0_0_0 I75 (L179_0r, L179_0a, L181_0r, L181_0a, L189_0r, L189_0a, L193_0r, L193_0a, L204_0r, L204_0a, L209_0r, L209_0a, L211_0r, L211_0a, reset);
  tko0m6_1nm6b0 I76 (L217_0r, L217_0a, L218_0r0[5:0], L218_0r1[5:0], L218_0a, reset);
  tkj7m6_1 I77 (L218_0r0[5:0], L218_0r1[5:0], L218_0a, L220_0r0, L220_0r1, L220_0a, L223_0r0[6:0], L223_0r1[6:0], L223_0a, reset);
  tkf0mo0w0_o0w0 I78 (L222_0r, L222_0a, L217_0r, L217_0a, L219_0r, L219_0a, reset);
  tkvaluResult32_wo0w32_ro0w32 I79 (L230_0r0[31:0], L230_0r1[31:0], L230_0a, L226_0r, L226_0a, L226_0r, L226_0a, L228_0r0[31:0], L228_0r1[31:0], L228_0a, reset);
  tko0m1_1nm1b1 I80 (L233_0r, L233_0a, L234_0r0, L234_0r1, L234_0a, reset);
  tkj3m1_2 I81 (L234_0r0, L234_0r1, L234_0a, L236_0r0[1:0], L236_0r1[1:0], L236_0a, L239_0r0[2:0], L239_0r1[2:0], L239_0a, reset);
  tkf0mo0w0_o0w0 I82 (L238_0r, L238_0a, L233_0r, L233_0a, L235_0r, L235_0a, reset);
  tkf4mo0w0 I83 (L242_0r0[3:0], L242_0r1[3:0], L242_0a, L241_0r, L241_0a, reset);
  tkvdread32_wo0w32_ro0w32 I84 (L249_0r0[31:0], L249_0r1[31:0], L249_0a, L245_0r, L245_0a, L245_0r, L245_0a, L247_0r0[31:0], L247_0r1[31:0], L247_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 I85 (L254_0r, L254_0a, L213_0r, L213_0a, L215_0r, L215_0a, L222_0r, L222_0a, L232_0r, L232_0a, L238_0r, L238_0a, L244_0r, L244_0a, L251_0r, L251_0a, L252_0r, L252_0a, reset);
  tkj0m0_0_0_0_0_0_0_0 I86 (L214_0r, L214_0a, L216_0r, L216_0a, L224_0r, L224_0a, L229_0r, L229_0a, L240_0r, L240_0a, L241_0r, L241_0a, L248_0r, L248_0a, L253_0r, L253_0a, L255_0r, L255_0a, reset);
  tko0m6_1nm6b0 I87 (L264_0r, L264_0a, L265_0r0[5:0], L265_0r1[5:0], L265_0a, reset);
  tkj7m6_1 I88 (L265_0r0[5:0], L265_0r1[5:0], L265_0a, L267_0r0, L267_0r1, L267_0a, L270_0r0[6:0], L270_0r1[6:0], L270_0a, reset);
  tkf0mo0w0_o0w0 I89 (L269_0r, L269_0a, L264_0r, L264_0a, L266_0r, L266_0a, reset);
  tkvaluResult32_wo0w32_ro0w32 I90 (L277_0r0[31:0], L277_0r1[31:0], L277_0a, L273_0r, L273_0a, L273_0r, L273_0a, L275_0r0[31:0], L275_0r1[31:0], L275_0a, reset);
  tko0m1_1nm1b0 I91 (L280_0r, L280_0a, L281_0r0, L281_0r1, L281_0a, reset);
  tkj3m1_2 I92 (L281_0r0, L281_0r1, L281_0a, L283_0r0[1:0], L283_0r1[1:0], L283_0a, L286_0r0[2:0], L286_0r1[2:0], L286_0a, reset);
  tkf0mo0w0_o0w0 I93 (L285_0r, L285_0a, L280_0r, L280_0a, L282_0r, L282_0a, reset);
  tkf4mo0w0 I94 (L289_0r0[3:0], L289_0r1[3:0], L289_0a, L288_0r, L288_0a, reset);
  tkvr232_wo0w32_ro0w32 I95 (L297_0r0[31:0], L297_0r1[31:0], L297_0a, L293_0r, L293_0a, L293_0r, L293_0a, L295_0r0[31:0], L295_0r1[31:0], L295_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 I96 (L302_0r, L302_0a, L260_0r, L260_0a, L262_0r, L262_0a, L269_0r, L269_0a, L279_0r, L279_0a, L285_0r, L285_0a, L291_0r, L291_0a, L299_0r, L299_0a, L300_0r, L300_0a, reset);
  tkj0m0_0_0_0_0_0_0_0 I97 (L261_0r, L261_0a, L263_0r, L263_0a, L271_0r, L271_0a, L276_0r, L276_0a, L287_0r, L287_0a, L288_0r, L288_0a, L296_0r, L296_0a, L301_0r, L301_0a, L303_0r, L303_0a, reset);
  tks3_o0w3_7o0w0_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0 I98 (L49_0r0[2:0], L49_0r1[2:0], L49_0a, L50_0r, L50_0a, L54_0r, L54_0a, L146_0r, L146_0a, L210_0r, L210_0a, L254_0r, L254_0a, L257_0r, L257_0a, L302_0r, L302_0a, L305_0r, L305_0a, reset);
  tkm8x0b I99 (L50_0r, L50_0a, L55_0r, L55_0a, L147_0r, L147_0a, L211_0r, L211_0a, L255_0r, L255_0a, L258_0r, L258_0a, L303_0r, L303_0a, L306_0r, L306_0a, L307_0r, L307_0a, reset);
  tkm2x0b I100 (L308_0r, L308_0a, L307_0r, L307_0a, L23_0r, L23_0a, reset);
  tkf0mo0w0_o0w0 I101 (L317_0r, L317_0a, L310_0r, L310_0a, L314_0r, L314_0a, reset);
  tkj0m0_0 I102 (L312_0r, L312_0a, L316_0r, L316_0a, L33_0r, L33_0a, reset);
  tko0m1_1nm1b0 I103 (L319_0r, L319_0a, L321_0r0, L321_0r1, L321_0a, reset);
  tkf0mo0w0_o0w0 I104 (L52_0r, L52_0a, L323_0r, L323_0a, L324_0r, L324_0a, reset);
  tkf0mo0w0_o0w0 I105 (L123_0r, L123_0a, L325_0r, L325_0a, L326_0r, L326_0a, reset);
  tkf0mo0w0_o0w0 I106 (L208_0r, L208_0a, L327_0r, L327_0a, L328_0r, L328_0a, reset);
  tkf0mo0w0_o0w0 I107 (L252_0r, L252_0a, L329_0r, L329_0a, L330_0r, L330_0a, reset);
  tkf0mo0w0_o0w0 I108 (L257_0r, L257_0a, L331_0r, L331_0a, L332_0r, L332_0a, reset);
  tkf0mo0w0_o0w0 I109 (L300_0r, L300_0a, L333_0r, L333_0a, L334_0r, L334_0a, reset);
  tkf0mo0w0_o0w0 I110 (L305_0r, L305_0a, L335_0r, L335_0a, L336_0r, L336_0a, reset);
  tkm7x0b I111 (L323_0r, L323_0a, L325_0r, L325_0a, L327_0r, L327_0a, L329_0r, L329_0a, L331_0r, L331_0a, L333_0r, L333_0a, L335_0r, L335_0a, L319_0r, L319_0a, reset);
  tko0m7_1nm7b1 I112 (L324_0r, L324_0a, L337_0r0[6:0], L337_0r1[6:0], L337_0a, reset);
  tko0m7_1nm7b2 I113 (L326_0r, L326_0a, L338_0r0[6:0], L338_0r1[6:0], L338_0a, reset);
  tko0m7_1nm7b4 I114 (L328_0r, L328_0a, L339_0r0[6:0], L339_0r1[6:0], L339_0a, reset);
  tko0m7_1nm7b8 I115 (L330_0r, L330_0a, L340_0r0[6:0], L340_0r1[6:0], L340_0a, reset);
  tko0m7_1nm7b10 I116 (L332_0r, L332_0a, L341_0r0[6:0], L341_0r1[6:0], L341_0a, reset);
  tko0m7_1nm7b20 I117 (L334_0r, L334_0a, L342_0r0[6:0], L342_0r1[6:0], L342_0a, reset);
  tko0m7_1nm7b40 I118 (L336_0r, L336_0a, L343_0r0[6:0], L343_0r1[6:0], L343_0a, reset);
  tkm7x7b I119 (L337_0r0[6:0], L337_0r1[6:0], L337_0a, L338_0r0[6:0], L338_0r1[6:0], L338_0a, L339_0r0[6:0], L339_0r1[6:0], L339_0a, L340_0r0[6:0], L340_0r1[6:0], L340_0a, L341_0r0[6:0], L341_0r1[6:0], L341_0a, L342_0r0[6:0], L342_0r1[6:0], L342_0a, L343_0r0[6:0], L343_0r1[6:0], L343_0a, L344_0r0[6:0], L344_0r1[6:0], L344_0a, reset);
  tkj7m0_7 I120 (L322_0r, L322_0a, L344_0r0[6:0], L344_0r1[6:0], L344_0a, L345_0r0[6:0], L345_0r1[6:0], L345_0a, reset);
  tks7_o0w7_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0_20o0w0_40o0w0 I121 (L345_0r0[6:0], L345_0r1[6:0], L345_0a, L53_0r, L53_0a, L124_0r, L124_0a, L209_0r, L209_0a, L253_0r, L253_0a, L258_0r, L258_0a, L301_0r, L301_0a, L306_0r, L306_0a, reset);
  tkvr132_wo0w32_ro0w32 I122 (L357_0r0[31:0], L357_0r1[31:0], L357_0a, L353_0r, L353_0a, L353_0r, L353_0a, L355_0r0[31:0], L355_0r1[31:0], L355_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I123 (L348_0r0, L348_0r1, L348_0a, L349_0r, L349_0a, L359_0r, L359_0a, reset);
  tkm2x0b I124 (L352_0r, L352_0a, L356_0r, L356_0a, L360_0r, L360_0a, reset);
  tkvr032_wo0w32_ro0w32 I125 (L365_0r0[31:0], L365_0r1[31:0], L365_0a, L361_0r, L361_0a, L361_0r, L361_0a, L363_0r0[31:0], L363_0r1[31:0], L363_0a, reset);
  tkf0mo0w0_o0w0 I126 (L368_0r, L368_0a, L347_0r, L347_0a, L367_0r, L367_0a, reset);
  tkj0m0_0 I127 (L360_0r, L360_0a, L364_0r, L364_0a, L369_0r, L369_0a, reset);
  tkf0mo0w0_o0w0 I128 (L180_0r, L180_0a, L370_0r, L370_0a, L371_0r, L371_0a, reset);
  tkf0mo0w0_o0w0 I129 (L215_0r, L215_0a, L372_0r, L372_0a, L373_0r, L373_0a, reset);
  tkf0mo0w0_o0w0 I130 (L262_0r, L262_0a, L374_0r, L374_0a, L375_0r, L375_0a, reset);
  tkm3x0b I131 (L370_0r, L370_0a, L372_0r, L372_0a, L374_0r, L374_0a, L368_0r, L368_0a, reset);
  tko0m3_1nm3b1 I132 (L371_0r, L371_0a, L376_0r0[2:0], L376_0r1[2:0], L376_0a, reset);
  tko0m3_1nm3b2 I133 (L373_0r, L373_0a, L377_0r0[2:0], L377_0r1[2:0], L377_0a, reset);
  tko0m3_1nm3b4 I134 (L375_0r, L375_0a, L378_0r0[2:0], L378_0r1[2:0], L378_0a, reset);
  tkm3x3b I135 (L376_0r0[2:0], L376_0r1[2:0], L376_0a, L377_0r0[2:0], L377_0r1[2:0], L377_0a, L378_0r0[2:0], L378_0r1[2:0], L378_0a, L379_0r0[2:0], L379_0r1[2:0], L379_0a, reset);
  tkj3m0_3 I136 (L369_0r, L369_0a, L379_0r0[2:0], L379_0r1[2:0], L379_0a, L380_0r0[2:0], L380_0r1[2:0], L380_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_4o0w0 I137 (L380_0r0[2:0], L380_0r1[2:0], L380_0a, L181_0r, L181_0a, L216_0r, L216_0a, L263_0r, L263_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I138 (L387_0r0, L387_0r1, L387_0a, L388_0r, L388_0a, L389_0r, L389_0a, reset);
  tkm2x0b I139 (L388_0r, L388_0a, L392_0r, L392_0a, L393_0r, L393_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I140 (L395_0r0, L395_0r1, L395_0a, L396_0r, L396_0a, L397_0r, L397_0a, reset);
  tkm2x0b I141 (L396_0r, L396_0a, L400_0r, L400_0a, L401_0r, L401_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I142 (L403_0r0, L403_0r1, L403_0a, L404_0r, L404_0a, L405_0r, L405_0a, reset);
  tkm2x0b I143 (L404_0r, L404_0a, L408_0r, L408_0a, L409_0r, L409_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I144 (L415_0r0, L415_0r1, L415_0a, L416_0r, L416_0a, L417_0r, L417_0a, reset);
  tkm2x0b I145 (L416_0r, L416_0a, L420_0r, L420_0a, L421_0r, L421_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0 I146 (L426_0r, L426_0a, L382_0r, L382_0a, L386_0r, L386_0a, L394_0r, L394_0a, L402_0r, L402_0a, L410_0r, L410_0a, L414_0r, L414_0a, L422_0r, L422_0a, reset);
  tkj0m0_0_0_0_0_0_0 I147 (L385_0r, L385_0a, L393_0r, L393_0a, L401_0r, L401_0a, L409_0r, L409_0a, L413_0r, L413_0a, L421_0r, L421_0a, L425_0r, L425_0a, L427_0r, L427_0a, reset);
  tkf0mo0w0_o0w0 I148 (L178_0r, L178_0a, L428_0r, L428_0a, L429_0r, L429_0a, reset);
  tkf0mo0w0_o0w0 I149 (L213_0r, L213_0a, L430_0r, L430_0a, L431_0r, L431_0a, reset);
  tkf0mo0w0_o0w0 I150 (L260_0r, L260_0a, L432_0r, L432_0a, L433_0r, L433_0a, reset);
  tkm3x0b I151 (L428_0r, L428_0a, L430_0r, L430_0a, L432_0r, L432_0a, L426_0r, L426_0a, reset);
  tko0m3_1nm3b1 I152 (L429_0r, L429_0a, L434_0r0[2:0], L434_0r1[2:0], L434_0a, reset);
  tko0m3_1nm3b2 I153 (L431_0r, L431_0a, L435_0r0[2:0], L435_0r1[2:0], L435_0a, reset);
  tko0m3_1nm3b4 I154 (L433_0r, L433_0a, L436_0r0[2:0], L436_0r1[2:0], L436_0a, reset);
  tkm3x3b I155 (L434_0r0[2:0], L434_0r1[2:0], L434_0a, L435_0r0[2:0], L435_0r1[2:0], L435_0a, L436_0r0[2:0], L436_0r1[2:0], L436_0a, L437_0r0[2:0], L437_0r1[2:0], L437_0a, reset);
  tkj3m0_3 I156 (L427_0r, L427_0a, L437_0r0[2:0], L437_0r1[2:0], L437_0a, L438_0r0[2:0], L438_0r1[2:0], L438_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_4o0w0 I157 (L438_0r0[2:0], L438_0r1[2:0], L438_0a, L179_0r, L179_0a, L214_0r, L214_0a, L261_0r, L261_0a, reset);
  tkf1mo0w0_o0w1 I158 (L36_0r0, L36_0r1, L36_0a, L441_0r, L441_0a, L442_0r0, L442_0r1, L442_0a, reset);
  tkf1mo0w0_o0w1 I159 (L16_0r0, L16_0r1, L16_0a, L443_0r, L443_0a, L444_0r0, L444_0r1, L444_0a, reset);
  tkm2x1b I160 (L442_0r0, L442_0r1, L442_0a, L444_0r0, L444_0r1, L444_0a, L439_0r0, L439_0r1, L439_0a, reset);
  tko0m2_1nm2b1 I161 (L441_0r, L441_0a, L445_0r0[1:0], L445_0r1[1:0], L445_0a, reset);
  tko0m2_1nm2b2 I162 (L443_0r, L443_0a, L446_0r0[1:0], L446_0r1[1:0], L446_0a, reset);
  tkm2x2b I163 (L445_0r0[1:0], L445_0r1[1:0], L445_0a, L446_0r0[1:0], L446_0r1[1:0], L446_0a, L447_0r0[1:0], L447_0r1[1:0], L447_0a, reset);
  tkj2m0_2 I164 (L440_0r, L440_0a, L447_0r0[1:0], L447_0r1[1:0], L447_0a, L448_0r0[1:0], L448_0r1[1:0], L448_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I165 (L448_0r0[1:0], L448_0r1[1:0], L448_0a, L37_0r, L37_0a, L17_0r, L17_0a, reset);
  tkvtakeBranch21_wo0w1_ro0w1 I166 (L439_0r0, L439_0r1, L439_0a, L440_0r, L440_0a, L26_0r, L26_0a, L27_0r0, L27_0r1, L27_0a, reset);
  tkf1mo0w0_o0w1 I167 (L119_0r0, L119_0r1, L119_0a, L451_0r, L451_0a, L452_0r0, L452_0r1, L452_0a, reset);
  tkf1mo0w0_o0w1 I168 (L46_0r0, L46_0r1, L46_0a, L453_0r, L453_0a, L454_0r0, L454_0r1, L454_0a, reset);
  tkf1mo0w0_o0w1 I169 (L12_0r0, L12_0r1, L12_0a, L455_0r, L455_0a, L456_0r0, L456_0r1, L456_0a, reset);
  tkm3x1b I170 (L452_0r0, L452_0r1, L452_0a, L454_0r0, L454_0r1, L454_0a, L456_0r0, L456_0r1, L456_0a, L449_0r0, L449_0r1, L449_0a, reset);
  tko0m3_1nm3b1 I171 (L451_0r, L451_0a, L457_0r0[2:0], L457_0r1[2:0], L457_0a, reset);
  tko0m3_1nm3b2 I172 (L453_0r, L453_0a, L458_0r0[2:0], L458_0r1[2:0], L458_0a, reset);
  tko0m3_1nm3b4 I173 (L455_0r, L455_0a, L459_0r0[2:0], L459_0r1[2:0], L459_0a, reset);
  tkm3x3b I174 (L457_0r0[2:0], L457_0r1[2:0], L457_0a, L458_0r0[2:0], L458_0r1[2:0], L458_0a, L459_0r0[2:0], L459_0r1[2:0], L459_0a, L460_0r0[2:0], L460_0r1[2:0], L460_0a, reset);
  tkj3m0_3 I175 (L450_0r, L450_0a, L460_0r0[2:0], L460_0r1[2:0], L460_0a, L461_0r0[2:0], L461_0r1[2:0], L461_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_4o0w0 I176 (L461_0r0[2:0], L461_0r1[2:0], L461_0a, L121_0r, L121_0a, L48_0r, L48_0a, L13_0r, L13_0a, reset);
  tkvtakeBranch1_wo0w1_ro0w1o0w1 I177 (L449_0r0, L449_0r1, L449_0a, L450_0r, L450_0a, L121_0r, L121_0a, L34_0r, L34_0a, L122_0r0, L122_0r1, L122_0a, L36_0r0, L36_0r1, L36_0a, reset);
  tkvcwp1_wo0w1_ro0w1 I178 (L4_0r0, L4_0r1, L4_0a, L5_0r, L5_0a, L422_0r, L422_0a, L424_0r0, L424_0r1, L424_0a, reset);
  tkvpreCarry1_wo0w1_ro0w1o0w1o0w1 I179 (L40_0r0, L40_0r1, L40_0a, L41_0r, L41_0a, L266_0r, L266_0a, L219_0r, L219_0a, L184_0r, L184_0a, L267_0r0, L267_0r1, L267_0a, L220_0r0, L220_0r1, L220_0a, L185_0r0, L185_0r1, L185_0a, reset);
  tkf4mo0w0_o0w4 I180 (L192_0r0[3:0], L192_0r1[3:0], L192_0a, L464_0r, L464_0a, L465_0r0[3:0], L465_0r1[3:0], L465_0a, reset);
  tkf4mo0w0_o0w4 I181 (L8_0r0[3:0], L8_0r1[3:0], L8_0a, L466_0r, L466_0a, L467_0r0[3:0], L467_0r1[3:0], L467_0a, reset);
  tkm2x4b I182 (L465_0r0[3:0], L465_0r1[3:0], L465_0a, L467_0r0[3:0], L467_0r1[3:0], L467_0a, L462_0r0[3:0], L462_0r1[3:0], L462_0a, reset);
  tko0m2_1nm2b1 I183 (L464_0r, L464_0a, L468_0r0[1:0], L468_0r1[1:0], L468_0a, reset);
  tko0m2_1nm2b2 I184 (L466_0r, L466_0a, L469_0r0[1:0], L469_0r1[1:0], L469_0a, reset);
  tkm2x2b I185 (L468_0r0[1:0], L468_0r1[1:0], L468_0a, L469_0r0[1:0], L469_0r1[1:0], L469_0a, L470_0r0[1:0], L470_0r1[1:0], L470_0a, reset);
  tkj2m0_2 I186 (L463_0r, L463_0a, L470_0r0[1:0], L470_0r1[1:0], L470_0a, L471_0r0[1:0], L471_0r1[1:0], L471_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I187 (L471_0r0[1:0], L471_0r1[1:0], L471_0a, L193_0r, L193_0a, L9_0r, L9_0a, reset);
  tkvflags4_wo0w4_ro2w1o1w1o3w1o0w1o3w1o2w1o1w1o2w1o1w1o0w1o0w1o3w1 I188 (L462_0r0[3:0], L462_0r1[3:0], L462_0a, L463_0r, L463_0a, L106_0r, L106_0a, L102_0r, L102_0a, L98_0r, L98_0a, L91_0r, L91_0a, L89_0r, L89_0a, L82_0r, L82_0a, L80_0r, L80_0a, L71_0r, L71_0a, L69_0r, L69_0a, L67_0r, L67_0a, L63_0r, L63_0a, L38_0r, L38_0a, L108_0r0, L108_0r1, L108_0a, L104_0r0, L104_0r1, L104_0a, L100_0r0, L100_0r1, L100_0a, L92_0r0, L92_0r1, L92_0a, L90_0r0, L90_0r1, L90_0a, L83_0r0, L83_0r1, L83_0a, L81_0r0, L81_0r1, L81_0a, L72_0r0, L72_0r1, L72_0a, L70_0r0, L70_0r1, L70_0a, L68_0r0, L68_0r1, L68_0a, L65_0r0, L65_0r1, L65_0a, L40_0r0, L40_0r1, L40_0a, reset);
  tkvpcr33_wo0w33_ro0w32o32w1 I189 (L315_0r0[32:0], L315_0r1[32:0], L315_0a, L316_0r, L316_0a, L127_0r, L127_0a, L29_0r, L29_0a, L128_0r0[31:0], L128_0r1[31:0], L128_0a, L30_0r0, L30_0r1, L30_0a, reset);
  tkvopr74_wo0w74_ro26w5o25w1o25w1o20w5o9w1o15w5o8w1o10w5o7w1o7w3o38w32o37w1o71w2o71w2o25w1o31w6o38w32o6w1o3w4o0w3 I190 (L311_0r0[73:0], L311_0r1[73:0], L311_0a, L312_0r, L312_0a, L417_0r, L417_0a, L414_0r, L414_0a, L410_0r, L410_0a, L405_0r, L405_0a, L402_0r, L402_0a, L397_0r, L397_0a, L394_0r, L394_0a, L389_0r, L389_0a, L386_0r, L386_0a, L382_0r, L382_0a, L349_0r, L349_0a, L347_0r, L347_0a, L282_0r, L282_0a, L235_0r, L235_0a, L195_0r, L195_0a, L182_0r, L182_0a, L129_0r, L129_0a, L114_0r, L114_0a, L57_0r, L57_0a, L48_0r, L48_0a, L419_0r0[4:0], L419_0r1[4:0], L419_0a, L415_0r0, L415_0r1, L415_0a, L412_0r0, L412_0r1, L412_0a, L407_0r0[4:0], L407_0r1[4:0], L407_0a, L403_0r0, L403_0r1, L403_0a, L399_0r0[4:0], L399_0r1[4:0], L399_0a, L395_0r0, L395_0r1, L395_0a, L391_0r0[4:0], L391_0r1[4:0], L391_0a, L387_0r0, L387_0r1, L387_0a, L384_0r0[2:0], L384_0r1[2:0], L384_0a, L351_0r0[31:0], L351_0r1[31:0], L351_0a, L348_0r0, L348_0r1, L348_0a, L283_0r0[1:0], L283_0r1[1:0], L283_0a, L236_0r0[1:0], L236_0r1[1:0], L236_0a, L196_0r0, L196_0r1, L196_0a, L183_0r0[5:0], L183_0r1[5:0], L183_0a, L130_0r0[31:0], L130_0r1[31:0], L130_0a, L115_0r0, L115_0r1, L115_0a, L58_0r0[3:0], L58_0r1[3:0], L58_0a, L49_0r0[2:0], L49_0r1[2:0], L49_0a, reset);
  tkj74m74_0 I191 (op_0r0[73:0], op_0r1[73:0], op_0a, L310_0r, L310_0a, L311_0r0[73:0], L311_0r1[73:0], L311_0a, reset);
  tkj33m33_0 I192 (pc_0r0[32:0], pc_0r1[32:0], pc_0a, L314_0r, L314_0a, L315_0r0[32:0], L315_0r1[32:0], L315_0a, reset);
  tkf1mo0w0_o0w1 I193 (L138_0r0, L138_0r1, L138_0a, L474_0r, L474_0a, L475_0r0, L475_0r1, L475_0a, reset);
  tkf1mo0w0_o0w1 I194 (L321_0r0, L321_0r1, L321_0a, L476_0r, L476_0a, L477_0r0, L477_0r1, L477_0a, reset);
  tkm2x1b I195 (L475_0r0, L475_0r1, L475_0a, L477_0r0, L477_0r1, L477_0a, L478_0r0, L478_0r1, L478_0a, reset);
  tkf1mo0w0_o0w1 I196 (L478_0r0, L478_0r1, L478_0a, L479_0r, L479_0a, doFetch_0r0, doFetch_0r1, doFetch_0a, reset);
  tko0m2_1nm2b1 I197 (L474_0r, L474_0a, L481_0r0[1:0], L481_0r1[1:0], L481_0a, reset);
  tko0m2_1nm2b2 I198 (L476_0r, L476_0a, L482_0r0[1:0], L482_0r1[1:0], L482_0a, reset);
  tkm2x2b I199 (L481_0r0[1:0], L481_0r1[1:0], L481_0a, L482_0r0[1:0], L482_0r1[1:0], L482_0a, L483_0r0[1:0], L483_0r1[1:0], L483_0a, reset);
  tkj2m0_2 I200 (L479_0r, L479_0a, L483_0r0[1:0], L483_0r1[1:0], L483_0a, L484_0r0[1:0], L484_0r1[1:0], L484_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I201 (L484_0r0[1:0], L484_0r1[1:0], L484_0a, L139_0r, L139_0a, L322_0r, L322_0a, reset);
  tkf32mo0w0_o0w32 I202 (L134_0r0[31:0], L134_0r1[31:0], L134_0a, L135_0r, L135_0a, newPc_0r0[31:0], newPc_0r1[31:0], newPc_0a, reset);
  tkf1mo0w0_o0w1 I203 (L412_0r0, L412_0r1, L412_0a, L413_0r, L413_0a, wEn_0r0, wEn_0r1, wEn_0a, reset);
  tkf3mo0w0_o0w3 I204 (L384_0r0[2:0], L384_0r1[2:0], L384_0a, L385_0r, L385_0a, rEn_0r0[2:0], rEn_0r1[2:0], rEn_0a, reset);
  tkf5mo0w0_o0w5 I205 (L419_0r0[4:0], L419_0r1[4:0], L419_0a, L420_0r, L420_0a, wSel_0r0[4:0], wSel_0r1[4:0], wSel_0a, reset);
  tkf5mo0w0_o0w5 I206 (L391_0r0[4:0], L391_0r1[4:0], L391_0a, L392_0r, L392_0a, r0Sel_0r0[4:0], r0Sel_0r1[4:0], r0Sel_0a, reset);
  tkf5mo0w0_o0w5 I207 (L399_0r0[4:0], L399_0r1[4:0], L399_0a, L400_0r, L400_0a, r1Sel_0r0[4:0], r1Sel_0r1[4:0], r1Sel_0a, reset);
  tkf5mo0w0_o0w5 I208 (L407_0r0[4:0], L407_0r1[4:0], L407_0a, L408_0r, L408_0a, r2Sel_0r0[4:0], r2Sel_0r1[4:0], r2Sel_0a, reset);
  tkf1mo0w0_o0w1 I209 (L424_0r0, L424_0r1, L424_0a, L425_0r, L425_0a, window_0r0, window_0r1, window_0a, reset);
  tkf32mo0w0_o0w32 I210 (L200_0r0[31:0], L200_0r1[31:0], L200_0a, L493_0r, L493_0a, L494_0r0[31:0], L494_0r1[31:0], L494_0a, reset);
  tkf32mo0w0_o0w32 I211 (L247_0r0[31:0], L247_0r1[31:0], L247_0a, L495_0r, L495_0a, L496_0r0[31:0], L496_0r1[31:0], L496_0a, reset);
  tkm2x32b I212 (L494_0r0[31:0], L494_0r1[31:0], L494_0a, L496_0r0[31:0], L496_0r1[31:0], L496_0a, L497_0r0[31:0], L497_0r1[31:0], L497_0a, reset);
  tkf32mo0w0_o0w32 I213 (L497_0r0[31:0], L497_0r1[31:0], L497_0a, L498_0r, L498_0a, w_0r0[31:0], w_0r1[31:0], w_0a, reset);
  tko0m2_1nm2b1 I214 (L493_0r, L493_0a, L500_0r0[1:0], L500_0r1[1:0], L500_0a, reset);
  tko0m2_1nm2b2 I215 (L495_0r, L495_0a, L501_0r0[1:0], L501_0r1[1:0], L501_0a, reset);
  tkm2x2b I216 (L500_0r0[1:0], L500_0r1[1:0], L500_0a, L501_0r0[1:0], L501_0r1[1:0], L501_0a, L502_0r0[1:0], L502_0r1[1:0], L502_0a, reset);
  tkj2m0_2 I217 (L498_0r, L498_0a, L502_0r0[1:0], L502_0r1[1:0], L502_0a, L503_0r0[1:0], L503_0r1[1:0], L503_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I218 (L503_0r0[1:0], L503_0r1[1:0], L503_0a, L201_0r, L201_0a, L248_0r, L248_0a, reset);
  tkj32m32_0 I219 (r0_0r0[31:0], r0_0r1[31:0], r0_0a, L367_0r, L367_0a, L365_0r0[31:0], L365_0r1[31:0], L365_0a, reset);
  tkj32m32_0 I220 (r1_0r0[31:0], r1_0r1[31:0], r1_0a, L359_0r, L359_0a, L357_0r0[31:0], L357_0r1[31:0], L357_0a, reset);
  tkj32m32_0 I221 (r2_0r0[31:0], r2_0r1[31:0], r2_0a, L299_0r, L299_0a, L297_0r0[31:0], L297_0r1[31:0], L297_0a, reset);
  tkf7mo0w0_o0w7 I222 (L188_0r0[6:0], L188_0r1[6:0], L188_0a, L507_0r, L507_0a, L508_0r0[6:0], L508_0r1[6:0], L508_0a, reset);
  tkf7mo0w0_o0w7 I223 (L223_0r0[6:0], L223_0r1[6:0], L223_0a, L509_0r, L509_0a, L510_0r0[6:0], L510_0r1[6:0], L510_0a, reset);
  tkf7mo0w0_o0w7 I224 (L270_0r0[6:0], L270_0r1[6:0], L270_0a, L511_0r, L511_0a, L512_0r0[6:0], L512_0r1[6:0], L512_0a, reset);
  tkm3x7b I225 (L508_0r0[6:0], L508_0r1[6:0], L508_0a, L510_0r0[6:0], L510_0r1[6:0], L510_0a, L512_0r0[6:0], L512_0r1[6:0], L512_0a, L513_0r0[6:0], L513_0r1[6:0], L513_0a, reset);
  tkf7mo0w0_o0w7 I226 (L513_0r0[6:0], L513_0r1[6:0], L513_0a, L514_0r, L514_0a, aluOp_0r0[6:0], aluOp_0r1[6:0], aluOp_0a, reset);
  tko0m3_1nm3b1 I227 (L507_0r, L507_0a, L516_0r0[2:0], L516_0r1[2:0], L516_0a, reset);
  tko0m3_1nm3b2 I228 (L509_0r, L509_0a, L517_0r0[2:0], L517_0r1[2:0], L517_0a, reset);
  tko0m3_1nm3b4 I229 (L511_0r, L511_0a, L518_0r0[2:0], L518_0r1[2:0], L518_0a, reset);
  tkm3x3b I230 (L516_0r0[2:0], L516_0r1[2:0], L516_0a, L517_0r0[2:0], L517_0r1[2:0], L517_0a, L518_0r0[2:0], L518_0r1[2:0], L518_0a, L519_0r0[2:0], L519_0r1[2:0], L519_0a, reset);
  tkj3m0_3 I231 (L514_0r, L514_0a, L519_0r0[2:0], L519_0r1[2:0], L519_0a, L520_0r0[2:0], L520_0r1[2:0], L520_0a, reset);
  tks3_o0w3_1o0w0_2o0w0_4o0w0 I232 (L520_0r0[2:0], L520_0r1[2:0], L520_0a, L189_0r, L189_0a, L224_0r, L224_0a, L271_0r, L271_0a, reset);
  tko0m3_1nm3b1 I233 (L207_0r, L207_0a, L522_0r0[2:0], L522_0r1[2:0], L522_0a, reset);
  tko0m3_1nm3b2 I234 (L232_0r, L232_0a, L523_0r0[2:0], L523_0r1[2:0], L523_0a, reset);
  tko0m3_1nm3b4 I235 (L279_0r, L279_0a, L524_0r0[2:0], L524_0r1[2:0], L524_0a, reset);
  tkm3x3b I236 (L522_0r0[2:0], L522_0r1[2:0], L522_0a, L523_0r0[2:0], L523_0r1[2:0], L523_0a, L524_0r0[2:0], L524_0r1[2:0], L524_0a, L525_0r0[2:0], L525_0r1[2:0], L525_0a, reset);
  tkj35m32_3 I237 (aluResult_0r0[31:0], aluResult_0r1[31:0], aluResult_0a, L525_0r0[2:0], L525_0r1[2:0], L525_0a, L526_0r0[34:0], L526_0r1[34:0], L526_0a, reset);
  tks35_o32w3_1o0w32_2o0w32_4o0w32 I238 (L526_0r0[34:0], L526_0r1[34:0], L526_0a, L205_0r0[31:0], L205_0r1[31:0], L205_0a, L230_0r0[31:0], L230_0r1[31:0], L230_0a, L277_0r0[31:0], L277_0r1[31:0], L277_0a, reset);
  tko0m3_1nm3b1 I239 (L191_0r, L191_0a, L528_0r0[2:0], L528_0r1[2:0], L528_0a, reset);
  tko0m3_1nm3b2 I240 (L244_0r, L244_0a, L529_0r0[2:0], L529_0r1[2:0], L529_0a, reset);
  tko0m3_1nm3b4 I241 (L291_0r, L291_0a, L530_0r0[2:0], L530_0r1[2:0], L530_0a, reset);
  tkm3x3b I242 (L528_0r0[2:0], L528_0r1[2:0], L528_0a, L529_0r0[2:0], L529_0r1[2:0], L529_0a, L530_0r0[2:0], L530_0r1[2:0], L530_0a, L531_0r0[2:0], L531_0r1[2:0], L531_0a, reset);
  tkj7m4_3 I243 (aluFlags_0r0[3:0], aluFlags_0r1[3:0], aluFlags_0a, L531_0r0[2:0], L531_0r1[2:0], L531_0a, L532_0r0[6:0], L532_0r1[6:0], L532_0a, reset);
  tks7_o4w3_1o0w4_2o0w4_4o0w4 I244 (L532_0r0[6:0], L532_0r1[6:0], L532_0a, L192_0r0[3:0], L192_0r1[3:0], L192_0a, L242_0r0[3:0], L242_0r1[3:0], L242_0a, L289_0r0[3:0], L289_0r1[3:0], L289_0a, reset);
  tkf32mo0w0_o0w32 I245 (L363_0r0[31:0], L363_0r1[31:0], L363_0a, L364_0r, L364_0a, aluLhs_0r0[31:0], aluLhs_0r1[31:0], aluLhs_0a, reset);
  tkf32mo0w0_o0w32 I246 (L351_0r0[31:0], L351_0r1[31:0], L351_0a, L534_0r, L534_0a, L535_0r0[31:0], L535_0r1[31:0], L535_0a, reset);
  tkf32mo0w0_o0w32 I247 (L355_0r0[31:0], L355_0r1[31:0], L355_0a, L536_0r, L536_0a, L537_0r0[31:0], L537_0r1[31:0], L537_0a, reset);
  tkm2x32b I248 (L535_0r0[31:0], L535_0r1[31:0], L535_0a, L537_0r0[31:0], L537_0r1[31:0], L537_0a, L538_0r0[31:0], L538_0r1[31:0], L538_0a, reset);
  tkf32mo0w0_o0w32 I249 (L538_0r0[31:0], L538_0r1[31:0], L538_0a, L539_0r, L539_0a, aluRhs_0r0[31:0], aluRhs_0r1[31:0], aluRhs_0a, reset);
  tko0m2_1nm2b1 I250 (L534_0r, L534_0a, L541_0r0[1:0], L541_0r1[1:0], L541_0a, reset);
  tko0m2_1nm2b2 I251 (L536_0r, L536_0a, L542_0r0[1:0], L542_0r1[1:0], L542_0a, reset);
  tkm2x2b I252 (L541_0r0[1:0], L541_0r1[1:0], L541_0a, L542_0r0[1:0], L542_0r1[1:0], L542_0a, L543_0r0[1:0], L543_0r1[1:0], L543_0a, reset);
  tkj2m0_2 I253 (L539_0r, L539_0a, L543_0r0[1:0], L543_0r1[1:0], L543_0a, L544_0r0[1:0], L544_0r1[1:0], L544_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I254 (L544_0r0[1:0], L544_0r1[1:0], L544_0a, L352_0r, L352_0a, L356_0r, L356_0a, reset);
  tkf32mo0w0_o0w32 I255 (L228_0r0[31:0], L228_0r1[31:0], L228_0a, L545_0r, L545_0a, L546_0r0[31:0], L546_0r1[31:0], L546_0a, reset);
  tkf32mo0w0_o0w32 I256 (L275_0r0[31:0], L275_0r1[31:0], L275_0a, L547_0r, L547_0a, L548_0r0[31:0], L548_0r1[31:0], L548_0a, reset);
  tkm2x32b I257 (L546_0r0[31:0], L546_0r1[31:0], L546_0a, L548_0r0[31:0], L548_0r1[31:0], L548_0a, L549_0r0[31:0], L549_0r1[31:0], L549_0a, reset);
  tkf32mo0w0_o0w32 I258 (L549_0r0[31:0], L549_0r1[31:0], L549_0a, L550_0r, L550_0a, daddr_0r0[31:0], daddr_0r1[31:0], daddr_0a, reset);
  tko0m2_1nm2b1 I259 (L545_0r, L545_0a, L552_0r0[1:0], L552_0r1[1:0], L552_0a, reset);
  tko0m2_1nm2b2 I260 (L547_0r, L547_0a, L553_0r0[1:0], L553_0r1[1:0], L553_0a, reset);
  tkm2x2b I261 (L552_0r0[1:0], L552_0r1[1:0], L552_0a, L553_0r0[1:0], L553_0r1[1:0], L553_0a, L554_0r0[1:0], L554_0r1[1:0], L554_0a, reset);
  tkj2m0_2 I262 (L550_0r, L550_0a, L554_0r0[1:0], L554_0r1[1:0], L554_0a, L555_0r0[1:0], L555_0r1[1:0], L555_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I263 (L555_0r0[1:0], L555_0r1[1:0], L555_0a, L229_0r, L229_0a, L276_0r, L276_0a, reset);
  tkf3mo0w0_o0w3 I264 (L239_0r0[2:0], L239_0r1[2:0], L239_0a, L556_0r, L556_0a, L557_0r0[2:0], L557_0r1[2:0], L557_0a, reset);
  tkf3mo0w0_o0w3 I265 (L286_0r0[2:0], L286_0r1[2:0], L286_0a, L558_0r, L558_0a, L559_0r0[2:0], L559_0r1[2:0], L559_0a, reset);
  tkm2x3b I266 (L557_0r0[2:0], L557_0r1[2:0], L557_0a, L559_0r0[2:0], L559_0r1[2:0], L559_0a, L560_0r0[2:0], L560_0r1[2:0], L560_0a, reset);
  tkf3mo0w0_o0w3 I267 (L560_0r0[2:0], L560_0r1[2:0], L560_0a, L561_0r, L561_0a, daccess_0r0[2:0], daccess_0r1[2:0], daccess_0a, reset);
  tko0m2_1nm2b1 I268 (L556_0r, L556_0a, L563_0r0[1:0], L563_0r1[1:0], L563_0a, reset);
  tko0m2_1nm2b2 I269 (L558_0r, L558_0a, L564_0r0[1:0], L564_0r1[1:0], L564_0a, reset);
  tkm2x2b I270 (L563_0r0[1:0], L563_0r1[1:0], L563_0a, L564_0r0[1:0], L564_0r1[1:0], L564_0a, L565_0r0[1:0], L565_0r1[1:0], L565_0a, reset);
  tkj2m0_2 I271 (L561_0r, L561_0a, L565_0r0[1:0], L565_0r1[1:0], L565_0a, L566_0r0[1:0], L566_0r1[1:0], L566_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I272 (L566_0r0[1:0], L566_0r1[1:0], L566_0a, L240_0r, L240_0a, L287_0r, L287_0a, reset);
  tkj32m32_0 I273 (dread_0r0[31:0], dread_0r1[31:0], dread_0a, L251_0r, L251_0a, L249_0r0[31:0], L249_0r1[31:0], L249_0a, reset);
  tkf32mo0w0_o0w32 I274 (L295_0r0[31:0], L295_0r1[31:0], L295_0a, L296_0r, L296_0a, dwrite_0r0[31:0], dwrite_0r1[31:0], dwrite_0a, reset);
  tkr I275 (L2_0r, L2_0a, reset);
  tkr I276 (L6_0r, L6_0a, reset);
  tkr I277 (L10_0r, L10_0a, reset);
  tkr I278 (L14_0r, L14_0a, reset);
endmodule

module teak_Execute (op_0r0, op_0r1, op_0a, pc_0r0, pc_0r1, pc_0a, doFetch_0r0, doFetch_0r1, doFetch_0a, newPc_0r0, newPc_0r1, newPc_0a, daddr_0r0, daddr_0r1, daddr_0a, daccess_0r0, daccess_0r1, daccess_0a, dread_0r0, dread_0r1, dread_0a, dwrite_0r0, dwrite_0r1, dwrite_0a, reset);
  input [73:0] op_0r0;
  input [73:0] op_0r1;
  output op_0a;
  input [32:0] pc_0r0;
  input [32:0] pc_0r1;
  output pc_0a;
  output doFetch_0r0;
  output doFetch_0r1;
  input doFetch_0a;
  output [31:0] newPc_0r0;
  output [31:0] newPc_0r1;
  input newPc_0a;
  output [31:0] daddr_0r0;
  output [31:0] daddr_0r1;
  input daddr_0a;
  output [2:0] daccess_0r0;
  output [2:0] daccess_0r1;
  input daccess_0a;
  input [31:0] dread_0r0;
  input [31:0] dread_0r1;
  output dread_0a;
  output [31:0] dwrite_0r0;
  output [31:0] dwrite_0r1;
  input dwrite_0a;
  input reset;
  wire L3_0r;
  wire L3_0a;
  wire [31:0] L4_0r0;
  wire [31:0] L4_0r1;
  wire L4_0a;
  wire L6_0r;
  wire L6_0a;
  wire [31:0] L8_0r0;
  wire [31:0] L8_0r1;
  wire L8_0a;
  wire L9_0r;
  wire L9_0a;
  wire [6:0] L11_0r0;
  wire [6:0] L11_0r1;
  wire L11_0a;
  wire [31:0] L14_0r0;
  wire [31:0] L14_0r1;
  wire L14_0a;
  wire [31:0] L15_0r0;
  wire [31:0] L15_0r1;
  wire L15_0a;
  wire L17_0r0;
  wire L17_0r1;
  wire L17_0a;
  wire [2:0] L18_0r0;
  wire [2:0] L18_0r1;
  wire L18_0a;
  wire [4:0] L19_0r0;
  wire [4:0] L19_0r1;
  wire L19_0a;
  wire [4:0] L20_0r0;
  wire [4:0] L20_0r1;
  wire L20_0a;
  wire [4:0] L21_0r0;
  wire [4:0] L21_0r1;
  wire L21_0a;
  wire [4:0] L22_0r0;
  wire [4:0] L22_0r1;
  wire L22_0a;
  wire L23_0r0;
  wire L23_0r1;
  wire L23_0a;
  wire [31:0] L24_0r0;
  wire [31:0] L24_0r1;
  wire L24_0a;
  wire [31:0] L40_0r0;
  wire [31:0] L40_0r1;
  wire L40_0a;
  wire [31:0] L41_0r0;
  wire [31:0] L41_0r1;
  wire L41_0a;
  wire [31:0] L42_0r0;
  wire [31:0] L42_0r1;
  wire L42_0a;
  wire [31:0] L43_0r0;
  wire [31:0] L43_0r1;
  wire L43_0a;
  wire [31:0] L45_0r0;
  wire [31:0] L45_0r1;
  wire L45_0a;
  wire [3:0] L46_0r0;
  wire [3:0] L46_0r1;
  wire L46_0a;
  tkvv32_wo0w32_ro0w32 I0 (L4_0r0[31:0], L4_0r1[31:0], L4_0a, L6_0r, L6_0a, L6_0r, L6_0a, L8_0r0[31:0], L8_0r1[31:0], L8_0a, reset);
  teak_Alu I1 (L11_0r0[6:0], L11_0r1[6:0], L11_0a, L45_0r0[31:0], L45_0r1[31:0], L45_0a, L46_0r0[3:0], L46_0r1[3:0], L46_0a, L14_0r0[31:0], L14_0r1[31:0], L14_0a, L15_0r0[31:0], L15_0r1[31:0], L15_0a, reset);
  teak_RegBank I2 (L17_0r0, L17_0r1, L17_0a, L18_0r0[2:0], L18_0r1[2:0], L18_0a, L19_0r0[4:0], L19_0r1[4:0], L19_0a, L20_0r0[4:0], L20_0r1[4:0], L20_0a, L21_0r0[4:0], L21_0r1[4:0], L21_0a, L22_0r0[4:0], L22_0r1[4:0], L22_0a, L23_0r0, L23_0r1, L23_0a, L24_0r0[31:0], L24_0r1[31:0], L24_0a, L41_0r0[31:0], L41_0r1[31:0], L41_0a, L42_0r0[31:0], L42_0r1[31:0], L42_0a, L43_0r0[31:0], L43_0r1[31:0], L43_0a, reset);
  teak_ExecuteCtrl I3 (op_0r0[73:0], op_0r1[73:0], op_0a, pc_0r0[32:0], pc_0r1[32:0], pc_0a, doFetch_0r0, doFetch_0r1, doFetch_0a, newPc_0r0[31:0], newPc_0r1[31:0], newPc_0a, L17_0r0, L17_0r1, L17_0a, L18_0r0[2:0], L18_0r1[2:0], L18_0a, L19_0r0[4:0], L19_0r1[4:0], L19_0a, L20_0r0[4:0], L20_0r1[4:0], L20_0a, L21_0r0[4:0], L21_0r1[4:0], L21_0a, L22_0r0[4:0], L22_0r1[4:0], L22_0a, L23_0r0, L23_0r1, L23_0a, L40_0r0[31:0], L40_0r1[31:0], L40_0a, L41_0r0[31:0], L41_0r1[31:0], L41_0a, L42_0r0[31:0], L42_0r1[31:0], L42_0a, L43_0r0[31:0], L43_0r1[31:0], L43_0a, L11_0r0[6:0], L11_0r1[6:0], L11_0a, L45_0r0[31:0], L45_0r1[31:0], L45_0a, L46_0r0[3:0], L46_0r1[3:0], L46_0a, L14_0r0[31:0], L14_0r1[31:0], L14_0a, L15_0r0[31:0], L15_0r1[31:0], L15_0a, daddr_0r0[31:0], daddr_0r1[31:0], daddr_0a, daccess_0r0[2:0], daccess_0r1[2:0], daccess_0a, dread_0r0[31:0], dread_0r1[31:0], dread_0a, dwrite_0r0[31:0], dwrite_0r1[31:0], dwrite_0a, reset);
  tkj32m32_0 I4 (L40_0r0[31:0], L40_0r1[31:0], L40_0a, L3_0r, L3_0a, L4_0r0[31:0], L4_0r1[31:0], L4_0a, reset);
  tkf32mo0w0_o0w32 I5 (L8_0r0[31:0], L8_0r1[31:0], L8_0a, L9_0r, L9_0a, L24_0r0[31:0], L24_0r1[31:0], L24_0a, reset);
  tki I6 (L9_0r, L9_0a, L3_0r, L3_0a, reset);
endmodule

module teak_MemArbiter (faddr_0r0, faddr_0r1, faddr_0a, finst_0r0, finst_0r1, finst_0a, daddr_0r0, daddr_0r1, daddr_0a, daccess_0r0, daccess_0r1, daccess_0a, dread_0r0, dread_0r1, dread_0a, dwrite_0r0, dwrite_0r1, dwrite_0a, maddr_0r0, maddr_0r1, maddr_0a, maccess_0r0, maccess_0r1, maccess_0a, mread_0r0, mread_0r1, mread_0a, mwrite_0r0, mwrite_0r1, mwrite_0a, reset);
  input [31:0] faddr_0r0;
  input [31:0] faddr_0r1;
  output faddr_0a;
  output [31:0] finst_0r0;
  output [31:0] finst_0r1;
  input finst_0a;
  input [31:0] daddr_0r0;
  input [31:0] daddr_0r1;
  output daddr_0a;
  input [2:0] daccess_0r0;
  input [2:0] daccess_0r1;
  output daccess_0a;
  output [31:0] dread_0r0;
  output [31:0] dread_0r1;
  input dread_0a;
  input [31:0] dwrite_0r0;
  input [31:0] dwrite_0r1;
  output dwrite_0a;
  output [31:0] maddr_0r0;
  output [31:0] maddr_0r1;
  input maddr_0a;
  output [2:0] maccess_0r0;
  output [2:0] maccess_0r1;
  input maccess_0a;
  input [31:0] mread_0r0;
  input [31:0] mread_0r1;
  output mread_0a;
  output [31:0] mwrite_0r0;
  output [31:0] mwrite_0r1;
  input mwrite_0a;
  input reset;
  wire L2_0r;
  wire L2_0a;
  wire L3_0r;
  wire L3_0a;
  wire [31:0] L5_0r0;
  wire [31:0] L5_0r1;
  wire L5_0a;
  wire L6_0r;
  wire L6_0a;
  wire L7_0r;
  wire L7_0a;
  wire [2:0] L9_0r0;
  wire [2:0] L9_0r1;
  wire L9_0a;
  wire L10_0r;
  wire L10_0a;
  wire L11_0r;
  wire L11_0a;
  wire [31:0] L13_0r0;
  wire [31:0] L13_0r1;
  wire L13_0a;
  wire L14_0r;
  wire L14_0a;
  wire [31:0] L15_0r0;
  wire [31:0] L15_0r1;
  wire L15_0a;
  wire L17_0r;
  wire L17_0a;
  wire L18_0r;
  wire L18_0a;
  wire L19_0r;
  wire L19_0a;
  wire [31:0] L20_0r0;
  wire [31:0] L20_0r1;
  wire L20_0a;
  wire L22_0r;
  wire L22_0a;
  wire [31:0] L24_0r0;
  wire [31:0] L24_0r1;
  wire L24_0a;
  wire L25_0r;
  wire L25_0a;
  wire L26_0r;
  wire L26_0a;
  wire L27_0r;
  wire L27_0a;
  wire [31:0] L29_0r0;
  wire [31:0] L29_0r1;
  wire L29_0a;
  wire L30_0r;
  wire L30_0a;
  wire L31_0r;
  wire L31_0a;
  wire [2:0] L33_0r0;
  wire [2:0] L33_0r1;
  wire L33_0a;
  wire L34_0r;
  wire L34_0a;
  wire L35_0r;
  wire L35_0a;
  wire L36_0r0;
  wire L36_0r1;
  wire L36_0a;
  wire L37_0r;
  wire L37_0a;
  wire [31:0] L39_0r0;
  wire [31:0] L39_0r1;
  wire L39_0a;
  wire L40_0r;
  wire L40_0a;
  wire [31:0] L41_0r0;
  wire [31:0] L41_0r1;
  wire L41_0a;
  wire L43_0r;
  wire L43_0a;
  wire L44_0r;
  wire L44_0a;
  wire [31:0] L46_0r0;
  wire [31:0] L46_0r1;
  wire L46_0a;
  wire L47_0r;
  wire L47_0a;
  wire [31:0] L48_0r0;
  wire [31:0] L48_0r1;
  wire L48_0a;
  wire L50_0r;
  wire L50_0a;
  wire L51_0r;
  wire L51_0a;
  wire L52_0r;
  wire L52_0a;
  wire L53_0r;
  wire L53_0a;
  wire [31:0] L54_0r0;
  wire [31:0] L54_0r1;
  wire L54_0a;
  wire L55_0r;
  wire L55_0a;
  wire [2:0] L56_0r0;
  wire [2:0] L56_0r1;
  wire L56_0a;
  wire L57_0r;
  wire L57_0a;
  wire L59_0r;
  wire L59_0a;
  wire [31:0] L61_0r0;
  wire [31:0] L61_0r1;
  wire L61_0a;
  wire L62_0r;
  wire L62_0a;
  wire L63_0r;
  wire L63_0a;
  wire [2:0] L65_0r0;
  wire [2:0] L65_0r1;
  wire L65_0a;
  wire L66_0r;
  wire L66_0a;
  wire L67_0r;
  wire L67_0a;
  wire L68_0r;
  wire L68_0a;
  wire L69_0r;
  wire L69_0a;
  wire [1:0] L70_0r0;
  wire [1:0] L70_0r1;
  wire L70_0a;
  wire [1:0] L71_0r0;
  wire [1:0] L71_0r1;
  wire L71_0a;
  wire [1:0] L72_0r0;
  wire [1:0] L72_0r1;
  wire L72_0a;
  wire [1:0] L73_0r0;
  wire [1:0] L73_0r1;
  wire L73_0a;
  wire L74_0r;
  wire L74_0a;
  wire L79_0r;
  wire L79_0a;
  wire [31:0] L80_0r0;
  wire [31:0] L80_0r1;
  wire L80_0a;
  wire L81_0r;
  wire L81_0a;
  wire [31:0] L82_0r0;
  wire [31:0] L82_0r1;
  wire L82_0a;
  wire [31:0] L83_0r0;
  wire [31:0] L83_0r1;
  wire L83_0a;
  wire L84_0r;
  wire L84_0a;
  wire [1:0] L86_0r0;
  wire [1:0] L86_0r1;
  wire L86_0a;
  wire [1:0] L87_0r0;
  wire [1:0] L87_0r1;
  wire L87_0a;
  wire [1:0] L88_0r0;
  wire [1:0] L88_0r1;
  wire L88_0a;
  wire [1:0] L89_0r0;
  wire [1:0] L89_0r1;
  wire L89_0a;
  wire L90_0r;
  wire L90_0a;
  wire [2:0] L91_0r0;
  wire [2:0] L91_0r1;
  wire L91_0a;
  wire L92_0r;
  wire L92_0a;
  wire [2:0] L93_0r0;
  wire [2:0] L93_0r1;
  wire L93_0a;
  wire [2:0] L94_0r0;
  wire [2:0] L94_0r1;
  wire L94_0a;
  wire L95_0r;
  wire L95_0a;
  wire [1:0] L97_0r0;
  wire [1:0] L97_0r1;
  wire L97_0a;
  wire [1:0] L98_0r0;
  wire [1:0] L98_0r1;
  wire L98_0a;
  wire [1:0] L99_0r0;
  wire [1:0] L99_0r1;
  wire L99_0a;
  wire [1:0] L100_0r0;
  wire [1:0] L100_0r1;
  wire L100_0a;
  wire [1:0] L102_0r0;
  wire [1:0] L102_0r1;
  wire L102_0a;
  wire [1:0] L103_0r0;
  wire [1:0] L103_0r1;
  wire L103_0a;
  wire [1:0] L104_0r0;
  wire [1:0] L104_0r1;
  wire L104_0a;
  wire [33:0] L105_0r0;
  wire [33:0] L105_0r1;
  wire L105_0a;
  tko0m3_1nm3b1 I0 (L7_0r, L7_0a, L9_0r0[2:0], L9_0r1[2:0], L9_0a, reset);
  tkvmread32_wo0w32_ro0w32 I1 (L15_0r0[31:0], L15_0r1[31:0], L15_0a, L11_0r, L11_0a, L11_0r, L11_0a, L13_0r0[31:0], L13_0r1[31:0], L13_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0 I2 (L18_0r, L18_0a, L2_0r, L2_0a, L3_0r, L3_0a, L7_0r, L7_0a, L17_0r, L17_0a, reset);
  tkj0m0_0_0_0 I3 (L2_0r, L2_0a, L6_0r, L6_0a, L10_0r, L10_0a, L14_0r, L14_0a, L19_0r, L19_0a, reset);
  tkvfaddr32_wo0w32_ro0w32 I4 (L20_0r0[31:0], L20_0r1[31:0], L20_0a, L18_0r, L18_0a, L3_0r, L3_0a, L5_0r0[31:0], L5_0r1[31:0], L5_0a, reset);
  tkf32mo0w0_o0w32 I5 (faddr_0r0[31:0], faddr_0r1[31:0], faddr_0a, L22_0r, L22_0a, L24_0r0[31:0], L24_0r1[31:0], L24_0a, reset);
  tkj32m0_32 I6 (L25_0r, L25_0a, L24_0r0[31:0], L24_0r1[31:0], L24_0a, L20_0r0[31:0], L20_0r1[31:0], L20_0a, reset);
  tkvdwrite32_wo0w32_ro0w32 I7 (L41_0r0[31:0], L41_0r1[31:0], L41_0a, L37_0r, L37_0a, L37_0r, L37_0a, L39_0r0[31:0], L39_0r1[31:0], L39_0a, reset);
  tkvmread32_wo0w32_ro0w32 I8 (L48_0r0[31:0], L48_0r1[31:0], L48_0a, L44_0r, L44_0a, L44_0r, L44_0a, L46_0r0[31:0], L46_0r1[31:0], L46_0a, reset);
  tks1_o0w1_0o0w0_1o0w0 I9 (L36_0r0, L36_0r1, L36_0a, L43_0r, L43_0a, L50_0r, L50_0a, reset);
  tkm2x0b I10 (L40_0r, L40_0a, L47_0r, L47_0a, L51_0r, L51_0a, reset);
  tkf0mo0w0_o0w0_o0w0_o0w0 I11 (L52_0r, L52_0a, L26_0r, L26_0a, L27_0r, L27_0a, L31_0r, L31_0a, L35_0r, L35_0a, reset);
  tkj0m0_0_0_0 I12 (L26_0r, L26_0a, L30_0r, L30_0a, L34_0r, L34_0a, L51_0r, L51_0a, L53_0r, L53_0a, reset);
  tkvdaddr32_wo0w32_ro0w32 I13 (L54_0r0[31:0], L54_0r1[31:0], L54_0a, L55_0r, L55_0a, L27_0r, L27_0a, L29_0r0[31:0], L29_0r1[31:0], L29_0a, reset);
  tkvdaccess3_wo0w3_ro0w3o0w1 I14 (L56_0r0[2:0], L56_0r1[2:0], L56_0a, L57_0r, L57_0a, L31_0r, L31_0a, L35_0r, L35_0a, L33_0r0[2:0], L33_0r1[2:0], L33_0a, L36_0r0, L36_0r1, L36_0a, reset);
  tkj0m0_0 I15 (L55_0r, L55_0a, L57_0r, L57_0a, L52_0r, L52_0a, reset);
  tkf32mo0w0_o0w32 I16 (daddr_0r0[31:0], daddr_0r1[31:0], daddr_0a, L59_0r, L59_0a, L61_0r0[31:0], L61_0r1[31:0], L61_0a, reset);
  tkj32m0_32 I17 (L62_0r, L62_0a, L61_0r0[31:0], L61_0r1[31:0], L61_0a, L54_0r0[31:0], L54_0r1[31:0], L54_0a, reset);
  tkf3mo0w0_o0w3 I18 (daccess_0r0[2:0], daccess_0r1[2:0], daccess_0a, L63_0r, L63_0a, L65_0r0[2:0], L65_0r1[2:0], L65_0a, reset);
  tkj3m0_3 I19 (L66_0r, L66_0a, L65_0r0[2:0], L65_0r1[2:0], L65_0a, L56_0r0[2:0], L56_0r1[2:0], L56_0a, reset);
  tkj0m0_0 I20 (L59_0r, L59_0a, L63_0r, L63_0a, L67_0r, L67_0a, reset);
  tkf0mo0w0_o0w0 I21 (L68_0r, L68_0a, L62_0r, L62_0a, L66_0r, L66_0a, reset);
  tko0m2_1nm2b1 I22 (L22_0r, L22_0a, L70_0r0[1:0], L70_0r1[1:0], L70_0a, reset);
  tko0m2_1nm2b2 I23 (L67_0r, L67_0a, L71_0r0[1:0], L71_0r1[1:0], L71_0a, reset);
  tka2x2b I24 (L70_0r0[1:0], L70_0r1[1:0], L70_0a, L71_0r0[1:0], L71_0r1[1:0], L71_0a, L72_0r0[1:0], L72_0r1[1:0], L72_0a, reset);
  tkj2m0_2 I25 (L69_0r, L69_0a, L72_0r0[1:0], L72_0r1[1:0], L72_0a, L73_0r0[1:0], L73_0r1[1:0], L73_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I26 (L73_0r0[1:0], L73_0r1[1:0], L73_0a, L25_0r, L25_0a, L68_0r, L68_0a, reset);
  tkm2x0b I27 (L19_0r, L19_0a, L53_0r, L53_0a, L74_0r, L74_0a, reset);
  tkf32mo0w0_o0w32 I28 (L13_0r0[31:0], L13_0r1[31:0], L13_0a, L14_0r, L14_0a, finst_0r0[31:0], finst_0r1[31:0], finst_0a, reset);
  tkf32mo0w0_o0w32 I29 (L46_0r0[31:0], L46_0r1[31:0], L46_0a, L47_0r, L47_0a, dread_0r0[31:0], dread_0r1[31:0], dread_0a, reset);
  tkj32m32_0 I30 (dwrite_0r0[31:0], dwrite_0r1[31:0], dwrite_0a, L43_0r, L43_0a, L41_0r0[31:0], L41_0r1[31:0], L41_0a, reset);
  tkf32mo0w0_o0w32 I31 (L5_0r0[31:0], L5_0r1[31:0], L5_0a, L79_0r, L79_0a, L80_0r0[31:0], L80_0r1[31:0], L80_0a, reset);
  tkf32mo0w0_o0w32 I32 (L29_0r0[31:0], L29_0r1[31:0], L29_0a, L81_0r, L81_0a, L82_0r0[31:0], L82_0r1[31:0], L82_0a, reset);
  tkm2x32b I33 (L80_0r0[31:0], L80_0r1[31:0], L80_0a, L82_0r0[31:0], L82_0r1[31:0], L82_0a, L83_0r0[31:0], L83_0r1[31:0], L83_0a, reset);
  tkf32mo0w0_o0w32 I34 (L83_0r0[31:0], L83_0r1[31:0], L83_0a, L84_0r, L84_0a, maddr_0r0[31:0], maddr_0r1[31:0], maddr_0a, reset);
  tko0m2_1nm2b1 I35 (L79_0r, L79_0a, L86_0r0[1:0], L86_0r1[1:0], L86_0a, reset);
  tko0m2_1nm2b2 I36 (L81_0r, L81_0a, L87_0r0[1:0], L87_0r1[1:0], L87_0a, reset);
  tkm2x2b I37 (L86_0r0[1:0], L86_0r1[1:0], L86_0a, L87_0r0[1:0], L87_0r1[1:0], L87_0a, L88_0r0[1:0], L88_0r1[1:0], L88_0a, reset);
  tkj2m0_2 I38 (L84_0r, L84_0a, L88_0r0[1:0], L88_0r1[1:0], L88_0a, L89_0r0[1:0], L89_0r1[1:0], L89_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I39 (L89_0r0[1:0], L89_0r1[1:0], L89_0a, L6_0r, L6_0a, L30_0r, L30_0a, reset);
  tkf3mo0w0_o0w3 I40 (L9_0r0[2:0], L9_0r1[2:0], L9_0a, L90_0r, L90_0a, L91_0r0[2:0], L91_0r1[2:0], L91_0a, reset);
  tkf3mo0w0_o0w3 I41 (L33_0r0[2:0], L33_0r1[2:0], L33_0a, L92_0r, L92_0a, L93_0r0[2:0], L93_0r1[2:0], L93_0a, reset);
  tkm2x3b I42 (L91_0r0[2:0], L91_0r1[2:0], L91_0a, L93_0r0[2:0], L93_0r1[2:0], L93_0a, L94_0r0[2:0], L94_0r1[2:0], L94_0a, reset);
  tkf3mo0w0_o0w3 I43 (L94_0r0[2:0], L94_0r1[2:0], L94_0a, L95_0r, L95_0a, maccess_0r0[2:0], maccess_0r1[2:0], maccess_0a, reset);
  tko0m2_1nm2b1 I44 (L90_0r, L90_0a, L97_0r0[1:0], L97_0r1[1:0], L97_0a, reset);
  tko0m2_1nm2b2 I45 (L92_0r, L92_0a, L98_0r0[1:0], L98_0r1[1:0], L98_0a, reset);
  tkm2x2b I46 (L97_0r0[1:0], L97_0r1[1:0], L97_0a, L98_0r0[1:0], L98_0r1[1:0], L98_0a, L99_0r0[1:0], L99_0r1[1:0], L99_0a, reset);
  tkj2m0_2 I47 (L95_0r, L95_0a, L99_0r0[1:0], L99_0r1[1:0], L99_0a, L100_0r0[1:0], L100_0r1[1:0], L100_0a, reset);
  tks2_o0w2_1o0w0_2o0w0 I48 (L100_0r0[1:0], L100_0r1[1:0], L100_0a, L10_0r, L10_0a, L34_0r, L34_0a, reset);
  tko0m2_1nm2b1 I49 (L17_0r, L17_0a, L102_0r0[1:0], L102_0r1[1:0], L102_0a, reset);
  tko0m2_1nm2b2 I50 (L50_0r, L50_0a, L103_0r0[1:0], L103_0r1[1:0], L103_0a, reset);
  tkm2x2b I51 (L102_0r0[1:0], L102_0r1[1:0], L102_0a, L103_0r0[1:0], L103_0r1[1:0], L103_0a, L104_0r0[1:0], L104_0r1[1:0], L104_0a, reset);
  tkj34m32_2 I52 (mread_0r0[31:0], mread_0r1[31:0], mread_0a, L104_0r0[1:0], L104_0r1[1:0], L104_0a, L105_0r0[33:0], L105_0r1[33:0], L105_0a, reset);
  tks34_o32w2_1o0w32_2o0w32 I53 (L105_0r0[33:0], L105_0r1[33:0], L105_0a, L15_0r0[31:0], L15_0r1[31:0], L15_0a, L48_0r0[31:0], L48_0r1[31:0], L48_0a, reset);
  tkf32mo0w0_o0w32 I54 (L39_0r0[31:0], L39_0r1[31:0], L39_0a, L40_0r, L40_0a, mwrite_0r0[31:0], mwrite_0r1[31:0], mwrite_0a, reset);
  tki I55 (L74_0r, L74_0a, L69_0r, L69_0a, reset);
endmodule

module teak_Sparkler2 (a_0r0, a_0r1, a_0a, access_0r0, access_0r1, access_0a, di_0r0, di_0r1, di_0a, do_0r0, do_0r1, do_0a, reset);
  output [31:0] a_0r0;
  output [31:0] a_0r1;
  input a_0a;
  output [2:0] access_0r0;
  output [2:0] access_0r1;
  input access_0a;
  input [31:0] di_0r0;
  input [31:0] di_0r1;
  output di_0a;
  output [31:0] do_0r0;
  output [31:0] do_0r1;
  input do_0a;
  input reset;
  wire L3_0r;
  wire L3_0a;
  wire [64:0] L4_0r0;
  wire [64:0] L4_0r1;
  wire L4_0a;
  wire L6_0r;
  wire L6_0a;
  wire [64:0] L8_0r0;
  wire [64:0] L8_0r1;
  wire L8_0a;
  wire L9_0r;
  wire L9_0a;
  wire L13_0r;
  wire L13_0a;
  wire [73:0] L14_0r0;
  wire [73:0] L14_0r1;
  wire L14_0a;
  wire L16_0r;
  wire L16_0a;
  wire [73:0] L18_0r0;
  wire [73:0] L18_0r1;
  wire L18_0a;
  wire L19_0r;
  wire L19_0a;
  wire L23_0r;
  wire L23_0a;
  wire [32:0] L24_0r0;
  wire [32:0] L24_0r1;
  wire L24_0a;
  wire L26_0r;
  wire L26_0a;
  wire [32:0] L28_0r0;
  wire [32:0] L28_0r1;
  wire L28_0a;
  wire L29_0r;
  wire L29_0a;
  wire L33_0r;
  wire L33_0a;
  wire L34_0r0;
  wire L34_0r1;
  wire L34_0a;
  wire L36_0r;
  wire L36_0a;
  wire L38_0r0;
  wire L38_0r1;
  wire L38_0a;
  wire L39_0r;
  wire L39_0a;
  wire L43_0r;
  wire L43_0a;
  wire L44_0r0;
  wire L44_0r1;
  wire L44_0a;
  wire L46_0r;
  wire L46_0a;
  wire L48_0r0;
  wire L48_0r1;
  wire L48_0a;
  wire L49_0r;
  wire L49_0a;
  wire L53_0r;
  wire L53_0a;
  wire [31:0] L54_0r0;
  wire [31:0] L54_0r1;
  wire L54_0a;
  wire L56_0r;
  wire L56_0a;
  wire [31:0] L58_0r0;
  wire [31:0] L58_0r1;
  wire L58_0a;
  wire L59_0r;
  wire L59_0a;
  wire L61_0r0;
  wire L61_0r1;
  wire L61_0a;
  wire L62_0r0;
  wire L62_0r1;
  wire L62_0a;
  wire L64_0r0;
  wire L64_0r1;
  wire L64_0a;
  wire [31:0] L65_0r0;
  wire [31:0] L65_0r1;
  wire L65_0a;
  wire [64:0] L66_0r0;
  wire [64:0] L66_0r1;
  wire L66_0a;
  wire [31:0] L68_0r0;
  wire [31:0] L68_0r1;
  wire L68_0a;
  wire [64:0] L70_0r0;
  wire [64:0] L70_0r1;
  wire L70_0a;
  wire [73:0] L71_0r0;
  wire [73:0] L71_0r1;
  wire L71_0a;
  wire [32:0] L72_0r0;
  wire [32:0] L72_0r1;
  wire L72_0a;
  wire [73:0] L74_0r0;
  wire [73:0] L74_0r1;
  wire L74_0a;
  wire [32:0] L75_0r0;
  wire [32:0] L75_0r1;
  wire L75_0a;
  wire L76_0r0;
  wire L76_0r1;
  wire L76_0a;
  wire [31:0] L77_0r0;
  wire [31:0] L77_0r1;
  wire L77_0a;
  wire [31:0] L80_0r0;
  wire [31:0] L80_0r1;
  wire L80_0a;
  wire [31:0] L83_0r0;
  wire [31:0] L83_0r1;
  wire L83_0a;
  wire [31:0] L85_0r0;
  wire [31:0] L85_0r1;
  wire L85_0a;
  wire [2:0] L86_0r0;
  wire [2:0] L86_0r1;
  wire L86_0a;
  wire [31:0] L88_0r0;
  wire [31:0] L88_0r1;
  wire L88_0a;
  tkvv65_wo0w65_ro0w65 I0 (L4_0r0[64:0], L4_0r1[64:0], L4_0a, L6_0r, L6_0a, L6_0r, L6_0a, L8_0r0[64:0], L8_0r1[64:0], L8_0a, reset);
  tkvv74_wo0w74_ro0w74 I1 (L14_0r0[73:0], L14_0r1[73:0], L14_0a, L16_0r, L16_0a, L16_0r, L16_0a, L18_0r0[73:0], L18_0r1[73:0], L18_0a, reset);
  tkvv33_wo0w33_ro0w33 I2 (L24_0r0[32:0], L24_0r1[32:0], L24_0a, L26_0r, L26_0a, L26_0r, L26_0a, L28_0r0[32:0], L28_0r1[32:0], L28_0a, reset);
  tkvv1_wo0w1_ro0w1 I3 (L34_0r0, L34_0r1, L34_0a, L36_0r, L36_0a, L36_0r, L36_0a, L38_0r0, L38_0r1, L38_0a, reset);
  tkvv1_wo0w1_ro0w1 I4 (L44_0r0, L44_0r1, L44_0a, L46_0r, L46_0a, L46_0r, L46_0a, L48_0r0, L48_0r1, L48_0a, reset);
  tkvv32_wo0w32_ro0w32 I5 (L54_0r0[31:0], L54_0r1[31:0], L54_0a, L56_0r, L56_0a, L56_0r, L56_0a, L58_0r0[31:0], L58_0r1[31:0], L58_0a, reset);
  teak_FetchInitial I6 (L61_0r0, L61_0r1, L61_0a, L62_0r0, L62_0r1, L62_0a, reset);
  teak_Fetch I7 (L64_0r0, L64_0r1, L64_0a, L65_0r0[31:0], L65_0r1[31:0], L65_0a, L66_0r0[64:0], L66_0r1[64:0], L66_0a, L83_0r0[31:0], L83_0r1[31:0], L83_0a, L68_0r0[31:0], L68_0r1[31:0], L68_0a, reset);
  teak_Decode I8 (L70_0r0[64:0], L70_0r1[64:0], L70_0a, L71_0r0[73:0], L71_0r1[73:0], L71_0a, L72_0r0[32:0], L72_0r1[32:0], L72_0a, reset);
  teak_Execute I9 (L74_0r0[73:0], L74_0r1[73:0], L74_0a, L75_0r0[32:0], L75_0r1[32:0], L75_0a, L76_0r0, L76_0r1, L76_0a, L77_0r0[31:0], L77_0r1[31:0], L77_0a, L85_0r0[31:0], L85_0r1[31:0], L85_0a, L86_0r0[2:0], L86_0r1[2:0], L86_0a, L80_0r0[31:0], L80_0r1[31:0], L80_0a, L88_0r0[31:0], L88_0r1[31:0], L88_0a, reset);
  teak_MemArbiter I10 (L83_0r0[31:0], L83_0r1[31:0], L83_0a, L68_0r0[31:0], L68_0r1[31:0], L68_0a, L85_0r0[31:0], L85_0r1[31:0], L85_0a, L86_0r0[2:0], L86_0r1[2:0], L86_0a, L80_0r0[31:0], L80_0r1[31:0], L80_0a, L88_0r0[31:0], L88_0r1[31:0], L88_0a, a_0r0[31:0], a_0r1[31:0], a_0a, access_0r0[2:0], access_0r1[2:0], access_0a, di_0r0[31:0], di_0r1[31:0], di_0a, do_0r0[31:0], do_0r1[31:0], do_0a, reset);
  tkf32mo0w0_o0w32 I11 (L58_0r0[31:0], L58_0r1[31:0], L58_0a, L59_0r, L59_0a, L65_0r0[31:0], L65_0r1[31:0], L65_0a, reset);
  tkj32m32_0 I12 (L77_0r0[31:0], L77_0r1[31:0], L77_0a, L53_0r, L53_0a, L54_0r0[31:0], L54_0r1[31:0], L54_0a, reset);
  tkf1mo0w0_o0w1 I13 (L48_0r0, L48_0r1, L48_0a, L49_0r, L49_0a, L64_0r0, L64_0r1, L64_0a, reset);
  tkj1m1_0 I14 (L62_0r0, L62_0r1, L62_0a, L43_0r, L43_0a, L44_0r0, L44_0r1, L44_0a, reset);
  tkf1mo0w0_o0w1 I15 (L38_0r0, L38_0r1, L38_0a, L39_0r, L39_0a, L61_0r0, L61_0r1, L61_0a, reset);
  tkj1m1_0 I16 (L76_0r0, L76_0r1, L76_0a, L33_0r, L33_0a, L34_0r0, L34_0r1, L34_0a, reset);
  tkf33mo0w0_o0w33 I17 (L28_0r0[32:0], L28_0r1[32:0], L28_0a, L29_0r, L29_0a, L75_0r0[32:0], L75_0r1[32:0], L75_0a, reset);
  tkj33m33_0 I18 (L72_0r0[32:0], L72_0r1[32:0], L72_0a, L23_0r, L23_0a, L24_0r0[32:0], L24_0r1[32:0], L24_0a, reset);
  tkf74mo0w0_o0w74 I19 (L18_0r0[73:0], L18_0r1[73:0], L18_0a, L19_0r, L19_0a, L74_0r0[73:0], L74_0r1[73:0], L74_0a, reset);
  tkj74m74_0 I20 (L71_0r0[73:0], L71_0r1[73:0], L71_0a, L13_0r, L13_0a, L14_0r0[73:0], L14_0r1[73:0], L14_0a, reset);
  tkf65mo0w0_o0w65 I21 (L8_0r0[64:0], L8_0r1[64:0], L8_0a, L9_0r, L9_0a, L70_0r0[64:0], L70_0r1[64:0], L70_0a, reset);
  tkj65m65_0 I22 (L66_0r0[64:0], L66_0r1[64:0], L66_0a, L3_0r, L3_0a, L4_0r0[64:0], L4_0r1[64:0], L4_0a, reset);
  tki I23 (L9_0r, L9_0a, L3_0r, L3_0a, reset);
  tki I24 (L19_0r, L19_0a, L13_0r, L13_0a, reset);
  tki I25 (L29_0r, L29_0a, L23_0r, L23_0a, reset);
  tki I26 (L39_0r, L39_0a, L33_0r, L33_0a, reset);
  tki I27 (L49_0r, L49_0a, L43_0r, L43_0a, reset);
  tki I28 (L59_0r, L59_0a, L53_0r, L53_0a, reset);
endmodule

// Netlist costs:
// teak_Alu: AND2*6339 AO22*423 AO222*66 BUFF*11497 C2*1275 C2R*234 C3*1371 GND*278 INV*494 NAND2*464 NAND3*20 NOR2*463 NOR3*917 OR2*1958 OR3*283
// teak_Decode: AND2*2266 AO22*84 BUFF*4840 C2*434 C2R*204 C3*711 GND*563 INV*91 NAND2*180 NAND3*78 NOR2*333 NOR3*491 OR2*1077 OR3*7
// teak_Execute: AND2*28408 AO22*1641 AO222*138 BUFF*23895 C2*4926 C2R*906 C3*5123 GND*715 INV*855 NAND2*798 NAND3*883 NOR2*2638 NOR3*4189 OR2*9098 OR3*365
// teak_ExecuteCtrl: AND2*3352 AO22*355 AO222*64 BUFF*4902 C2*609 C2R*244 C3*945 GND*222 INV*99 NAND2*70 NAND3*48 NOR2*432 NOR3*514 OR2*1312 OR3*73
// teak_Fetch: AND2*1280 AO22*136 AO222*64 BUFF*2095 C2*90 C2R*40 C3*455 GND*91 INV*70 NAND2*65 NOR2*150 NOR3*196 OR2*325 OR3*85
// teak_FetchInitial: AND2*31 AO22*2 BUFF*66 C2*9 C2R*16 C3*11 GND*11 INV*1 NOR2*8 NOR3*1 OR2*22 OR3*11
// teak_MemArbiter: AND2*1318 AO22*172 BUFF*1722 C2*218 C2R*30 C3*209 GND*19 INV*12 MUTEX*1 NAND2*1 NOR2*176 NOR3*164 OR2*406
// teak_RegBank: AND2*18492 AO22*827 AO222*8 BUFF*7200 C2*3035 C2R*428 C3*2777 GND*215 INV*258 NAND2*264 NAND3*815 NOR2*1710 NOR3*2726 OR2*5794 OR3*9
// teak_Shifter: AND2*3400 AO22*177 BUFF*5333 C2*288 C2R*130 C3*499 GND*173 INV*389 NAND2*375 NAND3*7 NOR2*199 NOR3*558 OR2*974 OR3*10
// teak_Sparkler2: AND2*34751 AO22*2265 AO222*202 BUFF*34519 C2*5703 C2R*1196 C3*6711 GND*1399 INV*1053 MUTEX*1 NAND2*1044 NAND3*961 NOR2*3517 NOR3*5247 OR2*11146 OR3*468
// tka2x2b: AND2*10 C2*2 C2R*2 INV*2 MUTEX*1 OR2*8
// tkf0mo0w0_o0w0: BUFF*2 C2*1
// tkf0mo0w0_o0w0_o0w0: BUFF*3 C3*1
// tkf0mo0w0_o0w0_o0w0_o0w0: BUFF*5 C2*1 C3*1
// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0: BUFF*6 C2*1 C3*2
// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0: BUFF*8 C3*3
// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0: BUFF*8 C2*1 C3*3
// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0: BUFF*12 C2*1 C3*4
// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0: BUFF*12 C2*2 C3*4
// tkf0mo0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0_o0w0: BUFF*14 C2*3 C3*5
// tkf1mo0w0_o0w1: BUFF*4 C3*1 OR2*1
// tkf2mo0w0_o0w2: BUFF*6 C3*1 OR2*1
// tkf2mo0w1: BUFF*1 C2*4 OR2*2
// tkf32mo0w0_o0w32: BUFF*66 C3*1 OR2*1
// tkf33mo0w0_o0w33: BUFF*68 C3*1 OR2*1
// tkf33mo0w32: BUFF*63 C2*4 OR2*2
// tkf34mo1w33: BUFF*65 C2*4 OR2*2
// tkf3mo0w0_o0w3: BUFF*8 C3*1 OR2*1
// tkf4mo0w0: BUFF*2 C2*3 C3*1 OR2*5
// tkf4mo0w0_o0w4: BUFF*10 C3*1 OR2*1
// tkf4mo0w3: BUFF*5 C2*4 OR2*2
// tkf5mo0w0_o0w5: BUFF*12 C3*1 OR2*1
// tkf65mo0w0_o0w65: BUFF*132 C3*1 OR2*1
// tkf74mo0w0_o0w74: BUFF*150 C3*1 OR2*1
// tkf7mo0w0_o0w7: BUFF*16 C3*1 OR2*1
// tki: AND2*1 AO22*3 INV*3
// tkj0m0_0: BUFF*2 C2*1
// tkj0m0_0_0: BUFF*3 C3*1
// tkj0m0_0_0_0: BUFF*5 C2*1 C3*1
// tkj0m0_0_0_0_0_0: BUFF*6 C2*1 C3*2
// tkj0m0_0_0_0_0_0_0: BUFF*8 C3*3
// tkj0m0_0_0_0_0_0_0_0: BUFF*8 C2*1 C3*3
// tkj11m0_11: BUFF*45 C2*2
// tkj12m6_6: BUFF*49 C2*2 OR2*1
// tkj15m5_5_5: BUFF*61 C2*3 OR2*2
// tkj1m1_0: BUFF*5 C2*2
// tkj24m2_22: BUFF*97 C2*2 OR2*1
// tkj2m0_2: BUFF*9 C2*2
// tkj2m1_1: BUFF*9 C2*2 OR2*1
// tkj2m2_0: BUFF*9 C2*2
// tkj32m0_32: BUFF*129 C2*2
// tkj32m10_22: BUFF*129 C2*2 OR2*1
// tkj32m16_16: BUFF*129 C2*2 OR2*1
// tkj32m1_31: BUFF*129 C2*2 OR2*1
// tkj32m24_8: BUFF*129 C2*2 OR2*1
// tkj32m28_4: BUFF*129 C2*2 OR2*1
// tkj32m2_30: BUFF*129 C2*2 OR2*1
// tkj32m30_2: BUFF*129 C2*2 OR2*1
// tkj32m31_1: BUFF*129 C2*2 OR2*1
// tkj32m32_0: BUFF*129 C2*2
// tkj32m4_28: BUFF*129 C2*2 OR2*1
// tkj32m8_24: BUFF*129 C2*2 OR2*1
// tkj33m0_33: BUFF*133 C2*2
// tkj33m1_32: BUFF*133 C2*2 OR2*1
// tkj33m32_1: BUFF*133 C2*2 OR2*1
// tkj33m33_0: BUFF*133 C2*2
// tkj34m32_2: BUFF*137 C2*2 OR2*1
// tkj35m32_3: BUFF*141 C2*2 OR2*1
// tkj3m0_3: BUFF*13 C2*2
// tkj3m1_1_1: BUFF*13 C2*3 OR2*2
// tkj3m1_2: BUFF*13 C2*2 OR2*1
// tkj3m3_0: BUFF*13 C2*2
// tkj4m0_4: BUFF*17 C2*2
// tkj4m1_1_1_1: BUFF*18 C2*2 C3*1 OR2*3
// tkj4m3_1: BUFF*17 C2*2 OR2*1
// tkj4m4_0: BUFF*17 C2*2
// tkj5m0_5: BUFF*21 C2*2
// tkj5m5_0: BUFF*21 C2*2
// tkj64m32_32: BUFF*257 C2*2 OR2*1
// tkj65m32_33: BUFF*261 C2*2 OR2*1
// tkj65m65_0: BUFF*261 C2*2
// tkj66m33_33: BUFF*265 C2*2 OR2*1
// tkj74m3_4_3_15_1_5_6_1_32_4: BUFF*304 C2*2 C3*4 OR2*9
// tkj74m74_0: BUFF*297 C2*2
// tkj7m0_7: BUFF*29 C2*2
// tkj7m4_3: BUFF*29 C2*2 OR2*1
// tkj7m6_1: BUFF*29 C2*2 OR2*1
// tkj7m7_0: BUFF*29 C2*2
// tkj8m0_8: BUFF*33 C2*2
// tkm11x0b: C2R*22 INV*1 NAND3*1 NOR2*2 NOR3*3 OR2*1
// tkm11x11b: AND2*242 BUFF*11 C2*22 C2R*22 C3*44 INV*23 NAND3*23 NOR2*24 NOR3*69 OR2*144
// tkm11x3b: AND2*66 C2R*22 C3*11 INV*7 NAND3*7 NOR2*8 NOR3*21 OR2*40
// tkm11x4b: AND2*88 BUFF*11 C2*11 C2R*22 C3*11 INV*9 NAND3*9 NOR2*10 NOR3*27 OR2*53
// tkm2x0b: C2R*4 NOR2*1 OR2*1
// tkm2x1b: AND2*4 BUFF*2 C2R*4 NOR2*1 OR2*5
// tkm2x2b: AND2*8 C2*2 C2R*4 NOR2*1 OR2*9
// tkm2x32b: AND2*128 BUFF*2 C2*6 C2R*4 C3*28 NOR2*1 OR2*129
// tkm2x3b: AND2*12 C2R*4 C3*2 NOR2*1 OR2*13
// tkm2x4b: AND2*16 BUFF*2 C2*2 C2R*4 C3*2 NOR2*1 OR2*17
// tkm3x0b: C2R*6 NOR2*1 OR3*1
// tkm3x1b: AND2*6 BUFF*3 C2R*6 NOR2*1 OR2*3 OR3*3
// tkm3x2b: AND2*12 C2*3 C2R*6 NOR2*1 OR2*6 OR3*5
// tkm3x32b: AND2*192 BUFF*3 C2*9 C2R*6 C3*42 NOR2*1 OR2*96 OR3*65
// tkm3x33b: AND2*198 BUFF*3 C2*6 C2R*6 C3*45 NOR2*1 OR2*99 OR3*67
// tkm3x3b: AND2*18 C2R*6 C3*3 NOR2*1 OR2*9 OR3*7
// tkm3x7b: AND2*42 BUFF*3 C2R*6 C3*9 NOR2*1 OR2*21 OR3*15
// tkm4x0b: C2R*8 INV*1 NAND2*1 NOR2*1 NOR3*1
// tkm4x1b: AND2*8 BUFF*4 C2R*8 INV*3 NAND2*3 NOR2*1 NOR3*3 OR2*4
// tkm4x32b: AND2*256 BUFF*4 C2*12 C2R*8 C3*56 INV*65 NAND2*65 NOR2*1 NOR3*65 OR2*128
// tkm4x4b: AND2*32 BUFF*4 C2*4 C2R*8 C3*4 INV*9 NAND2*9 NOR2*1 NOR3*9 OR2*16
// tkm5x0b: C2R*10 NAND2*1 NOR2*2 NOR3*1
// tkm5x32b: AND2*320 BUFF*5 C2*15 C2R*10 C3*70 NAND2*65 NOR2*66 NOR3*65 OR2*160
// tkm5x5b: AND2*50 C2*10 C2R*10 C3*5 NAND2*11 NOR2*12 NOR3*11 OR2*25
// tkm5x74b: AND2*740 BUFF*5 C2*5 C2R*10 C3*180 NAND2*149 NOR2*150 NOR3*149 OR2*370
// tkm7x0b: C2R*14 INV*1 NAND3*1 NOR2*1 NOR3*2
// tkm7x32b: AND2*448 BUFF*7 C2*21 C2R*14 C3*98 INV*65 NAND3*65 NOR2*1 NOR3*130 OR2*224
// tkm7x7b: AND2*98 BUFF*7 C2R*14 C3*21 INV*15 NAND3*15 NOR2*1 NOR3*30 OR2*49
// tkm8x0b: C2R*16 NAND3*1 NOR2*2 NOR3*2
// tkm8x1b: AND2*16 BUFF*8 C2R*16 NAND3*3 NOR2*4 NOR3*6 OR2*8
// tkm8x32b: AND2*512 BUFF*8 C2*24 C2R*16 C3*112 NAND3*65 NOR2*66 NOR3*130 OR2*256
// tkm8x8b: AND2*128 C2*8 C2R*16 C3*24 NAND3*17 NOR2*18 NOR3*34 OR2*64
// tko0m10_1nm10b0: BUFF*11 GND*10
// tko0m11_1nm11b1: BUFF*12 GND*11
// tko0m11_1nm11b10: BUFF*12 GND*11
// tko0m11_1nm11b100: BUFF*12 GND*11
// tko0m11_1nm11b2: BUFF*12 GND*11
// tko0m11_1nm11b20: BUFF*12 GND*11
// tko0m11_1nm11b200: BUFF*12 GND*11
// tko0m11_1nm11b4: BUFF*12 GND*11
// tko0m11_1nm11b40: BUFF*12 GND*11
// tko0m11_1nm11b400: BUFF*12 GND*11
// tko0m11_1nm11b8: BUFF*12 GND*11
// tko0m11_1nm11b80: BUFF*12 GND*11
// tko0m15_1nm15b0: BUFF*16 GND*15
// tko0m16_1nm16b0: BUFF*17 GND*16
// tko0m16_1nm16bffff: BUFF*17 GND*16
// tko0m1_1nm1b0: BUFF*2 GND*1
// tko0m1_1nm1b1: BUFF*2 GND*1
// tko0m2_1nm2b0: BUFF*3 GND*2
// tko0m2_1nm2b1: BUFF*3 GND*2
// tko0m2_1nm2b2: BUFF*3 GND*2
// tko0m2_1nm2b3: BUFF*3 GND*2
// tko0m32_1nm32b0: BUFF*33 GND*32
// tko0m3_1nm3b0: BUFF*4 GND*3
// tko0m3_1nm3b1: BUFF*4 GND*3
// tko0m3_1nm3b2: BUFF*4 GND*3
// tko0m3_1nm3b3: BUFF*4 GND*3
// tko0m3_1nm3b4: BUFF*4 GND*3
// tko0m3_1nm3b5: BUFF*4 GND*3
// tko0m4_1nm4b0: BUFF*5 GND*4
// tko0m4_1nm4b1: BUFF*5 GND*4
// tko0m4_1nm4b2: BUFF*5 GND*4
// tko0m4_1nm4b3: BUFF*5 GND*4
// tko0m4_1nm4b4: BUFF*5 GND*4
// tko0m4_1nm4b5: BUFF*5 GND*4
// tko0m4_1nm4b6: BUFF*5 GND*4
// tko0m4_1nm4b7: BUFF*5 GND*4
// tko0m4_1nm4b8: BUFF*5 GND*4
// tko0m4_1nm4bb: BUFF*5 GND*4
// tko0m4_1nm4bd: BUFF*5 GND*4
// tko0m4_1nm4bf: BUFF*5 GND*4
// tko0m5_1nm5b0: BUFF*6 GND*5
// tko0m5_1nm5b1: BUFF*6 GND*5
// tko0m5_1nm5b10: BUFF*6 GND*5
// tko0m5_1nm5b2: BUFF*6 GND*5
// tko0m5_1nm5b4: BUFF*6 GND*5
// tko0m5_1nm5b8: BUFF*6 GND*5
// tko0m6_1nm6b0: BUFF*7 GND*6
// tko0m6_1nm6b4: BUFF*7 GND*6
// tko0m74_1nm74b1c00000000000000040: BUFF*75 GND*74
// tko0m7_1nm7b1: BUFF*8 GND*7
// tko0m7_1nm7b10: BUFF*8 GND*7
// tko0m7_1nm7b2: BUFF*8 GND*7
// tko0m7_1nm7b20: BUFF*8 GND*7
// tko0m7_1nm7b4: BUFF*8 GND*7
// tko0m7_1nm7b40: BUFF*8 GND*7
// tko0m7_1nm7b8: BUFF*8 GND*7
// tko0m8_1nm8b0: BUFF*9 GND*8
// tko0m8_1nm8b1: BUFF*9 GND*8
// tko0m8_1nm8b10: BUFF*9 GND*8
// tko0m8_1nm8b2: BUFF*9 GND*8
// tko0m8_1nm8b20: BUFF*9 GND*8
// tko0m8_1nm8b4: BUFF*9 GND*8
// tko0m8_1nm8b40: BUFF*9 GND*8
// tko0m8_1nm8b8: BUFF*9 GND*8
// tko0m8_1nm8b80: BUFF*9 GND*8
// tko0m8_1nm8bff: BUFF*9 GND*8
// tko12m1_1api0w6b_2api6w6b_3eqt1o0w6bt2o0w6b: BUFF*32 C2*44 OR2*12 OR3*5
// tko13m32_1ap19xi12w1b_2api0w13bt1o0w19b: BUFF*103
// tko1m1_1noti0w1b: BUFF*3
// tko24m32_1ap8xi23w1b_2api0w24bt1o0w8b: BUFF*81
// tko2m1_1api0w1b_2api1w1b_3andt1o0w1bt2o0w1b: BUFF*6 C2*4 OR3*1
// tko2m1_1api0w1b_2api1w1b_3net1o0w1bt2o0w1b: BUFF*7 C2*4 OR2*2
// tko2m1_1api0w1b_2api1w1b_3ort1o0w1bt2o0w1b: BUFF*6 C2*4 OR3*1
// tko2m1_1api0w1b_2api1w1b_3xort1o0w1bt2o0w1b: BUFF*5 C2*4 OR2*2
// tko2m2_1api0w1b_2api1w1b_3nm1b0_4apt1o0w1bt3o0w1b_5nm1b0_6apt2o0w1bt5o0w1b_7addt4o0w2bt6o0w2b: AO222*2 BUFF*16 C2*5 C3*8 GND*2 INV*2 NAND2*2 NOR3*2 OR2*4 OR3*1
// tko32m32_1noti0w32b: BUFF*65
// tko33m1_1api0w32b_2api32w1b_3nm31b0_4apt2o0w1bt3o0w31b_5eqt1o0w32bt4o0w32b: BUFF*194 C2*254 C3*15 GND*31 OR2*97 OR3*31
// tko35m33_1api0w32b_2api32w3b_3nm1b0_4apt1o0w32bt3o0w1b_5nm30b0_6apt2o0w3bt5o0w30b_7addt4o0w33bt6o0w33b: AO222*64 BUFF*236 C2*6 C3*272 GND*31 INV*64 NAND2*64 NOR3*64 OR2*37 OR3*1
// tko64m32_1api0w32b_2api32w32b_3andt1o0w32bt2o0w32b: BUFF*161 C2*128 OR3*32
// tko64m32_1api0w32b_2api32w32b_3ort1o0w32bt2o0w32b: BUFF*161 C2*128 OR3*32
// tko64m32_1api0w32b_2api32w32b_3xort1o0w32bt2o0w32b: BUFF*129 C2*128 OR2*64
// tko64m33_1api0w32b_2api32w32b_3nm1b0_4apt1o0w32bt3o0w1b_5nm1b0_6apt2o0w32bt5o0w1b_7addt4o0w33bt6o0w33b: AO222*64 BUFF*266 C2*5 C3*287 GND*2 INV*64 NAND2*64 NOR3*64 OR2*66 OR3*1
// tko66m34_1api0w33b_2api33w33b_3nm1b0_4apt1o0w33bt3o0w1b_5nm1b0_6apt2o0w33bt5o0w1b_7addt4o0w34bt6o0w34b: AO222*66 BUFF*273 C2*5 C3*296 GND*2 INV*66 NAND2*66 NOR3*66 OR2*68 OR3*1
// tkr: NOR2*3
// tks11_o0w11_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0_20o0w0_40o0w0_80o0w0_100o0w0_200o0w0_400o0w0: BUFF*34 C2*36 C3*48 INV*1 NAND3*1 NOR2*1 NOR3*3 OR2*12
// tks1_o0w1_0o0w0_1o0w0: BUFF*7 C2*3 OR2*2
// tks1_o0w1_1o0w0_0o0w0: BUFF*7 C2*3 OR2*2
// tks2_o0w2_0c2o0w0_1o0w0_3o0w0: BUFF*7 C2*7 OR2*2 OR3*1
// tks2_o0w2_1o0w0_2o0w0: BUFF*4 C2*6 OR2*3
// tks2_o0w2_1o0w0_2o0w0_3o0w0_0o0w0: BUFF*8 C2*10 INV*1 NAND2*1 NOR3*1 OR2*2
// tks34_o32w2_1o0w32_2o0w32: BUFF*4 C2*134 C3*16 OR2*35
// tks35_o32w3_0o0w32_1o0w32_2o0w32_3o0w32_4o0w32_5o0w32_6o0w32_7o0w32: BUFF*9 C2*523 C3*24 NAND3*1 NOR2*1 NOR3*2 OR2*35
// tks35_o32w3_1o0w32_2o0w32_3o0w32_4o0w32_5o0w32_6o0w32_7o0w32: BUFF*8 C2*458 C3*23 INV*1 NAND3*1 NOR3*2 OR2*35
// tks35_o32w3_1o0w32_2o0w32_4o0w32: BUFF*4 C2*198 C3*19 OR2*35 OR3*1
// tks3_o0w3_0c4m1m2m3c4o0w0_5m6o0w0: BUFF*2 C2*5 C3*5 INV*1 NAND2*1 NOR3*1 OR2*5
// tks3_o0w3_0m1c6m6o0w0_2o0w0_4o0w0: BUFF*6 C2*4 C3*5 OR2*3 OR3*2
// tks3_o0w3_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0: BUFF*16 C2*9 C3*9 NAND3*1 NOR2*1 NOR3*2 OR2*3
// tks3_o0w3_1c6m2c4m4o0w0_0o0w0: BUFF*4 C2*4 C3*3 OR2*4 OR3*1
// tks3_o0w3_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0: BUFF*14 C2*8 C3*8 INV*1 NAND3*1 NOR3*2 OR2*3
// tks3_o0w3_1o0w0_2o0w0_4o0w0: BUFF*6 C2*4 C3*4 OR2*3 OR3*1
// tks3_o0w3_7o0w0_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0: BUFF*16 C2*9 C3*9 NAND3*1 NOR2*1 NOR3*2 OR2*3
// tks4_o0w4_0m8o0w0_1m9o0w0_2mao0w0_3mbo0w0_4mco0w0_5mdo0w0_6meo0w0_7mfo0w0: BUFF*25 C2*26 C3*17 NAND3*1 NOR2*1 NOR3*2 OR2*12
// tks4_o0w4_1o0w0_2o0w0_4o0w0_8o0w0: BUFF*13 C2*10 C3*5 INV*1 NAND2*1 NOR3*1 OR2*4
// tks5_o0w5_0o0w0_1m2c1m4c3o0w0_8c7o0w0_10c7o0w0_18c7o0w0: BUFF*10 C2*16 C3*5 NAND2*1 NOR2*1 NOR3*1 OR2*5 OR3*1
// tks5_o0w5_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0: BUFF*10 C2*18 C3*6 NAND2*1 NOR2*1 NOR3*1 OR2*5
// tks6_o0w6_0c30m1c3em2c3cm24m28m2cm34m38m3co0w0_4m14o0w0_8m18o0w0_cm1co0w0: BUFF*6 C2*20 C3*27 INV*1 NAND2*1 NAND3*1 NOR3*4 OR2*9
// tks6_o0w6_0c38m1c3em2c3cm24m2cm34m3co0w0_4mcm14m1co0w0: BUFF*3 C2*13 C3*19 INV*2 NAND2*1 NAND3*1 NOR3*3 OR2*7
// tks6_o0w6_0c3cm1c38m2c38m3c38m5m6m7mdc30mec30mfc30m15c20m16c20m17c20o0w0_25m26m27o0w0: BUFF*5 C2*20 C3*23 INV*1 NAND2*1 NAND3*1 NOR3*4 OR2*8 OR3*1
// tks6_o0w6_4c20m9c30mac30mbc30mdc30mec30mfc30m20m21m22m23m28m2cm30m31m32m33m34m35m36m37m38m3co0w0_0m8mcm10m14m18m1co0w0_1m5m11m15o0w0_2m6m12m16o0w0_3m7m13m17o0w0_25o0w0_26o0w0_27o0w0: BUFF*17 C2*56 C3*85 INV*4 NAND2*4 NAND3*4 NOR2*2 NOR3*14 OR2*6 OR3*1
// tks6_o0w6_8c30mbc30mcc30mdc30mec30mfc30m10c20m11c20m12c20m13c20m14c20m15c20m16c20m17c20m19c20m1ac20m20m21m22m23m24m25m26m27m29m2ao0w0_0o0w0_1o0w0_2o0w0_3o0w0_4o0w0_5o0w0_6o0w0_7o0w0_9o0w0_ao0w0: BUFF*27 C2*59 C3*58 INV*1 NAND3*4 NOR2*2 NOR3*11 OR2*7 OR3*1
// tks6_o0w6_9c30mac30mbc30mdc30mec30mfc30m20m21m22m23m24m28m2cm30m31m32m33m34m35m36m37m38m3co0w0_0m1m2m3m4m5m6m7m8mcm10m11m12m13m14m15m16m17m18m1cm25m26m27o0w0: BUFF*8 C2*50 C3*88 NAND2*2 NAND3*4 NOR2*2 NOR3*14 OR2*7 OR3*2
// tks7_o0w7_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0_20o0w0_40o0w0: BUFF*22 C2*8 C3*24 INV*1 NAND3*1 NOR3*2 OR2*7
// tks7_o4w3_1o0w4_2o0w4_4o0w4: BUFF*4 C2*28 C3*6 OR2*7 OR3*1
// tks8_o0w8_1o0w0_2o0w0_4o0w0_8o0w0_10o0w0_20o0w0_40o0w0_80o0w0: BUFF*16 C2*18 C3*27 NAND3*1 NOR2*1 NOR3*2 OR2*8
// tkvaddCarryIn1_wo0w1_ro0w1o0w1: AND2*9 AO22*2 BUFF*8 C2*1 INV*2 NAND2*1 NOR2*2 NOR3*2 OR2*1
// tkvaddResult33_wo0w33_ro0w33: AND2*231 AO22*34 BUFF*105 C2*3 C3*31 INV*1 NOR2*34 NOR3*33 OR2*34
// tkvaluResult32_wo0w32_ro0w32: AND2*224 AO22*33 BUFF*101 C2*5 C3*29 INV*1 NOR2*33 NOR3*32 OR2*33
// tkvcwp1_wo0w1_ro0w1: AND2*7 AO22*2 BUFF*7 C2*1 INV*1 NOR2*2 NOR3*1 OR2*2
// tkvdaccess3_wo0w3_ro0w3o0w1: AND2*23 AO22*4 BUFF*14 C2*1 C3*2 INV*2 NAND2*1 NOR2*4 NOR3*4 OR2*3
// tkvdaddr32_wo0w32_ro0w32: AND2*224 AO22*33 BUFF*101 C2*5 C3*29 INV*1 NOR2*33 NOR3*32 OR2*33
// tkvdistanceI5_wo0w5_ro0w1o1w1o2w1o3w1o4w1: AND2*35 AO22*6 BUFF*22 C2*3 C3*3 INV*3 NAND3*1 NOR2*6 NOR3*8 OR2*6
// tkvdoFetch1_wo0w1_ro0w1: AND2*7 AO22*2 BUFF*7 C2*1 INV*1 NOR2*2 NOR3*1 OR2*2
// tkvdoFetchI1_wo0w1_ro0w1: AND2*7 AO22*2 BUFF*7 C2*1 INV*1 NOR2*2 NOR3*1 OR2*2
// tkvdread32_wo0w32_ro0w32: AND2*224 AO22*33 BUFF*101 C2*5 C3*29 INV*1 NOR2*33 NOR3*32 OR2*33
// tkvdwrite32_wo0w32_ro0w32: AND2*224 AO22*33 BUFF*101 C2*5 C3*29 INV*1 NOR2*33 NOR3*32 OR2*33
// tkvfaddr32_wo0w32_ro0w32: AND2*224 AO22*33 BUFF*101 C2*5 C3*29 INV*1 NOR2*33 NOR3*32 OR2*33
// tkvfinst32_wo0w32_ro0w32: AND2*224 AO22*33 BUFF*101 C2*5 C3*29 INV*1 NOR2*33 NOR3*32 OR2*33
// tkvflags4_wo0w4_ro2w1o1w1o3w1o0w1o3w1o2w1o1w1o2w1o1w1o0w1o0w1o3w1: AND2*44 AO22*5 BUFF*27 C2*3 C3*2 INV*1 NAND2*1 NAND3*2 NOR2*5 NOR3*12 OR2*4 OR3*1
// tkvglobals_1279632_wo0w32_ro0w32o0w32o0w32: AND2*352 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvglobals_15912832_wo0w32_ro0w32o0w32o0w32: AND2*352 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvglobals_19116032_wo0w32_ro0w32o0w32o0w32: AND2*352 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvglobals_22319232_wo0w32_ro0w32o0w32o0w32: AND2*352 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvglobals_31032_wo0w32_ro0w32o0w32o0w32: AND2*352 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvglobals_633232_wo0w32_ro0w32o0w32o0w32: AND2*352 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvglobals_956432_wo0w32_ro0w32o0w32o0w32: AND2*352 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvi32_wo0w32_ro0w32o0w16o16w16o16w16: AND2*320 AO22*33 BUFF*104 C2*5 C3*29 INV*1 NAND3*1 NOR2*34 NOR3*34 OR2*32
// tkvi32_wo0w32_ro0w32o0w24o8w24o8w24: AND2*368 AO22*33 BUFF*104 C2*5 C3*29 INV*1 NAND3*1 NOR2*34 NOR3*34 OR2*32
// tkvi32_wo0w32_ro0w32o0w28o4w28o4w28: AND2*392 AO22*33 BUFF*104 C2*5 C3*29 INV*1 NAND3*1 NOR2*34 NOR3*34 OR2*32
// tkvi32_wo0w32_ro0w32o0w30o2w30o2w30: AND2*404 AO22*33 BUFF*104 C2*5 C3*29 INV*1 NAND3*1 NOR2*34 NOR3*34 OR2*32
// tkvi32_wo0w32_ro0w32o0w31o1w31o1w31: AND2*410 AO22*33 BUFF*104 C2*5 C3*29 INV*1 NAND3*1 NOR2*34 NOR3*34 OR2*32
// tkvimmOrReg1_wo0w1_ro0w1: AND2*7 AO22*2 BUFF*7 C2*1 INV*1 NOR2*2 NOR3*1 OR2*2
// tkvinouts_1279632_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32: AND2*544 AO22*33 BUFF*106 C2*5 C3*29 INV*2 NAND3*1 NOR2*33 NOR3*36 OR2*33
// tkvinouts_15912832_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32: AND2*544 AO22*33 BUFF*106 C2*5 C3*29 INV*2 NAND3*1 NOR2*33 NOR3*36 OR2*33
// tkvinouts_19116032_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32: AND2*544 AO22*33 BUFF*106 C2*5 C3*29 INV*2 NAND3*1 NOR2*33 NOR3*36 OR2*33
// tkvinouts_22319232_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32: AND2*544 AO22*33 BUFF*106 C2*5 C3*29 INV*2 NAND3*1 NOR2*33 NOR3*36 OR2*33
// tkvinouts_25522432_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32: AND2*544 AO22*33 BUFF*106 C2*5 C3*29 INV*2 NAND3*1 NOR2*33 NOR3*36 OR2*33
// tkvinouts_31032_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32: AND2*544 AO22*33 BUFF*106 C2*5 C3*29 INV*2 NAND3*1 NOR2*33 NOR3*36 OR2*33
// tkvinouts_633232_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32: AND2*544 AO22*33 BUFF*106 C2*5 C3*29 INV*2 NAND3*1 NOR2*33 NOR3*36 OR2*33
// tkvinouts_956432_wo0w32_ro0w32o0w32o0w32o0w32o0w32o0w32: AND2*544 AO22*33 BUFF*106 C2*5 C3*29 INV*2 NAND3*1 NOR2*33 NOR3*36 OR2*33
// tkvinstKind3_wo0w3_ro0w3o0w3o0w3: AND2*33 AO22*4 BUFF*15 C2*1 C3*2 INV*1 NAND2*1 NOR2*4 NOR3*5 OR2*3
// tkvir65_wo0w65_ro0w22o25w5o0w22o25w4o22w3o19w6o13w1o0w13o19w6o25w5o25w5o0w5o14w5o13w1o13w1o0w13o19w6o25w5o0w5o14w5o13w1o19w6o30w2o32w33: AND2*685 AO22*66 BUFF*223 C2*3 C3*63 INV*2 NAND2*1 NAND3*5 NOR2*66 NOR3*83 OR2*65
// tkvlhs32_wo0w32_ro0w32o0w32o0w32o0w32o0w32o31w1: AND2*482 AO22*33 BUFF*106 C2*5 C3*29 INV*2 NAND3*1 NOR2*33 NOR3*36 OR2*33
// tkvlocals_1279632_wo0w32_ro0w32o0w32o0w32: AND2*352 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvlocals_15912832_wo0w32_ro0w32o0w32o0w32: AND2*352 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvlocals_19116032_wo0w32_ro0w32o0w32o0w32: AND2*352 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvlocals_22319232_wo0w32_ro0w32o0w32o0w32: AND2*352 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvlocals_25522432_wo0w32_ro0w32o0w32o0w32: AND2*352 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvlocals_31032_wo0w32_ro0w32o0w32o0w32: AND2*352 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvlocals_633232_wo0w32_ro0w32o0w32o0w32: AND2*352 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvlocals_956432_wo0w32_ro0w32o0w32o0w32: AND2*352 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvlogicResult32_wo0w32_ro0w32: AND2*224 AO22*33 BUFF*101 C2*5 C3*29 INV*1 NOR2*33 NOR3*32 OR2*33
// tkvmemAccess4_wo0w4_ro0w4: AND2*28 AO22*5 BUFF*16 C2*3 C3*2 INV*1 NOR2*5 NOR3*4 OR2*5
// tkvmergedResult33_wo0w33_ro0w32o0w32o31w1o32w1o31w1o32w1: AND2*301 AO22*34 BUFF*110 C2*3 C3*31 INV*2 NAND3*1 NOR2*34 NOR3*37 OR2*34
// tkvmread32_wo0w32_ro0w32: AND2*224 AO22*33 BUFF*101 C2*5 C3*29 INV*1 NOR2*33 NOR3*32 OR2*33
// tkvnewPc32_wo0w32_ro0w32: AND2*224 AO22*33 BUFF*101 C2*5 C3*29 INV*1 NOR2*33 NOR3*32 OR2*33
// tkvnewStream1_wo0w1_ro0w1: AND2*7 AO22*2 BUFF*7 C2*1 INV*1 NOR2*2 NOR3*1 OR2*2
// tkvop7_wo0w7_ro0w6o0w6o6w1o6w1o0w6o0w6o0w6: AND2*99 AO22*8 BUFF*31 C2*1 C3*6 INV*1 NAND2*1 NAND3*1 NOR2*9 NOR3*11 OR2*8
// tkvopr74_wo0w74_ro26w5o25w1o25w1o20w5o9w1o15w5o8w1o10w5o7w1o7w3o38w32o37w1o71w2o71w2o25w1o31w6o38w32o6w1o3w4o0w3: AND2*594 AO22*75 BUFF*246 C2*1 C3*73 INV*2 NAND2*2 NAND3*4 NOR2*76 NOR3*88 OR2*74
// tkvpc32_wo0w32_ro0w32o0w32o0w32: AND2*352 AO22*33 BUFF*103 C2*5 C3*29 INV*1 NAND2*1 NOR2*33 NOR3*34 OR2*32
// tkvpcTemp32_wo0w32_ro0w32: AND2*224 AO22*33 BUFF*101 C2*5 C3*29 INV*1 NOR2*33 NOR3*32 OR2*33
// tkvpcr33_wo0w33_ro0w32o32w1: AND2*231 AO22*34 BUFF*106 C2*3 C3*31 INV*2 NAND2*1 NOR2*34 NOR3*34 OR2*33
// tkvpostRhs32_wo0w32_ro0w32o31w1o0w5o31w1: AND2*238 AO22*33 BUFF*104 C2*5 C3*29 INV*1 NAND3*1 NOR2*34 NOR3*34 OR2*32
// tkvpreCarry1_wo0w1_ro0w1o0w1o0w1: AND2*11 AO22*2 BUFF*9 C2*1 INV*1 NAND2*1 NOR2*2 NOR3*3 OR2*1
// tkvr032_wo0w32_ro0w32: AND2*224 AO22*33 BUFF*101 C2*5 C3*29 INV*1 NOR2*33 NOR3*32 OR2*33
// tkvr132_wo0w32_ro0w32: AND2*224 AO22*33 BUFF*101 C2*5 C3*29 INV*1 NOR2*33 NOR3*32 OR2*33
// tkvr232_wo0w32_ro0w32: AND2*224 AO22*33 BUFF*101 C2*5 C3*29 INV*1 NOR2*33 NOR3*32 OR2*33
// tkvrEn3_wo0w3_ro0w1o1w1o2w1: AND2*21 AO22*4 BUFF*15 C2*1 C3*2 INV*1 NAND2*1 NOR2*4 NOR3*5 OR2*3
// tkvrhs32_wo0w32_ro0w32o0w32o0w32o0w32o0w32: AND2*480 AO22*33 BUFF*105 C2*5 C3*29 INV*3 NAND3*1 NOR2*33 NOR3*35 OR2*33
// tkvsel5_wo0w5_ro0w5o0w3o0w3o0w3o0w3: AND2*59 AO22*6 BUFF*22 C2*3 C3*3 INV*3 NAND3*1 NOR2*6 NOR3*8 OR2*6
// tkvshift2_wo0w2_ro0w2o0w2o0w2o0w2o0w2: AND2*30 AO22*3 BUFF*13 C2*1 C3*1 INV*3 NAND3*1 NOR2*3 NOR3*5 OR2*3
// tkvshiftResult32_wo0w32_ro0w32: AND2*224 AO22*33 BUFF*101 C2*5 C3*29 INV*1 NOR2*33 NOR3*32 OR2*33
// tkvstore1_wo0w1_ro0w1o0w1: AND2*9 AO22*2 BUFF*8 C2*1 INV*2 NAND2*1 NOR2*2 NOR3*2 OR2*1
// tkvtake1_wo0w1_ro0w1: AND2*7 AO22*2 BUFF*7 C2*1 INV*1 NOR2*2 NOR3*1 OR2*2
// tkvtakeBranch1_wo0w1_ro0w1o0w1: AND2*9 AO22*2 BUFF*8 C2*1 INV*2 NAND2*1 NOR2*2 NOR3*2 OR2*1
// tkvtakeBranch21_wo0w1_ro0w1: AND2*7 AO22*2 BUFF*7 C2*1 INV*1 NOR2*2 NOR3*1 OR2*2
// tkvv1_wo0w1_ro0w1: AND2*7 AO22*2 BUFF*7 C2*1 INV*1 NOR2*2 NOR3*1 OR2*2
// tkvv32_wo0w32_ro0w32: AND2*224 AO22*33 BUFF*101 C2*5 C3*29 INV*1 NOR2*33 NOR3*32 OR2*33
// tkvv33_wo0w33_ro0w33: AND2*231 AO22*34 BUFF*105 C2*3 C3*31 INV*1 NOR2*34 NOR3*33 OR2*34
// tkvv65_wo0w65_ro0w65: AND2*455 AO22*66 BUFF*200 C2*3 C3*63 INV*1 NOR2*66 NOR3*65 OR2*66
// tkvv74_wo0w74_ro0w74: AND2*518 AO22*75 BUFF*227 C2*1 C3*73 INV*1 NOR2*75 NOR3*74 OR2*75
// tkvw32_wo0w32_ro0w32o0w32o0w32o0w32: AND2*416 AO22*33 BUFF*104 C2*5 C3*29 INV*1 NAND3*1 NOR2*34 NOR3*34 OR2*32
// tkvwEn1_wo0w1_ro0w1: AND2*7 AO22*2 BUFF*7 C2*1 INV*1 NOR2*2 NOR3*1 OR2*2
// tkvwindow1_wo0w1_ro0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1o0w1: AND2*29 AO22*2 BUFF*18 C2*1 INV*1 NAND2*1 NAND3*2 NOR2*2 NOR3*9 OR2*1 OR3*1
